module real_aes_2833_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_185;
wire n_285;
wire n_624;
wire n_800;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_822;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_792;
wire n_386;
wire n_635;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_817;
wire n_443;
wire n_565;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_449;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_756;
wire n_735;
wire n_713;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_765;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_809;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_798;
wire n_797;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_SL g565 ( .A(n_0), .B(n_510), .Y(n_565) );
AOI21xp5_ASAP7_75t_L g511 ( .A1(n_1), .A2(n_512), .B(n_513), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g817 ( .A(n_2), .B(n_818), .Y(n_817) );
AOI22xp5_ASAP7_75t_L g123 ( .A1(n_3), .A2(n_4), .B1(n_124), .B2(n_125), .Y(n_123) );
CKINVDCx20_ASAP7_75t_R g125 ( .A(n_3), .Y(n_125) );
CKINVDCx20_ASAP7_75t_R g124 ( .A(n_4), .Y(n_124) );
NAND2xp5_ASAP7_75t_SL g547 ( .A(n_5), .B(n_228), .Y(n_547) );
INVx1_ASAP7_75t_L g160 ( .A(n_6), .Y(n_160) );
NAND2xp5_ASAP7_75t_SL g216 ( .A(n_7), .B(n_217), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_8), .B(n_228), .Y(n_596) );
INVx1_ASAP7_75t_L g198 ( .A(n_9), .Y(n_198) );
CKINVDCx16_ASAP7_75t_R g818 ( .A(n_10), .Y(n_818) );
CKINVDCx5p33_ASAP7_75t_R g166 ( .A(n_11), .Y(n_166) );
NAND2xp33_ASAP7_75t_L g588 ( .A(n_12), .B(n_225), .Y(n_588) );
INVx2_ASAP7_75t_L g142 ( .A(n_13), .Y(n_142) );
OAI22xp5_ASAP7_75t_SL g121 ( .A1(n_14), .A2(n_122), .B1(n_123), .B2(n_126), .Y(n_121) );
CKINVDCx20_ASAP7_75t_R g126 ( .A(n_14), .Y(n_126) );
AOI221x1_ASAP7_75t_L g532 ( .A1(n_15), .A2(n_29), .B1(n_510), .B2(n_512), .C(n_533), .Y(n_532) );
CKINVDCx16_ASAP7_75t_R g499 ( .A(n_16), .Y(n_499) );
NOR3xp33_ASAP7_75t_L g816 ( .A(n_16), .B(n_817), .C(n_819), .Y(n_816) );
NAND2xp5_ASAP7_75t_SL g584 ( .A(n_17), .B(n_510), .Y(n_584) );
AOI22xp5_ASAP7_75t_SL g119 ( .A1(n_18), .A2(n_120), .B1(n_121), .B2(n_127), .Y(n_119) );
CKINVDCx20_ASAP7_75t_R g127 ( .A(n_18), .Y(n_127) );
INVx1_ASAP7_75t_L g226 ( .A(n_19), .Y(n_226) );
AO21x2_ASAP7_75t_L g582 ( .A1(n_20), .A2(n_195), .B(n_583), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_21), .B(n_190), .Y(n_536) );
OAI22xp5_ASAP7_75t_L g806 ( .A1(n_22), .A2(n_83), .B1(n_807), .B2(n_808), .Y(n_806) );
INVx1_ASAP7_75t_L g807 ( .A(n_22), .Y(n_807) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_23), .B(n_228), .Y(n_521) );
AO21x1_ASAP7_75t_L g542 ( .A1(n_24), .A2(n_510), .B(n_543), .Y(n_542) );
INVx1_ASAP7_75t_L g116 ( .A(n_25), .Y(n_116) );
INVx1_ASAP7_75t_L g223 ( .A(n_26), .Y(n_223) );
INVx1_ASAP7_75t_SL g210 ( .A(n_27), .Y(n_210) );
NAND2xp5_ASAP7_75t_SL g268 ( .A(n_28), .B(n_153), .Y(n_268) );
AOI33xp33_ASAP7_75t_L g248 ( .A1(n_30), .A2(n_55), .A3(n_146), .B1(n_171), .B2(n_249), .B3(n_250), .Y(n_248) );
NAND2x1_ASAP7_75t_L g563 ( .A(n_31), .B(n_228), .Y(n_563) );
NAND2x1_ASAP7_75t_L g595 ( .A(n_32), .B(n_225), .Y(n_595) );
INVx1_ASAP7_75t_L g151 ( .A(n_33), .Y(n_151) );
OA21x2_ASAP7_75t_L g141 ( .A1(n_34), .A2(n_90), .B(n_142), .Y(n_141) );
OR2x2_ASAP7_75t_L g192 ( .A(n_34), .B(n_90), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_35), .B(n_175), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_36), .B(n_225), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_37), .B(n_228), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_38), .B(n_225), .Y(n_546) );
AOI21xp5_ASAP7_75t_L g552 ( .A1(n_39), .A2(n_512), .B(n_553), .Y(n_552) );
AND2x2_ASAP7_75t_L g159 ( .A(n_40), .B(n_160), .Y(n_159) );
INVx1_ASAP7_75t_L g170 ( .A(n_40), .Y(n_170) );
AND2x2_ASAP7_75t_L g179 ( .A(n_40), .B(n_149), .Y(n_179) );
OR2x6_ASAP7_75t_L g114 ( .A(n_41), .B(n_115), .Y(n_114) );
INVxp67_ASAP7_75t_L g819 ( .A(n_41), .Y(n_819) );
CKINVDCx20_ASAP7_75t_R g161 ( .A(n_42), .Y(n_161) );
NAND2xp5_ASAP7_75t_SL g556 ( .A(n_43), .B(n_510), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_44), .B(n_175), .Y(n_183) );
AOI22xp5_ASAP7_75t_L g261 ( .A1(n_45), .A2(n_140), .B1(n_217), .B2(n_262), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_46), .B(n_270), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_47), .B(n_153), .Y(n_211) );
CKINVDCx20_ASAP7_75t_R g525 ( .A(n_48), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_49), .B(n_225), .Y(n_554) );
NAND2xp5_ASAP7_75t_SL g200 ( .A(n_50), .B(n_195), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_51), .B(n_153), .Y(n_199) );
AOI21xp5_ASAP7_75t_L g593 ( .A1(n_52), .A2(n_512), .B(n_594), .Y(n_593) );
CKINVDCx5p33_ASAP7_75t_R g265 ( .A(n_53), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_54), .B(n_225), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_56), .B(n_153), .Y(n_187) );
INVx1_ASAP7_75t_L g147 ( .A(n_57), .Y(n_147) );
INVx1_ASAP7_75t_L g155 ( .A(n_57), .Y(n_155) );
AND2x2_ASAP7_75t_L g189 ( .A(n_58), .B(n_190), .Y(n_189) );
AOI221xp5_ASAP7_75t_L g196 ( .A1(n_59), .A2(n_78), .B1(n_168), .B2(n_175), .C(n_197), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_60), .B(n_175), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_61), .B(n_228), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_62), .B(n_140), .Y(n_173) );
AOI21xp5_ASAP7_75t_SL g235 ( .A1(n_63), .A2(n_168), .B(n_236), .Y(n_235) );
AOI21xp5_ASAP7_75t_L g561 ( .A1(n_64), .A2(n_512), .B(n_562), .Y(n_561) );
CKINVDCx20_ASAP7_75t_R g794 ( .A(n_65), .Y(n_794) );
INVx1_ASAP7_75t_L g220 ( .A(n_66), .Y(n_220) );
AO21x1_ASAP7_75t_L g544 ( .A1(n_67), .A2(n_512), .B(n_545), .Y(n_544) );
NAND2xp5_ASAP7_75t_SL g509 ( .A(n_68), .B(n_510), .Y(n_509) );
INVx1_ASAP7_75t_L g186 ( .A(n_69), .Y(n_186) );
XOR2xp5_ASAP7_75t_L g803 ( .A(n_70), .B(n_86), .Y(n_803) );
NAND2xp5_ASAP7_75t_SL g597 ( .A(n_71), .B(n_510), .Y(n_597) );
AOI21xp5_ASAP7_75t_L g184 ( .A1(n_72), .A2(n_168), .B(n_185), .Y(n_184) );
AND2x2_ASAP7_75t_L g557 ( .A(n_73), .B(n_191), .Y(n_557) );
INVx1_ASAP7_75t_L g149 ( .A(n_74), .Y(n_149) );
INVx1_ASAP7_75t_L g157 ( .A(n_74), .Y(n_157) );
AND2x2_ASAP7_75t_L g598 ( .A(n_75), .B(n_139), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_76), .B(n_175), .Y(n_251) );
CKINVDCx20_ASAP7_75t_R g821 ( .A(n_77), .Y(n_821) );
AND2x2_ASAP7_75t_L g212 ( .A(n_79), .B(n_139), .Y(n_212) );
INVx1_ASAP7_75t_L g221 ( .A(n_80), .Y(n_221) );
AOI21xp5_ASAP7_75t_L g208 ( .A1(n_81), .A2(n_168), .B(n_209), .Y(n_208) );
A2O1A1Ixp33_ASAP7_75t_L g266 ( .A1(n_82), .A2(n_168), .B(n_243), .C(n_267), .Y(n_266) );
INVx1_ASAP7_75t_L g808 ( .A(n_83), .Y(n_808) );
INVx1_ASAP7_75t_L g117 ( .A(n_84), .Y(n_117) );
AND2x2_ASAP7_75t_L g507 ( .A(n_85), .B(n_139), .Y(n_507) );
AND2x2_ASAP7_75t_SL g233 ( .A(n_86), .B(n_139), .Y(n_233) );
NAND2xp5_ASAP7_75t_SL g523 ( .A(n_87), .B(n_510), .Y(n_523) );
AOI22xp5_ASAP7_75t_L g245 ( .A1(n_88), .A2(n_168), .B1(n_246), .B2(n_247), .Y(n_245) );
AND2x2_ASAP7_75t_L g543 ( .A(n_89), .B(n_217), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_91), .B(n_225), .Y(n_522) );
AND2x2_ASAP7_75t_L g566 ( .A(n_92), .B(n_139), .Y(n_566) );
INVx1_ASAP7_75t_L g237 ( .A(n_93), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_94), .B(n_228), .Y(n_555) );
AOI21xp5_ASAP7_75t_L g519 ( .A1(n_95), .A2(n_512), .B(n_520), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_96), .B(n_225), .Y(n_534) );
AND2x2_ASAP7_75t_L g252 ( .A(n_97), .B(n_139), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g809 ( .A(n_98), .B(n_810), .Y(n_809) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_99), .B(n_228), .Y(n_514) );
A2O1A1Ixp33_ASAP7_75t_L g143 ( .A1(n_100), .A2(n_144), .B(n_150), .C(n_158), .Y(n_143) );
BUFx2_ASAP7_75t_L g111 ( .A(n_101), .Y(n_111) );
AOI21xp5_ASAP7_75t_L g585 ( .A1(n_102), .A2(n_512), .B(n_586), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_103), .B(n_153), .Y(n_238) );
AOI21xp33_ASAP7_75t_L g104 ( .A1(n_105), .A2(n_812), .B(n_820), .Y(n_104) );
AO21x2_ASAP7_75t_L g105 ( .A1(n_106), .A2(n_112), .B(n_797), .Y(n_105) );
HB1xp67_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g107 ( .A(n_108), .Y(n_107) );
BUFx3_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
CKINVDCx20_ASAP7_75t_R g109 ( .A(n_110), .Y(n_109) );
HB1xp67_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
NOR2x1_ASAP7_75t_R g799 ( .A(n_111), .B(n_800), .Y(n_799) );
OAI22xp5_ASAP7_75t_L g112 ( .A1(n_113), .A2(n_118), .B1(n_794), .B2(n_795), .Y(n_112) );
NAND2xp5_ASAP7_75t_L g801 ( .A(n_113), .B(n_499), .Y(n_801) );
CKINVDCx5p33_ASAP7_75t_R g113 ( .A(n_114), .Y(n_113) );
OR2x2_ASAP7_75t_L g796 ( .A(n_114), .B(n_499), .Y(n_796) );
INVx1_ASAP7_75t_L g815 ( .A(n_115), .Y(n_815) );
NAND2xp5_ASAP7_75t_L g115 ( .A(n_116), .B(n_117), .Y(n_115) );
XOR2xp5_ASAP7_75t_L g118 ( .A(n_119), .B(n_128), .Y(n_118) );
INVxp33_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
INVx1_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
OAI22xp5_ASAP7_75t_L g128 ( .A1(n_129), .A2(n_497), .B1(n_498), .B2(n_500), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
NAND3x1_ASAP7_75t_L g130 ( .A(n_131), .B(n_376), .C(n_443), .Y(n_130) );
AND2x2_ASAP7_75t_L g131 ( .A(n_132), .B(n_336), .Y(n_131) );
NOR3x1_ASAP7_75t_L g132 ( .A(n_133), .B(n_287), .C(n_316), .Y(n_132) );
OAI221xp5_ASAP7_75t_L g133 ( .A1(n_134), .A2(n_201), .B1(n_240), .B2(n_255), .C(n_272), .Y(n_133) );
A2O1A1Ixp33_ASAP7_75t_SL g450 ( .A1(n_134), .A2(n_214), .B(n_451), .C(n_452), .Y(n_450) );
INVx1_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
AOI22xp5_ASAP7_75t_L g421 ( .A1(n_135), .A2(n_422), .B1(n_425), .B2(n_427), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_135), .B(n_241), .Y(n_496) );
AND2x2_ASAP7_75t_L g135 ( .A(n_136), .B(n_180), .Y(n_135) );
BUFx2_ASAP7_75t_L g415 ( .A(n_136), .Y(n_415) );
INVx1_ASAP7_75t_SL g428 ( .A(n_136), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_136), .B(n_283), .Y(n_470) );
INVx1_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
AND2x4_ASAP7_75t_L g253 ( .A(n_137), .B(n_254), .Y(n_253) );
AND2x2_ASAP7_75t_L g298 ( .A(n_137), .B(n_194), .Y(n_298) );
INVx1_ASAP7_75t_L g309 ( .A(n_137), .Y(n_309) );
INVx2_ASAP7_75t_L g313 ( .A(n_137), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_137), .B(n_284), .Y(n_440) );
OR2x2_ASAP7_75t_L g137 ( .A(n_138), .B(n_163), .Y(n_137) );
OAI22xp5_ASAP7_75t_L g138 ( .A1(n_139), .A2(n_143), .B1(n_161), .B2(n_162), .Y(n_138) );
INVx3_ASAP7_75t_L g162 ( .A(n_139), .Y(n_162) );
INVx4_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_140), .B(n_165), .Y(n_164) );
INVx3_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
BUFx4f_ASAP7_75t_L g195 ( .A(n_141), .Y(n_195) );
AND2x2_ASAP7_75t_SL g191 ( .A(n_142), .B(n_192), .Y(n_191) );
AND2x4_ASAP7_75t_L g217 ( .A(n_142), .B(n_192), .Y(n_217) );
INVxp67_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
O2A1O1Ixp33_ASAP7_75t_L g185 ( .A1(n_145), .A2(n_186), .B(n_187), .C(n_188), .Y(n_185) );
O2A1O1Ixp33_ASAP7_75t_SL g197 ( .A1(n_145), .A2(n_188), .B(n_198), .C(n_199), .Y(n_197) );
O2A1O1Ixp33_ASAP7_75t_SL g209 ( .A1(n_145), .A2(n_188), .B(n_210), .C(n_211), .Y(n_209) );
OAI22xp5_ASAP7_75t_L g219 ( .A1(n_145), .A2(n_152), .B1(n_220), .B2(n_221), .Y(n_219) );
O2A1O1Ixp33_ASAP7_75t_L g236 ( .A1(n_145), .A2(n_188), .B(n_237), .C(n_238), .Y(n_236) );
INVx2_ASAP7_75t_L g270 ( .A(n_145), .Y(n_270) );
OR2x6_ASAP7_75t_L g145 ( .A(n_146), .B(n_148), .Y(n_145) );
AND2x2_ASAP7_75t_L g176 ( .A(n_146), .B(n_177), .Y(n_176) );
INVxp33_ASAP7_75t_L g249 ( .A(n_146), .Y(n_249) );
INVx2_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
AND2x2_ASAP7_75t_L g172 ( .A(n_147), .B(n_160), .Y(n_172) );
AND2x4_ASAP7_75t_L g228 ( .A(n_147), .B(n_156), .Y(n_228) );
INVx3_ASAP7_75t_L g171 ( .A(n_148), .Y(n_171) );
INVx2_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
AND2x6_ASAP7_75t_L g225 ( .A(n_149), .B(n_154), .Y(n_225) );
NOR2xp33_ASAP7_75t_L g150 ( .A(n_151), .B(n_152), .Y(n_150) );
INVx1_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
AND2x4_ASAP7_75t_L g510 ( .A(n_153), .B(n_159), .Y(n_510) );
AND2x4_ASAP7_75t_L g153 ( .A(n_154), .B(n_156), .Y(n_153) );
INVx2_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx2_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
HB1xp67_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
INVx5_ASAP7_75t_L g188 ( .A(n_159), .Y(n_188) );
HB1xp67_ASAP7_75t_L g177 ( .A(n_160), .Y(n_177) );
AO21x2_ASAP7_75t_L g181 ( .A1(n_162), .A2(n_182), .B(n_189), .Y(n_181) );
AO21x2_ASAP7_75t_L g284 ( .A1(n_162), .A2(n_182), .B(n_189), .Y(n_284) );
AO21x2_ASAP7_75t_L g550 ( .A1(n_162), .A2(n_551), .B(n_557), .Y(n_550) );
AO21x2_ASAP7_75t_L g559 ( .A1(n_162), .A2(n_560), .B(n_566), .Y(n_559) );
AO21x2_ASAP7_75t_L g572 ( .A1(n_162), .A2(n_560), .B(n_566), .Y(n_572) );
AO21x2_ASAP7_75t_L g575 ( .A1(n_162), .A2(n_551), .B(n_557), .Y(n_575) );
OAI22xp5_ASAP7_75t_L g163 ( .A1(n_164), .A2(n_167), .B1(n_173), .B2(n_174), .Y(n_163) );
INVx1_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
INVxp67_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
AND2x4_ASAP7_75t_L g168 ( .A(n_169), .B(n_172), .Y(n_168) );
NOR2x1p5_ASAP7_75t_L g169 ( .A(n_170), .B(n_171), .Y(n_169) );
INVx1_ASAP7_75t_L g250 ( .A(n_171), .Y(n_250) );
AND2x6_ASAP7_75t_L g512 ( .A(n_172), .B(n_179), .Y(n_512) );
INVx1_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
AND2x4_ASAP7_75t_L g175 ( .A(n_176), .B(n_178), .Y(n_175) );
INVx1_ASAP7_75t_L g263 ( .A(n_176), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_178), .Y(n_264) );
BUFx3_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
AND2x2_ASAP7_75t_L g389 ( .A(n_180), .B(n_390), .Y(n_389) );
NOR2x1_ASAP7_75t_L g180 ( .A(n_181), .B(n_193), .Y(n_180) );
INVx2_ASAP7_75t_L g292 ( .A(n_181), .Y(n_292) );
AND2x2_ASAP7_75t_L g312 ( .A(n_181), .B(n_313), .Y(n_312) );
NOR2xp67_ASAP7_75t_L g437 ( .A(n_181), .B(n_313), .Y(n_437) );
AND2x2_ASAP7_75t_L g462 ( .A(n_181), .B(n_305), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_183), .B(n_184), .Y(n_182) );
NOR2xp33_ASAP7_75t_L g229 ( .A(n_188), .B(n_217), .Y(n_229) );
INVx1_ASAP7_75t_L g246 ( .A(n_188), .Y(n_246) );
AOI21xp5_ASAP7_75t_L g267 ( .A1(n_188), .A2(n_268), .B(n_269), .Y(n_267) );
AOI21xp5_ASAP7_75t_L g513 ( .A1(n_188), .A2(n_514), .B(n_515), .Y(n_513) );
AOI21xp5_ASAP7_75t_L g520 ( .A1(n_188), .A2(n_521), .B(n_522), .Y(n_520) );
AOI21xp5_ASAP7_75t_L g533 ( .A1(n_188), .A2(n_534), .B(n_535), .Y(n_533) );
AOI21xp5_ASAP7_75t_L g545 ( .A1(n_188), .A2(n_546), .B(n_547), .Y(n_545) );
AOI21xp5_ASAP7_75t_L g553 ( .A1(n_188), .A2(n_554), .B(n_555), .Y(n_553) );
AOI21xp5_ASAP7_75t_L g562 ( .A1(n_188), .A2(n_563), .B(n_564), .Y(n_562) );
AOI21xp5_ASAP7_75t_L g586 ( .A1(n_188), .A2(n_587), .B(n_588), .Y(n_586) );
AOI21xp5_ASAP7_75t_L g594 ( .A1(n_188), .A2(n_595), .B(n_596), .Y(n_594) );
CKINVDCx5p33_ASAP7_75t_R g205 ( .A(n_190), .Y(n_205) );
AOI21xp5_ASAP7_75t_L g508 ( .A1(n_190), .A2(n_509), .B(n_511), .Y(n_508) );
OA21x2_ASAP7_75t_L g531 ( .A1(n_190), .A2(n_532), .B(n_536), .Y(n_531) );
OA21x2_ASAP7_75t_L g602 ( .A1(n_190), .A2(n_532), .B(n_536), .Y(n_602) );
BUFx6f_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
INVx1_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
INVx2_ASAP7_75t_L g254 ( .A(n_194), .Y(n_254) );
INVx1_ASAP7_75t_L g276 ( .A(n_194), .Y(n_276) );
INVxp67_ASAP7_75t_L g315 ( .A(n_194), .Y(n_315) );
AND2x4_ASAP7_75t_L g355 ( .A(n_194), .B(n_356), .Y(n_355) );
HB1xp67_ASAP7_75t_L g410 ( .A(n_194), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_194), .B(n_306), .Y(n_441) );
OA21x2_ASAP7_75t_L g194 ( .A1(n_195), .A2(n_196), .B(n_200), .Y(n_194) );
INVx2_ASAP7_75t_SL g243 ( .A(n_195), .Y(n_243) );
INVx1_ASAP7_75t_SL g201 ( .A(n_202), .Y(n_201) );
AND2x2_ASAP7_75t_L g202 ( .A(n_203), .B(n_213), .Y(n_202) );
AND2x2_ASAP7_75t_L g329 ( .A(n_203), .B(n_301), .Y(n_329) );
INVx1_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
HB1xp67_ASAP7_75t_L g257 ( .A(n_204), .Y(n_257) );
AND2x2_ASAP7_75t_L g285 ( .A(n_204), .B(n_286), .Y(n_285) );
INVx2_ASAP7_75t_L g296 ( .A(n_204), .Y(n_296) );
INVx1_ASAP7_75t_L g320 ( .A(n_204), .Y(n_320) );
AND2x2_ASAP7_75t_L g323 ( .A(n_204), .B(n_215), .Y(n_323) );
HB1xp67_ASAP7_75t_L g345 ( .A(n_204), .Y(n_345) );
AO21x2_ASAP7_75t_L g204 ( .A1(n_205), .A2(n_206), .B(n_212), .Y(n_204) );
AO21x2_ASAP7_75t_L g591 ( .A1(n_205), .A2(n_592), .B(n_598), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_207), .B(n_208), .Y(n_206) );
NOR2x1_ASAP7_75t_L g213 ( .A(n_214), .B(n_230), .Y(n_213) );
AND2x2_ASAP7_75t_L g310 ( .A(n_214), .B(n_232), .Y(n_310) );
NAND2x1_ASAP7_75t_L g343 ( .A(n_214), .B(n_344), .Y(n_343) );
INVx1_ASAP7_75t_L g446 ( .A(n_214), .Y(n_446) );
INVx2_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
INVx3_ASAP7_75t_L g286 ( .A(n_215), .Y(n_286) );
AND2x2_ASAP7_75t_L g301 ( .A(n_215), .B(n_260), .Y(n_301) );
NOR2x1_ASAP7_75t_SL g370 ( .A(n_215), .B(n_232), .Y(n_370) );
AND2x4_ASAP7_75t_L g215 ( .A(n_216), .B(n_218), .Y(n_215) );
AOI21xp5_ASAP7_75t_L g234 ( .A1(n_217), .A2(n_235), .B(n_239), .Y(n_234) );
INVx1_ASAP7_75t_SL g517 ( .A(n_217), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_217), .B(n_549), .Y(n_548) );
AOI21xp5_ASAP7_75t_L g583 ( .A1(n_217), .A2(n_584), .B(n_585), .Y(n_583) );
OAI21xp5_ASAP7_75t_L g218 ( .A1(n_219), .A2(n_222), .B(n_229), .Y(n_218) );
OAI22xp5_ASAP7_75t_L g222 ( .A1(n_223), .A2(n_224), .B1(n_226), .B2(n_227), .Y(n_222) );
INVxp67_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
INVxp67_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
NOR2x1_ASAP7_75t_L g407 ( .A(n_230), .B(n_394), .Y(n_407) );
INVx1_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
AND2x2_ASAP7_75t_L g332 ( .A(n_231), .B(n_333), .Y(n_332) );
INVx2_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
INVx4_ASAP7_75t_L g271 ( .A(n_232), .Y(n_271) );
AND2x4_ASAP7_75t_L g278 ( .A(n_232), .B(n_279), .Y(n_278) );
BUFx6f_ASAP7_75t_L g302 ( .A(n_232), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_232), .B(n_295), .Y(n_395) );
AND2x2_ASAP7_75t_L g423 ( .A(n_232), .B(n_260), .Y(n_423) );
OR2x6_ASAP7_75t_L g232 ( .A(n_233), .B(n_234), .Y(n_232) );
NAND2x1_ASAP7_75t_SL g240 ( .A(n_241), .B(n_253), .Y(n_240) );
OR2x2_ASAP7_75t_L g451 ( .A(n_241), .B(n_363), .Y(n_451) );
INVx1_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
AND2x4_ASAP7_75t_L g291 ( .A(n_242), .B(n_292), .Y(n_291) );
INVx2_ASAP7_75t_L g356 ( .A(n_242), .Y(n_356) );
AND2x2_ASAP7_75t_L g390 ( .A(n_242), .B(n_313), .Y(n_390) );
AO21x2_ASAP7_75t_L g242 ( .A1(n_243), .A2(n_244), .B(n_252), .Y(n_242) );
AO21x2_ASAP7_75t_L g306 ( .A1(n_243), .A2(n_244), .B(n_252), .Y(n_306) );
NAND2xp5_ASAP7_75t_SL g244 ( .A(n_245), .B(n_251), .Y(n_244) );
INVx1_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
INVx3_ASAP7_75t_L g363 ( .A(n_253), .Y(n_363) );
AND2x2_ASAP7_75t_L g371 ( .A(n_253), .B(n_304), .Y(n_371) );
AND2x2_ASAP7_75t_L g488 ( .A(n_253), .B(n_291), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_256), .B(n_258), .Y(n_255) );
BUFx2_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
AND2x2_ASAP7_75t_L g442 ( .A(n_257), .B(n_383), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_257), .B(n_282), .Y(n_477) );
AOI21xp5_ASAP7_75t_L g318 ( .A1(n_258), .A2(n_319), .B(n_322), .Y(n_318) );
AND2x2_ASAP7_75t_L g388 ( .A(n_258), .B(n_294), .Y(n_388) );
INVx2_ASAP7_75t_SL g475 ( .A(n_258), .Y(n_475) );
AND2x4_ASAP7_75t_SL g258 ( .A(n_259), .B(n_271), .Y(n_258) );
HB1xp67_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
INVx1_ASAP7_75t_L g279 ( .A(n_260), .Y(n_279) );
INVx2_ASAP7_75t_L g326 ( .A(n_260), .Y(n_326) );
AND2x4_ASAP7_75t_L g333 ( .A(n_260), .B(n_286), .Y(n_333) );
AND2x2_ASAP7_75t_L g260 ( .A(n_261), .B(n_266), .Y(n_260) );
NOR3xp33_ASAP7_75t_L g262 ( .A(n_263), .B(n_264), .C(n_265), .Y(n_262) );
HB1xp67_ASAP7_75t_L g289 ( .A(n_271), .Y(n_289) );
AND2x4_ASAP7_75t_L g365 ( .A(n_271), .B(n_279), .Y(n_365) );
OR2x2_ASAP7_75t_L g491 ( .A(n_271), .B(n_492), .Y(n_491) );
NAND4xp25_ASAP7_75t_L g272 ( .A(n_273), .B(n_277), .C(n_280), .D(n_285), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
OR2x2_ASAP7_75t_L g338 ( .A(n_274), .B(n_339), .Y(n_338) );
INVx2_ASAP7_75t_L g435 ( .A(n_274), .Y(n_435) );
INVx3_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
NAND2x1p5_ASAP7_75t_L g335 ( .A(n_275), .B(n_283), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_275), .B(n_340), .Y(n_469) );
BUFx3_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
HB1xp67_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_278), .B(n_294), .Y(n_347) );
INVx2_ASAP7_75t_L g449 ( .A(n_278), .Y(n_449) );
AND2x2_ASAP7_75t_SL g459 ( .A(n_278), .B(n_319), .Y(n_459) );
NOR2xp33_ASAP7_75t_L g484 ( .A(n_278), .B(n_485), .Y(n_484) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
AND2x2_ASAP7_75t_L g351 ( .A(n_282), .B(n_298), .Y(n_351) );
AND2x2_ASAP7_75t_L g419 ( .A(n_282), .B(n_355), .Y(n_419) );
INVx3_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
AND2x4_ASAP7_75t_L g304 ( .A(n_283), .B(n_305), .Y(n_304) );
INVx3_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
HB1xp67_ASAP7_75t_L g358 ( .A(n_284), .Y(n_358) );
AND2x2_ASAP7_75t_L g409 ( .A(n_284), .B(n_410), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_284), .B(n_306), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_285), .B(n_449), .Y(n_456) );
INVx1_ASAP7_75t_SL g492 ( .A(n_285), .Y(n_492) );
INVx1_ASAP7_75t_L g321 ( .A(n_286), .Y(n_321) );
AND2x2_ASAP7_75t_L g383 ( .A(n_286), .B(n_326), .Y(n_383) );
OAI21xp5_ASAP7_75t_L g287 ( .A1(n_288), .A2(n_297), .B(n_299), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_289), .B(n_290), .Y(n_288) );
AND2x2_ASAP7_75t_L g290 ( .A(n_291), .B(n_293), .Y(n_290) );
AND2x2_ASAP7_75t_L g349 ( .A(n_291), .B(n_298), .Y(n_349) );
AND2x2_ASAP7_75t_L g457 ( .A(n_291), .B(n_308), .Y(n_457) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
INVx1_ASAP7_75t_L g331 ( .A(n_294), .Y(n_331) );
AND2x2_ASAP7_75t_L g364 ( .A(n_294), .B(n_365), .Y(n_364) );
AND2x2_ASAP7_75t_L g369 ( .A(n_294), .B(n_370), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_294), .B(n_333), .Y(n_418) );
NOR3xp33_ASAP7_75t_L g468 ( .A(n_294), .B(n_469), .C(n_470), .Y(n_468) );
INVx3_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
INVx2_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
INVxp67_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
AOI22xp33_ASAP7_75t_L g299 ( .A1(n_300), .A2(n_303), .B1(n_310), .B2(n_311), .Y(n_299) );
AND2x2_ASAP7_75t_L g300 ( .A(n_301), .B(n_302), .Y(n_300) );
INVx2_ASAP7_75t_L g394 ( .A(n_301), .Y(n_394) );
AND2x2_ASAP7_75t_L g328 ( .A(n_302), .B(n_329), .Y(n_328) );
AND2x2_ASAP7_75t_L g350 ( .A(n_302), .B(n_323), .Y(n_350) );
AND2x2_ASAP7_75t_SL g382 ( .A(n_302), .B(n_383), .Y(n_382) );
AND2x2_ASAP7_75t_L g303 ( .A(n_304), .B(n_307), .Y(n_303) );
INVx1_ASAP7_75t_L g361 ( .A(n_304), .Y(n_361) );
AND2x2_ASAP7_75t_L g314 ( .A(n_305), .B(n_315), .Y(n_314) );
INVx1_ASAP7_75t_L g340 ( .A(n_305), .Y(n_340) );
INVx2_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
INVx2_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
AND2x2_ASAP7_75t_L g403 ( .A(n_309), .B(n_355), .Y(n_403) );
INVx1_ASAP7_75t_L g461 ( .A(n_309), .Y(n_461) );
INVx1_ASAP7_75t_L g317 ( .A(n_311), .Y(n_317) );
AND2x2_ASAP7_75t_L g311 ( .A(n_312), .B(n_314), .Y(n_311) );
NAND2x1p5_ASAP7_75t_L g339 ( .A(n_312), .B(n_340), .Y(n_339) );
AND2x2_ASAP7_75t_L g448 ( .A(n_312), .B(n_355), .Y(n_448) );
AND2x2_ASAP7_75t_L g414 ( .A(n_314), .B(n_415), .Y(n_414) );
NAND2x1p5_ASAP7_75t_L g482 ( .A(n_314), .B(n_483), .Y(n_482) );
OAI21xp5_ASAP7_75t_L g316 ( .A1(n_317), .A2(n_318), .B(n_327), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_319), .B(n_354), .Y(n_353) );
AND2x4_ASAP7_75t_L g375 ( .A(n_319), .B(n_324), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_319), .B(n_365), .Y(n_426) );
AND2x4_ASAP7_75t_SL g319 ( .A(n_320), .B(n_321), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_320), .B(n_383), .Y(n_413) );
HB1xp67_ASAP7_75t_L g433 ( .A(n_320), .Y(n_433) );
AOI22xp5_ASAP7_75t_L g348 ( .A1(n_322), .A2(n_349), .B1(n_350), .B2(n_351), .Y(n_348) );
AND2x2_ASAP7_75t_SL g322 ( .A(n_323), .B(n_324), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_323), .B(n_365), .Y(n_384) );
INVx1_ASAP7_75t_L g485 ( .A(n_323), .Y(n_485) );
INVx2_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
OAI21xp5_ASAP7_75t_L g327 ( .A1(n_328), .A2(n_330), .B(n_334), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_329), .B(n_488), .Y(n_487) );
AND2x2_ASAP7_75t_L g330 ( .A(n_331), .B(n_332), .Y(n_330) );
INVx1_ASAP7_75t_L g466 ( .A(n_332), .Y(n_466) );
INVx4_ASAP7_75t_L g368 ( .A(n_333), .Y(n_368) );
INVxp33_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
OR2x2_ASAP7_75t_L g396 ( .A(n_335), .B(n_397), .Y(n_396) );
NOR2x1_ASAP7_75t_L g336 ( .A(n_337), .B(n_352), .Y(n_336) );
OAI21xp5_ASAP7_75t_L g337 ( .A1(n_338), .A2(n_341), .B(n_348), .Y(n_337) );
INVx1_ASAP7_75t_L g386 ( .A(n_339), .Y(n_386) );
NOR2xp33_ASAP7_75t_L g341 ( .A(n_342), .B(n_346), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
INVx1_ASAP7_75t_L g391 ( .A(n_343), .Y(n_391) );
INVx1_ASAP7_75t_L g424 ( .A(n_344), .Y(n_424) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
AOI22xp5_ASAP7_75t_L g387 ( .A1(n_349), .A2(n_388), .B1(n_389), .B2(n_391), .Y(n_387) );
INVx1_ASAP7_75t_L g401 ( .A(n_350), .Y(n_401) );
NAND4xp25_ASAP7_75t_SL g352 ( .A(n_353), .B(n_359), .C(n_366), .D(n_372), .Y(n_352) );
AND2x2_ASAP7_75t_L g354 ( .A(n_355), .B(n_357), .Y(n_354) );
INVx1_ASAP7_75t_L g374 ( .A(n_355), .Y(n_374) );
AND2x2_ASAP7_75t_L g486 ( .A(n_355), .B(n_483), .Y(n_486) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_360), .B(n_364), .Y(n_359) );
NOR2xp33_ASAP7_75t_L g360 ( .A(n_361), .B(n_362), .Y(n_360) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
OR2x2_ASAP7_75t_L g493 ( .A(n_363), .B(n_430), .Y(n_493) );
INVx1_ASAP7_75t_L g490 ( .A(n_364), .Y(n_490) );
HB1xp67_ASAP7_75t_L g399 ( .A(n_365), .Y(n_399) );
OAI21xp5_ASAP7_75t_L g366 ( .A1(n_367), .A2(n_369), .B(n_371), .Y(n_366) );
INVx2_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_373), .B(n_375), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
AND2x2_ASAP7_75t_L g376 ( .A(n_377), .B(n_404), .Y(n_376) );
NOR3xp33_ASAP7_75t_L g377 ( .A(n_378), .B(n_392), .C(n_400), .Y(n_377) );
OAI21xp5_ASAP7_75t_L g378 ( .A1(n_379), .A2(n_385), .B(n_387), .Y(n_378) );
INVxp67_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_381), .B(n_384), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
AOI22xp5_ASAP7_75t_L g416 ( .A1(n_382), .A2(n_414), .B1(n_417), .B2(n_419), .Y(n_416) );
OAI22xp33_ASAP7_75t_L g392 ( .A1(n_385), .A2(n_393), .B1(n_396), .B2(n_398), .Y(n_392) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g397 ( .A(n_390), .Y(n_397) );
AND2x4_ASAP7_75t_L g408 ( .A(n_390), .B(n_409), .Y(n_408) );
OR2x2_ASAP7_75t_L g393 ( .A(n_394), .B(n_395), .Y(n_393) );
HB1xp67_ASAP7_75t_L g495 ( .A(n_395), .Y(n_495) );
AOI31xp33_ASAP7_75t_L g494 ( .A1(n_398), .A2(n_471), .A3(n_495), .B(n_496), .Y(n_494) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
NOR2xp33_ASAP7_75t_L g400 ( .A(n_401), .B(n_402), .Y(n_400) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
NOR2xp33_ASAP7_75t_L g404 ( .A(n_405), .B(n_420), .Y(n_404) );
NAND2xp5_ASAP7_75t_SL g405 ( .A(n_406), .B(n_416), .Y(n_405) );
AOI22xp5_ASAP7_75t_L g406 ( .A1(n_407), .A2(n_408), .B1(n_411), .B2(n_414), .Y(n_406) );
HB1xp67_ASAP7_75t_L g474 ( .A(n_410), .Y(n_474) );
INVx2_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
BUFx2_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_418), .B(n_466), .Y(n_465) );
NAND2xp5_ASAP7_75t_SL g420 ( .A(n_421), .B(n_431), .Y(n_420) );
AND2x2_ASAP7_75t_L g422 ( .A(n_423), .B(n_424), .Y(n_422) );
AND2x2_ASAP7_75t_L g432 ( .A(n_423), .B(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g471 ( .A(n_423), .Y(n_471) );
AOI22xp33_ASAP7_75t_SL g480 ( .A1(n_423), .A2(n_481), .B1(n_484), .B2(n_486), .Y(n_480) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
AND2x2_ASAP7_75t_L g427 ( .A(n_428), .B(n_429), .Y(n_427) );
NOR2xp33_ASAP7_75t_L g476 ( .A(n_428), .B(n_477), .Y(n_476) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
AOI22xp5_ASAP7_75t_L g431 ( .A1(n_432), .A2(n_434), .B1(n_438), .B2(n_442), .Y(n_431) );
NOR2xp33_ASAP7_75t_SL g434 ( .A(n_435), .B(n_436), .Y(n_434) );
INVxp67_ASAP7_75t_SL g436 ( .A(n_437), .Y(n_436) );
INVx1_ASAP7_75t_SL g438 ( .A(n_439), .Y(n_438) );
OR2x2_ASAP7_75t_L g439 ( .A(n_440), .B(n_441), .Y(n_439) );
INVx2_ASAP7_75t_SL g483 ( .A(n_440), .Y(n_483) );
INVx2_ASAP7_75t_L g464 ( .A(n_441), .Y(n_464) );
AND2x2_ASAP7_75t_L g443 ( .A(n_444), .B(n_478), .Y(n_443) );
AOI211xp5_ASAP7_75t_L g444 ( .A1(n_445), .A2(n_450), .B(n_453), .C(n_467), .Y(n_444) );
OAI21xp33_ASAP7_75t_L g445 ( .A1(n_446), .A2(n_447), .B(n_449), .Y(n_445) );
INVx1_ASAP7_75t_SL g447 ( .A(n_448), .Y(n_447) );
INVx1_ASAP7_75t_L g452 ( .A(n_449), .Y(n_452) );
NAND2xp5_ASAP7_75t_SL g453 ( .A(n_454), .B(n_458), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_455), .B(n_457), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
AOI22xp5_ASAP7_75t_L g458 ( .A1(n_459), .A2(n_460), .B1(n_463), .B2(n_465), .Y(n_458) );
AND2x2_ASAP7_75t_L g460 ( .A(n_461), .B(n_462), .Y(n_460) );
AND2x2_ASAP7_75t_L g463 ( .A(n_461), .B(n_464), .Y(n_463) );
AO22x1_ASAP7_75t_L g467 ( .A1(n_468), .A2(n_471), .B1(n_472), .B2(n_476), .Y(n_467) );
NOR2xp33_ASAP7_75t_L g472 ( .A(n_473), .B(n_475), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
NOR3xp33_ASAP7_75t_L g478 ( .A(n_479), .B(n_489), .C(n_494), .Y(n_478) );
NAND2xp5_ASAP7_75t_SL g479 ( .A(n_480), .B(n_487), .Y(n_479) );
INVx3_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
AOI21xp33_ASAP7_75t_R g489 ( .A1(n_490), .A2(n_491), .B(n_493), .Y(n_489) );
CKINVDCx5p33_ASAP7_75t_R g497 ( .A(n_498), .Y(n_497) );
CKINVDCx16_ASAP7_75t_R g498 ( .A(n_499), .Y(n_498) );
INVx3_ASAP7_75t_SL g805 ( .A(n_500), .Y(n_805) );
NOR2x2_ASAP7_75t_L g500 ( .A(n_501), .B(n_681), .Y(n_500) );
AO211x2_ASAP7_75t_L g501 ( .A1(n_502), .A2(n_526), .B(n_576), .C(n_649), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
INVxp67_ASAP7_75t_SL g503 ( .A(n_504), .Y(n_503) );
AND3x2_ASAP7_75t_L g730 ( .A(n_504), .B(n_611), .C(n_627), .Y(n_730) );
AND2x4_ASAP7_75t_L g733 ( .A(n_504), .B(n_734), .Y(n_733) );
AND2x2_ASAP7_75t_L g504 ( .A(n_505), .B(n_516), .Y(n_504) );
NAND2x1p5_ASAP7_75t_L g589 ( .A(n_505), .B(n_590), .Y(n_589) );
INVx4_ASAP7_75t_L g642 ( .A(n_505), .Y(n_642) );
AND2x2_ASAP7_75t_SL g727 ( .A(n_505), .B(n_636), .Y(n_727) );
AND2x2_ASAP7_75t_L g770 ( .A(n_505), .B(n_591), .Y(n_770) );
INVx5_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
BUFx2_ASAP7_75t_L g619 ( .A(n_506), .Y(n_619) );
AND2x2_ASAP7_75t_L g638 ( .A(n_506), .B(n_582), .Y(n_638) );
AND2x2_ASAP7_75t_L g656 ( .A(n_506), .B(n_591), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_506), .B(n_590), .Y(n_716) );
NOR2x1_ASAP7_75t_SL g743 ( .A(n_506), .B(n_516), .Y(n_743) );
OR2x6_ASAP7_75t_L g506 ( .A(n_507), .B(n_508), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_516), .B(n_582), .Y(n_581) );
AO21x2_ASAP7_75t_L g516 ( .A1(n_517), .A2(n_518), .B(n_524), .Y(n_516) );
NOR2xp33_ASAP7_75t_L g524 ( .A(n_517), .B(n_525), .Y(n_524) );
AO21x2_ASAP7_75t_L g615 ( .A1(n_517), .A2(n_518), .B(n_524), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_519), .B(n_523), .Y(n_518) );
AO21x1_ASAP7_75t_L g526 ( .A1(n_527), .A2(n_558), .B(n_567), .Y(n_526) );
INVx2_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
OAI22xp33_ASAP7_75t_L g624 ( .A1(n_528), .A2(n_625), .B1(n_629), .B2(n_630), .Y(n_624) );
OR2x2_ASAP7_75t_L g528 ( .A(n_529), .B(n_537), .Y(n_528) );
AND2x2_ASAP7_75t_L g685 ( .A(n_529), .B(n_573), .Y(n_685) );
BUFx2_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
AND2x4_ASAP7_75t_L g618 ( .A(n_530), .B(n_601), .Y(n_618) );
AND2x2_ASAP7_75t_L g690 ( .A(n_530), .B(n_575), .Y(n_690) );
AND2x2_ASAP7_75t_L g709 ( .A(n_530), .B(n_675), .Y(n_709) );
INVx2_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
INVx2_ASAP7_75t_L g568 ( .A(n_531), .Y(n_568) );
HB1xp67_ASAP7_75t_L g696 ( .A(n_531), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_537), .B(n_679), .Y(n_678) );
INVx2_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
AND2x2_ASAP7_75t_L g669 ( .A(n_538), .B(n_570), .Y(n_669) );
AND2x4_ASAP7_75t_L g538 ( .A(n_539), .B(n_550), .Y(n_538) );
AND2x2_ASAP7_75t_L g573 ( .A(n_539), .B(n_574), .Y(n_573) );
OR2x2_ASAP7_75t_L g606 ( .A(n_539), .B(n_607), .Y(n_606) );
AND2x2_ASAP7_75t_SL g666 ( .A(n_539), .B(n_602), .Y(n_666) );
INVx2_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
BUFx2_ASAP7_75t_L g759 ( .A(n_540), .Y(n_759) );
INVx2_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
INVx2_ASAP7_75t_L g601 ( .A(n_541), .Y(n_601) );
OAI21x1_ASAP7_75t_SL g541 ( .A1(n_542), .A2(n_544), .B(n_548), .Y(n_541) );
INVx1_ASAP7_75t_L g549 ( .A(n_543), .Y(n_549) );
INVx2_ASAP7_75t_L g607 ( .A(n_550), .Y(n_607) );
HB1xp67_ASAP7_75t_L g707 ( .A(n_550), .Y(n_707) );
NAND2xp5_ASAP7_75t_SL g551 ( .A(n_552), .B(n_556), .Y(n_551) );
INVx2_ASAP7_75t_L g603 ( .A(n_558), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g761 ( .A(n_558), .B(n_735), .Y(n_761) );
AND2x2_ASAP7_75t_L g780 ( .A(n_558), .B(n_770), .Y(n_780) );
BUFx2_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
AND2x4_ASAP7_75t_SL g648 ( .A(n_559), .B(n_607), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_561), .B(n_565), .Y(n_560) );
AND2x2_ASAP7_75t_SL g567 ( .A(n_568), .B(n_569), .Y(n_567) );
AND2x2_ASAP7_75t_L g647 ( .A(n_568), .B(n_648), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_568), .B(n_617), .Y(n_652) );
INVx1_ASAP7_75t_SL g779 ( .A(n_568), .Y(n_779) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_569), .B(n_730), .Y(n_729) );
AND2x2_ASAP7_75t_L g569 ( .A(n_570), .B(n_573), .Y(n_569) );
INVx1_ASAP7_75t_L g605 ( .A(n_570), .Y(n_605) );
AND2x2_ASAP7_75t_L g791 ( .A(n_570), .B(n_792), .Y(n_791) );
BUFx2_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
AND2x2_ASAP7_75t_L g667 ( .A(n_571), .B(n_574), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_571), .B(n_680), .Y(n_679) );
AND2x2_ASAP7_75t_L g721 ( .A(n_571), .B(n_575), .Y(n_721) );
AND2x2_ASAP7_75t_L g752 ( .A(n_571), .B(n_753), .Y(n_752) );
INVx2_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
AND2x2_ASAP7_75t_L g617 ( .A(n_572), .B(n_575), .Y(n_617) );
INVxp67_ASAP7_75t_L g634 ( .A(n_572), .Y(n_634) );
BUFx3_ASAP7_75t_L g675 ( .A(n_572), .Y(n_675) );
AND2x2_ASAP7_75t_L g695 ( .A(n_573), .B(n_696), .Y(n_695) );
NAND2xp33_ASAP7_75t_L g708 ( .A(n_573), .B(n_709), .Y(n_708) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_574), .B(n_601), .Y(n_664) );
AND2x2_ASAP7_75t_L g753 ( .A(n_574), .B(n_602), .Y(n_753) );
INVx2_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
AND2x2_ASAP7_75t_L g680 ( .A(n_575), .B(n_602), .Y(n_680) );
OR3x1_ASAP7_75t_L g576 ( .A(n_577), .B(n_624), .C(n_639), .Y(n_576) );
OAI321xp33_ASAP7_75t_L g577 ( .A1(n_578), .A2(n_589), .A3(n_599), .B1(n_604), .B2(n_608), .C(n_616), .Y(n_577) );
INVx1_ASAP7_75t_SL g578 ( .A(n_579), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
INVxp67_ASAP7_75t_SL g655 ( .A(n_581), .Y(n_655) );
INVxp67_ASAP7_75t_SL g673 ( .A(n_581), .Y(n_673) );
OR2x2_ASAP7_75t_L g677 ( .A(n_581), .B(n_589), .Y(n_677) );
BUFx3_ASAP7_75t_L g611 ( .A(n_582), .Y(n_611) );
AND2x2_ASAP7_75t_L g628 ( .A(n_582), .B(n_614), .Y(n_628) );
INVx1_ASAP7_75t_L g645 ( .A(n_582), .Y(n_645) );
INVx2_ASAP7_75t_L g661 ( .A(n_582), .Y(n_661) );
OR2x2_ASAP7_75t_L g700 ( .A(n_582), .B(n_590), .Y(n_700) );
INVx2_ASAP7_75t_L g688 ( .A(n_589), .Y(n_688) );
AND2x2_ASAP7_75t_L g612 ( .A(n_590), .B(n_613), .Y(n_612) );
INVx2_ASAP7_75t_L g627 ( .A(n_590), .Y(n_627) );
AND2x4_ASAP7_75t_L g636 ( .A(n_590), .B(n_637), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_590), .B(n_613), .Y(n_659) );
AND2x2_ASAP7_75t_L g766 ( .A(n_590), .B(n_661), .Y(n_766) );
INVx4_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
HB1xp67_ASAP7_75t_L g725 ( .A(n_591), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_593), .B(n_597), .Y(n_592) );
INVx1_ASAP7_75t_L g653 ( .A(n_599), .Y(n_653) );
NAND2xp5_ASAP7_75t_SL g599 ( .A(n_600), .B(n_603), .Y(n_599) );
AND2x2_ASAP7_75t_L g740 ( .A(n_600), .B(n_667), .Y(n_740) );
INVx1_ASAP7_75t_SL g757 ( .A(n_600), .Y(n_757) );
NAND2xp5_ASAP7_75t_L g786 ( .A(n_600), .B(n_733), .Y(n_786) );
AND2x4_ASAP7_75t_L g600 ( .A(n_601), .B(n_602), .Y(n_600) );
OR2x2_ASAP7_75t_L g629 ( .A(n_601), .B(n_602), .Y(n_629) );
AND2x2_ASAP7_75t_L g722 ( .A(n_603), .B(n_618), .Y(n_722) );
OR2x2_ASAP7_75t_L g604 ( .A(n_605), .B(n_606), .Y(n_604) );
NAND2xp5_ASAP7_75t_SL g745 ( .A(n_607), .B(n_618), .Y(n_745) );
INVx2_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
AOI22xp33_ASAP7_75t_L g762 ( .A1(n_609), .A2(n_758), .B1(n_763), .B2(n_765), .Y(n_762) );
AND2x4_ASAP7_75t_L g609 ( .A(n_610), .B(n_612), .Y(n_609) );
AND2x2_ASAP7_75t_L g687 ( .A(n_610), .B(n_688), .Y(n_687) );
OR2x2_ASAP7_75t_L g782 ( .A(n_610), .B(n_783), .Y(n_782) );
INVx2_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
AND2x2_ASAP7_75t_L g738 ( .A(n_611), .B(n_656), .Y(n_738) );
AND2x4_ASAP7_75t_L g692 ( .A(n_612), .B(n_638), .Y(n_692) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
HB1xp67_ASAP7_75t_L g790 ( .A(n_614), .Y(n_790) );
INVx2_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
INVx1_ASAP7_75t_L g623 ( .A(n_615), .Y(n_623) );
INVx1_ASAP7_75t_L g637 ( .A(n_615), .Y(n_637) );
NAND4xp25_ASAP7_75t_L g616 ( .A(n_617), .B(n_618), .C(n_619), .D(n_620), .Y(n_616) );
AND2x2_ASAP7_75t_L g774 ( .A(n_617), .B(n_759), .Y(n_774) );
NAND2xp5_ASAP7_75t_L g784 ( .A(n_617), .B(n_785), .Y(n_784) );
NOR2xp33_ASAP7_75t_L g693 ( .A(n_618), .B(n_694), .Y(n_693) );
OAI322xp33_ASAP7_75t_L g701 ( .A1(n_618), .A2(n_702), .A3(n_706), .B1(n_708), .B2(n_710), .C1(n_712), .C2(n_717), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_618), .B(n_667), .Y(n_717) );
INVx1_ASAP7_75t_L g785 ( .A(n_618), .Y(n_785) );
INVx2_ASAP7_75t_L g631 ( .A(n_619), .Y(n_631) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
INVx2_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_622), .B(n_725), .Y(n_724) );
INVx2_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_623), .B(n_642), .Y(n_699) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_626), .B(n_669), .Y(n_668) );
AND2x2_ASAP7_75t_L g626 ( .A(n_627), .B(n_628), .Y(n_626) );
INVx1_ASAP7_75t_L g672 ( .A(n_627), .Y(n_672) );
AND2x2_ASAP7_75t_L g744 ( .A(n_627), .B(n_655), .Y(n_744) );
AOI31xp33_ASAP7_75t_L g630 ( .A1(n_628), .A2(n_631), .A3(n_632), .B(n_635), .Y(n_630) );
AND2x2_ASAP7_75t_L g641 ( .A(n_628), .B(n_642), .Y(n_641) );
AND2x2_ASAP7_75t_L g769 ( .A(n_628), .B(n_770), .Y(n_769) );
AND2x2_ASAP7_75t_SL g776 ( .A(n_628), .B(n_656), .Y(n_776) );
INVx1_ASAP7_75t_L g777 ( .A(n_628), .Y(n_777) );
INVx1_ASAP7_75t_SL g735 ( .A(n_629), .Y(n_735) );
NAND3xp33_ASAP7_75t_SL g763 ( .A(n_629), .B(n_757), .C(n_764), .Y(n_763) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
OR2x2_ASAP7_75t_L g663 ( .A(n_634), .B(n_664), .Y(n_663) );
AND2x2_ASAP7_75t_L g635 ( .A(n_636), .B(n_638), .Y(n_635) );
AND2x2_ASAP7_75t_L g644 ( .A(n_636), .B(n_645), .Y(n_644) );
INVx2_ASAP7_75t_L g705 ( .A(n_636), .Y(n_705) );
AOI322xp5_ASAP7_75t_L g787 ( .A1(n_636), .A2(n_666), .A3(n_669), .B1(n_788), .B2(n_789), .C1(n_791), .C2(n_793), .Y(n_787) );
AND2x2_ASAP7_75t_L g793 ( .A(n_636), .B(n_642), .Y(n_793) );
AOI21xp5_ASAP7_75t_L g639 ( .A1(n_640), .A2(n_643), .B(n_646), .Y(n_639) );
INVx1_ASAP7_75t_SL g640 ( .A(n_641), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_642), .B(n_661), .Y(n_660) );
AND2x4_ASAP7_75t_L g788 ( .A(n_642), .B(n_675), .Y(n_788) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
INVx1_ASAP7_75t_L g714 ( .A(n_645), .Y(n_714) );
AND2x2_ASAP7_75t_L g742 ( .A(n_645), .B(n_743), .Y(n_742) );
AND2x2_ASAP7_75t_L g789 ( .A(n_645), .B(n_790), .Y(n_789) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
INVx1_ASAP7_75t_L g694 ( .A(n_648), .Y(n_694) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
O2A1O1Ixp5_ASAP7_75t_L g650 ( .A1(n_651), .A2(n_653), .B(n_654), .C(n_657), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
AND2x2_ASAP7_75t_L g654 ( .A(n_655), .B(n_656), .Y(n_654) );
AND2x2_ASAP7_75t_L g711 ( .A(n_656), .B(n_661), .Y(n_711) );
OAI211xp5_ASAP7_75t_L g657 ( .A1(n_658), .A2(n_662), .B(n_668), .C(n_670), .Y(n_657) );
OAI221xp5_ASAP7_75t_L g683 ( .A1(n_658), .A2(n_684), .B1(n_686), .B2(n_689), .C(n_691), .Y(n_683) );
OR2x2_ASAP7_75t_L g658 ( .A(n_659), .B(n_660), .Y(n_658) );
INVx1_ASAP7_75t_L g703 ( .A(n_660), .Y(n_703) );
OR2x2_ASAP7_75t_L g723 ( .A(n_660), .B(n_724), .Y(n_723) );
AND2x2_ASAP7_75t_L g662 ( .A(n_663), .B(n_665), .Y(n_662) );
INVx1_ASAP7_75t_L g768 ( .A(n_663), .Y(n_768) );
INVx1_ASAP7_75t_L g792 ( .A(n_664), .Y(n_792) );
NAND2xp5_ASAP7_75t_SL g665 ( .A(n_666), .B(n_667), .Y(n_665) );
AND2x2_ASAP7_75t_L g674 ( .A(n_666), .B(n_675), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g748 ( .A(n_666), .B(n_736), .Y(n_748) );
INVx1_ASAP7_75t_L g728 ( .A(n_667), .Y(n_728) );
AOI22xp5_ASAP7_75t_L g670 ( .A1(n_671), .A2(n_674), .B1(n_676), .B2(n_678), .Y(n_670) );
AND2x2_ASAP7_75t_L g671 ( .A(n_672), .B(n_673), .Y(n_671) );
INVx1_ASAP7_75t_SL g736 ( .A(n_675), .Y(n_736) );
INVx2_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
NAND4xp75_ASAP7_75t_L g681 ( .A(n_682), .B(n_718), .C(n_746), .D(n_771), .Y(n_681) );
NOR2xp67_ASAP7_75t_L g682 ( .A(n_683), .B(n_701), .Y(n_682) );
INVx1_ASAP7_75t_SL g684 ( .A(n_685), .Y(n_684) );
INVx2_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
AND2x2_ASAP7_75t_SL g758 ( .A(n_690), .B(n_759), .Y(n_758) );
AOI22xp5_ASAP7_75t_L g691 ( .A1(n_692), .A2(n_693), .B1(n_695), .B2(n_697), .Y(n_691) );
NOR2xp33_ASAP7_75t_L g756 ( .A(n_694), .B(n_757), .Y(n_756) );
INVx2_ASAP7_75t_SL g697 ( .A(n_698), .Y(n_697) );
OR2x2_ASAP7_75t_L g698 ( .A(n_699), .B(n_700), .Y(n_698) );
INVx2_ASAP7_75t_L g734 ( .A(n_700), .Y(n_734) );
OR2x2_ASAP7_75t_L g749 ( .A(n_700), .B(n_750), .Y(n_749) );
NAND2xp5_ASAP7_75t_SL g702 ( .A(n_703), .B(n_704), .Y(n_702) );
INVx1_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
INVx1_ASAP7_75t_L g764 ( .A(n_709), .Y(n_764) );
INVx1_ASAP7_75t_SL g710 ( .A(n_711), .Y(n_710) );
OAI21xp5_ASAP7_75t_SL g755 ( .A1(n_711), .A2(n_756), .B(n_758), .Y(n_755) );
INVxp67_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
AND2x2_ASAP7_75t_L g713 ( .A(n_714), .B(n_715), .Y(n_713) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
NOR2x1_ASAP7_75t_L g718 ( .A(n_719), .B(n_731), .Y(n_718) );
OAI221xp5_ASAP7_75t_L g719 ( .A1(n_720), .A2(n_723), .B1(n_726), .B2(n_728), .C(n_729), .Y(n_719) );
NOR2xp33_ASAP7_75t_L g720 ( .A(n_721), .B(n_722), .Y(n_720) );
OAI21xp33_ASAP7_75t_L g767 ( .A1(n_721), .A2(n_768), .B(n_769), .Y(n_767) );
INVx3_ASAP7_75t_SL g726 ( .A(n_727), .Y(n_726) );
OAI322xp33_ASAP7_75t_L g731 ( .A1(n_732), .A2(n_735), .A3(n_736), .B1(n_737), .B2(n_739), .C1(n_741), .C2(n_745), .Y(n_731) );
INVx1_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
INVx1_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
INVx1_ASAP7_75t_SL g739 ( .A(n_740), .Y(n_739) );
NOR2x1_ASAP7_75t_L g741 ( .A(n_742), .B(n_744), .Y(n_741) );
INVx1_ASAP7_75t_L g754 ( .A(n_742), .Y(n_754) );
INVx1_ASAP7_75t_L g750 ( .A(n_743), .Y(n_750) );
AND2x2_ASAP7_75t_L g765 ( .A(n_743), .B(n_766), .Y(n_765) );
NOR2x1_ASAP7_75t_L g746 ( .A(n_747), .B(n_760), .Y(n_746) );
OAI221xp5_ASAP7_75t_L g747 ( .A1(n_748), .A2(n_749), .B1(n_751), .B2(n_754), .C(n_755), .Y(n_747) );
INVx1_ASAP7_75t_SL g751 ( .A(n_752), .Y(n_751) );
OAI211xp5_ASAP7_75t_SL g760 ( .A1(n_754), .A2(n_761), .B(n_762), .C(n_767), .Y(n_760) );
INVx2_ASAP7_75t_SL g783 ( .A(n_770), .Y(n_783) );
NOR2x1_ASAP7_75t_L g771 ( .A(n_772), .B(n_781), .Y(n_771) );
OAI22xp33_ASAP7_75t_L g772 ( .A1(n_773), .A2(n_775), .B1(n_777), .B2(n_778), .Y(n_772) );
INVx1_ASAP7_75t_SL g773 ( .A(n_774), .Y(n_773) );
INVx2_ASAP7_75t_SL g775 ( .A(n_776), .Y(n_775) );
NAND2xp5_ASAP7_75t_L g778 ( .A(n_779), .B(n_780), .Y(n_778) );
OAI211xp5_ASAP7_75t_SL g781 ( .A1(n_782), .A2(n_784), .B(n_786), .C(n_787), .Y(n_781) );
BUFx2_ASAP7_75t_L g795 ( .A(n_796), .Y(n_795) );
OAI21xp5_ASAP7_75t_L g797 ( .A1(n_798), .A2(n_802), .B(n_809), .Y(n_797) );
INVx2_ASAP7_75t_L g798 ( .A(n_799), .Y(n_798) );
INVxp67_ASAP7_75t_SL g800 ( .A(n_801), .Y(n_800) );
BUFx2_ASAP7_75t_L g811 ( .A(n_801), .Y(n_811) );
XNOR2xp5_ASAP7_75t_L g802 ( .A(n_803), .B(n_804), .Y(n_802) );
XOR2x2_ASAP7_75t_L g804 ( .A(n_805), .B(n_806), .Y(n_804) );
INVx1_ASAP7_75t_L g810 ( .A(n_811), .Y(n_810) );
INVx3_ASAP7_75t_SL g812 ( .A(n_813), .Y(n_812) );
INVx1_ASAP7_75t_SL g822 ( .A(n_813), .Y(n_822) );
INVx2_ASAP7_75t_SL g813 ( .A(n_814), .Y(n_813) );
AND2x2_ASAP7_75t_SL g814 ( .A(n_815), .B(n_816), .Y(n_814) );
NOR2xp33_ASAP7_75t_L g820 ( .A(n_821), .B(n_822), .Y(n_820) );
endmodule