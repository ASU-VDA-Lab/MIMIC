module real_jpeg_7329_n_13 (n_8, n_0, n_95, n_2, n_10, n_9, n_12, n_97, n_6, n_104, n_100, n_11, n_7, n_3, n_99, n_5, n_4, n_102, n_98, n_101, n_1, n_96, n_103, n_13);

input n_8;
input n_0;
input n_95;
input n_2;
input n_10;
input n_9;
input n_12;
input n_97;
input n_6;
input n_104;
input n_100;
input n_11;
input n_7;
input n_3;
input n_99;
input n_5;
input n_4;
input n_102;
input n_98;
input n_101;
input n_1;
input n_96;
input n_103;

output n_13;

wire n_54;
wire n_37;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_68;
wire n_78;
wire n_83;
wire n_64;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_27;
wire n_56;
wire n_48;
wire n_93;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_45;
wire n_42;
wire n_18;
wire n_77;
wire n_39;
wire n_26;
wire n_19;
wire n_17;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_24;
wire n_92;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_81;
wire n_85;
wire n_89;
wire n_16;

INVx1_ASAP7_75t_L g76 ( 
.A(n_0),
.Y(n_76)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_1),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_1),
.B(n_61),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g16 ( 
.A(n_2),
.B(n_17),
.Y(n_16)
);

AND2x2_ASAP7_75t_L g23 ( 
.A(n_2),
.B(n_17),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_3),
.B(n_38),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_3),
.B(n_38),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_4),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_5),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_6),
.B(n_79),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_6),
.B(n_79),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_7),
.B(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_7),
.B(n_65),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_8),
.B(n_87),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_8),
.B(n_87),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_9),
.B(n_41),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_9),
.B(n_41),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_10),
.B(n_27),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_10),
.B(n_27),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_11),
.B(n_55),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_12),
.Y(n_18)
);

XNOR2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_24),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_SL g14 ( 
.A(n_15),
.B(n_22),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_19),
.Y(n_17)
);

BUFx2_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_21),
.B(n_39),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_21),
.B(n_66),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_85),
.B(n_91),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_32),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_29),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_31),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_31),
.Y(n_90)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

OAI21x1_ASAP7_75t_L g33 ( 
.A1(n_34),
.A2(n_78),
.B(n_84),
.Y(n_33)
);

AOI21xp5_ASAP7_75t_L g34 ( 
.A1(n_35),
.A2(n_72),
.B(n_77),
.Y(n_34)
);

AO221x1_ASAP7_75t_L g35 ( 
.A1(n_36),
.A2(n_44),
.B1(n_69),
.B2(n_70),
.C(n_71),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_40),
.Y(n_36)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_40),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_43),
.Y(n_41)
);

AO21x1_ASAP7_75t_L g44 ( 
.A1(n_45),
.A2(n_52),
.B(n_68),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_46),
.B(n_51),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_46),
.B(n_51),
.Y(n_68)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_49),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_49),
.B(n_75),
.Y(n_74)
);

BUFx12_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

OAI21xp5_ASAP7_75t_SL g52 ( 
.A1(n_53),
.A2(n_64),
.B(n_67),
.Y(n_52)
);

AOI21xp5_ASAP7_75t_L g53 ( 
.A1(n_54),
.A2(n_58),
.B(n_63),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_57),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_59),
.B(n_62),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_59),
.B(n_62),
.Y(n_63)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_73),
.B(n_76),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_73),
.B(n_76),
.Y(n_77)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_81),
.Y(n_79)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g91 ( 
.A1(n_86),
.A2(n_92),
.B(n_93),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_89),
.Y(n_87)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_95),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_96),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_97),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_98),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_99),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_100),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_101),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_102),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_103),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_104),
.Y(n_88)
);


endmodule