module fake_jpeg_8049_n_341 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_341);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_341;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_260;
wire n_199;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_0),
.B(n_3),
.Y(n_21)
);

BUFx4f_ASAP7_75t_SL g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_15),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_14),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_4),
.B(n_1),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_11),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_36),
.Y(n_77)
);

OR2x2_ASAP7_75t_L g37 ( 
.A(n_28),
.B(n_1),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_37),
.B(n_39),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_35),
.Y(n_38)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_21),
.Y(n_39)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_40),
.Y(n_70)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

INVx1_ASAP7_75t_SL g56 ( 
.A(n_41),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

BUFx10_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_21),
.B(n_15),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_43),
.B(n_48),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_28),
.B(n_1),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_45),
.B(n_32),
.Y(n_57)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_46),
.B(n_30),
.Y(n_59)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_23),
.Y(n_47)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_22),
.Y(n_48)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_26),
.Y(n_49)
);

BUFx2_ASAP7_75t_L g78 ( 
.A(n_49),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_34),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_51),
.B(n_54),
.Y(n_105)
);

INVx13_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_52),
.B(n_62),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_49),
.A2(n_30),
.B1(n_32),
.B2(n_18),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_53),
.A2(n_16),
.B1(n_20),
.B2(n_24),
.Y(n_83)
);

NAND2xp67_ASAP7_75t_SL g54 ( 
.A(n_37),
.B(n_31),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_55),
.B(n_64),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_57),
.B(n_71),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_49),
.A2(n_30),
.B1(n_18),
.B2(n_19),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_58),
.A2(n_60),
.B1(n_54),
.B2(n_27),
.Y(n_89)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_59),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_40),
.A2(n_19),
.B1(n_27),
.B2(n_24),
.Y(n_60)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_37),
.B(n_34),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_45),
.B(n_33),
.Y(n_65)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_65),
.Y(n_109)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_66),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_37),
.B(n_33),
.Y(n_67)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_67),
.Y(n_114)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_36),
.Y(n_68)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_68),
.Y(n_82)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_69),
.B(n_56),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_43),
.B(n_16),
.Y(n_71)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_36),
.Y(n_74)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_74),
.Y(n_90)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_36),
.Y(n_76)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_76),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_77),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_79),
.B(n_80),
.Y(n_124)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_63),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_63),
.Y(n_81)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_81),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_83),
.A2(n_87),
.B1(n_97),
.B2(n_104),
.Y(n_118)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_70),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_84),
.B(n_96),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_61),
.Y(n_86)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_86),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_53),
.A2(n_73),
.B1(n_72),
.B2(n_47),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_89),
.A2(n_91),
.B(n_75),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_70),
.A2(n_20),
.B1(n_47),
.B2(n_48),
.Y(n_91)
);

OR2x2_ASAP7_75t_L g92 ( 
.A(n_72),
.B(n_25),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_92),
.B(n_93),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_51),
.B(n_57),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_73),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_95),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_51),
.B(n_25),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_64),
.A2(n_29),
.B1(n_26),
.B2(n_22),
.Y(n_97)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_75),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_98),
.B(n_101),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_55),
.B(n_48),
.C(n_44),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_99),
.B(n_44),
.C(n_61),
.Y(n_131)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_74),
.Y(n_101)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_62),
.Y(n_102)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_102),
.Y(n_133)
);

OR2x2_ASAP7_75t_L g103 ( 
.A(n_71),
.B(n_12),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_103),
.B(n_108),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_50),
.A2(n_29),
.B1(n_26),
.B2(n_38),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_77),
.A2(n_46),
.B1(n_29),
.B2(n_26),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_107),
.A2(n_76),
.B1(n_23),
.B2(n_17),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_69),
.B(n_10),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_66),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_110),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_66),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_111),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_50),
.A2(n_29),
.B1(n_38),
.B2(n_17),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_112),
.A2(n_56),
.B1(n_52),
.B2(n_68),
.Y(n_122)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_78),
.Y(n_113)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_113),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_78),
.B(n_17),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_116),
.B(n_66),
.Y(n_121)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_117),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_121),
.B(n_108),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_122),
.A2(n_142),
.B1(n_118),
.B2(n_134),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_99),
.B(n_52),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_126),
.A2(n_129),
.B(n_136),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_95),
.B(n_78),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_127),
.B(n_130),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_94),
.B(n_106),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_131),
.B(n_88),
.C(n_102),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_132),
.A2(n_84),
.B1(n_104),
.B2(n_112),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_94),
.B(n_2),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_134),
.B(n_137),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_90),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_135),
.B(n_144),
.Y(n_164)
);

O2A1O1Ixp33_ASAP7_75t_L g136 ( 
.A1(n_97),
.A2(n_44),
.B(n_17),
.C(n_61),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_106),
.B(n_2),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_105),
.A2(n_44),
.B(n_61),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_138),
.A2(n_141),
.B(n_127),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_105),
.B(n_87),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_83),
.A2(n_23),
.B1(n_8),
.B2(n_9),
.Y(n_142)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_85),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_117),
.Y(n_148)
);

INVx1_ASAP7_75t_SL g173 ( 
.A(n_148),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_149),
.A2(n_154),
.B1(n_146),
.B2(n_115),
.Y(n_190)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_124),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_150),
.B(n_151),
.Y(n_212)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_124),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_140),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_152),
.B(n_155),
.Y(n_196)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_143),
.Y(n_153)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_153),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_118),
.A2(n_105),
.B1(n_116),
.B2(n_79),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_140),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_156),
.A2(n_163),
.B(n_169),
.Y(n_198)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_121),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_157),
.B(n_158),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_128),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_160),
.A2(n_113),
.B1(n_115),
.B2(n_82),
.Y(n_187)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_122),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_161),
.B(n_166),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_128),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_142),
.Y(n_165)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_165),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_130),
.B(n_92),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_167),
.B(n_170),
.Y(n_194)
);

MAJx2_ASAP7_75t_L g168 ( 
.A(n_141),
.B(n_103),
.C(n_100),
.Y(n_168)
);

MAJx2_ASAP7_75t_L g185 ( 
.A(n_168),
.B(n_126),
.C(n_138),
.Y(n_185)
);

O2A1O1Ixp33_ASAP7_75t_L g169 ( 
.A1(n_132),
.A2(n_120),
.B(n_141),
.C(n_136),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_137),
.B(n_100),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_171),
.B(n_133),
.C(n_86),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_125),
.B(n_114),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_172),
.B(n_174),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_119),
.B(n_109),
.Y(n_174)
);

INVx11_ASAP7_75t_L g175 ( 
.A(n_139),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_175),
.Y(n_200)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_136),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_176),
.B(n_180),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_129),
.A2(n_114),
.B1(n_109),
.B2(n_90),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_178),
.A2(n_23),
.B(n_145),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_143),
.B(n_98),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_179),
.Y(n_199)
);

OR2x2_ASAP7_75t_L g180 ( 
.A(n_146),
.B(n_82),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_125),
.B(n_80),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_181),
.B(n_182),
.Y(n_206)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_131),
.Y(n_182)
);

OAI21xp33_ASAP7_75t_SL g183 ( 
.A1(n_177),
.A2(n_158),
.B(n_163),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_183),
.A2(n_185),
.B(n_208),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_156),
.B(n_126),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_186),
.B(n_201),
.C(n_202),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_187),
.A2(n_188),
.B1(n_213),
.B2(n_175),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_165),
.A2(n_119),
.B1(n_144),
.B2(n_135),
.Y(n_188)
);

NAND2xp33_ASAP7_75t_SL g189 ( 
.A(n_177),
.B(n_101),
.Y(n_189)
);

AOI32xp33_ASAP7_75t_L g229 ( 
.A1(n_189),
.A2(n_172),
.A3(n_162),
.B1(n_180),
.B2(n_153),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_190),
.A2(n_167),
.B1(n_170),
.B2(n_166),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_182),
.A2(n_133),
.B1(n_139),
.B2(n_123),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_191),
.A2(n_197),
.B1(n_215),
.B2(n_149),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_164),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_192),
.B(n_180),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_161),
.A2(n_133),
.B1(n_147),
.B2(n_81),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_171),
.B(n_145),
.C(n_81),
.Y(n_202)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_181),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_205),
.B(n_210),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_169),
.A2(n_23),
.B(n_3),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_209),
.A2(n_176),
.B(n_150),
.Y(n_219)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_164),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_159),
.Y(n_211)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_211),
.Y(n_235)
);

OAI22x1_ASAP7_75t_L g213 ( 
.A1(n_169),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_159),
.Y(n_214)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_214),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_160),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_204),
.A2(n_178),
.B(n_151),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_SL g250 ( 
.A1(n_218),
.A2(n_219),
.B(n_229),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g258 ( 
.A(n_220),
.Y(n_258)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_196),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_221),
.B(n_223),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_193),
.A2(n_154),
.B1(n_157),
.B2(n_152),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_222),
.A2(n_226),
.B1(n_227),
.B2(n_237),
.Y(n_264)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_212),
.Y(n_223)
);

INVx2_ASAP7_75t_SL g224 ( 
.A(n_195),
.Y(n_224)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_224),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_207),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_225),
.B(n_232),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_193),
.A2(n_155),
.B1(n_173),
.B2(n_168),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_213),
.A2(n_173),
.B1(n_168),
.B2(n_174),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_228),
.A2(n_234),
.B1(n_231),
.B2(n_235),
.Y(n_256)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_230),
.Y(n_266)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_204),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_231),
.B(n_234),
.Y(n_262)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_184),
.Y(n_234)
);

BUFx2_ASAP7_75t_L g236 ( 
.A(n_200),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_236),
.B(n_240),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_215),
.A2(n_162),
.B1(n_5),
.B2(n_6),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_186),
.B(n_206),
.C(n_202),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_239),
.B(n_241),
.C(n_198),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_206),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_201),
.B(n_4),
.C(n_5),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_203),
.Y(n_242)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_242),
.Y(n_245)
);

BUFx3_ASAP7_75t_L g243 ( 
.A(n_195),
.Y(n_243)
);

INVxp33_ASAP7_75t_L g248 ( 
.A(n_243),
.Y(n_248)
);

NOR2xp67_ASAP7_75t_SL g247 ( 
.A(n_218),
.B(n_198),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_SL g268 ( 
.A(n_247),
.B(n_263),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_249),
.B(n_252),
.C(n_257),
.Y(n_272)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_233),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_251),
.B(n_253),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_238),
.B(n_214),
.C(n_211),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_233),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_238),
.B(n_190),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_255),
.B(n_260),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_256),
.A2(n_220),
.B1(n_222),
.B2(n_227),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_239),
.B(n_185),
.C(n_191),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_217),
.B(n_226),
.C(n_216),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_217),
.B(n_184),
.C(n_194),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_261),
.B(n_228),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_219),
.A2(n_209),
.B(n_208),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_216),
.B(n_194),
.Y(n_265)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_265),
.Y(n_276)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_267),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_270),
.B(n_280),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_254),
.B(n_199),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_273),
.B(n_274),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_248),
.B(n_224),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_259),
.B(n_221),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_275),
.B(n_278),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_258),
.A2(n_197),
.B1(n_223),
.B2(n_210),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_277),
.A2(n_245),
.B1(n_262),
.B2(n_246),
.Y(n_300)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_256),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_254),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_279),
.B(n_284),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_255),
.B(n_241),
.Y(n_280)
);

MAJx2_ASAP7_75t_L g281 ( 
.A(n_247),
.B(n_203),
.C(n_205),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_SL g299 ( 
.A(n_281),
.B(n_261),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_257),
.B(n_237),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_282),
.B(n_285),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_SL g283 ( 
.A(n_250),
.B(n_199),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_SL g298 ( 
.A(n_283),
.B(n_250),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_266),
.B(n_236),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_260),
.B(n_224),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_280),
.B(n_252),
.C(n_249),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_288),
.B(n_269),
.C(n_272),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_271),
.A2(n_263),
.B(n_258),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_289),
.A2(n_291),
.B(n_262),
.Y(n_303)
);

INVx13_ASAP7_75t_L g290 ( 
.A(n_281),
.Y(n_290)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_290),
.Y(n_305)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_276),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_268),
.A2(n_253),
.B1(n_251),
.B2(n_264),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_292),
.A2(n_299),
.B1(n_300),
.B2(n_290),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_285),
.B(n_265),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_293),
.B(n_269),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_298),
.B(n_289),
.Y(n_314)
);

AOI322xp5_ASAP7_75t_SL g301 ( 
.A1(n_283),
.A2(n_266),
.A3(n_264),
.B1(n_245),
.B2(n_270),
.C1(n_272),
.C2(n_268),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_301),
.B(n_9),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_302),
.B(n_311),
.C(n_313),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_303),
.B(n_310),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_287),
.B(n_282),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_304),
.B(n_298),
.C(n_292),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_306),
.B(n_307),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_300),
.B(n_244),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_293),
.B(n_244),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_308),
.B(n_309),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_291),
.B(n_243),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_287),
.B(n_200),
.C(n_10),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_312),
.B(n_314),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_286),
.B(n_9),
.C(n_11),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_302),
.B(n_288),
.C(n_286),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_319),
.B(n_320),
.C(n_321),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_L g320 ( 
.A1(n_305),
.A2(n_297),
.B(n_295),
.Y(n_320)
);

NOR2xp67_ASAP7_75t_R g323 ( 
.A(n_314),
.B(n_299),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_323),
.B(n_304),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_L g332 ( 
.A1(n_324),
.A2(n_325),
.B(n_328),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_322),
.B(n_318),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_317),
.B(n_311),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_327),
.B(n_330),
.Y(n_333)
);

MAJx2_ASAP7_75t_L g328 ( 
.A(n_322),
.B(n_319),
.C(n_313),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g329 ( 
.A(n_316),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_329),
.B(n_326),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_317),
.B(n_294),
.Y(n_330)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_331),
.Y(n_336)
);

BUFx24_ASAP7_75t_SL g334 ( 
.A(n_328),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_L g335 ( 
.A1(n_334),
.A2(n_332),
.B1(n_329),
.B2(n_296),
.Y(n_335)
);

INVxp67_ASAP7_75t_L g337 ( 
.A(n_335),
.Y(n_337)
);

OAI221xp5_ASAP7_75t_L g338 ( 
.A1(n_337),
.A2(n_333),
.B1(n_336),
.B2(n_315),
.C(n_11),
.Y(n_338)
);

OAI321xp33_ASAP7_75t_L g339 ( 
.A1(n_338),
.A2(n_14),
.A3(n_13),
.B1(n_7),
.B2(n_6),
.C(n_5),
.Y(n_339)
);

AOI21xp5_ASAP7_75t_L g340 ( 
.A1(n_339),
.A2(n_13),
.B(n_14),
.Y(n_340)
);

AOI21xp5_ASAP7_75t_L g341 ( 
.A1(n_340),
.A2(n_13),
.B(n_6),
.Y(n_341)
);


endmodule