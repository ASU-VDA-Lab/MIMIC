module fake_jpeg_31219_n_168 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_168);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_168;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_12),
.Y(n_49)
);

BUFx4f_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_27),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_28),
.Y(n_53)
);

INVx6_ASAP7_75t_SL g54 ( 
.A(n_39),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_3),
.B(n_42),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_25),
.Y(n_57)
);

BUFx16f_ASAP7_75t_L g58 ( 
.A(n_22),
.Y(n_58)
);

INVx6_ASAP7_75t_SL g59 ( 
.A(n_37),
.Y(n_59)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_29),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_33),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_20),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_23),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_13),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_19),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_34),
.Y(n_67)
);

BUFx10_ASAP7_75t_L g68 ( 
.A(n_21),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_1),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_61),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_70),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_61),
.Y(n_71)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_71),
.Y(n_90)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_58),
.Y(n_72)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_72),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_64),
.Y(n_73)
);

BUFx2_ASAP7_75t_L g79 ( 
.A(n_73),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_68),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_74),
.B(n_51),
.Y(n_91)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_58),
.Y(n_75)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_75),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_65),
.Y(n_76)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_76),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_65),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g88 ( 
.A(n_77),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_64),
.Y(n_78)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_78),
.Y(n_83)
);

INVx6_ASAP7_75t_SL g80 ( 
.A(n_72),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_80),
.B(n_68),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_70),
.A2(n_78),
.B1(n_73),
.B2(n_71),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_85),
.A2(n_92),
.B1(n_83),
.B2(n_82),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_72),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_86),
.B(n_91),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_74),
.B(n_57),
.C(n_49),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_87),
.A2(n_89),
.B(n_0),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_72),
.B(n_56),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_76),
.A2(n_52),
.B1(n_49),
.B2(n_50),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_92),
.A2(n_50),
.B1(n_79),
.B2(n_90),
.Y(n_95)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_93),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_95),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_96),
.A2(n_97),
.B1(n_103),
.B2(n_2),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_85),
.A2(n_52),
.B1(n_60),
.B2(n_67),
.Y(n_97)
);

OAI32xp33_ASAP7_75t_L g98 ( 
.A1(n_81),
.A2(n_52),
.A3(n_56),
.B1(n_63),
.B2(n_53),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_98),
.B(n_104),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_99),
.Y(n_122)
);

OR2x6_ASAP7_75t_SL g100 ( 
.A(n_89),
.B(n_68),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_100),
.B(n_101),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_79),
.B(n_69),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_82),
.A2(n_60),
.B1(n_55),
.B2(n_66),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_88),
.Y(n_104)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_84),
.Y(n_105)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_105),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_106),
.B(n_0),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_88),
.B(n_62),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_107),
.B(n_111),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_88),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_91),
.Y(n_109)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_109),
.Y(n_117)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_91),
.Y(n_110)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_110),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_91),
.B(n_48),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_100),
.A2(n_48),
.B1(n_59),
.B2(n_54),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_112),
.A2(n_114),
.B1(n_116),
.B2(n_120),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_100),
.A2(n_14),
.B1(n_44),
.B2(n_41),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_96),
.A2(n_11),
.B1(n_40),
.B2(n_38),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_118),
.B(n_126),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_102),
.B(n_1),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_119),
.B(n_7),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_98),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_120)
);

INVxp33_ASAP7_75t_L g126 ( 
.A(n_94),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_108),
.Y(n_127)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_127),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_128),
.A2(n_131),
.B1(n_5),
.B2(n_6),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_109),
.B(n_4),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_129),
.B(n_130),
.Y(n_137)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_101),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_100),
.A2(n_17),
.B1(n_36),
.B2(n_32),
.Y(n_131)
);

XOR2x1_ASAP7_75t_L g132 ( 
.A(n_115),
.B(n_5),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_132),
.B(n_134),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_133),
.B(n_139),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_122),
.B(n_16),
.C(n_31),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_113),
.A2(n_6),
.B(n_7),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_135),
.B(n_138),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_121),
.B(n_124),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_117),
.B(n_8),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_140),
.B(n_141),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_114),
.B(n_8),
.Y(n_141)
);

XNOR2x1_ASAP7_75t_L g144 ( 
.A(n_131),
.B(n_9),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_144),
.A2(n_147),
.B1(n_9),
.B2(n_10),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_123),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_145),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_126),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_146),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_125),
.B(n_18),
.C(n_30),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_152),
.A2(n_137),
.B(n_147),
.Y(n_157)
);

OA21x2_ASAP7_75t_L g155 ( 
.A1(n_149),
.A2(n_132),
.B(n_143),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_155),
.B(n_157),
.Y(n_160)
);

AOI322xp5_ASAP7_75t_L g156 ( 
.A1(n_148),
.A2(n_150),
.A3(n_153),
.B1(n_154),
.B2(n_136),
.C1(n_135),
.C2(n_125),
.Y(n_156)
);

BUFx24_ASAP7_75t_SL g159 ( 
.A(n_156),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_151),
.B(n_142),
.Y(n_158)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_160),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_161),
.B(n_158),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_162),
.B(n_153),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_163),
.B(n_159),
.Y(n_164)
);

AOI21x1_ASAP7_75t_L g165 ( 
.A1(n_164),
.A2(n_144),
.B(n_134),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_165),
.B(n_116),
.Y(n_166)
);

NOR3xp33_ASAP7_75t_SL g167 ( 
.A(n_166),
.B(n_47),
.C(n_26),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_167),
.B(n_24),
.Y(n_168)
);


endmodule