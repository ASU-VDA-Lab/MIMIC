module fake_netlist_5_2446_n_1706 (n_137, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_109, n_112, n_85, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1706);

input n_137;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_109;
input n_112;
input n_85;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1706;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1166;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_155;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_173;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1580;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_1107;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_171;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_156;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_157;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1598;
wire n_955;
wire n_163;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1036;
wire n_1097;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_475;
wire n_422;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_164;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1672;
wire n_675;
wire n_888;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1623;
wire n_1565;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_857;
wire n_832;
wire n_207;
wire n_561;
wire n_1319;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1199;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1660;
wire n_887;
wire n_154;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1662;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_759;
wire n_806;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_843;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1647;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_284;
wire n_1128;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_372;
wire n_293;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_314;
wire n_433;
wire n_368;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_448;
wire n_259;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_168;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1612;
wire n_1416;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_261;
wire n_174;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_572;
wire n_366;
wire n_815;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_162;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_280;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_153;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1400;
wire n_1342;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_661;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_1638;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_165;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1685;
wire n_601;
wire n_917;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_206;
wire n_172;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_818;
wire n_861;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1059;
wire n_1345;
wire n_176;
wire n_1133;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1440;
wire n_177;
wire n_421;
wire n_1356;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_435;
wire n_159;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_198;
wire n_714;
wire n_1683;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1564;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_1675;
wire n_1554;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_167;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_158;
wire n_704;
wire n_787;
wire n_961;
wire n_771;
wire n_276;
wire n_1225;
wire n_1520;
wire n_169;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_432;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_685;
wire n_598;
wire n_608;
wire n_928;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_413;
wire n_402;
wire n_1086;
wire n_796;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_170;
wire n_161;
wire n_273;
wire n_585;
wire n_270;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_160;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_175;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_166;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_100),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_23),
.Y(n_154)
);

BUFx2_ASAP7_75t_L g155 ( 
.A(n_66),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_121),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_69),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_23),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_147),
.Y(n_159)
);

INVx1_ASAP7_75t_SL g160 ( 
.A(n_9),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_112),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_76),
.Y(n_162)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_139),
.Y(n_163)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_5),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_138),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_77),
.Y(n_166)
);

BUFx3_ASAP7_75t_L g167 ( 
.A(n_10),
.Y(n_167)
);

INVx2_ASAP7_75t_SL g168 ( 
.A(n_75),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_120),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_54),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_10),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_2),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_129),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_47),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_26),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_102),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_71),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_99),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_80),
.Y(n_179)
);

BUFx3_ASAP7_75t_L g180 ( 
.A(n_2),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_89),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_37),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_63),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_114),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_25),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_108),
.Y(n_186)
);

BUFx10_ASAP7_75t_L g187 ( 
.A(n_118),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_87),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_149),
.Y(n_189)
);

INVx1_ASAP7_75t_SL g190 ( 
.A(n_130),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_128),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_95),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_78),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_65),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_148),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_115),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_85),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_1),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_49),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_42),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_5),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_24),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_96),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_41),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_90),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_3),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_124),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_110),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_127),
.Y(n_209)
);

INVx2_ASAP7_75t_SL g210 ( 
.A(n_58),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_144),
.Y(n_211)
);

BUFx2_ASAP7_75t_L g212 ( 
.A(n_28),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_21),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_17),
.Y(n_214)
);

BUFx3_ASAP7_75t_L g215 ( 
.A(n_37),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_64),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_131),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_22),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_19),
.Y(n_219)
);

INVx2_ASAP7_75t_SL g220 ( 
.A(n_56),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_39),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_134),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_70),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_53),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_42),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_27),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_72),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_32),
.Y(n_228)
);

INVx1_ASAP7_75t_SL g229 ( 
.A(n_86),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_143),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_126),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_40),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_41),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_13),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_21),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_116),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_40),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_9),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_22),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_19),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_38),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_97),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_46),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_106),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_103),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_11),
.Y(n_246)
);

BUFx10_ASAP7_75t_L g247 ( 
.A(n_48),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_24),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_32),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_123),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_151),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_104),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_31),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_38),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_4),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_67),
.Y(n_256)
);

INVx2_ASAP7_75t_SL g257 ( 
.A(n_98),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_132),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_31),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_30),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_133),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_101),
.Y(n_262)
);

BUFx3_ASAP7_75t_L g263 ( 
.A(n_30),
.Y(n_263)
);

INVx2_ASAP7_75t_SL g264 ( 
.A(n_35),
.Y(n_264)
);

CKINVDCx16_ASAP7_75t_R g265 ( 
.A(n_36),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_35),
.Y(n_266)
);

CKINVDCx14_ASAP7_75t_R g267 ( 
.A(n_7),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_18),
.Y(n_268)
);

INVx3_ASAP7_75t_L g269 ( 
.A(n_73),
.Y(n_269)
);

BUFx2_ASAP7_75t_SL g270 ( 
.A(n_6),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_84),
.Y(n_271)
);

BUFx10_ASAP7_75t_L g272 ( 
.A(n_8),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_12),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_20),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_55),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_117),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_61),
.Y(n_277)
);

CKINVDCx14_ASAP7_75t_R g278 ( 
.A(n_135),
.Y(n_278)
);

INVx1_ASAP7_75t_SL g279 ( 
.A(n_92),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_20),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_51),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_119),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_68),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_105),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_142),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_57),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_145),
.Y(n_287)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_43),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_140),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_60),
.Y(n_290)
);

INVx2_ASAP7_75t_SL g291 ( 
.A(n_14),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_25),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_94),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_34),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_18),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_33),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_62),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_83),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_29),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_29),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_33),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_93),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_109),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_196),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_167),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_233),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_223),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_212),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_267),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_233),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_233),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_167),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_233),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_233),
.Y(n_314)
);

INVx3_ASAP7_75t_L g315 ( 
.A(n_163),
.Y(n_315)
);

CKINVDCx16_ASAP7_75t_R g316 ( 
.A(n_265),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_164),
.Y(n_317)
);

INVxp67_ASAP7_75t_SL g318 ( 
.A(n_155),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_164),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_239),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_239),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_200),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_253),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_253),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_180),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_201),
.Y(n_326)
);

BUFx2_ASAP7_75t_L g327 ( 
.A(n_180),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_245),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_215),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_171),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_202),
.Y(n_331)
);

HB1xp67_ASAP7_75t_L g332 ( 
.A(n_154),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_215),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_263),
.Y(n_334)
);

INVxp67_ASAP7_75t_SL g335 ( 
.A(n_269),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_263),
.Y(n_336)
);

HB1xp67_ASAP7_75t_L g337 ( 
.A(n_154),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_182),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_251),
.Y(n_339)
);

HB1xp67_ASAP7_75t_L g340 ( 
.A(n_158),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_185),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_198),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_206),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_204),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_219),
.Y(n_345)
);

INVxp67_ASAP7_75t_L g346 ( 
.A(n_272),
.Y(n_346)
);

INVxp67_ASAP7_75t_SL g347 ( 
.A(n_269),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_213),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_226),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_237),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_214),
.Y(n_351)
);

INVxp67_ASAP7_75t_SL g352 ( 
.A(n_269),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_218),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_282),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_221),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_238),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_249),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_268),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_284),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_274),
.Y(n_360)
);

INVxp67_ASAP7_75t_L g361 ( 
.A(n_272),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_225),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_278),
.Y(n_363)
);

INVxp67_ASAP7_75t_SL g364 ( 
.A(n_174),
.Y(n_364)
);

INVxp67_ASAP7_75t_SL g365 ( 
.A(n_179),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_280),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_177),
.Y(n_367)
);

INVxp67_ASAP7_75t_L g368 ( 
.A(n_272),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_228),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_232),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_178),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_300),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_183),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_256),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_193),
.Y(n_375)
);

BUFx6f_ASAP7_75t_L g376 ( 
.A(n_256),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_264),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_199),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_304),
.Y(n_379)
);

INVx3_ASAP7_75t_L g380 ( 
.A(n_376),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_306),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_306),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_307),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_374),
.Y(n_384)
);

XNOR2x2_ASAP7_75t_L g385 ( 
.A(n_377),
.B(n_160),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_335),
.B(n_168),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_374),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_310),
.Y(n_388)
);

HB1xp67_ASAP7_75t_L g389 ( 
.A(n_322),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_310),
.Y(n_390)
);

INVx3_ASAP7_75t_L g391 ( 
.A(n_376),
.Y(n_391)
);

BUFx6f_ASAP7_75t_L g392 ( 
.A(n_376),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_367),
.Y(n_393)
);

BUFx6f_ASAP7_75t_L g394 ( 
.A(n_376),
.Y(n_394)
);

AND2x4_ASAP7_75t_L g395 ( 
.A(n_347),
.B(n_168),
.Y(n_395)
);

INVx4_ASAP7_75t_L g396 ( 
.A(n_376),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_352),
.B(n_210),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_311),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_316),
.A2(n_241),
.B1(n_295),
.B2(n_301),
.Y(n_399)
);

HB1xp67_ASAP7_75t_L g400 ( 
.A(n_322),
.Y(n_400)
);

BUFx6f_ASAP7_75t_L g401 ( 
.A(n_311),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_371),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_313),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_313),
.Y(n_404)
);

BUFx6f_ASAP7_75t_L g405 ( 
.A(n_314),
.Y(n_405)
);

BUFx2_ASAP7_75t_L g406 ( 
.A(n_309),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_314),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_321),
.Y(n_408)
);

AND2x2_ASAP7_75t_L g409 ( 
.A(n_325),
.B(n_264),
.Y(n_409)
);

NAND2x1_ASAP7_75t_L g410 ( 
.A(n_315),
.B(n_210),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_315),
.Y(n_411)
);

AND2x2_ASAP7_75t_L g412 ( 
.A(n_325),
.B(n_291),
.Y(n_412)
);

BUFx6f_ASAP7_75t_L g413 ( 
.A(n_321),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_364),
.B(n_220),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_315),
.Y(n_415)
);

AND2x2_ASAP7_75t_L g416 ( 
.A(n_329),
.B(n_291),
.Y(n_416)
);

INVx6_ASAP7_75t_L g417 ( 
.A(n_365),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_330),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_328),
.A2(n_172),
.B1(n_158),
.B2(n_301),
.Y(n_419)
);

AND2x4_ASAP7_75t_L g420 ( 
.A(n_375),
.B(n_220),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_330),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_317),
.Y(n_422)
);

INVx4_ASAP7_75t_L g423 ( 
.A(n_357),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_357),
.Y(n_424)
);

INVx3_ASAP7_75t_L g425 ( 
.A(n_317),
.Y(n_425)
);

BUFx6f_ASAP7_75t_L g426 ( 
.A(n_319),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_356),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_356),
.Y(n_428)
);

AND2x4_ASAP7_75t_L g429 ( 
.A(n_378),
.B(n_257),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_358),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_373),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_358),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_360),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_360),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_319),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_326),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_320),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_320),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_L g439 ( 
.A1(n_318),
.A2(n_292),
.B1(n_172),
.B2(n_299),
.Y(n_439)
);

BUFx3_ASAP7_75t_L g440 ( 
.A(n_305),
.Y(n_440)
);

CKINVDCx8_ASAP7_75t_R g441 ( 
.A(n_309),
.Y(n_441)
);

BUFx6f_ASAP7_75t_L g442 ( 
.A(n_323),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_323),
.Y(n_443)
);

BUFx6f_ASAP7_75t_L g444 ( 
.A(n_324),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_326),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_324),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_382),
.Y(n_447)
);

BUFx6f_ASAP7_75t_SL g448 ( 
.A(n_395),
.Y(n_448)
);

NAND2xp33_ASAP7_75t_SL g449 ( 
.A(n_419),
.B(n_363),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_381),
.Y(n_450)
);

INVx5_ASAP7_75t_L g451 ( 
.A(n_392),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_381),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_388),
.Y(n_453)
);

AND2x2_ASAP7_75t_L g454 ( 
.A(n_395),
.B(n_420),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_417),
.B(n_331),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_SL g456 ( 
.A(n_441),
.B(n_343),
.Y(n_456)
);

INVx3_ASAP7_75t_L g457 ( 
.A(n_392),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_382),
.Y(n_458)
);

INVx3_ASAP7_75t_L g459 ( 
.A(n_392),
.Y(n_459)
);

INVx3_ASAP7_75t_L g460 ( 
.A(n_392),
.Y(n_460)
);

BUFx3_ASAP7_75t_L g461 ( 
.A(n_440),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_388),
.Y(n_462)
);

AOI22xp33_ASAP7_75t_L g463 ( 
.A1(n_395),
.A2(n_308),
.B1(n_270),
.B2(n_288),
.Y(n_463)
);

AND2x2_ASAP7_75t_L g464 ( 
.A(n_395),
.B(n_329),
.Y(n_464)
);

CKINVDCx20_ASAP7_75t_R g465 ( 
.A(n_379),
.Y(n_465)
);

OAI22xp33_ASAP7_75t_L g466 ( 
.A1(n_414),
.A2(n_255),
.B1(n_234),
.B2(n_260),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_SL g467 ( 
.A(n_441),
.B(n_343),
.Y(n_467)
);

AOI22xp5_ASAP7_75t_L g468 ( 
.A1(n_399),
.A2(n_175),
.B1(n_292),
.B2(n_294),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_SL g469 ( 
.A(n_436),
.B(n_348),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_413),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_417),
.B(n_348),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_390),
.Y(n_472)
);

INVx3_ASAP7_75t_L g473 ( 
.A(n_392),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_413),
.Y(n_474)
);

BUFx2_ASAP7_75t_L g475 ( 
.A(n_385),
.Y(n_475)
);

INVx2_ASAP7_75t_SL g476 ( 
.A(n_417),
.Y(n_476)
);

BUFx6f_ASAP7_75t_L g477 ( 
.A(n_392),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_390),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_398),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_413),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_417),
.B(n_351),
.Y(n_481)
);

NOR3xp33_ASAP7_75t_L g482 ( 
.A(n_439),
.B(n_361),
.C(n_346),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_413),
.Y(n_483)
);

AND2x2_ASAP7_75t_L g484 ( 
.A(n_420),
.B(n_312),
.Y(n_484)
);

INVx1_ASAP7_75t_SL g485 ( 
.A(n_383),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_386),
.B(n_351),
.Y(n_486)
);

BUFx10_ASAP7_75t_L g487 ( 
.A(n_445),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_397),
.B(n_353),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_SL g489 ( 
.A(n_406),
.B(n_353),
.Y(n_489)
);

BUFx10_ASAP7_75t_L g490 ( 
.A(n_389),
.Y(n_490)
);

INVx4_ASAP7_75t_L g491 ( 
.A(n_401),
.Y(n_491)
);

INVx3_ASAP7_75t_L g492 ( 
.A(n_394),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_413),
.Y(n_493)
);

BUFx6f_ASAP7_75t_L g494 ( 
.A(n_394),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_413),
.Y(n_495)
);

BUFx10_ASAP7_75t_L g496 ( 
.A(n_400),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_398),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_403),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_423),
.B(n_355),
.Y(n_499)
);

AND2x4_ASAP7_75t_L g500 ( 
.A(n_420),
.B(n_163),
.Y(n_500)
);

INVx2_ASAP7_75t_SL g501 ( 
.A(n_409),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_393),
.Y(n_502)
);

BUFx6f_ASAP7_75t_L g503 ( 
.A(n_394),
.Y(n_503)
);

AOI22xp33_ASAP7_75t_L g504 ( 
.A1(n_420),
.A2(n_181),
.B1(n_298),
.B2(n_189),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_402),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_431),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_403),
.Y(n_507)
);

INVx3_ASAP7_75t_L g508 ( 
.A(n_394),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_404),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_440),
.B(n_355),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_384),
.Y(n_511)
);

AO21x2_ASAP7_75t_L g512 ( 
.A1(n_404),
.A2(n_208),
.B(n_203),
.Y(n_512)
);

INVx3_ASAP7_75t_L g513 ( 
.A(n_394),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_387),
.Y(n_514)
);

BUFx3_ASAP7_75t_L g515 ( 
.A(n_440),
.Y(n_515)
);

BUFx3_ASAP7_75t_L g516 ( 
.A(n_380),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_387),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_406),
.B(n_362),
.Y(n_518)
);

NOR2x1p5_ASAP7_75t_L g519 ( 
.A(n_410),
.B(n_175),
.Y(n_519)
);

INVx3_ASAP7_75t_L g520 ( 
.A(n_394),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_387),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_407),
.Y(n_522)
);

AND2x6_ASAP7_75t_L g523 ( 
.A(n_429),
.B(n_181),
.Y(n_523)
);

INVx4_ASAP7_75t_L g524 ( 
.A(n_401),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_407),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_423),
.B(n_362),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_426),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_426),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_426),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_423),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_423),
.B(n_369),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_427),
.Y(n_532)
);

NAND3xp33_ASAP7_75t_L g533 ( 
.A(n_409),
.B(n_416),
.C(n_412),
.Y(n_533)
);

INVx3_ASAP7_75t_L g534 ( 
.A(n_396),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_429),
.B(n_369),
.Y(n_535)
);

AND2x2_ASAP7_75t_L g536 ( 
.A(n_429),
.B(n_333),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_SL g537 ( 
.A(n_429),
.B(n_370),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_380),
.B(n_370),
.Y(n_538)
);

INVx1_ASAP7_75t_SL g539 ( 
.A(n_412),
.Y(n_539)
);

INVx3_ASAP7_75t_L g540 ( 
.A(n_396),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_426),
.Y(n_541)
);

INVx1_ASAP7_75t_SL g542 ( 
.A(n_416),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_427),
.Y(n_543)
);

BUFx3_ASAP7_75t_L g544 ( 
.A(n_410),
.Y(n_544)
);

INVx3_ASAP7_75t_L g545 ( 
.A(n_396),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_426),
.Y(n_546)
);

HB1xp67_ASAP7_75t_L g547 ( 
.A(n_385),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_380),
.B(n_190),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_426),
.Y(n_549)
);

AO22x2_ASAP7_75t_L g550 ( 
.A1(n_428),
.A2(n_189),
.B1(n_211),
.B2(n_288),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_442),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_428),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_430),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_442),
.Y(n_554)
);

INVx2_ASAP7_75t_SL g555 ( 
.A(n_430),
.Y(n_555)
);

BUFx3_ASAP7_75t_L g556 ( 
.A(n_380),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_442),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_432),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_442),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_432),
.B(n_332),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_433),
.Y(n_561)
);

NOR2xp33_ASAP7_75t_SL g562 ( 
.A(n_433),
.B(n_339),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_434),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_434),
.Y(n_564)
);

BUFx3_ASAP7_75t_L g565 ( 
.A(n_391),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_442),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_442),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_444),
.Y(n_568)
);

INVx3_ASAP7_75t_L g569 ( 
.A(n_396),
.Y(n_569)
);

BUFx4f_ASAP7_75t_L g570 ( 
.A(n_401),
.Y(n_570)
);

AOI22xp5_ASAP7_75t_L g571 ( 
.A1(n_418),
.A2(n_299),
.B1(n_296),
.B2(n_294),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_435),
.Y(n_572)
);

AO22x2_ASAP7_75t_L g573 ( 
.A1(n_435),
.A2(n_211),
.B1(n_298),
.B2(n_236),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_444),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_444),
.Y(n_575)
);

INVx3_ASAP7_75t_L g576 ( 
.A(n_401),
.Y(n_576)
);

INVx4_ASAP7_75t_L g577 ( 
.A(n_401),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_444),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_425),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_391),
.B(n_229),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_443),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_391),
.B(n_279),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_444),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_444),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_SL g585 ( 
.A(n_418),
.B(n_368),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_443),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_401),
.Y(n_587)
);

BUFx2_ASAP7_75t_L g588 ( 
.A(n_425),
.Y(n_588)
);

INVx2_ASAP7_75t_SL g589 ( 
.A(n_411),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_411),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_405),
.Y(n_591)
);

OR2x6_ASAP7_75t_L g592 ( 
.A(n_438),
.B(n_222),
.Y(n_592)
);

AND2x2_ASAP7_75t_L g593 ( 
.A(n_438),
.B(n_334),
.Y(n_593)
);

CKINVDCx20_ASAP7_75t_R g594 ( 
.A(n_465),
.Y(n_594)
);

XNOR2xp5_ASAP7_75t_L g595 ( 
.A(n_502),
.B(n_354),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_588),
.Y(n_596)
);

NOR2xp33_ASAP7_75t_L g597 ( 
.A(n_486),
.B(n_337),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_SL g598 ( 
.A(n_476),
.B(n_256),
.Y(n_598)
);

BUFx3_ASAP7_75t_L g599 ( 
.A(n_502),
.Y(n_599)
);

AOI22xp33_ASAP7_75t_L g600 ( 
.A1(n_475),
.A2(n_261),
.B1(n_256),
.B2(n_242),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_L g601 ( 
.A(n_488),
.B(n_340),
.Y(n_601)
);

OAI22xp33_ASAP7_75t_L g602 ( 
.A1(n_475),
.A2(n_296),
.B1(n_235),
.B2(n_266),
.Y(n_602)
);

INVx3_ASAP7_75t_L g603 ( 
.A(n_516),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_588),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_454),
.B(n_425),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_454),
.B(n_425),
.Y(n_606)
);

OAI22xp33_ASAP7_75t_L g607 ( 
.A1(n_547),
.A2(n_273),
.B1(n_240),
.B2(n_246),
.Y(n_607)
);

AOI22xp33_ASAP7_75t_L g608 ( 
.A1(n_512),
.A2(n_256),
.B1(n_261),
.B2(n_290),
.Y(n_608)
);

BUFx6f_ASAP7_75t_SL g609 ( 
.A(n_487),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_476),
.B(n_391),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_L g611 ( 
.A(n_539),
.B(n_153),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_532),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_579),
.B(n_405),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_SL g614 ( 
.A(n_501),
.B(n_261),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_579),
.B(n_405),
.Y(n_615)
);

AND2x4_ASAP7_75t_L g616 ( 
.A(n_461),
.B(n_338),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_555),
.B(n_405),
.Y(n_617)
);

AND2x2_ASAP7_75t_L g618 ( 
.A(n_542),
.B(n_327),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_L g619 ( 
.A(n_471),
.B(n_153),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_555),
.B(n_405),
.Y(n_620)
);

AOI21xp5_ASAP7_75t_L g621 ( 
.A1(n_530),
.A2(n_415),
.B(n_437),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_SL g622 ( 
.A(n_501),
.B(n_455),
.Y(n_622)
);

INVx2_ASAP7_75t_SL g623 ( 
.A(n_484),
.Y(n_623)
);

OAI22x1_ASAP7_75t_L g624 ( 
.A1(n_468),
.A2(n_518),
.B1(n_571),
.B2(n_505),
.Y(n_624)
);

INVx2_ASAP7_75t_SL g625 ( 
.A(n_484),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_532),
.Y(n_626)
);

AOI22xp5_ASAP7_75t_L g627 ( 
.A1(n_448),
.A2(n_359),
.B1(n_216),
.B2(n_244),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_543),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_543),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_481),
.B(n_405),
.Y(n_630)
);

A2O1A1Ixp33_ASAP7_75t_L g631 ( 
.A1(n_533),
.A2(n_250),
.B(n_297),
.C(n_446),
.Y(n_631)
);

INVx5_ASAP7_75t_L g632 ( 
.A(n_523),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_530),
.B(n_415),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_589),
.B(n_415),
.Y(n_634)
);

INVxp67_ASAP7_75t_L g635 ( 
.A(n_560),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_552),
.Y(n_636)
);

INVx8_ASAP7_75t_L g637 ( 
.A(n_448),
.Y(n_637)
);

NAND2x1p5_ASAP7_75t_L g638 ( 
.A(n_544),
.B(n_261),
.Y(n_638)
);

NOR2xp33_ASAP7_75t_L g639 ( 
.A(n_499),
.B(n_156),
.Y(n_639)
);

AOI22xp33_ASAP7_75t_L g640 ( 
.A1(n_512),
.A2(n_261),
.B1(n_344),
.B2(n_349),
.Y(n_640)
);

AOI22xp33_ASAP7_75t_L g641 ( 
.A1(n_512),
.A2(n_341),
.B1(n_342),
.B2(n_372),
.Y(n_641)
);

AOI22xp5_ASAP7_75t_L g642 ( 
.A1(n_448),
.A2(n_464),
.B1(n_562),
.B2(n_531),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_SL g643 ( 
.A(n_533),
.B(n_184),
.Y(n_643)
);

AOI22xp5_ASAP7_75t_L g644 ( 
.A1(n_464),
.A2(n_186),
.B1(n_188),
.B2(n_191),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_553),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_589),
.B(n_422),
.Y(n_646)
);

INVxp67_ASAP7_75t_L g647 ( 
.A(n_510),
.Y(n_647)
);

AND2x2_ASAP7_75t_L g648 ( 
.A(n_536),
.B(n_327),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_SL g649 ( 
.A(n_526),
.B(n_192),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_558),
.B(n_422),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_558),
.B(n_422),
.Y(n_651)
);

INVx4_ASAP7_75t_L g652 ( 
.A(n_461),
.Y(n_652)
);

O2A1O1Ixp5_ASAP7_75t_L g653 ( 
.A1(n_500),
.A2(n_446),
.B(n_437),
.C(n_336),
.Y(n_653)
);

AND2x2_ASAP7_75t_L g654 ( 
.A(n_536),
.B(n_377),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_SL g655 ( 
.A(n_535),
.B(n_561),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_561),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_563),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_563),
.B(n_437),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_564),
.B(n_446),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_564),
.Y(n_660)
);

BUFx6f_ASAP7_75t_L g661 ( 
.A(n_461),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_SL g662 ( 
.A(n_544),
.B(n_194),
.Y(n_662)
);

O2A1O1Ixp33_ASAP7_75t_L g663 ( 
.A1(n_537),
.A2(n_366),
.B(n_350),
.C(n_345),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_572),
.B(n_408),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_572),
.B(n_581),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_593),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_511),
.Y(n_667)
);

AND2x2_ASAP7_75t_L g668 ( 
.A(n_490),
.B(n_421),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_593),
.Y(n_669)
);

AND2x2_ASAP7_75t_L g670 ( 
.A(n_490),
.B(n_421),
.Y(n_670)
);

INVx1_ASAP7_75t_SL g671 ( 
.A(n_485),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_511),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_581),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_586),
.B(n_408),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_586),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_514),
.Y(n_676)
);

AND2x2_ASAP7_75t_L g677 ( 
.A(n_490),
.B(n_424),
.Y(n_677)
);

INVx2_ASAP7_75t_SL g678 ( 
.A(n_538),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_SL g679 ( 
.A(n_500),
.B(n_195),
.Y(n_679)
);

INVx2_ASAP7_75t_SL g680 ( 
.A(n_519),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_514),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_450),
.Y(n_682)
);

INVx2_ASAP7_75t_SL g683 ( 
.A(n_519),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_450),
.B(n_424),
.Y(n_684)
);

OR2x2_ASAP7_75t_L g685 ( 
.A(n_489),
.B(n_248),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_452),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_517),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_517),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_452),
.B(n_197),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_SL g690 ( 
.A(n_500),
.B(n_515),
.Y(n_690)
);

INVxp67_ASAP7_75t_L g691 ( 
.A(n_585),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_521),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_SL g693 ( 
.A(n_500),
.B(n_205),
.Y(n_693)
);

NAND2xp33_ASAP7_75t_L g694 ( 
.A(n_523),
.B(n_207),
.Y(n_694)
);

NOR2xp33_ASAP7_75t_L g695 ( 
.A(n_515),
.B(n_156),
.Y(n_695)
);

AND2x2_ASAP7_75t_L g696 ( 
.A(n_490),
.B(n_254),
.Y(n_696)
);

AOI22xp33_ASAP7_75t_L g697 ( 
.A1(n_550),
.A2(n_573),
.B1(n_523),
.B2(n_504),
.Y(n_697)
);

XOR2xp5_ASAP7_75t_L g698 ( 
.A(n_506),
.B(n_209),
.Y(n_698)
);

AND2x2_ASAP7_75t_L g699 ( 
.A(n_496),
.B(n_259),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_453),
.B(n_462),
.Y(n_700)
);

NOR2xp33_ASAP7_75t_L g701 ( 
.A(n_515),
.B(n_157),
.Y(n_701)
);

INVx2_ASAP7_75t_SL g702 ( 
.A(n_496),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_453),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_462),
.B(n_217),
.Y(n_704)
);

AO22x2_ASAP7_75t_L g705 ( 
.A1(n_482),
.A2(n_469),
.B1(n_467),
.B2(n_456),
.Y(n_705)
);

AO22x2_ASAP7_75t_L g706 ( 
.A1(n_468),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_706)
);

AND2x2_ASAP7_75t_L g707 ( 
.A(n_496),
.B(n_187),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_472),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_472),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_L g710 ( 
.A(n_466),
.B(n_157),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_478),
.B(n_224),
.Y(n_711)
);

BUFx12f_ASAP7_75t_SL g712 ( 
.A(n_592),
.Y(n_712)
);

A2O1A1Ixp33_ASAP7_75t_L g713 ( 
.A1(n_463),
.A2(n_252),
.B(n_227),
.C(n_230),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_479),
.B(n_497),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_521),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_479),
.B(n_231),
.Y(n_716)
);

NOR2xp33_ASAP7_75t_L g717 ( 
.A(n_497),
.B(n_159),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_498),
.B(n_243),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_498),
.B(n_258),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_447),
.Y(n_720)
);

INVxp67_ASAP7_75t_L g721 ( 
.A(n_571),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_507),
.B(n_262),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_507),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_SL g724 ( 
.A(n_534),
.B(n_271),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_509),
.B(n_275),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_509),
.B(n_522),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_SL g727 ( 
.A(n_487),
.B(n_303),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_522),
.B(n_276),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_447),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_525),
.Y(n_730)
);

OAI21xp5_ASAP7_75t_L g731 ( 
.A1(n_534),
.A2(n_277),
.B(n_281),
.Y(n_731)
);

OAI221xp5_ASAP7_75t_L g732 ( 
.A1(n_525),
.A2(n_303),
.B1(n_302),
.B2(n_293),
.C(n_289),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_458),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_548),
.B(n_283),
.Y(n_734)
);

INVx1_ASAP7_75t_SL g735 ( 
.A(n_506),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_SL g736 ( 
.A(n_534),
.B(n_285),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_580),
.B(n_286),
.Y(n_737)
);

INVx2_ASAP7_75t_SL g738 ( 
.A(n_496),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_458),
.Y(n_739)
);

HB1xp67_ASAP7_75t_L g740 ( 
.A(n_592),
.Y(n_740)
);

NOR2xp33_ASAP7_75t_SL g741 ( 
.A(n_487),
.B(n_187),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_SL g742 ( 
.A(n_487),
.B(n_293),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_582),
.B(n_287),
.Y(n_743)
);

NOR2xp67_ASAP7_75t_L g744 ( 
.A(n_590),
.B(n_289),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_540),
.B(n_169),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_540),
.B(n_169),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_SL g747 ( 
.A(n_540),
.B(n_166),
.Y(n_747)
);

OAI22xp5_ASAP7_75t_L g748 ( 
.A1(n_592),
.A2(n_166),
.B1(n_161),
.B2(n_176),
.Y(n_748)
);

AOI21xp5_ASAP7_75t_L g749 ( 
.A1(n_540),
.A2(n_170),
.B(n_161),
.Y(n_749)
);

NOR2xp67_ASAP7_75t_L g750 ( 
.A(n_590),
.B(n_159),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_SL g751 ( 
.A(n_545),
.B(n_176),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_SL g752 ( 
.A(n_545),
.B(n_173),
.Y(n_752)
);

OAI22xp5_ASAP7_75t_L g753 ( 
.A1(n_592),
.A2(n_173),
.B1(n_170),
.B2(n_165),
.Y(n_753)
);

OR2x2_ASAP7_75t_L g754 ( 
.A(n_449),
.B(n_162),
.Y(n_754)
);

INVx2_ASAP7_75t_SL g755 ( 
.A(n_592),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_545),
.B(n_165),
.Y(n_756)
);

NOR2xp33_ASAP7_75t_L g757 ( 
.A(n_647),
.B(n_545),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_612),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_626),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_720),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_729),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_594),
.Y(n_762)
);

BUFx2_ASAP7_75t_L g763 ( 
.A(n_618),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_733),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_628),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_739),
.Y(n_766)
);

AOI22xp33_ASAP7_75t_L g767 ( 
.A1(n_710),
.A2(n_523),
.B1(n_516),
.B2(n_556),
.Y(n_767)
);

AND2x4_ASAP7_75t_L g768 ( 
.A(n_623),
.B(n_556),
.Y(n_768)
);

BUFx3_ASAP7_75t_L g769 ( 
.A(n_599),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_629),
.Y(n_770)
);

AND2x4_ASAP7_75t_L g771 ( 
.A(n_625),
.B(n_556),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_636),
.Y(n_772)
);

AND2x4_ASAP7_75t_L g773 ( 
.A(n_616),
.B(n_565),
.Y(n_773)
);

AND2x4_ASAP7_75t_L g774 ( 
.A(n_616),
.B(n_565),
.Y(n_774)
);

INVx1_ASAP7_75t_SL g775 ( 
.A(n_671),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_678),
.B(n_647),
.Y(n_776)
);

AOI22xp33_ASAP7_75t_L g777 ( 
.A1(n_710),
.A2(n_523),
.B1(n_565),
.B2(n_573),
.Y(n_777)
);

AND2x2_ASAP7_75t_L g778 ( 
.A(n_635),
.B(n_573),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_665),
.B(n_523),
.Y(n_779)
);

INVx2_ASAP7_75t_SL g780 ( 
.A(n_648),
.Y(n_780)
);

INVx4_ASAP7_75t_L g781 ( 
.A(n_661),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_700),
.B(n_523),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_645),
.Y(n_783)
);

NAND2xp33_ASAP7_75t_SL g784 ( 
.A(n_609),
.B(n_162),
.Y(n_784)
);

AOI22xp33_ASAP7_75t_L g785 ( 
.A1(n_600),
.A2(n_573),
.B1(n_550),
.B2(n_584),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_656),
.Y(n_786)
);

BUFx6f_ASAP7_75t_L g787 ( 
.A(n_661),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_657),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_635),
.B(n_569),
.Y(n_789)
);

AND2x4_ASAP7_75t_L g790 ( 
.A(n_680),
.B(n_587),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_639),
.B(n_569),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_SL g792 ( 
.A(n_642),
.B(n_570),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_660),
.Y(n_793)
);

NAND3xp33_ASAP7_75t_SL g794 ( 
.A(n_741),
.B(n_247),
.C(n_557),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_714),
.B(n_527),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_SL g796 ( 
.A(n_619),
.B(n_570),
.Y(n_796)
);

BUFx5_ASAP7_75t_L g797 ( 
.A(n_673),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_675),
.Y(n_798)
);

AOI22xp5_ASAP7_75t_L g799 ( 
.A1(n_639),
.A2(n_554),
.B1(n_527),
.B2(n_584),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_682),
.Y(n_800)
);

INVx3_ASAP7_75t_SL g801 ( 
.A(n_735),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_686),
.Y(n_802)
);

AND2x2_ASAP7_75t_L g803 ( 
.A(n_597),
.B(n_550),
.Y(n_803)
);

AND2x6_ASAP7_75t_L g804 ( 
.A(n_668),
.B(n_470),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_619),
.B(n_457),
.Y(n_805)
);

NOR2xp33_ASAP7_75t_R g806 ( 
.A(n_595),
.B(n_457),
.Y(n_806)
);

AOI22xp33_ASAP7_75t_L g807 ( 
.A1(n_600),
.A2(n_550),
.B1(n_529),
.B2(n_583),
.Y(n_807)
);

INVx1_ASAP7_75t_SL g808 ( 
.A(n_670),
.Y(n_808)
);

INVx2_ASAP7_75t_SL g809 ( 
.A(n_654),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_703),
.Y(n_810)
);

NOR2xp33_ASAP7_75t_L g811 ( 
.A(n_597),
.B(n_491),
.Y(n_811)
);

AND2x2_ASAP7_75t_L g812 ( 
.A(n_601),
.B(n_247),
.Y(n_812)
);

BUFx3_ASAP7_75t_L g813 ( 
.A(n_637),
.Y(n_813)
);

BUFx6f_ASAP7_75t_L g814 ( 
.A(n_661),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_726),
.B(n_528),
.Y(n_815)
);

INVxp67_ASAP7_75t_SL g816 ( 
.A(n_661),
.Y(n_816)
);

OR2x6_ASAP7_75t_L g817 ( 
.A(n_637),
.B(n_528),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_605),
.B(n_529),
.Y(n_818)
);

OAI22xp5_ASAP7_75t_L g819 ( 
.A1(n_608),
.A2(n_470),
.B1(n_474),
.B2(n_480),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_SL g820 ( 
.A(n_622),
.B(n_570),
.Y(n_820)
);

AND2x4_ASAP7_75t_L g821 ( 
.A(n_683),
.B(n_587),
.Y(n_821)
);

AOI22xp5_ASAP7_75t_L g822 ( 
.A1(n_622),
.A2(n_559),
.B1(n_583),
.B2(n_578),
.Y(n_822)
);

INVx5_ASAP7_75t_L g823 ( 
.A(n_637),
.Y(n_823)
);

INVxp67_ASAP7_75t_L g824 ( 
.A(n_611),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_SL g825 ( 
.A(n_677),
.B(n_477),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_708),
.Y(n_826)
);

BUFx4f_ASAP7_75t_L g827 ( 
.A(n_702),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_709),
.Y(n_828)
);

INVx8_ASAP7_75t_L g829 ( 
.A(n_609),
.Y(n_829)
);

AOI21xp5_ASAP7_75t_L g830 ( 
.A1(n_630),
.A2(n_491),
.B(n_524),
.Y(n_830)
);

AOI22xp5_ASAP7_75t_L g831 ( 
.A1(n_655),
.A2(n_557),
.B1(n_578),
.B2(n_541),
.Y(n_831)
);

OAI22xp5_ASAP7_75t_SL g832 ( 
.A1(n_721),
.A2(n_0),
.B1(n_4),
.B2(n_6),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_606),
.B(n_541),
.Y(n_833)
);

NAND2x1p5_ASAP7_75t_L g834 ( 
.A(n_632),
.B(n_491),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_SL g835 ( 
.A(n_601),
.B(n_477),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_667),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_723),
.Y(n_837)
);

AOI22xp33_ASAP7_75t_L g838 ( 
.A1(n_655),
.A2(n_559),
.B1(n_546),
.B2(n_549),
.Y(n_838)
);

OAI21xp5_ASAP7_75t_L g839 ( 
.A1(n_653),
.A2(n_495),
.B(n_474),
.Y(n_839)
);

INVxp67_ASAP7_75t_L g840 ( 
.A(n_611),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_672),
.Y(n_841)
);

INVx3_ASAP7_75t_L g842 ( 
.A(n_603),
.Y(n_842)
);

INVx2_ASAP7_75t_SL g843 ( 
.A(n_696),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_676),
.Y(n_844)
);

CKINVDCx5p33_ASAP7_75t_R g845 ( 
.A(n_698),
.Y(n_845)
);

INVx3_ASAP7_75t_L g846 ( 
.A(n_603),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_730),
.B(n_457),
.Y(n_847)
);

INVx5_ASAP7_75t_L g848 ( 
.A(n_738),
.Y(n_848)
);

AND2x4_ASAP7_75t_L g849 ( 
.A(n_666),
.B(n_591),
.Y(n_849)
);

BUFx6f_ASAP7_75t_L g850 ( 
.A(n_652),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_646),
.Y(n_851)
);

BUFx4f_ASAP7_75t_L g852 ( 
.A(n_596),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_669),
.B(n_546),
.Y(n_853)
);

INVx1_ASAP7_75t_SL g854 ( 
.A(n_604),
.Y(n_854)
);

AND2x2_ASAP7_75t_L g855 ( 
.A(n_699),
.B(n_707),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_641),
.B(n_549),
.Y(n_856)
);

NOR2xp33_ASAP7_75t_L g857 ( 
.A(n_721),
.B(n_691),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_681),
.Y(n_858)
);

AND2x2_ASAP7_75t_L g859 ( 
.A(n_691),
.B(n_551),
.Y(n_859)
);

INVx1_ASAP7_75t_SL g860 ( 
.A(n_685),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_634),
.Y(n_861)
);

CKINVDCx5p33_ASAP7_75t_R g862 ( 
.A(n_624),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_664),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_641),
.B(n_551),
.Y(n_864)
);

AOI21xp5_ASAP7_75t_L g865 ( 
.A1(n_690),
.A2(n_491),
.B(n_577),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_674),
.Y(n_866)
);

INVx2_ASAP7_75t_SL g867 ( 
.A(n_705),
.Y(n_867)
);

NAND2xp33_ASAP7_75t_L g868 ( 
.A(n_632),
.B(n_477),
.Y(n_868)
);

NOR2xp33_ASAP7_75t_L g869 ( 
.A(n_754),
.B(n_524),
.Y(n_869)
);

INVxp67_ASAP7_75t_L g870 ( 
.A(n_705),
.Y(n_870)
);

HB1xp67_ASAP7_75t_L g871 ( 
.A(n_712),
.Y(n_871)
);

NAND2x1p5_ASAP7_75t_L g872 ( 
.A(n_632),
.B(n_524),
.Y(n_872)
);

BUFx8_ASAP7_75t_L g873 ( 
.A(n_755),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_684),
.Y(n_874)
);

AND2x4_ASAP7_75t_L g875 ( 
.A(n_740),
.B(n_591),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_687),
.Y(n_876)
);

INVx2_ASAP7_75t_SL g877 ( 
.A(n_662),
.Y(n_877)
);

AOI22xp5_ASAP7_75t_L g878 ( 
.A1(n_643),
.A2(n_567),
.B1(n_575),
.B2(n_574),
.Y(n_878)
);

BUFx6f_ASAP7_75t_L g879 ( 
.A(n_652),
.Y(n_879)
);

HB1xp67_ASAP7_75t_L g880 ( 
.A(n_740),
.Y(n_880)
);

BUFx2_ASAP7_75t_L g881 ( 
.A(n_706),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_608),
.B(n_567),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_650),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_651),
.B(n_658),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_659),
.Y(n_885)
);

BUFx2_ASAP7_75t_L g886 ( 
.A(n_706),
.Y(n_886)
);

OR2x2_ASAP7_75t_L g887 ( 
.A(n_727),
.B(n_495),
.Y(n_887)
);

AND2x2_ASAP7_75t_L g888 ( 
.A(n_742),
.B(n_575),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_SL g889 ( 
.A(n_632),
.B(n_494),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_688),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_692),
.Y(n_891)
);

INVx3_ASAP7_75t_L g892 ( 
.A(n_715),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_613),
.B(n_568),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_633),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_690),
.Y(n_895)
);

NAND2x1p5_ASAP7_75t_L g896 ( 
.A(n_614),
.B(n_577),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_617),
.Y(n_897)
);

INVx5_ASAP7_75t_L g898 ( 
.A(n_694),
.Y(n_898)
);

INVx2_ASAP7_75t_SL g899 ( 
.A(n_662),
.Y(n_899)
);

INVx2_ASAP7_75t_L g900 ( 
.A(n_610),
.Y(n_900)
);

CKINVDCx5p33_ASAP7_75t_R g901 ( 
.A(n_627),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_615),
.B(n_566),
.Y(n_902)
);

CKINVDCx5p33_ASAP7_75t_R g903 ( 
.A(n_644),
.Y(n_903)
);

BUFx3_ASAP7_75t_L g904 ( 
.A(n_689),
.Y(n_904)
);

BUFx3_ASAP7_75t_L g905 ( 
.A(n_704),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_SL g906 ( 
.A(n_711),
.B(n_503),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_631),
.B(n_554),
.Y(n_907)
);

AND2x2_ASAP7_75t_L g908 ( 
.A(n_717),
.B(n_493),
.Y(n_908)
);

BUFx6f_ASAP7_75t_L g909 ( 
.A(n_638),
.Y(n_909)
);

INVx3_ASAP7_75t_L g910 ( 
.A(n_638),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_SL g911 ( 
.A(n_716),
.B(n_494),
.Y(n_911)
);

AOI22xp5_ASAP7_75t_L g912 ( 
.A1(n_649),
.A2(n_736),
.B1(n_724),
.B2(n_679),
.Y(n_912)
);

NAND2x1p5_ASAP7_75t_L g913 ( 
.A(n_614),
.B(n_577),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_640),
.B(n_480),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_717),
.B(n_492),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_620),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_598),
.Y(n_917)
);

INVx2_ASAP7_75t_L g918 ( 
.A(n_598),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_734),
.B(n_492),
.Y(n_919)
);

OAI21xp5_ASAP7_75t_L g920 ( 
.A1(n_621),
.A2(n_483),
.B(n_493),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_640),
.B(n_737),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_743),
.B(n_483),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_663),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_718),
.Y(n_924)
);

AND2x4_ASAP7_75t_L g925 ( 
.A(n_679),
.B(n_576),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_719),
.Y(n_926)
);

OAI22xp5_ASAP7_75t_SL g927 ( 
.A1(n_732),
.A2(n_7),
.B1(n_8),
.B2(n_11),
.Y(n_927)
);

AOI22xp5_ASAP7_75t_L g928 ( 
.A1(n_649),
.A2(n_576),
.B1(n_492),
.B2(n_520),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_722),
.Y(n_929)
);

BUFx6f_ASAP7_75t_L g930 ( 
.A(n_693),
.Y(n_930)
);

INVx2_ASAP7_75t_SL g931 ( 
.A(n_725),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_SL g932 ( 
.A(n_728),
.B(n_695),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_745),
.B(n_576),
.Y(n_933)
);

BUFx3_ASAP7_75t_L g934 ( 
.A(n_769),
.Y(n_934)
);

OAI22xp5_ASAP7_75t_SL g935 ( 
.A1(n_901),
.A2(n_862),
.B1(n_903),
.B2(n_845),
.Y(n_935)
);

OAI22xp5_ASAP7_75t_L g936 ( 
.A1(n_870),
.A2(n_697),
.B1(n_706),
.B2(n_695),
.Y(n_936)
);

AOI21xp5_ASAP7_75t_L g937 ( 
.A1(n_791),
.A2(n_731),
.B(n_724),
.Y(n_937)
);

INVx2_ASAP7_75t_L g938 ( 
.A(n_849),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_SL g939 ( 
.A(n_824),
.B(n_701),
.Y(n_939)
);

A2O1A1Ixp33_ASAP7_75t_L g940 ( 
.A1(n_924),
.A2(n_701),
.B(n_713),
.C(n_693),
.Y(n_940)
);

AOI21xp5_ASAP7_75t_L g941 ( 
.A1(n_868),
.A2(n_736),
.B(n_752),
.Y(n_941)
);

INVx2_ASAP7_75t_L g942 ( 
.A(n_849),
.Y(n_942)
);

OR2x2_ASAP7_75t_L g943 ( 
.A(n_763),
.B(n_607),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_863),
.B(n_756),
.Y(n_944)
);

NOR2xp33_ASAP7_75t_R g945 ( 
.A(n_762),
.B(n_746),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_758),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_892),
.Y(n_947)
);

AOI21x1_ASAP7_75t_L g948 ( 
.A1(n_796),
.A2(n_752),
.B(n_751),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_759),
.Y(n_949)
);

A2O1A1Ixp33_ASAP7_75t_L g950 ( 
.A1(n_926),
.A2(n_747),
.B(n_751),
.C(n_750),
.Y(n_950)
);

HB1xp67_ASAP7_75t_L g951 ( 
.A(n_775),
.Y(n_951)
);

NOR2xp33_ASAP7_75t_L g952 ( 
.A(n_840),
.B(n_602),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_SL g953 ( 
.A(n_808),
.B(n_744),
.Y(n_953)
);

OR2x6_ASAP7_75t_SL g954 ( 
.A(n_776),
.B(n_753),
.Y(n_954)
);

INVx2_ASAP7_75t_SL g955 ( 
.A(n_775),
.Y(n_955)
);

CKINVDCx5p33_ASAP7_75t_R g956 ( 
.A(n_801),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_765),
.Y(n_957)
);

AOI22xp33_ASAP7_75t_L g958 ( 
.A1(n_867),
.A2(n_697),
.B1(n_748),
.B2(n_749),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_770),
.Y(n_959)
);

AOI21xp5_ASAP7_75t_L g960 ( 
.A1(n_834),
.A2(n_477),
.B(n_494),
.Y(n_960)
);

AO22x1_ASAP7_75t_L g961 ( 
.A1(n_857),
.A2(n_12),
.B1(n_14),
.B2(n_15),
.Y(n_961)
);

O2A1O1Ixp5_ASAP7_75t_L g962 ( 
.A1(n_932),
.A2(n_520),
.B(n_513),
.C(n_508),
.Y(n_962)
);

NAND2xp33_ASAP7_75t_L g963 ( 
.A(n_797),
.B(n_477),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_772),
.Y(n_964)
);

HB1xp67_ASAP7_75t_L g965 ( 
.A(n_880),
.Y(n_965)
);

AOI21xp5_ASAP7_75t_L g966 ( 
.A1(n_872),
.A2(n_494),
.B(n_503),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_866),
.B(n_874),
.Y(n_967)
);

AOI21xp5_ASAP7_75t_L g968 ( 
.A1(n_872),
.A2(n_494),
.B(n_503),
.Y(n_968)
);

BUFx2_ASAP7_75t_SL g969 ( 
.A(n_823),
.Y(n_969)
);

CKINVDCx20_ASAP7_75t_R g970 ( 
.A(n_806),
.Y(n_970)
);

AOI21xp5_ASAP7_75t_L g971 ( 
.A1(n_884),
.A2(n_503),
.B(n_451),
.Y(n_971)
);

AOI22xp5_ASAP7_75t_L g972 ( 
.A1(n_855),
.A2(n_520),
.B1(n_513),
.B2(n_508),
.Y(n_972)
);

AOI33xp33_ASAP7_75t_L g973 ( 
.A1(n_860),
.A2(n_854),
.A3(n_780),
.B1(n_809),
.B2(n_843),
.B3(n_808),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_783),
.Y(n_974)
);

AOI21xp5_ASAP7_75t_L g975 ( 
.A1(n_884),
.A2(n_503),
.B(n_451),
.Y(n_975)
);

AOI21xp5_ASAP7_75t_L g976 ( 
.A1(n_779),
.A2(n_782),
.B(n_830),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_786),
.Y(n_977)
);

NOR2xp33_ASAP7_75t_L g978 ( 
.A(n_929),
.B(n_513),
.Y(n_978)
);

OAI22xp33_ASAP7_75t_L g979 ( 
.A1(n_860),
.A2(n_508),
.B1(n_492),
.B2(n_473),
.Y(n_979)
);

OAI22xp5_ASAP7_75t_L g980 ( 
.A1(n_921),
.A2(n_508),
.B1(n_473),
.B2(n_460),
.Y(n_980)
);

NAND2xp33_ASAP7_75t_L g981 ( 
.A(n_797),
.B(n_460),
.Y(n_981)
);

AO21x1_ASAP7_75t_L g982 ( 
.A1(n_912),
.A2(n_15),
.B(n_16),
.Y(n_982)
);

BUFx6f_ASAP7_75t_L g983 ( 
.A(n_787),
.Y(n_983)
);

O2A1O1Ixp33_ASAP7_75t_L g984 ( 
.A1(n_877),
.A2(n_473),
.B(n_460),
.C(n_459),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_851),
.B(n_459),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_894),
.B(n_459),
.Y(n_986)
);

OAI22xp5_ASAP7_75t_L g987 ( 
.A1(n_921),
.A2(n_457),
.B1(n_451),
.B2(n_26),
.Y(n_987)
);

NOR2xp33_ASAP7_75t_L g988 ( 
.A(n_931),
.B(n_16),
.Y(n_988)
);

BUFx3_ASAP7_75t_L g989 ( 
.A(n_813),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_SL g990 ( 
.A(n_899),
.B(n_451),
.Y(n_990)
);

O2A1O1Ixp33_ASAP7_75t_SL g991 ( 
.A1(n_820),
.A2(n_82),
.B(n_152),
.C(n_150),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_788),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_793),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_883),
.B(n_451),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_885),
.B(n_79),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_798),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_SL g997 ( 
.A(n_930),
.B(n_74),
.Y(n_997)
);

AND2x4_ASAP7_75t_L g998 ( 
.A(n_823),
.B(n_81),
.Y(n_998)
);

INVxp67_ASAP7_75t_L g999 ( 
.A(n_854),
.Y(n_999)
);

NOR2xp33_ASAP7_75t_L g1000 ( 
.A(n_904),
.B(n_17),
.Y(n_1000)
);

AND2x2_ASAP7_75t_L g1001 ( 
.A(n_852),
.B(n_27),
.Y(n_1001)
);

BUFx3_ASAP7_75t_L g1002 ( 
.A(n_829),
.Y(n_1002)
);

AOI21xp5_ASAP7_75t_L g1003 ( 
.A1(n_782),
.A2(n_88),
.B(n_141),
.Y(n_1003)
);

O2A1O1Ixp33_ASAP7_75t_L g1004 ( 
.A1(n_792),
.A2(n_28),
.B(n_34),
.C(n_36),
.Y(n_1004)
);

INVx1_ASAP7_75t_SL g1005 ( 
.A(n_859),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_800),
.Y(n_1006)
);

INVx3_ASAP7_75t_L g1007 ( 
.A(n_787),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_802),
.Y(n_1008)
);

AOI21xp5_ASAP7_75t_L g1009 ( 
.A1(n_893),
.A2(n_107),
.B(n_44),
.Y(n_1009)
);

AOI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_893),
.A2(n_902),
.B(n_933),
.Y(n_1010)
);

BUFx12f_ASAP7_75t_L g1011 ( 
.A(n_873),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_810),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_861),
.B(n_897),
.Y(n_1013)
);

O2A1O1Ixp33_ASAP7_75t_L g1014 ( 
.A1(n_794),
.A2(n_45),
.B(n_50),
.C(n_52),
.Y(n_1014)
);

OR2x2_ASAP7_75t_L g1015 ( 
.A(n_881),
.B(n_59),
.Y(n_1015)
);

BUFx2_ASAP7_75t_L g1016 ( 
.A(n_871),
.Y(n_1016)
);

OAI22x1_ASAP7_75t_L g1017 ( 
.A1(n_886),
.A2(n_91),
.B1(n_111),
.B2(n_113),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_916),
.B(n_122),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_757),
.B(n_125),
.Y(n_1019)
);

OAI22xp5_ASAP7_75t_L g1020 ( 
.A1(n_807),
.A2(n_146),
.B1(n_136),
.B2(n_137),
.Y(n_1020)
);

AOI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_902),
.A2(n_933),
.B(n_922),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_826),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_789),
.B(n_895),
.Y(n_1023)
);

BUFx6f_ASAP7_75t_L g1024 ( 
.A(n_787),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_905),
.B(n_828),
.Y(n_1025)
);

AOI22xp5_ASAP7_75t_L g1026 ( 
.A1(n_930),
.A2(n_888),
.B1(n_804),
.B2(n_803),
.Y(n_1026)
);

INVx3_ASAP7_75t_L g1027 ( 
.A(n_814),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_837),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_908),
.B(n_869),
.Y(n_1029)
);

HB1xp67_ASAP7_75t_L g1030 ( 
.A(n_875),
.Y(n_1030)
);

A2O1A1Ixp33_ASAP7_75t_L g1031 ( 
.A1(n_923),
.A2(n_925),
.B(n_887),
.C(n_900),
.Y(n_1031)
);

INVx3_ASAP7_75t_L g1032 ( 
.A(n_814),
.Y(n_1032)
);

NOR3xp33_ASAP7_75t_SL g1033 ( 
.A(n_832),
.B(n_927),
.C(n_784),
.Y(n_1033)
);

AOI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_922),
.A2(n_898),
.B(n_865),
.Y(n_1034)
);

NOR2xp33_ASAP7_75t_L g1035 ( 
.A(n_768),
.B(n_771),
.Y(n_1035)
);

AND2x4_ASAP7_75t_L g1036 ( 
.A(n_773),
.B(n_774),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_804),
.B(n_778),
.Y(n_1037)
);

OR2x6_ASAP7_75t_L g1038 ( 
.A(n_829),
.B(n_817),
.Y(n_1038)
);

BUFx2_ASAP7_75t_L g1039 ( 
.A(n_873),
.Y(n_1039)
);

AOI21xp5_ASAP7_75t_L g1040 ( 
.A1(n_898),
.A2(n_919),
.B(n_795),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_853),
.Y(n_1041)
);

O2A1O1Ixp5_ASAP7_75t_L g1042 ( 
.A1(n_835),
.A2(n_911),
.B(n_906),
.C(n_805),
.Y(n_1042)
);

NAND3xp33_ASAP7_75t_SL g1043 ( 
.A(n_767),
.B(n_777),
.C(n_915),
.Y(n_1043)
);

AOI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_898),
.A2(n_815),
.B(n_795),
.Y(n_1044)
);

NOR2xp33_ASAP7_75t_SL g1045 ( 
.A(n_927),
.B(n_832),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_SL g1046 ( 
.A(n_797),
.B(n_879),
.Y(n_1046)
);

A2O1A1Ixp33_ASAP7_75t_L g1047 ( 
.A1(n_925),
.A2(n_864),
.B(n_856),
.C(n_918),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_804),
.B(n_815),
.Y(n_1048)
);

BUFx12f_ASAP7_75t_L g1049 ( 
.A(n_848),
.Y(n_1049)
);

A2O1A1Ixp33_ASAP7_75t_L g1050 ( 
.A1(n_856),
.A2(n_864),
.B(n_917),
.C(n_907),
.Y(n_1050)
);

CKINVDCx6p67_ASAP7_75t_R g1051 ( 
.A(n_829),
.Y(n_1051)
);

BUFx6f_ASAP7_75t_L g1052 ( 
.A(n_814),
.Y(n_1052)
);

AND2x2_ASAP7_75t_SL g1053 ( 
.A(n_827),
.B(n_850),
.Y(n_1053)
);

NAND2x1p5_ASAP7_75t_L g1054 ( 
.A(n_850),
.B(n_879),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_853),
.Y(n_1055)
);

A2O1A1Ixp33_ASAP7_75t_L g1056 ( 
.A1(n_882),
.A2(n_833),
.B(n_818),
.C(n_878),
.Y(n_1056)
);

A2O1A1Ixp33_ASAP7_75t_L g1057 ( 
.A1(n_914),
.A2(n_891),
.B(n_890),
.C(n_822),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_SL g1058 ( 
.A(n_797),
.B(n_879),
.Y(n_1058)
);

CKINVDCx11_ASAP7_75t_R g1059 ( 
.A(n_817),
.Y(n_1059)
);

AOI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_816),
.A2(n_889),
.B(n_825),
.Y(n_1060)
);

AOI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_842),
.A2(n_846),
.B(n_896),
.Y(n_1061)
);

AOI21xp5_ASAP7_75t_L g1062 ( 
.A1(n_842),
.A2(n_846),
.B(n_896),
.Y(n_1062)
);

AOI21xp5_ASAP7_75t_L g1063 ( 
.A1(n_913),
.A2(n_819),
.B(n_920),
.Y(n_1063)
);

O2A1O1Ixp5_ASAP7_75t_SL g1064 ( 
.A1(n_819),
.A2(n_839),
.B(n_920),
.C(n_910),
.Y(n_1064)
);

AND2x4_ASAP7_75t_L g1065 ( 
.A(n_1036),
.B(n_774),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_946),
.Y(n_1066)
);

NAND2xp33_ASAP7_75t_L g1067 ( 
.A(n_967),
.B(n_797),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_949),
.Y(n_1068)
);

AOI21xp33_ASAP7_75t_L g1069 ( 
.A1(n_952),
.A2(n_799),
.B(n_847),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_957),
.Y(n_1070)
);

INVx2_ASAP7_75t_L g1071 ( 
.A(n_959),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_964),
.Y(n_1072)
);

OA21x2_ASAP7_75t_L g1073 ( 
.A1(n_1063),
.A2(n_839),
.B(n_831),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_967),
.B(n_768),
.Y(n_1074)
);

NOR2xp33_ASAP7_75t_L g1075 ( 
.A(n_939),
.B(n_771),
.Y(n_1075)
);

INVx4_ASAP7_75t_L g1076 ( 
.A(n_934),
.Y(n_1076)
);

A2O1A1Ixp33_ASAP7_75t_L g1077 ( 
.A1(n_940),
.A2(n_827),
.B(n_910),
.C(n_821),
.Y(n_1077)
);

OR2x2_ASAP7_75t_L g1078 ( 
.A(n_951),
.B(n_821),
.Y(n_1078)
);

OAI21x1_ASAP7_75t_L g1079 ( 
.A1(n_976),
.A2(n_838),
.B(n_928),
.Y(n_1079)
);

AOI221xp5_ASAP7_75t_L g1080 ( 
.A1(n_1045),
.A2(n_790),
.B1(n_773),
.B2(n_785),
.C(n_875),
.Y(n_1080)
);

OAI21xp5_ASAP7_75t_SL g1081 ( 
.A1(n_1001),
.A2(n_790),
.B(n_909),
.Y(n_1081)
);

AOI21xp5_ASAP7_75t_L g1082 ( 
.A1(n_937),
.A2(n_781),
.B(n_909),
.Y(n_1082)
);

AO31x2_ASAP7_75t_L g1083 ( 
.A1(n_1031),
.A2(n_858),
.A3(n_844),
.B(n_841),
.Y(n_1083)
);

OAI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_1064),
.A2(n_804),
.B(n_876),
.Y(n_1084)
);

OAI21x1_ASAP7_75t_L g1085 ( 
.A1(n_1061),
.A2(n_836),
.B(n_761),
.Y(n_1085)
);

NOR2xp33_ASAP7_75t_L g1086 ( 
.A(n_999),
.B(n_760),
.Y(n_1086)
);

OR2x2_ASAP7_75t_L g1087 ( 
.A(n_943),
.B(n_764),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_1005),
.B(n_766),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_974),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_SL g1090 ( 
.A(n_955),
.B(n_909),
.Y(n_1090)
);

OAI21x1_ASAP7_75t_L g1091 ( 
.A1(n_1062),
.A2(n_817),
.B(n_781),
.Y(n_1091)
);

AO21x1_ASAP7_75t_L g1092 ( 
.A1(n_987),
.A2(n_1029),
.B(n_1019),
.Y(n_1092)
);

AO21x2_ASAP7_75t_L g1093 ( 
.A1(n_1044),
.A2(n_1040),
.B(n_1021),
.Y(n_1093)
);

AOI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_1010),
.A2(n_981),
.B(n_941),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_1005),
.B(n_1013),
.Y(n_1095)
);

BUFx12f_ASAP7_75t_L g1096 ( 
.A(n_956),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_1041),
.B(n_1055),
.Y(n_1097)
);

AOI22xp5_ASAP7_75t_L g1098 ( 
.A1(n_1045),
.A2(n_970),
.B1(n_935),
.B2(n_953),
.Y(n_1098)
);

BUFx3_ASAP7_75t_L g1099 ( 
.A(n_989),
.Y(n_1099)
);

INVx2_ASAP7_75t_L g1100 ( 
.A(n_977),
.Y(n_1100)
);

O2A1O1Ixp33_ASAP7_75t_L g1101 ( 
.A1(n_1033),
.A2(n_950),
.B(n_1000),
.C(n_988),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_SL g1102 ( 
.A(n_1053),
.B(n_1025),
.Y(n_1102)
);

CKINVDCx5p33_ASAP7_75t_R g1103 ( 
.A(n_945),
.Y(n_1103)
);

OAI21x1_ASAP7_75t_L g1104 ( 
.A1(n_960),
.A2(n_968),
.B(n_966),
.Y(n_1104)
);

OAI21xp5_ASAP7_75t_L g1105 ( 
.A1(n_1047),
.A2(n_1050),
.B(n_1043),
.Y(n_1105)
);

AOI22x1_ASAP7_75t_L g1106 ( 
.A1(n_1017),
.A2(n_1003),
.B1(n_1060),
.B2(n_1009),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_1013),
.B(n_944),
.Y(n_1107)
);

OA21x2_ASAP7_75t_L g1108 ( 
.A1(n_1042),
.A2(n_962),
.B(n_1057),
.Y(n_1108)
);

AOI21xp5_ASAP7_75t_L g1109 ( 
.A1(n_1019),
.A2(n_1023),
.B(n_1048),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_1035),
.B(n_1023),
.Y(n_1110)
);

OAI21x1_ASAP7_75t_L g1111 ( 
.A1(n_980),
.A2(n_975),
.B(n_971),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_1030),
.B(n_992),
.Y(n_1112)
);

AO21x2_ASAP7_75t_L g1113 ( 
.A1(n_948),
.A2(n_980),
.B(n_987),
.Y(n_1113)
);

AO31x2_ASAP7_75t_L g1114 ( 
.A1(n_982),
.A2(n_936),
.A3(n_1020),
.B(n_1018),
.Y(n_1114)
);

OA21x2_ASAP7_75t_L g1115 ( 
.A1(n_1018),
.A2(n_995),
.B(n_994),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_993),
.Y(n_1116)
);

NAND3xp33_ASAP7_75t_L g1117 ( 
.A(n_973),
.B(n_1004),
.C(n_961),
.Y(n_1117)
);

A2O1A1Ixp33_ASAP7_75t_L g1118 ( 
.A1(n_995),
.A2(n_1020),
.B(n_1026),
.C(n_978),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_996),
.Y(n_1119)
);

NOR2xp67_ASAP7_75t_SL g1120 ( 
.A(n_969),
.B(n_1049),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_1006),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_1008),
.Y(n_1122)
);

OAI21xp5_ASAP7_75t_L g1123 ( 
.A1(n_984),
.A2(n_936),
.B(n_986),
.Y(n_1123)
);

OAI22xp5_ASAP7_75t_L g1124 ( 
.A1(n_958),
.A2(n_954),
.B1(n_1028),
.B2(n_1022),
.Y(n_1124)
);

OA21x2_ASAP7_75t_L g1125 ( 
.A1(n_994),
.A2(n_1037),
.B(n_985),
.Y(n_1125)
);

OAI21x1_ASAP7_75t_L g1126 ( 
.A1(n_1046),
.A2(n_1058),
.B(n_990),
.Y(n_1126)
);

OAI21xp5_ASAP7_75t_L g1127 ( 
.A1(n_972),
.A2(n_1014),
.B(n_979),
.Y(n_1127)
);

OAI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_997),
.A2(n_1012),
.B(n_991),
.Y(n_1128)
);

OAI21x1_ASAP7_75t_L g1129 ( 
.A1(n_1054),
.A2(n_1032),
.B(n_1027),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_1036),
.B(n_938),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_942),
.B(n_947),
.Y(n_1131)
);

OR2x4_ASAP7_75t_L g1132 ( 
.A(n_1015),
.B(n_983),
.Y(n_1132)
);

INVx1_ASAP7_75t_SL g1133 ( 
.A(n_965),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_1007),
.B(n_1032),
.Y(n_1134)
);

OAI21x1_ASAP7_75t_L g1135 ( 
.A1(n_1007),
.A2(n_1027),
.B(n_1038),
.Y(n_1135)
);

CKINVDCx11_ASAP7_75t_R g1136 ( 
.A(n_1011),
.Y(n_1136)
);

AO31x2_ASAP7_75t_L g1137 ( 
.A1(n_1016),
.A2(n_1039),
.A3(n_1052),
.B(n_983),
.Y(n_1137)
);

OAI21x1_ASAP7_75t_L g1138 ( 
.A1(n_1038),
.A2(n_1059),
.B(n_983),
.Y(n_1138)
);

INVx3_ASAP7_75t_L g1139 ( 
.A(n_1024),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_998),
.B(n_1024),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_1024),
.Y(n_1141)
);

AOI21xp5_ASAP7_75t_L g1142 ( 
.A1(n_1052),
.A2(n_1002),
.B(n_1051),
.Y(n_1142)
);

NOR2xp67_ASAP7_75t_L g1143 ( 
.A(n_1052),
.B(n_823),
.Y(n_1143)
);

OAI21xp5_ASAP7_75t_L g1144 ( 
.A1(n_1063),
.A2(n_1064),
.B(n_1056),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_946),
.Y(n_1145)
);

OAI21x1_ASAP7_75t_L g1146 ( 
.A1(n_976),
.A2(n_1062),
.B(n_1061),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_967),
.B(n_824),
.Y(n_1147)
);

NOR2xp33_ASAP7_75t_L g1148 ( 
.A(n_967),
.B(n_824),
.Y(n_1148)
);

NAND2x1p5_ASAP7_75t_L g1149 ( 
.A(n_1053),
.B(n_850),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_SL g1150 ( 
.A(n_955),
.B(n_824),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_967),
.B(n_1041),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_967),
.B(n_824),
.Y(n_1152)
);

O2A1O1Ixp5_ASAP7_75t_L g1153 ( 
.A1(n_1029),
.A2(n_796),
.B(n_811),
.C(n_937),
.Y(n_1153)
);

BUFx4_ASAP7_75t_R g1154 ( 
.A(n_934),
.Y(n_1154)
);

INVxp67_ASAP7_75t_SL g1155 ( 
.A(n_999),
.Y(n_1155)
);

INVx2_ASAP7_75t_SL g1156 ( 
.A(n_934),
.Y(n_1156)
);

AOI21xp5_ASAP7_75t_L g1157 ( 
.A1(n_963),
.A2(n_937),
.B(n_1034),
.Y(n_1157)
);

AO31x2_ASAP7_75t_L g1158 ( 
.A1(n_1063),
.A2(n_937),
.A3(n_1031),
.B(n_987),
.Y(n_1158)
);

INVx2_ASAP7_75t_L g1159 ( 
.A(n_946),
.Y(n_1159)
);

OAI21x1_ASAP7_75t_L g1160 ( 
.A1(n_976),
.A2(n_1062),
.B(n_1061),
.Y(n_1160)
);

AOI22xp5_ASAP7_75t_L g1161 ( 
.A1(n_1045),
.A2(n_307),
.B1(n_328),
.B2(n_304),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_967),
.B(n_1041),
.Y(n_1162)
);

AO21x2_ASAP7_75t_L g1163 ( 
.A1(n_1063),
.A2(n_937),
.B(n_1034),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_L g1164 ( 
.A(n_967),
.B(n_824),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_SL g1165 ( 
.A(n_955),
.B(n_824),
.Y(n_1165)
);

CKINVDCx11_ASAP7_75t_R g1166 ( 
.A(n_1011),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_SL g1167 ( 
.A(n_955),
.B(n_824),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_946),
.Y(n_1168)
);

AND2x4_ASAP7_75t_L g1169 ( 
.A(n_1036),
.B(n_1038),
.Y(n_1169)
);

OAI21xp5_ASAP7_75t_L g1170 ( 
.A1(n_1063),
.A2(n_1064),
.B(n_1056),
.Y(n_1170)
);

INVxp67_ASAP7_75t_L g1171 ( 
.A(n_951),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_L g1172 ( 
.A(n_967),
.B(n_1041),
.Y(n_1172)
);

A2O1A1Ixp33_ASAP7_75t_L g1173 ( 
.A1(n_952),
.A2(n_912),
.B(n_811),
.C(n_924),
.Y(n_1173)
);

NAND3xp33_ASAP7_75t_SL g1174 ( 
.A(n_1045),
.B(n_741),
.C(n_812),
.Y(n_1174)
);

INVx2_ASAP7_75t_L g1175 ( 
.A(n_946),
.Y(n_1175)
);

OAI21xp5_ASAP7_75t_L g1176 ( 
.A1(n_1063),
.A2(n_1064),
.B(n_1056),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_967),
.B(n_824),
.Y(n_1177)
);

INVx3_ASAP7_75t_SL g1178 ( 
.A(n_956),
.Y(n_1178)
);

O2A1O1Ixp33_ASAP7_75t_L g1179 ( 
.A1(n_939),
.A2(n_812),
.B(n_840),
.C(n_824),
.Y(n_1179)
);

BUFx3_ASAP7_75t_L g1180 ( 
.A(n_934),
.Y(n_1180)
);

OAI21xp5_ASAP7_75t_L g1181 ( 
.A1(n_1063),
.A2(n_1064),
.B(n_1056),
.Y(n_1181)
);

AO31x2_ASAP7_75t_L g1182 ( 
.A1(n_1063),
.A2(n_937),
.A3(n_1031),
.B(n_987),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_946),
.Y(n_1183)
);

AO21x1_ASAP7_75t_L g1184 ( 
.A1(n_987),
.A2(n_1029),
.B(n_1019),
.Y(n_1184)
);

OAI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_1063),
.A2(n_1064),
.B(n_1056),
.Y(n_1185)
);

INVx3_ASAP7_75t_L g1186 ( 
.A(n_1054),
.Y(n_1186)
);

NOR2xp33_ASAP7_75t_L g1187 ( 
.A(n_967),
.B(n_824),
.Y(n_1187)
);

OAI22xp5_ASAP7_75t_L g1188 ( 
.A1(n_967),
.A2(n_600),
.B1(n_608),
.B2(n_1013),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_967),
.B(n_1041),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_946),
.Y(n_1190)
);

AOI21xp5_ASAP7_75t_L g1191 ( 
.A1(n_963),
.A2(n_937),
.B(n_1034),
.Y(n_1191)
);

AOI21xp33_ASAP7_75t_L g1192 ( 
.A1(n_952),
.A2(n_812),
.B(n_811),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_946),
.Y(n_1193)
);

AOI21xp5_ASAP7_75t_L g1194 ( 
.A1(n_963),
.A2(n_937),
.B(n_1034),
.Y(n_1194)
);

HB1xp67_ASAP7_75t_L g1195 ( 
.A(n_951),
.Y(n_1195)
);

INVx2_ASAP7_75t_L g1196 ( 
.A(n_946),
.Y(n_1196)
);

BUFx6f_ASAP7_75t_L g1197 ( 
.A(n_1053),
.Y(n_1197)
);

OAI221xp5_ASAP7_75t_L g1198 ( 
.A1(n_1192),
.A2(n_1173),
.B1(n_1101),
.B2(n_1174),
.C(n_1179),
.Y(n_1198)
);

AOI22xp33_ASAP7_75t_L g1199 ( 
.A1(n_1192),
.A2(n_1117),
.B1(n_1184),
.B2(n_1092),
.Y(n_1199)
);

INVx2_ASAP7_75t_L g1200 ( 
.A(n_1071),
.Y(n_1200)
);

O2A1O1Ixp33_ASAP7_75t_L g1201 ( 
.A1(n_1124),
.A2(n_1118),
.B(n_1102),
.C(n_1107),
.Y(n_1201)
);

O2A1O1Ixp33_ASAP7_75t_SL g1202 ( 
.A1(n_1077),
.A2(n_1188),
.B(n_1069),
.C(n_1128),
.Y(n_1202)
);

AOI21xp5_ASAP7_75t_L g1203 ( 
.A1(n_1094),
.A2(n_1191),
.B(n_1157),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_1100),
.Y(n_1204)
);

A2O1A1Ixp33_ASAP7_75t_L g1205 ( 
.A1(n_1188),
.A2(n_1105),
.B(n_1148),
.C(n_1187),
.Y(n_1205)
);

AND2x6_ASAP7_75t_SL g1206 ( 
.A(n_1086),
.B(n_1075),
.Y(n_1206)
);

BUFx2_ASAP7_75t_L g1207 ( 
.A(n_1195),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_1151),
.B(n_1162),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_1151),
.B(n_1162),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1159),
.Y(n_1210)
);

OR2x2_ASAP7_75t_L g1211 ( 
.A(n_1095),
.B(n_1087),
.Y(n_1211)
);

INVx2_ASAP7_75t_SL g1212 ( 
.A(n_1180),
.Y(n_1212)
);

OR2x2_ASAP7_75t_L g1213 ( 
.A(n_1110),
.B(n_1147),
.Y(n_1213)
);

AO31x2_ASAP7_75t_L g1214 ( 
.A1(n_1194),
.A2(n_1109),
.A3(n_1124),
.B(n_1082),
.Y(n_1214)
);

OAI22xp5_ASAP7_75t_L g1215 ( 
.A1(n_1172),
.A2(n_1189),
.B1(n_1164),
.B2(n_1177),
.Y(n_1215)
);

INVx2_ASAP7_75t_L g1216 ( 
.A(n_1175),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1196),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1066),
.Y(n_1218)
);

BUFx2_ASAP7_75t_SL g1219 ( 
.A(n_1076),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1068),
.Y(n_1220)
);

OR2x2_ASAP7_75t_L g1221 ( 
.A(n_1152),
.B(n_1133),
.Y(n_1221)
);

BUFx6f_ASAP7_75t_L g1222 ( 
.A(n_1197),
.Y(n_1222)
);

AND2x2_ASAP7_75t_L g1223 ( 
.A(n_1197),
.B(n_1065),
.Y(n_1223)
);

INVxp67_ASAP7_75t_L g1224 ( 
.A(n_1155),
.Y(n_1224)
);

AOI22xp33_ASAP7_75t_L g1225 ( 
.A1(n_1117),
.A2(n_1105),
.B1(n_1189),
.B2(n_1172),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_1097),
.B(n_1074),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_1070),
.Y(n_1227)
);

BUFx8_ASAP7_75t_L g1228 ( 
.A(n_1096),
.Y(n_1228)
);

OAI21x1_ASAP7_75t_L g1229 ( 
.A1(n_1111),
.A2(n_1079),
.B(n_1085),
.Y(n_1229)
);

OAI21x1_ASAP7_75t_L g1230 ( 
.A1(n_1091),
.A2(n_1106),
.B(n_1126),
.Y(n_1230)
);

INVx1_ASAP7_75t_SL g1231 ( 
.A(n_1154),
.Y(n_1231)
);

INVx2_ASAP7_75t_SL g1232 ( 
.A(n_1099),
.Y(n_1232)
);

NOR2xp33_ASAP7_75t_SL g1233 ( 
.A(n_1076),
.B(n_1103),
.Y(n_1233)
);

NAND2x1p5_ASAP7_75t_L g1234 ( 
.A(n_1138),
.B(n_1135),
.Y(n_1234)
);

OA21x2_ASAP7_75t_L g1235 ( 
.A1(n_1144),
.A2(n_1185),
.B(n_1181),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1072),
.Y(n_1236)
);

OAI21x1_ASAP7_75t_L g1237 ( 
.A1(n_1144),
.A2(n_1176),
.B(n_1170),
.Y(n_1237)
);

AOI221xp5_ASAP7_75t_L g1238 ( 
.A1(n_1069),
.A2(n_1170),
.B1(n_1185),
.B2(n_1127),
.C(n_1171),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_1089),
.Y(n_1239)
);

INVx1_ASAP7_75t_SL g1240 ( 
.A(n_1133),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_1116),
.Y(n_1241)
);

OAI21x1_ASAP7_75t_L g1242 ( 
.A1(n_1084),
.A2(n_1073),
.B(n_1123),
.Y(n_1242)
);

NAND2x1p5_ASAP7_75t_L g1243 ( 
.A(n_1186),
.B(n_1197),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1119),
.Y(n_1244)
);

OAI21x1_ASAP7_75t_L g1245 ( 
.A1(n_1084),
.A2(n_1073),
.B(n_1123),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1121),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_L g1247 ( 
.A(n_1097),
.B(n_1114),
.Y(n_1247)
);

A2O1A1Ixp33_ASAP7_75t_L g1248 ( 
.A1(n_1127),
.A2(n_1080),
.B(n_1067),
.C(n_1081),
.Y(n_1248)
);

OR2x6_ASAP7_75t_L g1249 ( 
.A(n_1081),
.B(n_1149),
.Y(n_1249)
);

INVx2_ASAP7_75t_L g1250 ( 
.A(n_1122),
.Y(n_1250)
);

OAI21x1_ASAP7_75t_L g1251 ( 
.A1(n_1108),
.A2(n_1115),
.B(n_1125),
.Y(n_1251)
);

BUFx6f_ASAP7_75t_L g1252 ( 
.A(n_1169),
.Y(n_1252)
);

CKINVDCx20_ASAP7_75t_R g1253 ( 
.A(n_1136),
.Y(n_1253)
);

NOR2x1p5_ASAP7_75t_L g1254 ( 
.A(n_1140),
.B(n_1130),
.Y(n_1254)
);

OA21x2_ASAP7_75t_L g1255 ( 
.A1(n_1145),
.A2(n_1193),
.B(n_1168),
.Y(n_1255)
);

AOI221x1_ASAP7_75t_L g1256 ( 
.A1(n_1183),
.A2(n_1190),
.B1(n_1134),
.B2(n_1088),
.C(n_1112),
.Y(n_1256)
);

OAI21x1_ASAP7_75t_L g1257 ( 
.A1(n_1108),
.A2(n_1115),
.B(n_1125),
.Y(n_1257)
);

AND2x2_ASAP7_75t_L g1258 ( 
.A(n_1065),
.B(n_1078),
.Y(n_1258)
);

AOI22x1_ASAP7_75t_L g1259 ( 
.A1(n_1186),
.A2(n_1142),
.B1(n_1141),
.B2(n_1139),
.Y(n_1259)
);

OAI21x1_ASAP7_75t_L g1260 ( 
.A1(n_1129),
.A2(n_1134),
.B(n_1131),
.Y(n_1260)
);

INVx2_ASAP7_75t_SL g1261 ( 
.A(n_1156),
.Y(n_1261)
);

O2A1O1Ixp33_ASAP7_75t_SL g1262 ( 
.A1(n_1090),
.A2(n_1131),
.B(n_1114),
.C(n_1098),
.Y(n_1262)
);

INVxp67_ASAP7_75t_SL g1263 ( 
.A(n_1150),
.Y(n_1263)
);

AOI22xp33_ASAP7_75t_L g1264 ( 
.A1(n_1161),
.A2(n_1113),
.B1(n_1165),
.B2(n_1167),
.Y(n_1264)
);

HB1xp67_ASAP7_75t_L g1265 ( 
.A(n_1137),
.Y(n_1265)
);

OAI21x1_ASAP7_75t_L g1266 ( 
.A1(n_1093),
.A2(n_1163),
.B(n_1143),
.Y(n_1266)
);

AOI21x1_ASAP7_75t_L g1267 ( 
.A1(n_1120),
.A2(n_1113),
.B(n_1083),
.Y(n_1267)
);

AOI22xp33_ASAP7_75t_L g1268 ( 
.A1(n_1178),
.A2(n_1166),
.B1(n_1132),
.B2(n_1158),
.Y(n_1268)
);

OR2x6_ASAP7_75t_L g1269 ( 
.A(n_1132),
.B(n_1137),
.Y(n_1269)
);

OAI21x1_ASAP7_75t_L g1270 ( 
.A1(n_1158),
.A2(n_1182),
.B(n_1137),
.Y(n_1270)
);

OA21x2_ASAP7_75t_L g1271 ( 
.A1(n_1182),
.A2(n_1170),
.B(n_1144),
.Y(n_1271)
);

BUFx3_ASAP7_75t_L g1272 ( 
.A(n_1180),
.Y(n_1272)
);

NAND3xp33_ASAP7_75t_L g1273 ( 
.A(n_1192),
.B(n_812),
.C(n_741),
.Y(n_1273)
);

OA21x2_ASAP7_75t_L g1274 ( 
.A1(n_1144),
.A2(n_1176),
.B(n_1170),
.Y(n_1274)
);

CKINVDCx5p33_ASAP7_75t_R g1275 ( 
.A(n_1154),
.Y(n_1275)
);

O2A1O1Ixp33_ASAP7_75t_L g1276 ( 
.A1(n_1192),
.A2(n_1101),
.B(n_1174),
.C(n_1173),
.Y(n_1276)
);

OAI21xp5_ASAP7_75t_L g1277 ( 
.A1(n_1173),
.A2(n_1192),
.B(n_1153),
.Y(n_1277)
);

BUFx3_ASAP7_75t_L g1278 ( 
.A(n_1180),
.Y(n_1278)
);

INVx3_ASAP7_75t_L g1279 ( 
.A(n_1149),
.Y(n_1279)
);

INVx3_ASAP7_75t_L g1280 ( 
.A(n_1149),
.Y(n_1280)
);

BUFx6f_ASAP7_75t_L g1281 ( 
.A(n_1197),
.Y(n_1281)
);

INVx4_ASAP7_75t_L g1282 ( 
.A(n_1154),
.Y(n_1282)
);

OR2x2_ASAP7_75t_L g1283 ( 
.A(n_1095),
.B(n_1087),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1071),
.Y(n_1284)
);

INVx2_ASAP7_75t_L g1285 ( 
.A(n_1071),
.Y(n_1285)
);

OAI21xp33_ASAP7_75t_SL g1286 ( 
.A1(n_1107),
.A2(n_600),
.B(n_1151),
.Y(n_1286)
);

OAI21xp5_ASAP7_75t_L g1287 ( 
.A1(n_1173),
.A2(n_1192),
.B(n_1153),
.Y(n_1287)
);

OA21x2_ASAP7_75t_L g1288 ( 
.A1(n_1144),
.A2(n_1176),
.B(n_1170),
.Y(n_1288)
);

NOR2xp67_ASAP7_75t_L g1289 ( 
.A(n_1171),
.B(n_999),
.Y(n_1289)
);

INVx2_ASAP7_75t_L g1290 ( 
.A(n_1071),
.Y(n_1290)
);

AO31x2_ASAP7_75t_L g1291 ( 
.A1(n_1092),
.A2(n_1184),
.A3(n_1191),
.B(n_1157),
.Y(n_1291)
);

AO31x2_ASAP7_75t_L g1292 ( 
.A1(n_1092),
.A2(n_1184),
.A3(n_1191),
.B(n_1157),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_L g1293 ( 
.A(n_1151),
.B(n_1162),
.Y(n_1293)
);

A2O1A1Ixp33_ASAP7_75t_L g1294 ( 
.A1(n_1101),
.A2(n_1173),
.B(n_1045),
.C(n_1192),
.Y(n_1294)
);

BUFx3_ASAP7_75t_L g1295 ( 
.A(n_1180),
.Y(n_1295)
);

INVx2_ASAP7_75t_SL g1296 ( 
.A(n_1180),
.Y(n_1296)
);

INVx2_ASAP7_75t_SL g1297 ( 
.A(n_1180),
.Y(n_1297)
);

AOI211xp5_ASAP7_75t_L g1298 ( 
.A1(n_1174),
.A2(n_812),
.B(n_597),
.C(n_601),
.Y(n_1298)
);

OAI22xp5_ASAP7_75t_L g1299 ( 
.A1(n_1107),
.A2(n_600),
.B1(n_1033),
.B2(n_1151),
.Y(n_1299)
);

NOR2xp33_ASAP7_75t_L g1300 ( 
.A(n_1174),
.B(n_1045),
.Y(n_1300)
);

OAI21x1_ASAP7_75t_L g1301 ( 
.A1(n_1104),
.A2(n_1160),
.B(n_1146),
.Y(n_1301)
);

OAI21x1_ASAP7_75t_L g1302 ( 
.A1(n_1104),
.A2(n_1160),
.B(n_1146),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_L g1303 ( 
.A(n_1151),
.B(n_1162),
.Y(n_1303)
);

OAI21x1_ASAP7_75t_L g1304 ( 
.A1(n_1104),
.A2(n_1160),
.B(n_1146),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1071),
.Y(n_1305)
);

BUFx3_ASAP7_75t_L g1306 ( 
.A(n_1180),
.Y(n_1306)
);

BUFx3_ASAP7_75t_L g1307 ( 
.A(n_1180),
.Y(n_1307)
);

INVxp67_ASAP7_75t_L g1308 ( 
.A(n_1195),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_1151),
.B(n_1162),
.Y(n_1309)
);

INVx1_ASAP7_75t_SL g1310 ( 
.A(n_1154),
.Y(n_1310)
);

CKINVDCx20_ASAP7_75t_R g1311 ( 
.A(n_1136),
.Y(n_1311)
);

CKINVDCx5p33_ASAP7_75t_R g1312 ( 
.A(n_1154),
.Y(n_1312)
);

INVx2_ASAP7_75t_L g1313 ( 
.A(n_1071),
.Y(n_1313)
);

INVx3_ASAP7_75t_L g1314 ( 
.A(n_1149),
.Y(n_1314)
);

AOI21xp5_ASAP7_75t_L g1315 ( 
.A1(n_1094),
.A2(n_1191),
.B(n_1157),
.Y(n_1315)
);

AO21x2_ASAP7_75t_L g1316 ( 
.A1(n_1157),
.A2(n_1194),
.B(n_1191),
.Y(n_1316)
);

AND2x4_ASAP7_75t_L g1317 ( 
.A(n_1169),
.B(n_1065),
.Y(n_1317)
);

AOI22xp5_ASAP7_75t_L g1318 ( 
.A1(n_1174),
.A2(n_307),
.B1(n_328),
.B2(n_304),
.Y(n_1318)
);

BUFx3_ASAP7_75t_L g1319 ( 
.A(n_1180),
.Y(n_1319)
);

O2A1O1Ixp33_ASAP7_75t_L g1320 ( 
.A1(n_1192),
.A2(n_1101),
.B(n_1174),
.C(n_1173),
.Y(n_1320)
);

AO31x2_ASAP7_75t_L g1321 ( 
.A1(n_1092),
.A2(n_1184),
.A3(n_1191),
.B(n_1157),
.Y(n_1321)
);

NOR2xp67_ASAP7_75t_L g1322 ( 
.A(n_1171),
.B(n_999),
.Y(n_1322)
);

AOI221x1_ASAP7_75t_SL g1323 ( 
.A1(n_1298),
.A2(n_1300),
.B1(n_1273),
.B2(n_1215),
.C(n_1299),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1255),
.Y(n_1324)
);

AND2x2_ASAP7_75t_L g1325 ( 
.A(n_1300),
.B(n_1258),
.Y(n_1325)
);

INVx2_ASAP7_75t_L g1326 ( 
.A(n_1200),
.Y(n_1326)
);

NOR2xp67_ASAP7_75t_L g1327 ( 
.A(n_1282),
.B(n_1224),
.Y(n_1327)
);

HB1xp67_ASAP7_75t_L g1328 ( 
.A(n_1265),
.Y(n_1328)
);

NAND2xp5_ASAP7_75t_L g1329 ( 
.A(n_1213),
.B(n_1215),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1218),
.Y(n_1330)
);

AND2x2_ASAP7_75t_SL g1331 ( 
.A(n_1199),
.B(n_1238),
.Y(n_1331)
);

AOI221x1_ASAP7_75t_SL g1332 ( 
.A1(n_1299),
.A2(n_1322),
.B1(n_1289),
.B2(n_1239),
.C(n_1241),
.Y(n_1332)
);

AND2x2_ASAP7_75t_L g1333 ( 
.A(n_1223),
.B(n_1211),
.Y(n_1333)
);

OAI22xp5_ASAP7_75t_L g1334 ( 
.A1(n_1294),
.A2(n_1318),
.B1(n_1205),
.B2(n_1264),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1220),
.Y(n_1335)
);

CKINVDCx16_ASAP7_75t_R g1336 ( 
.A(n_1253),
.Y(n_1336)
);

HB1xp67_ASAP7_75t_L g1337 ( 
.A(n_1265),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_L g1338 ( 
.A(n_1283),
.B(n_1226),
.Y(n_1338)
);

AOI21x1_ASAP7_75t_SL g1339 ( 
.A1(n_1247),
.A2(n_1226),
.B(n_1293),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1227),
.Y(n_1340)
);

NAND2xp33_ASAP7_75t_SL g1341 ( 
.A(n_1275),
.B(n_1312),
.Y(n_1341)
);

CKINVDCx5p33_ASAP7_75t_R g1342 ( 
.A(n_1253),
.Y(n_1342)
);

AND2x4_ASAP7_75t_L g1343 ( 
.A(n_1249),
.B(n_1222),
.Y(n_1343)
);

AND2x2_ASAP7_75t_L g1344 ( 
.A(n_1254),
.B(n_1317),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_L g1345 ( 
.A(n_1208),
.B(n_1209),
.Y(n_1345)
);

OAI22xp5_ASAP7_75t_L g1346 ( 
.A1(n_1205),
.A2(n_1264),
.B1(n_1225),
.B2(n_1198),
.Y(n_1346)
);

AOI211xp5_ASAP7_75t_L g1347 ( 
.A1(n_1198),
.A2(n_1276),
.B(n_1320),
.C(n_1277),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_L g1348 ( 
.A(n_1208),
.B(n_1209),
.Y(n_1348)
);

HB1xp67_ASAP7_75t_L g1349 ( 
.A(n_1270),
.Y(n_1349)
);

AOI21x1_ASAP7_75t_SL g1350 ( 
.A1(n_1247),
.A2(n_1309),
.B(n_1303),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_L g1351 ( 
.A(n_1293),
.B(n_1303),
.Y(n_1351)
);

OAI22xp5_ASAP7_75t_L g1352 ( 
.A1(n_1225),
.A2(n_1268),
.B1(n_1263),
.B2(n_1248),
.Y(n_1352)
);

AND2x4_ASAP7_75t_L g1353 ( 
.A(n_1249),
.B(n_1222),
.Y(n_1353)
);

O2A1O1Ixp33_ASAP7_75t_L g1354 ( 
.A1(n_1276),
.A2(n_1320),
.B(n_1248),
.C(n_1202),
.Y(n_1354)
);

O2A1O1Ixp5_ASAP7_75t_L g1355 ( 
.A1(n_1287),
.A2(n_1267),
.B(n_1315),
.C(n_1203),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1236),
.Y(n_1356)
);

OA21x2_ASAP7_75t_L g1357 ( 
.A1(n_1237),
.A2(n_1257),
.B(n_1251),
.Y(n_1357)
);

AOI21xp5_ASAP7_75t_SL g1358 ( 
.A1(n_1201),
.A2(n_1256),
.B(n_1221),
.Y(n_1358)
);

OAI22xp5_ASAP7_75t_SL g1359 ( 
.A1(n_1311),
.A2(n_1231),
.B1(n_1310),
.B2(n_1268),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1244),
.Y(n_1360)
);

AND2x2_ASAP7_75t_L g1361 ( 
.A(n_1252),
.B(n_1222),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_L g1362 ( 
.A(n_1240),
.B(n_1207),
.Y(n_1362)
);

OA21x2_ASAP7_75t_L g1363 ( 
.A1(n_1242),
.A2(n_1245),
.B(n_1229),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1246),
.Y(n_1364)
);

AOI21xp5_ASAP7_75t_L g1365 ( 
.A1(n_1316),
.A2(n_1201),
.B(n_1286),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1250),
.Y(n_1366)
);

HB1xp67_ASAP7_75t_L g1367 ( 
.A(n_1291),
.Y(n_1367)
);

A2O1A1Ixp33_ASAP7_75t_L g1368 ( 
.A1(n_1199),
.A2(n_1217),
.B(n_1204),
.C(n_1305),
.Y(n_1368)
);

BUFx2_ASAP7_75t_L g1369 ( 
.A(n_1281),
.Y(n_1369)
);

NOR2xp67_ASAP7_75t_L g1370 ( 
.A(n_1261),
.B(n_1308),
.Y(n_1370)
);

OR2x2_ASAP7_75t_L g1371 ( 
.A(n_1308),
.B(n_1284),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_L g1372 ( 
.A(n_1216),
.B(n_1313),
.Y(n_1372)
);

OAI22xp5_ASAP7_75t_L g1373 ( 
.A1(n_1269),
.A2(n_1243),
.B1(n_1279),
.B2(n_1280),
.Y(n_1373)
);

BUFx3_ASAP7_75t_L g1374 ( 
.A(n_1272),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1210),
.Y(n_1375)
);

AND2x2_ASAP7_75t_L g1376 ( 
.A(n_1285),
.B(n_1290),
.Y(n_1376)
);

AOI21xp5_ASAP7_75t_SL g1377 ( 
.A1(n_1272),
.A2(n_1295),
.B(n_1306),
.Y(n_1377)
);

BUFx3_ASAP7_75t_L g1378 ( 
.A(n_1278),
.Y(n_1378)
);

AOI221xp5_ASAP7_75t_L g1379 ( 
.A1(n_1262),
.A2(n_1232),
.B1(n_1212),
.B2(n_1296),
.C(n_1297),
.Y(n_1379)
);

NAND2x1_ASAP7_75t_L g1380 ( 
.A(n_1269),
.B(n_1279),
.Y(n_1380)
);

AND2x2_ASAP7_75t_L g1381 ( 
.A(n_1314),
.B(n_1243),
.Y(n_1381)
);

AOI21x1_ASAP7_75t_SL g1382 ( 
.A1(n_1235),
.A2(n_1288),
.B(n_1274),
.Y(n_1382)
);

BUFx12f_ASAP7_75t_L g1383 ( 
.A(n_1228),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1260),
.Y(n_1384)
);

AOI21xp5_ASAP7_75t_SL g1385 ( 
.A1(n_1278),
.A2(n_1295),
.B(n_1306),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1234),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_L g1387 ( 
.A(n_1206),
.B(n_1314),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_L g1388 ( 
.A(n_1233),
.B(n_1319),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_L g1389 ( 
.A(n_1307),
.B(n_1319),
.Y(n_1389)
);

AND2x2_ASAP7_75t_L g1390 ( 
.A(n_1307),
.B(n_1288),
.Y(n_1390)
);

AOI21xp5_ASAP7_75t_SL g1391 ( 
.A1(n_1219),
.A2(n_1271),
.B(n_1274),
.Y(n_1391)
);

O2A1O1Ixp5_ASAP7_75t_L g1392 ( 
.A1(n_1291),
.A2(n_1321),
.B(n_1292),
.C(n_1235),
.Y(n_1392)
);

AND2x2_ASAP7_75t_L g1393 ( 
.A(n_1271),
.B(n_1321),
.Y(n_1393)
);

CKINVDCx5p33_ASAP7_75t_R g1394 ( 
.A(n_1311),
.Y(n_1394)
);

AOI21xp5_ASAP7_75t_SL g1395 ( 
.A1(n_1259),
.A2(n_1228),
.B(n_1214),
.Y(n_1395)
);

AND2x2_ASAP7_75t_L g1396 ( 
.A(n_1321),
.B(n_1292),
.Y(n_1396)
);

NAND2xp5_ASAP7_75t_L g1397 ( 
.A(n_1214),
.B(n_1292),
.Y(n_1397)
);

OA21x2_ASAP7_75t_L g1398 ( 
.A1(n_1301),
.A2(n_1302),
.B(n_1304),
.Y(n_1398)
);

NOR2xp33_ASAP7_75t_L g1399 ( 
.A(n_1266),
.B(n_1230),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_L g1400 ( 
.A(n_1213),
.B(n_1215),
.Y(n_1400)
);

BUFx3_ASAP7_75t_L g1401 ( 
.A(n_1272),
.Y(n_1401)
);

O2A1O1Ixp33_ASAP7_75t_L g1402 ( 
.A1(n_1298),
.A2(n_1174),
.B(n_1192),
.C(n_1101),
.Y(n_1402)
);

CKINVDCx5p33_ASAP7_75t_R g1403 ( 
.A(n_1275),
.Y(n_1403)
);

AOI221x1_ASAP7_75t_SL g1404 ( 
.A1(n_1298),
.A2(n_602),
.B1(n_607),
.B2(n_952),
.C(n_1300),
.Y(n_1404)
);

A2O1A1Ixp33_ASAP7_75t_L g1405 ( 
.A1(n_1201),
.A2(n_1294),
.B(n_1298),
.C(n_1276),
.Y(n_1405)
);

AOI211xp5_ASAP7_75t_L g1406 ( 
.A1(n_1298),
.A2(n_1174),
.B(n_812),
.C(n_741),
.Y(n_1406)
);

OA21x2_ASAP7_75t_L g1407 ( 
.A1(n_1237),
.A2(n_1257),
.B(n_1251),
.Y(n_1407)
);

AOI21xp5_ASAP7_75t_SL g1408 ( 
.A1(n_1248),
.A2(n_1173),
.B(n_609),
.Y(n_1408)
);

NAND2xp5_ASAP7_75t_L g1409 ( 
.A(n_1213),
.B(n_1215),
.Y(n_1409)
);

A2O1A1Ixp33_ASAP7_75t_SL g1410 ( 
.A1(n_1298),
.A2(n_1287),
.B(n_1277),
.C(n_1198),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1255),
.Y(n_1411)
);

INVx2_ASAP7_75t_L g1412 ( 
.A(n_1324),
.Y(n_1412)
);

AND2x2_ASAP7_75t_L g1413 ( 
.A(n_1393),
.B(n_1396),
.Y(n_1413)
);

OA21x2_ASAP7_75t_L g1414 ( 
.A1(n_1355),
.A2(n_1392),
.B(n_1365),
.Y(n_1414)
);

OR2x6_ASAP7_75t_L g1415 ( 
.A(n_1391),
.B(n_1395),
.Y(n_1415)
);

NOR2xp33_ASAP7_75t_L g1416 ( 
.A(n_1387),
.B(n_1333),
.Y(n_1416)
);

AND2x4_ASAP7_75t_L g1417 ( 
.A(n_1386),
.B(n_1390),
.Y(n_1417)
);

BUFx6f_ASAP7_75t_L g1418 ( 
.A(n_1357),
.Y(n_1418)
);

OR2x2_ASAP7_75t_L g1419 ( 
.A(n_1397),
.B(n_1411),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_L g1420 ( 
.A(n_1329),
.B(n_1400),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1409),
.B(n_1347),
.Y(n_1421)
);

AND2x4_ASAP7_75t_L g1422 ( 
.A(n_1384),
.B(n_1380),
.Y(n_1422)
);

HB1xp67_ASAP7_75t_L g1423 ( 
.A(n_1328),
.Y(n_1423)
);

INVx2_ASAP7_75t_L g1424 ( 
.A(n_1357),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1330),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1335),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1340),
.Y(n_1427)
);

AND2x2_ASAP7_75t_L g1428 ( 
.A(n_1367),
.B(n_1407),
.Y(n_1428)
);

OR2x6_ASAP7_75t_L g1429 ( 
.A(n_1408),
.B(n_1358),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1356),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1360),
.Y(n_1431)
);

AND2x2_ASAP7_75t_L g1432 ( 
.A(n_1363),
.B(n_1349),
.Y(n_1432)
);

BUFx2_ASAP7_75t_L g1433 ( 
.A(n_1337),
.Y(n_1433)
);

INVxp67_ASAP7_75t_L g1434 ( 
.A(n_1364),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_L g1435 ( 
.A(n_1331),
.B(n_1345),
.Y(n_1435)
);

AND2x4_ASAP7_75t_L g1436 ( 
.A(n_1343),
.B(n_1353),
.Y(n_1436)
);

OR2x2_ASAP7_75t_L g1437 ( 
.A(n_1338),
.B(n_1346),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1375),
.Y(n_1438)
);

AO21x1_ASAP7_75t_L g1439 ( 
.A1(n_1334),
.A2(n_1354),
.B(n_1352),
.Y(n_1439)
);

AO21x2_ASAP7_75t_L g1440 ( 
.A1(n_1410),
.A2(n_1399),
.B(n_1368),
.Y(n_1440)
);

HB1xp67_ASAP7_75t_L g1441 ( 
.A(n_1399),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1366),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1326),
.Y(n_1443)
);

OA21x2_ASAP7_75t_L g1444 ( 
.A1(n_1368),
.A2(n_1405),
.B(n_1382),
.Y(n_1444)
);

AND2x2_ASAP7_75t_L g1445 ( 
.A(n_1331),
.B(n_1325),
.Y(n_1445)
);

AO21x2_ASAP7_75t_L g1446 ( 
.A1(n_1410),
.A2(n_1405),
.B(n_1402),
.Y(n_1446)
);

NOR2xp33_ASAP7_75t_L g1447 ( 
.A(n_1344),
.B(n_1403),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1372),
.Y(n_1448)
);

OR2x2_ASAP7_75t_L g1449 ( 
.A(n_1371),
.B(n_1362),
.Y(n_1449)
);

AND2x2_ASAP7_75t_L g1450 ( 
.A(n_1398),
.B(n_1376),
.Y(n_1450)
);

AO21x2_ASAP7_75t_L g1451 ( 
.A1(n_1373),
.A2(n_1351),
.B(n_1348),
.Y(n_1451)
);

AO21x2_ASAP7_75t_L g1452 ( 
.A1(n_1339),
.A2(n_1350),
.B(n_1327),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1412),
.Y(n_1453)
);

OR2x2_ASAP7_75t_L g1454 ( 
.A(n_1419),
.B(n_1441),
.Y(n_1454)
);

AND2x2_ASAP7_75t_L g1455 ( 
.A(n_1450),
.B(n_1413),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1412),
.Y(n_1456)
);

OAI221xp5_ASAP7_75t_L g1457 ( 
.A1(n_1421),
.A2(n_1406),
.B1(n_1404),
.B2(n_1323),
.C(n_1332),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_L g1458 ( 
.A(n_1420),
.B(n_1451),
.Y(n_1458)
);

BUFx6f_ASAP7_75t_L g1459 ( 
.A(n_1418),
.Y(n_1459)
);

NOR2x1_ASAP7_75t_L g1460 ( 
.A(n_1429),
.B(n_1385),
.Y(n_1460)
);

INVx2_ASAP7_75t_L g1461 ( 
.A(n_1424),
.Y(n_1461)
);

OR2x2_ASAP7_75t_L g1462 ( 
.A(n_1419),
.B(n_1369),
.Y(n_1462)
);

AND2x2_ASAP7_75t_L g1463 ( 
.A(n_1413),
.B(n_1361),
.Y(n_1463)
);

AND2x2_ASAP7_75t_L g1464 ( 
.A(n_1413),
.B(n_1381),
.Y(n_1464)
);

BUFx2_ASAP7_75t_L g1465 ( 
.A(n_1422),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_L g1466 ( 
.A(n_1420),
.B(n_1379),
.Y(n_1466)
);

NAND2xp5_ASAP7_75t_L g1467 ( 
.A(n_1451),
.B(n_1370),
.Y(n_1467)
);

OR2x2_ASAP7_75t_L g1468 ( 
.A(n_1441),
.B(n_1433),
.Y(n_1468)
);

INVxp67_ASAP7_75t_SL g1469 ( 
.A(n_1423),
.Y(n_1469)
);

AND2x2_ASAP7_75t_L g1470 ( 
.A(n_1432),
.B(n_1401),
.Y(n_1470)
);

NOR2xp33_ASAP7_75t_SL g1471 ( 
.A(n_1429),
.B(n_1336),
.Y(n_1471)
);

BUFx3_ASAP7_75t_L g1472 ( 
.A(n_1422),
.Y(n_1472)
);

OR2x2_ASAP7_75t_L g1473 ( 
.A(n_1428),
.B(n_1389),
.Y(n_1473)
);

AND2x4_ASAP7_75t_L g1474 ( 
.A(n_1422),
.B(n_1374),
.Y(n_1474)
);

BUFx2_ASAP7_75t_L g1475 ( 
.A(n_1433),
.Y(n_1475)
);

AOI22xp33_ASAP7_75t_SL g1476 ( 
.A1(n_1471),
.A2(n_1446),
.B1(n_1429),
.B2(n_1421),
.Y(n_1476)
);

INVx2_ASAP7_75t_L g1477 ( 
.A(n_1461),
.Y(n_1477)
);

AOI33xp33_ASAP7_75t_L g1478 ( 
.A1(n_1470),
.A2(n_1445),
.A3(n_1431),
.B1(n_1430),
.B2(n_1426),
.B3(n_1425),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_L g1479 ( 
.A(n_1458),
.B(n_1451),
.Y(n_1479)
);

AND2x4_ASAP7_75t_L g1480 ( 
.A(n_1472),
.B(n_1415),
.Y(n_1480)
);

OAI22xp5_ASAP7_75t_L g1481 ( 
.A1(n_1457),
.A2(n_1429),
.B1(n_1435),
.B2(n_1437),
.Y(n_1481)
);

INVx3_ASAP7_75t_L g1482 ( 
.A(n_1459),
.Y(n_1482)
);

AOI33xp33_ASAP7_75t_L g1483 ( 
.A1(n_1470),
.A2(n_1445),
.A3(n_1431),
.B1(n_1430),
.B2(n_1426),
.B3(n_1425),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1453),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_L g1485 ( 
.A(n_1458),
.B(n_1451),
.Y(n_1485)
);

OAI211xp5_ASAP7_75t_L g1486 ( 
.A1(n_1457),
.A2(n_1435),
.B(n_1437),
.C(n_1445),
.Y(n_1486)
);

BUFx8_ASAP7_75t_L g1487 ( 
.A(n_1475),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1453),
.Y(n_1488)
);

INVxp67_ASAP7_75t_SL g1489 ( 
.A(n_1467),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1453),
.Y(n_1490)
);

AOI211xp5_ASAP7_75t_SL g1491 ( 
.A1(n_1471),
.A2(n_1377),
.B(n_1359),
.C(n_1439),
.Y(n_1491)
);

AND2x2_ASAP7_75t_L g1492 ( 
.A(n_1455),
.B(n_1417),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1456),
.Y(n_1493)
);

NAND2xp33_ASAP7_75t_R g1494 ( 
.A(n_1466),
.B(n_1342),
.Y(n_1494)
);

NOR2x1_ASAP7_75t_L g1495 ( 
.A(n_1460),
.B(n_1429),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1456),
.Y(n_1496)
);

AND2x4_ASAP7_75t_L g1497 ( 
.A(n_1472),
.B(n_1415),
.Y(n_1497)
);

OAI221xp5_ASAP7_75t_L g1498 ( 
.A1(n_1466),
.A2(n_1416),
.B1(n_1388),
.B2(n_1449),
.C(n_1415),
.Y(n_1498)
);

AOI22xp33_ASAP7_75t_L g1499 ( 
.A1(n_1460),
.A2(n_1439),
.B1(n_1446),
.B2(n_1440),
.Y(n_1499)
);

OAI33xp33_ASAP7_75t_L g1500 ( 
.A1(n_1454),
.A2(n_1434),
.A3(n_1449),
.B1(n_1427),
.B2(n_1438),
.B3(n_1442),
.Y(n_1500)
);

BUFx3_ASAP7_75t_L g1501 ( 
.A(n_1474),
.Y(n_1501)
);

AOI221xp5_ASAP7_75t_L g1502 ( 
.A1(n_1469),
.A2(n_1446),
.B1(n_1440),
.B2(n_1434),
.C(n_1448),
.Y(n_1502)
);

AND2x2_ASAP7_75t_L g1503 ( 
.A(n_1455),
.B(n_1417),
.Y(n_1503)
);

OAI321xp33_ASAP7_75t_L g1504 ( 
.A1(n_1473),
.A2(n_1446),
.A3(n_1415),
.B1(n_1442),
.B2(n_1448),
.C(n_1443),
.Y(n_1504)
);

NOR2xp33_ASAP7_75t_R g1505 ( 
.A(n_1462),
.B(n_1394),
.Y(n_1505)
);

INVx5_ASAP7_75t_SL g1506 ( 
.A(n_1459),
.Y(n_1506)
);

BUFx3_ASAP7_75t_L g1507 ( 
.A(n_1474),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1484),
.Y(n_1508)
);

AND2x2_ASAP7_75t_L g1509 ( 
.A(n_1492),
.B(n_1455),
.Y(n_1509)
);

INVx3_ASAP7_75t_L g1510 ( 
.A(n_1506),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_L g1511 ( 
.A(n_1479),
.B(n_1454),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1484),
.Y(n_1512)
);

HB1xp67_ASAP7_75t_L g1513 ( 
.A(n_1488),
.Y(n_1513)
);

OAI21xp5_ASAP7_75t_SL g1514 ( 
.A1(n_1491),
.A2(n_1447),
.B(n_1436),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1488),
.Y(n_1515)
);

INVx2_ASAP7_75t_L g1516 ( 
.A(n_1477),
.Y(n_1516)
);

NAND3xp33_ASAP7_75t_L g1517 ( 
.A(n_1502),
.B(n_1444),
.C(n_1414),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1490),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1490),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1493),
.Y(n_1520)
);

BUFx3_ASAP7_75t_L g1521 ( 
.A(n_1487),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1492),
.B(n_1503),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_SL g1523 ( 
.A(n_1476),
.B(n_1474),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_L g1524 ( 
.A(n_1485),
.B(n_1454),
.Y(n_1524)
);

AND2x2_ASAP7_75t_L g1525 ( 
.A(n_1503),
.B(n_1455),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1493),
.Y(n_1526)
);

INVx4_ASAP7_75t_L g1527 ( 
.A(n_1480),
.Y(n_1527)
);

AOI21xp5_ASAP7_75t_L g1528 ( 
.A1(n_1504),
.A2(n_1444),
.B(n_1440),
.Y(n_1528)
);

BUFx2_ASAP7_75t_L g1529 ( 
.A(n_1487),
.Y(n_1529)
);

OAI21xp5_ASAP7_75t_SL g1530 ( 
.A1(n_1491),
.A2(n_1436),
.B(n_1474),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1496),
.Y(n_1531)
);

NAND3xp33_ASAP7_75t_L g1532 ( 
.A(n_1499),
.B(n_1444),
.C(n_1414),
.Y(n_1532)
);

OR2x2_ASAP7_75t_L g1533 ( 
.A(n_1511),
.B(n_1524),
.Y(n_1533)
);

AND2x2_ASAP7_75t_L g1534 ( 
.A(n_1522),
.B(n_1501),
.Y(n_1534)
);

AND2x2_ASAP7_75t_L g1535 ( 
.A(n_1522),
.B(n_1501),
.Y(n_1535)
);

AND2x2_ASAP7_75t_L g1536 ( 
.A(n_1522),
.B(n_1507),
.Y(n_1536)
);

INVx2_ASAP7_75t_L g1537 ( 
.A(n_1516),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1513),
.Y(n_1538)
);

HB1xp67_ASAP7_75t_L g1539 ( 
.A(n_1513),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1508),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1508),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1512),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1512),
.Y(n_1543)
);

CKINVDCx5p33_ASAP7_75t_R g1544 ( 
.A(n_1529),
.Y(n_1544)
);

AND2x2_ASAP7_75t_L g1545 ( 
.A(n_1527),
.B(n_1507),
.Y(n_1545)
);

AND2x2_ASAP7_75t_L g1546 ( 
.A(n_1527),
.B(n_1489),
.Y(n_1546)
);

BUFx2_ASAP7_75t_L g1547 ( 
.A(n_1529),
.Y(n_1547)
);

INVx2_ASAP7_75t_L g1548 ( 
.A(n_1516),
.Y(n_1548)
);

AND2x4_ASAP7_75t_SL g1549 ( 
.A(n_1510),
.B(n_1527),
.Y(n_1549)
);

OR2x2_ASAP7_75t_L g1550 ( 
.A(n_1511),
.B(n_1468),
.Y(n_1550)
);

AOI221xp5_ASAP7_75t_L g1551 ( 
.A1(n_1523),
.A2(n_1481),
.B1(n_1486),
.B2(n_1498),
.C(n_1500),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_L g1552 ( 
.A(n_1529),
.B(n_1478),
.Y(n_1552)
);

AND2x4_ASAP7_75t_L g1553 ( 
.A(n_1527),
.B(n_1480),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1515),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1527),
.B(n_1509),
.Y(n_1555)
);

AND2x2_ASAP7_75t_L g1556 ( 
.A(n_1509),
.B(n_1480),
.Y(n_1556)
);

AND2x2_ASAP7_75t_L g1557 ( 
.A(n_1509),
.B(n_1525),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1525),
.B(n_1480),
.Y(n_1558)
);

NAND4xp25_ASAP7_75t_L g1559 ( 
.A(n_1517),
.B(n_1494),
.C(n_1495),
.D(n_1483),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1525),
.B(n_1497),
.Y(n_1560)
);

AND2x2_ASAP7_75t_L g1561 ( 
.A(n_1510),
.B(n_1497),
.Y(n_1561)
);

AND2x2_ASAP7_75t_L g1562 ( 
.A(n_1510),
.B(n_1497),
.Y(n_1562)
);

INVx2_ASAP7_75t_L g1563 ( 
.A(n_1516),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1515),
.Y(n_1564)
);

AOI22xp33_ASAP7_75t_L g1565 ( 
.A1(n_1523),
.A2(n_1495),
.B1(n_1440),
.B2(n_1497),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1518),
.Y(n_1566)
);

AND3x1_ASAP7_75t_L g1567 ( 
.A(n_1514),
.B(n_1482),
.C(n_1505),
.Y(n_1567)
);

NOR3xp33_ASAP7_75t_L g1568 ( 
.A(n_1514),
.B(n_1341),
.C(n_1482),
.Y(n_1568)
);

NAND2xp5_ASAP7_75t_L g1569 ( 
.A(n_1524),
.B(n_1464),
.Y(n_1569)
);

AOI22xp5_ASAP7_75t_L g1570 ( 
.A1(n_1530),
.A2(n_1444),
.B1(n_1415),
.B2(n_1452),
.Y(n_1570)
);

OAI221xp5_ASAP7_75t_SL g1571 ( 
.A1(n_1530),
.A2(n_1517),
.B1(n_1528),
.B2(n_1532),
.C(n_1521),
.Y(n_1571)
);

NAND4xp25_ASAP7_75t_L g1572 ( 
.A(n_1528),
.B(n_1374),
.C(n_1378),
.D(n_1473),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_L g1573 ( 
.A(n_1521),
.B(n_1464),
.Y(n_1573)
);

NOR2xp33_ASAP7_75t_L g1574 ( 
.A(n_1521),
.B(n_1383),
.Y(n_1574)
);

INVx3_ASAP7_75t_SL g1575 ( 
.A(n_1544),
.Y(n_1575)
);

AND2x4_ASAP7_75t_L g1576 ( 
.A(n_1547),
.B(n_1521),
.Y(n_1576)
);

OR2x2_ASAP7_75t_L g1577 ( 
.A(n_1533),
.B(n_1518),
.Y(n_1577)
);

HB1xp67_ASAP7_75t_L g1578 ( 
.A(n_1547),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_L g1579 ( 
.A(n_1551),
.B(n_1464),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1540),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1540),
.Y(n_1581)
);

AND2x2_ASAP7_75t_L g1582 ( 
.A(n_1567),
.B(n_1510),
.Y(n_1582)
);

AND2x4_ASAP7_75t_L g1583 ( 
.A(n_1549),
.B(n_1510),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1552),
.B(n_1464),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1541),
.Y(n_1585)
);

OR2x2_ASAP7_75t_L g1586 ( 
.A(n_1533),
.B(n_1519),
.Y(n_1586)
);

INVx2_ASAP7_75t_L g1587 ( 
.A(n_1557),
.Y(n_1587)
);

AND2x2_ASAP7_75t_L g1588 ( 
.A(n_1567),
.B(n_1506),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1541),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1559),
.B(n_1463),
.Y(n_1590)
);

NOR2x1_ASAP7_75t_L g1591 ( 
.A(n_1559),
.B(n_1378),
.Y(n_1591)
);

OR2x6_ASAP7_75t_L g1592 ( 
.A(n_1574),
.B(n_1415),
.Y(n_1592)
);

OAI21xp33_ASAP7_75t_L g1593 ( 
.A1(n_1571),
.A2(n_1532),
.B(n_1473),
.Y(n_1593)
);

OR2x2_ASAP7_75t_L g1594 ( 
.A(n_1550),
.B(n_1569),
.Y(n_1594)
);

AOI221xp5_ASAP7_75t_L g1595 ( 
.A1(n_1565),
.A2(n_1526),
.B1(n_1519),
.B2(n_1520),
.C(n_1531),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_L g1596 ( 
.A(n_1573),
.B(n_1546),
.Y(n_1596)
);

INVx2_ASAP7_75t_L g1597 ( 
.A(n_1557),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1561),
.B(n_1506),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1542),
.Y(n_1599)
);

AND2x4_ASAP7_75t_L g1600 ( 
.A(n_1549),
.B(n_1520),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1542),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1543),
.Y(n_1602)
);

AND2x2_ASAP7_75t_L g1603 ( 
.A(n_1561),
.B(n_1506),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1543),
.Y(n_1604)
);

INVx2_ASAP7_75t_L g1605 ( 
.A(n_1537),
.Y(n_1605)
);

AND2x2_ASAP7_75t_L g1606 ( 
.A(n_1562),
.B(n_1465),
.Y(n_1606)
);

INVx3_ASAP7_75t_L g1607 ( 
.A(n_1549),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_L g1608 ( 
.A(n_1546),
.B(n_1463),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1554),
.Y(n_1609)
);

CKINVDCx16_ASAP7_75t_R g1610 ( 
.A(n_1576),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_L g1611 ( 
.A(n_1578),
.B(n_1568),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1582),
.B(n_1562),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1580),
.Y(n_1613)
);

INVx2_ASAP7_75t_L g1614 ( 
.A(n_1587),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1581),
.Y(n_1615)
);

BUFx2_ASAP7_75t_L g1616 ( 
.A(n_1607),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1585),
.Y(n_1617)
);

OAI21x1_ASAP7_75t_L g1618 ( 
.A1(n_1591),
.A2(n_1538),
.B(n_1537),
.Y(n_1618)
);

INVx2_ASAP7_75t_SL g1619 ( 
.A(n_1607),
.Y(n_1619)
);

INVx1_ASAP7_75t_SL g1620 ( 
.A(n_1575),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1589),
.Y(n_1621)
);

AND2x4_ASAP7_75t_L g1622 ( 
.A(n_1607),
.B(n_1555),
.Y(n_1622)
);

BUFx3_ASAP7_75t_L g1623 ( 
.A(n_1575),
.Y(n_1623)
);

OR2x2_ASAP7_75t_L g1624 ( 
.A(n_1587),
.B(n_1550),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1599),
.Y(n_1625)
);

INVx2_ASAP7_75t_L g1626 ( 
.A(n_1600),
.Y(n_1626)
);

INVx2_ASAP7_75t_L g1627 ( 
.A(n_1597),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1579),
.B(n_1534),
.Y(n_1628)
);

AOI22xp33_ASAP7_75t_L g1629 ( 
.A1(n_1593),
.A2(n_1572),
.B1(n_1553),
.B2(n_1570),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1582),
.B(n_1555),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1601),
.Y(n_1631)
);

OR2x2_ASAP7_75t_L g1632 ( 
.A(n_1597),
.B(n_1539),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1576),
.B(n_1556),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1602),
.Y(n_1634)
);

A2O1A1Ixp33_ASAP7_75t_L g1635 ( 
.A1(n_1618),
.A2(n_1595),
.B(n_1590),
.C(n_1588),
.Y(n_1635)
);

HB1xp67_ASAP7_75t_L g1636 ( 
.A(n_1616),
.Y(n_1636)
);

OAI211xp5_ASAP7_75t_L g1637 ( 
.A1(n_1629),
.A2(n_1572),
.B(n_1570),
.C(n_1588),
.Y(n_1637)
);

OAI22xp33_ASAP7_75t_L g1638 ( 
.A1(n_1610),
.A2(n_1592),
.B1(n_1596),
.B2(n_1584),
.Y(n_1638)
);

OAI31xp33_ASAP7_75t_L g1639 ( 
.A1(n_1620),
.A2(n_1576),
.A3(n_1583),
.B(n_1600),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1614),
.Y(n_1640)
);

OAI322xp33_ASAP7_75t_L g1641 ( 
.A1(n_1611),
.A2(n_1609),
.A3(n_1604),
.B1(n_1577),
.B2(n_1586),
.C1(n_1594),
.C2(n_1538),
.Y(n_1641)
);

NOR2x1_ASAP7_75t_L g1642 ( 
.A(n_1623),
.B(n_1583),
.Y(n_1642)
);

AND2x2_ASAP7_75t_SL g1643 ( 
.A(n_1610),
.B(n_1583),
.Y(n_1643)
);

OAI221xp5_ASAP7_75t_L g1644 ( 
.A1(n_1623),
.A2(n_1592),
.B1(n_1603),
.B2(n_1598),
.C(n_1594),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_L g1645 ( 
.A(n_1616),
.B(n_1608),
.Y(n_1645)
);

OR2x2_ASAP7_75t_L g1646 ( 
.A(n_1628),
.B(n_1577),
.Y(n_1646)
);

AND2x2_ASAP7_75t_SL g1647 ( 
.A(n_1626),
.B(n_1600),
.Y(n_1647)
);

AOI22xp33_ASAP7_75t_L g1648 ( 
.A1(n_1623),
.A2(n_1592),
.B1(n_1603),
.B2(n_1598),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1614),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1614),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1627),
.Y(n_1651)
);

NOR2x1_ASAP7_75t_L g1652 ( 
.A(n_1626),
.B(n_1605),
.Y(n_1652)
);

CKINVDCx20_ASAP7_75t_R g1653 ( 
.A(n_1633),
.Y(n_1653)
);

INVx1_ASAP7_75t_SL g1654 ( 
.A(n_1643),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1636),
.Y(n_1655)
);

AND2x4_ASAP7_75t_L g1656 ( 
.A(n_1642),
.B(n_1619),
.Y(n_1656)
);

NAND2x1_ASAP7_75t_SL g1657 ( 
.A(n_1636),
.B(n_1622),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1640),
.Y(n_1658)
);

HB1xp67_ASAP7_75t_L g1659 ( 
.A(n_1652),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_L g1660 ( 
.A(n_1643),
.B(n_1612),
.Y(n_1660)
);

INVx1_ASAP7_75t_SL g1661 ( 
.A(n_1653),
.Y(n_1661)
);

NOR2xp33_ASAP7_75t_SL g1662 ( 
.A(n_1639),
.B(n_1619),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1649),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1650),
.Y(n_1664)
);

AOI22xp33_ASAP7_75t_L g1665 ( 
.A1(n_1662),
.A2(n_1644),
.B1(n_1641),
.B2(n_1612),
.Y(n_1665)
);

AOI211xp5_ASAP7_75t_L g1666 ( 
.A1(n_1662),
.A2(n_1654),
.B(n_1637),
.C(n_1659),
.Y(n_1666)
);

AOI21xp33_ASAP7_75t_L g1667 ( 
.A1(n_1661),
.A2(n_1638),
.B(n_1648),
.Y(n_1667)
);

OAI211xp5_ASAP7_75t_L g1668 ( 
.A1(n_1657),
.A2(n_1635),
.B(n_1618),
.C(n_1645),
.Y(n_1668)
);

AOI221xp5_ASAP7_75t_L g1669 ( 
.A1(n_1655),
.A2(n_1625),
.B1(n_1613),
.B2(n_1615),
.C(n_1631),
.Y(n_1669)
);

AOI221xp5_ASAP7_75t_L g1670 ( 
.A1(n_1660),
.A2(n_1625),
.B1(n_1613),
.B2(n_1615),
.C(n_1631),
.Y(n_1670)
);

INVx2_ASAP7_75t_L g1671 ( 
.A(n_1656),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1656),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_SL g1673 ( 
.A(n_1658),
.B(n_1647),
.Y(n_1673)
);

OAI21xp5_ASAP7_75t_L g1674 ( 
.A1(n_1668),
.A2(n_1647),
.B(n_1646),
.Y(n_1674)
);

HB1xp67_ASAP7_75t_L g1675 ( 
.A(n_1671),
.Y(n_1675)
);

AOI22xp5_ASAP7_75t_L g1676 ( 
.A1(n_1666),
.A2(n_1630),
.B1(n_1622),
.B2(n_1633),
.Y(n_1676)
);

O2A1O1Ixp33_ASAP7_75t_L g1677 ( 
.A1(n_1673),
.A2(n_1664),
.B(n_1663),
.C(n_1651),
.Y(n_1677)
);

NOR2xp33_ASAP7_75t_SL g1678 ( 
.A(n_1672),
.B(n_1630),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_L g1679 ( 
.A(n_1678),
.B(n_1665),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_L g1680 ( 
.A(n_1676),
.B(n_1667),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1675),
.Y(n_1681)
);

INVx3_ASAP7_75t_L g1682 ( 
.A(n_1677),
.Y(n_1682)
);

BUFx3_ASAP7_75t_L g1683 ( 
.A(n_1674),
.Y(n_1683)
);

NOR2x1_ASAP7_75t_SL g1684 ( 
.A(n_1678),
.B(n_1627),
.Y(n_1684)
);

A2O1A1Ixp33_ASAP7_75t_L g1685 ( 
.A1(n_1683),
.A2(n_1670),
.B(n_1669),
.C(n_1617),
.Y(n_1685)
);

HB1xp67_ASAP7_75t_L g1686 ( 
.A(n_1684),
.Y(n_1686)
);

OAI22xp5_ASAP7_75t_SL g1687 ( 
.A1(n_1679),
.A2(n_1622),
.B1(n_1617),
.B2(n_1634),
.Y(n_1687)
);

INVx3_ASAP7_75t_L g1688 ( 
.A(n_1681),
.Y(n_1688)
);

AOI322xp5_ASAP7_75t_L g1689 ( 
.A1(n_1680),
.A2(n_1682),
.A3(n_1634),
.B1(n_1621),
.B2(n_1622),
.C1(n_1627),
.C2(n_1605),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1686),
.Y(n_1690)
);

INVx2_ASAP7_75t_L g1691 ( 
.A(n_1688),
.Y(n_1691)
);

OR2x2_ASAP7_75t_L g1692 ( 
.A(n_1685),
.B(n_1682),
.Y(n_1692)
);

AOI22xp5_ASAP7_75t_L g1693 ( 
.A1(n_1691),
.A2(n_1687),
.B1(n_1621),
.B2(n_1632),
.Y(n_1693)
);

AOI322xp5_ASAP7_75t_L g1694 ( 
.A1(n_1693),
.A2(n_1690),
.A3(n_1692),
.B1(n_1689),
.B2(n_1606),
.C1(n_1553),
.C2(n_1545),
.Y(n_1694)
);

OR2x2_ASAP7_75t_L g1695 ( 
.A(n_1694),
.B(n_1632),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1694),
.Y(n_1696)
);

INVxp67_ASAP7_75t_SL g1697 ( 
.A(n_1695),
.Y(n_1697)
);

INVx2_ASAP7_75t_L g1698 ( 
.A(n_1696),
.Y(n_1698)
);

CKINVDCx20_ASAP7_75t_R g1699 ( 
.A(n_1698),
.Y(n_1699)
);

OAI22x1_ASAP7_75t_L g1700 ( 
.A1(n_1697),
.A2(n_1624),
.B1(n_1586),
.B2(n_1553),
.Y(n_1700)
);

OAI21x1_ASAP7_75t_L g1701 ( 
.A1(n_1699),
.A2(n_1624),
.B(n_1548),
.Y(n_1701)
);

OAI322xp33_ASAP7_75t_L g1702 ( 
.A1(n_1701),
.A2(n_1700),
.A3(n_1548),
.B1(n_1563),
.B2(n_1566),
.C1(n_1564),
.C2(n_1554),
.Y(n_1702)
);

OAI21xp5_ASAP7_75t_SL g1703 ( 
.A1(n_1702),
.A2(n_1606),
.B(n_1553),
.Y(n_1703)
);

AOI322xp5_ASAP7_75t_L g1704 ( 
.A1(n_1703),
.A2(n_1545),
.A3(n_1563),
.B1(n_1564),
.B2(n_1566),
.C1(n_1536),
.C2(n_1535),
.Y(n_1704)
);

AOI22xp5_ASAP7_75t_L g1705 ( 
.A1(n_1704),
.A2(n_1592),
.B1(n_1560),
.B2(n_1558),
.Y(n_1705)
);

AOI211xp5_ASAP7_75t_L g1706 ( 
.A1(n_1705),
.A2(n_1560),
.B(n_1558),
.C(n_1556),
.Y(n_1706)
);


endmodule