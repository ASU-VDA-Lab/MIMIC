module fake_jpeg_2267_n_289 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_289);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_289;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_270;
wire n_199;
wire n_112;
wire n_260;
wire n_176;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx6f_ASAP7_75t_SL g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_14),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_4),
.B(n_7),
.Y(n_35)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

CKINVDCx14_ASAP7_75t_R g37 ( 
.A(n_12),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_3),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_9),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_6),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_7),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_4),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_37),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_45),
.B(n_46),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_35),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_22),
.Y(n_47)
);

INVx8_ASAP7_75t_L g121 ( 
.A(n_47),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_25),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_48),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g49 ( 
.A(n_25),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_49),
.B(n_57),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_21),
.B(n_16),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_50),
.B(n_52),
.Y(n_93)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_29),
.Y(n_51)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_51),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_16),
.Y(n_52)
);

INVx1_ASAP7_75t_SL g53 ( 
.A(n_24),
.Y(n_53)
);

NAND2xp33_ASAP7_75t_SL g96 ( 
.A(n_53),
.B(n_66),
.Y(n_96)
);

INVx13_ASAP7_75t_L g54 ( 
.A(n_22),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g110 ( 
.A(n_54),
.Y(n_110)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

INVx5_ASAP7_75t_L g119 ( 
.A(n_55),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_30),
.Y(n_56)
);

INVx6_ASAP7_75t_L g130 ( 
.A(n_56),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_30),
.Y(n_57)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_24),
.Y(n_58)
);

INVx3_ASAP7_75t_SL g133 ( 
.A(n_58),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

INVx8_ASAP7_75t_L g122 ( 
.A(n_59),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx8_ASAP7_75t_L g124 ( 
.A(n_60),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g107 ( 
.A(n_61),
.Y(n_107)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_22),
.Y(n_62)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_62),
.Y(n_116)
);

BUFx10_ASAP7_75t_L g63 ( 
.A(n_29),
.Y(n_63)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_63),
.Y(n_104)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_19),
.Y(n_64)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_64),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_31),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_65),
.B(n_73),
.Y(n_112)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_19),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_28),
.B(n_0),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_67),
.B(n_71),
.Y(n_97)
);

BUFx12_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_68),
.Y(n_105)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_20),
.Y(n_69)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_69),
.Y(n_89)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_70),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_31),
.B(n_15),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_26),
.Y(n_72)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_72),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_20),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_33),
.Y(n_74)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_74),
.Y(n_98)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_28),
.Y(n_75)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_75),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_33),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_76),
.B(n_82),
.Y(n_118)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_40),
.Y(n_77)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_77),
.Y(n_111)
);

INVx13_ASAP7_75t_L g78 ( 
.A(n_42),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_78),
.Y(n_90)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_42),
.Y(n_79)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_79),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_17),
.B(n_11),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_80),
.B(n_84),
.Y(n_128)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_44),
.Y(n_81)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_81),
.Y(n_117)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_26),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_43),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_83),
.B(n_86),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_18),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_84),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_18),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_85),
.Y(n_129)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_27),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_27),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_87),
.Y(n_132)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_32),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_88),
.B(n_1),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_48),
.A2(n_34),
.B1(n_32),
.B2(n_43),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g167 ( 
.A1(n_95),
.A2(n_102),
.B1(n_129),
.B2(n_115),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_53),
.A2(n_38),
.B1(n_17),
.B2(n_23),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_100),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_72),
.A2(n_38),
.B1(n_36),
.B2(n_23),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_101),
.A2(n_108),
.B(n_125),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_56),
.A2(n_36),
.B1(n_34),
.B2(n_2),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_72),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_109),
.B(n_97),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_54),
.A2(n_9),
.B(n_3),
.Y(n_113)
);

AOI21xp33_ASAP7_75t_L g168 ( 
.A1(n_113),
.A2(n_128),
.B(n_108),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_87),
.B(n_3),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_123),
.B(n_133),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_82),
.A2(n_7),
.B1(n_9),
.B2(n_85),
.Y(n_125)
);

OA22x2_ASAP7_75t_SL g127 ( 
.A1(n_78),
.A2(n_63),
.B1(n_81),
.B2(n_70),
.Y(n_127)
);

A2O1A1Ixp33_ASAP7_75t_L g152 ( 
.A1(n_127),
.A2(n_63),
.B(n_68),
.C(n_96),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_59),
.B(n_61),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_134),
.B(n_47),
.Y(n_145)
);

INVx2_ASAP7_75t_SL g135 ( 
.A(n_114),
.Y(n_135)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_135),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_96),
.B(n_55),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_137),
.B(n_145),
.Y(n_184)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_103),
.Y(n_138)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_138),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_139),
.B(n_140),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_112),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_118),
.B(n_89),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_SL g196 ( 
.A(n_141),
.B(n_148),
.Y(n_196)
);

BUFx3_ASAP7_75t_L g142 ( 
.A(n_121),
.Y(n_142)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_142),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_93),
.B(n_60),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_143),
.B(n_147),
.Y(n_182)
);

AND2x6_ASAP7_75t_L g144 ( 
.A(n_127),
.B(n_47),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_144),
.B(n_150),
.Y(n_180)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_130),
.Y(n_146)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_146),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_92),
.B(n_79),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_98),
.B(n_62),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_126),
.B(n_62),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_149),
.B(n_153),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_106),
.Y(n_150)
);

INVx13_ASAP7_75t_L g151 ( 
.A(n_110),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_151),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g195 ( 
.A(n_152),
.B(n_161),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_90),
.B(n_68),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_99),
.B(n_131),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_154),
.B(n_162),
.Y(n_173)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_133),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_155),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_116),
.B(n_111),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_156),
.B(n_157),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_105),
.B(n_117),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_107),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_158),
.B(n_160),
.Y(n_190)
);

OR2x2_ASAP7_75t_SL g159 ( 
.A(n_127),
.B(n_116),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_159),
.B(n_163),
.C(n_91),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_94),
.Y(n_160)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_119),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_132),
.B(n_95),
.Y(n_162)
);

OR2x2_ASAP7_75t_SL g163 ( 
.A(n_100),
.B(n_105),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_110),
.B(n_120),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_164),
.B(n_165),
.Y(n_178)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_130),
.Y(n_165)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_94),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_166),
.B(n_168),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_167),
.A2(n_104),
.B1(n_107),
.B2(n_91),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_170),
.B(n_119),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_136),
.A2(n_101),
.B(n_125),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_181),
.A2(n_194),
.B(n_169),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_183),
.A2(n_186),
.B1(n_158),
.B2(n_155),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_136),
.A2(n_124),
.B1(n_122),
.B2(n_104),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_148),
.B(n_110),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_188),
.B(n_137),
.C(n_159),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_189),
.B(n_161),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_191),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_154),
.B(n_122),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_192),
.B(n_162),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_152),
.A2(n_121),
.B(n_124),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_198),
.A2(n_204),
.B(n_210),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_SL g222 ( 
.A(n_199),
.B(n_217),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_182),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_200),
.B(n_203),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_201),
.B(n_207),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_196),
.B(n_141),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_202),
.B(n_203),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_175),
.B(n_150),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_194),
.A2(n_163),
.B(n_169),
.Y(n_204)
);

INVx13_ASAP7_75t_L g205 ( 
.A(n_172),
.Y(n_205)
);

INVx4_ASAP7_75t_L g228 ( 
.A(n_205),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_179),
.A2(n_137),
.B(n_144),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g232 ( 
.A1(n_206),
.A2(n_215),
.B(n_216),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_187),
.B(n_135),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_193),
.B(n_189),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_208),
.B(n_178),
.Y(n_226)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_209),
.Y(n_223)
);

O2A1O1Ixp33_ASAP7_75t_L g210 ( 
.A1(n_181),
.A2(n_142),
.B(n_138),
.C(n_151),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_174),
.Y(n_211)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_211),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_173),
.A2(n_146),
.B1(n_165),
.B2(n_166),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_212),
.A2(n_219),
.B1(n_188),
.B2(n_184),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_213),
.B(n_185),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_186),
.A2(n_135),
.B1(n_160),
.B2(n_191),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_214),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_195),
.A2(n_179),
.B(n_180),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_195),
.A2(n_184),
.B1(n_173),
.B2(n_192),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_196),
.B(n_184),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_174),
.Y(n_218)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_218),
.Y(n_231)
);

OAI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_195),
.A2(n_178),
.B1(n_190),
.B2(n_183),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_207),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_220),
.B(n_218),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_221),
.A2(n_201),
.B1(n_212),
.B2(n_209),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_226),
.B(n_233),
.Y(n_246)
);

INVx1_ASAP7_75t_SL g248 ( 
.A(n_230),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_213),
.B(n_185),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_234),
.B(n_235),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_208),
.B(n_177),
.Y(n_235)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_229),
.Y(n_237)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_237),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_236),
.A2(n_198),
.B(n_204),
.Y(n_238)
);

CKINVDCx14_ASAP7_75t_R g262 ( 
.A(n_238),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_222),
.B(n_197),
.C(n_232),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_239),
.B(n_241),
.C(n_249),
.Y(n_261)
);

A2O1A1O1Ixp25_ASAP7_75t_L g240 ( 
.A1(n_232),
.A2(n_199),
.B(n_202),
.C(n_216),
.D(n_215),
.Y(n_240)
);

HB1xp67_ASAP7_75t_L g255 ( 
.A(n_240),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_222),
.B(n_217),
.C(n_206),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_242),
.B(n_243),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_230),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_244),
.A2(n_223),
.B1(n_224),
.B2(n_220),
.Y(n_254)
);

CKINVDCx16_ASAP7_75t_R g245 ( 
.A(n_234),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_245),
.B(n_251),
.Y(n_260)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_229),
.Y(n_247)
);

INVx2_ASAP7_75t_SL g252 ( 
.A(n_247),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_224),
.B(n_219),
.C(n_211),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_235),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_237),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_253),
.B(n_256),
.Y(n_263)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_254),
.Y(n_267)
);

OAI22xp33_ASAP7_75t_L g256 ( 
.A1(n_243),
.A2(n_223),
.B1(n_225),
.B2(n_236),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_239),
.B(n_226),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_258),
.B(n_261),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_260),
.B(n_227),
.Y(n_264)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_264),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_262),
.A2(n_238),
.B(n_240),
.Y(n_265)
);

AOI21xp33_ASAP7_75t_L g277 ( 
.A1(n_265),
.A2(n_269),
.B(n_221),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_L g266 ( 
.A1(n_254),
.A2(n_248),
.B(n_249),
.Y(n_266)
);

AND2x2_ASAP7_75t_L g276 ( 
.A(n_266),
.B(n_270),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_268),
.B(n_261),
.C(n_258),
.Y(n_274)
);

AOI322xp5_ASAP7_75t_L g269 ( 
.A1(n_259),
.A2(n_246),
.A3(n_250),
.B1(n_248),
.B2(n_251),
.C1(n_227),
.C2(n_241),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_253),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_252),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_271),
.A2(n_252),
.B1(n_257),
.B2(n_247),
.Y(n_273)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_273),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_274),
.B(n_275),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_268),
.B(n_255),
.C(n_256),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_277),
.A2(n_266),
.B(n_267),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_278),
.A2(n_279),
.B1(n_276),
.B2(n_263),
.Y(n_282)
);

OAI21xp33_ASAP7_75t_SL g279 ( 
.A1(n_276),
.A2(n_265),
.B(n_267),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_282),
.B(n_283),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_281),
.B(n_280),
.C(n_272),
.Y(n_283)
);

AO22x1_ASAP7_75t_L g284 ( 
.A1(n_279),
.A2(n_263),
.B1(n_231),
.B2(n_210),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_284),
.B(n_231),
.C(n_228),
.Y(n_286)
);

AOI322xp5_ASAP7_75t_L g287 ( 
.A1(n_286),
.A2(n_205),
.A3(n_284),
.B1(n_210),
.B2(n_172),
.C1(n_228),
.C2(n_176),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_287),
.B(n_285),
.C(n_205),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_288),
.B(n_171),
.Y(n_289)
);


endmodule