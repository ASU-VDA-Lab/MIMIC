module real_aes_8478_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_659;
wire n_547;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_417;
wire n_363;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_502;
wire n_434;
wire n_527;
wire n_600;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_713;
wire n_288;
wire n_404;
wire n_598;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_217;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_717;
wire n_359;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_719;
wire n_473;
wire n_465;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND3xp33_ASAP7_75t_SL g107 ( .A(n_0), .B(n_108), .C(n_109), .Y(n_107) );
INVx1_ASAP7_75t_L g124 ( .A(n_0), .Y(n_124) );
A2O1A1Ixp33_ASAP7_75t_L g502 ( .A1(n_1), .A2(n_148), .B(n_153), .C(n_503), .Y(n_502) );
INVx1_ASAP7_75t_L g260 ( .A(n_2), .Y(n_260) );
AOI21xp5_ASAP7_75t_L g459 ( .A1(n_3), .A2(n_143), .B(n_460), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_4), .B(n_220), .Y(n_465) );
CKINVDCx20_ASAP7_75t_R g126 ( .A(n_5), .Y(n_126) );
AOI21xp33_ASAP7_75t_L g221 ( .A1(n_6), .A2(n_143), .B(n_222), .Y(n_221) );
AND2x6_ASAP7_75t_L g148 ( .A(n_7), .B(n_149), .Y(n_148) );
AOI21xp5_ASAP7_75t_L g141 ( .A1(n_8), .A2(n_142), .B(n_150), .Y(n_141) );
INVx1_ASAP7_75t_L g105 ( .A(n_9), .Y(n_105) );
NOR2xp33_ASAP7_75t_L g125 ( .A(n_9), .B(n_40), .Y(n_125) );
INVx1_ASAP7_75t_L g554 ( .A(n_10), .Y(n_554) );
NAND2xp5_ASAP7_75t_SL g505 ( .A(n_11), .B(n_192), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_12), .B(n_208), .Y(n_207) );
INVx1_ASAP7_75t_L g227 ( .A(n_13), .Y(n_227) );
INVx1_ASAP7_75t_L g140 ( .A(n_14), .Y(n_140) );
INVx1_ASAP7_75t_L g160 ( .A(n_15), .Y(n_160) );
A2O1A1Ixp33_ASAP7_75t_L g513 ( .A1(n_16), .A2(n_161), .B(n_175), .C(n_514), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_17), .B(n_220), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_18), .B(n_177), .Y(n_193) );
NAND2xp5_ASAP7_75t_SL g170 ( .A(n_19), .B(n_143), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_20), .B(n_478), .Y(n_477) );
A2O1A1Ixp33_ASAP7_75t_L g521 ( .A1(n_21), .A2(n_208), .B(n_234), .C(n_522), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_22), .B(n_220), .Y(n_250) );
NAND2xp5_ASAP7_75t_SL g487 ( .A(n_23), .B(n_192), .Y(n_487) );
A2O1A1Ixp33_ASAP7_75t_L g156 ( .A1(n_24), .A2(n_157), .B(n_159), .C(n_161), .Y(n_156) );
NAND2xp5_ASAP7_75t_SL g451 ( .A(n_25), .B(n_192), .Y(n_451) );
CKINVDCx16_ASAP7_75t_R g482 ( .A(n_26), .Y(n_482) );
INVx1_ASAP7_75t_L g450 ( .A(n_27), .Y(n_450) );
BUFx6f_ASAP7_75t_L g147 ( .A(n_28), .Y(n_147) );
CKINVDCx20_ASAP7_75t_R g501 ( .A(n_29), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_30), .B(n_192), .Y(n_261) );
INVx1_ASAP7_75t_L g475 ( .A(n_31), .Y(n_475) );
INVx1_ASAP7_75t_L g239 ( .A(n_32), .Y(n_239) );
INVx2_ASAP7_75t_L g146 ( .A(n_33), .Y(n_146) );
CKINVDCx20_ASAP7_75t_R g507 ( .A(n_34), .Y(n_507) );
A2O1A1Ixp33_ASAP7_75t_L g462 ( .A1(n_35), .A2(n_208), .B(n_228), .C(n_463), .Y(n_462) );
INVxp67_ASAP7_75t_L g476 ( .A(n_36), .Y(n_476) );
A2O1A1Ixp33_ASAP7_75t_L g171 ( .A1(n_37), .A2(n_148), .B(n_153), .C(n_172), .Y(n_171) );
A2O1A1Ixp33_ASAP7_75t_L g448 ( .A1(n_38), .A2(n_153), .B(n_449), .C(n_454), .Y(n_448) );
CKINVDCx14_ASAP7_75t_R g461 ( .A(n_39), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g104 ( .A(n_40), .B(n_105), .Y(n_104) );
INVx1_ASAP7_75t_L g237 ( .A(n_41), .Y(n_237) );
A2O1A1Ixp33_ASAP7_75t_L g552 ( .A1(n_42), .A2(n_179), .B(n_225), .C(n_553), .Y(n_552) );
NAND2xp5_ASAP7_75t_SL g191 ( .A(n_43), .B(n_192), .Y(n_191) );
OAI22xp5_ASAP7_75t_L g715 ( .A1(n_44), .A2(n_438), .B1(n_707), .B2(n_716), .Y(n_715) );
CKINVDCx20_ASAP7_75t_R g716 ( .A(n_44), .Y(n_716) );
CKINVDCx20_ASAP7_75t_R g456 ( .A(n_45), .Y(n_456) );
CKINVDCx20_ASAP7_75t_R g472 ( .A(n_46), .Y(n_472) );
INVx1_ASAP7_75t_L g520 ( .A(n_47), .Y(n_520) );
CKINVDCx16_ASAP7_75t_R g240 ( .A(n_48), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_49), .B(n_143), .Y(n_211) );
AOI22xp5_ASAP7_75t_L g233 ( .A1(n_50), .A2(n_153), .B1(n_234), .B2(n_236), .Y(n_233) );
CKINVDCx20_ASAP7_75t_R g183 ( .A(n_51), .Y(n_183) );
CKINVDCx16_ASAP7_75t_R g257 ( .A(n_52), .Y(n_257) );
AOI22xp33_ASAP7_75t_L g99 ( .A1(n_53), .A2(n_100), .B1(n_112), .B2(n_719), .Y(n_99) );
A2O1A1Ixp33_ASAP7_75t_L g224 ( .A1(n_54), .A2(n_225), .B(n_226), .C(n_228), .Y(n_224) );
CKINVDCx14_ASAP7_75t_R g551 ( .A(n_55), .Y(n_551) );
CKINVDCx20_ASAP7_75t_R g196 ( .A(n_56), .Y(n_196) );
INVx1_ASAP7_75t_L g223 ( .A(n_57), .Y(n_223) );
INVx1_ASAP7_75t_L g149 ( .A(n_58), .Y(n_149) );
INVx1_ASAP7_75t_L g139 ( .A(n_59), .Y(n_139) );
INVx1_ASAP7_75t_SL g464 ( .A(n_60), .Y(n_464) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_61), .Y(n_117) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_62), .B(n_220), .Y(n_524) );
INVx1_ASAP7_75t_L g485 ( .A(n_63), .Y(n_485) );
A2O1A1Ixp33_ASAP7_75t_SL g247 ( .A1(n_64), .A2(n_177), .B(n_228), .C(n_248), .Y(n_247) );
INVxp67_ASAP7_75t_L g249 ( .A(n_65), .Y(n_249) );
AOI222xp33_ASAP7_75t_SL g127 ( .A1(n_66), .A2(n_68), .B1(n_128), .B2(n_702), .C1(n_703), .C2(n_710), .Y(n_127) );
INVx1_ASAP7_75t_L g111 ( .A(n_67), .Y(n_111) );
INVx1_ASAP7_75t_L g702 ( .A(n_68), .Y(n_702) );
AOI21xp5_ASAP7_75t_L g549 ( .A1(n_69), .A2(n_143), .B(n_550), .Y(n_549) );
CKINVDCx20_ASAP7_75t_R g490 ( .A(n_70), .Y(n_490) );
CKINVDCx20_ASAP7_75t_R g242 ( .A(n_71), .Y(n_242) );
AOI21xp5_ASAP7_75t_L g510 ( .A1(n_72), .A2(n_143), .B(n_511), .Y(n_510) );
INVx1_ASAP7_75t_L g187 ( .A(n_73), .Y(n_187) );
AOI21xp5_ASAP7_75t_L g470 ( .A1(n_74), .A2(n_142), .B(n_471), .Y(n_470) );
CKINVDCx16_ASAP7_75t_R g447 ( .A(n_75), .Y(n_447) );
INVx1_ASAP7_75t_L g512 ( .A(n_76), .Y(n_512) );
A2O1A1Ixp33_ASAP7_75t_L g189 ( .A1(n_77), .A2(n_148), .B(n_153), .C(n_190), .Y(n_189) );
AOI21xp5_ASAP7_75t_L g518 ( .A1(n_78), .A2(n_143), .B(n_519), .Y(n_518) );
INVx1_ASAP7_75t_L g515 ( .A(n_79), .Y(n_515) );
NAND2xp5_ASAP7_75t_SL g173 ( .A(n_80), .B(n_174), .Y(n_173) );
INVx2_ASAP7_75t_L g137 ( .A(n_81), .Y(n_137) );
INVx1_ASAP7_75t_L g504 ( .A(n_82), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_83), .B(n_177), .Y(n_176) );
A2O1A1Ixp33_ASAP7_75t_L g258 ( .A1(n_84), .A2(n_148), .B(n_153), .C(n_259), .Y(n_258) );
INVx2_ASAP7_75t_L g108 ( .A(n_85), .Y(n_108) );
OR2x2_ASAP7_75t_L g121 ( .A(n_85), .B(n_122), .Y(n_121) );
OR2x2_ASAP7_75t_L g701 ( .A(n_85), .B(n_123), .Y(n_701) );
A2O1A1Ixp33_ASAP7_75t_L g483 ( .A1(n_86), .A2(n_153), .B(n_484), .C(n_488), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_87), .B(n_136), .Y(n_229) );
CKINVDCx20_ASAP7_75t_R g264 ( .A(n_88), .Y(n_264) );
A2O1A1Ixp33_ASAP7_75t_L g204 ( .A1(n_89), .A2(n_148), .B(n_153), .C(n_205), .Y(n_204) );
CKINVDCx20_ASAP7_75t_R g213 ( .A(n_90), .Y(n_213) );
INVx1_ASAP7_75t_L g246 ( .A(n_91), .Y(n_246) );
CKINVDCx16_ASAP7_75t_R g151 ( .A(n_92), .Y(n_151) );
NAND2xp5_ASAP7_75t_SL g206 ( .A(n_93), .B(n_174), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_94), .B(n_165), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_95), .B(n_165), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g110 ( .A(n_96), .B(n_111), .Y(n_110) );
AOI21xp5_ASAP7_75t_L g244 ( .A1(n_97), .A2(n_143), .B(n_245), .Y(n_244) );
INVx2_ASAP7_75t_L g523 ( .A(n_98), .Y(n_523) );
INVx1_ASAP7_75t_L g100 ( .A(n_101), .Y(n_100) );
INVx2_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
INVx2_ASAP7_75t_SL g719 ( .A(n_102), .Y(n_719) );
AND2x2_ASAP7_75t_L g102 ( .A(n_103), .B(n_106), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
INVx1_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
OR2x2_ASAP7_75t_L g437 ( .A(n_108), .B(n_123), .Y(n_437) );
NOR2x2_ASAP7_75t_L g712 ( .A(n_108), .B(n_122), .Y(n_712) );
INVx1_ASAP7_75t_SL g109 ( .A(n_110), .Y(n_109) );
AOI22x1_ASAP7_75t_L g112 ( .A1(n_113), .A2(n_127), .B1(n_713), .B2(n_714), .Y(n_112) );
NOR2xp33_ASAP7_75t_L g113 ( .A(n_114), .B(n_118), .Y(n_113) );
INVx1_ASAP7_75t_SL g114 ( .A(n_115), .Y(n_114) );
BUFx2_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
INVx2_ASAP7_75t_SL g713 ( .A(n_116), .Y(n_713) );
INVx2_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
AOI21xp5_ASAP7_75t_L g714 ( .A1(n_118), .A2(n_715), .B(n_717), .Y(n_714) );
NOR2xp33_ASAP7_75t_SL g118 ( .A(n_119), .B(n_126), .Y(n_118) );
INVx1_ASAP7_75t_SL g119 ( .A(n_120), .Y(n_119) );
INVx1_ASAP7_75t_SL g120 ( .A(n_121), .Y(n_120) );
INVx1_ASAP7_75t_SL g718 ( .A(n_121), .Y(n_718) );
INVx2_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
AND2x2_ASAP7_75t_L g123 ( .A(n_124), .B(n_125), .Y(n_123) );
OAI22xp5_ASAP7_75t_SL g128 ( .A1(n_129), .A2(n_437), .B1(n_438), .B2(n_701), .Y(n_128) );
INVx2_ASAP7_75t_SL g704 ( .A(n_129), .Y(n_704) );
OR4x2_ASAP7_75t_L g129 ( .A(n_130), .B(n_333), .C(n_392), .D(n_419), .Y(n_129) );
NAND3xp33_ASAP7_75t_SL g130 ( .A(n_131), .B(n_275), .C(n_300), .Y(n_130) );
O2A1O1Ixp33_ASAP7_75t_L g131 ( .A1(n_132), .A2(n_198), .B(n_218), .C(n_251), .Y(n_131) );
AOI211xp5_ASAP7_75t_SL g423 ( .A1(n_132), .A2(n_424), .B(n_426), .C(n_429), .Y(n_423) );
AND2x2_ASAP7_75t_L g132 ( .A(n_133), .B(n_167), .Y(n_132) );
INVx1_ASAP7_75t_L g298 ( .A(n_133), .Y(n_298) );
INVx1_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
OR2x2_ASAP7_75t_L g273 ( .A(n_134), .B(n_274), .Y(n_273) );
INVx2_ASAP7_75t_L g305 ( .A(n_134), .Y(n_305) );
AND2x2_ASAP7_75t_L g360 ( .A(n_134), .B(n_329), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_134), .B(n_216), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_134), .B(n_217), .Y(n_418) );
INVx2_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
INVx1_ASAP7_75t_L g279 ( .A(n_135), .Y(n_279) );
AND2x2_ASAP7_75t_L g322 ( .A(n_135), .B(n_185), .Y(n_322) );
AND2x2_ASAP7_75t_L g340 ( .A(n_135), .B(n_217), .Y(n_340) );
OA21x2_ASAP7_75t_L g135 ( .A1(n_136), .A2(n_141), .B(n_164), .Y(n_135) );
INVx1_ASAP7_75t_L g197 ( .A(n_136), .Y(n_197) );
INVx2_ASAP7_75t_L g202 ( .A(n_136), .Y(n_202) );
O2A1O1Ixp33_ASAP7_75t_L g446 ( .A1(n_136), .A2(n_188), .B(n_447), .C(n_448), .Y(n_446) );
OA21x2_ASAP7_75t_L g548 ( .A1(n_136), .A2(n_549), .B(n_555), .Y(n_548) );
AND2x2_ASAP7_75t_SL g136 ( .A(n_137), .B(n_138), .Y(n_136) );
AND2x2_ASAP7_75t_L g166 ( .A(n_137), .B(n_138), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g138 ( .A(n_139), .B(n_140), .Y(n_138) );
BUFx2_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
AND2x4_ASAP7_75t_L g143 ( .A(n_144), .B(n_148), .Y(n_143) );
NAND2x1p5_ASAP7_75t_L g188 ( .A(n_144), .B(n_148), .Y(n_188) );
AND2x2_ASAP7_75t_L g144 ( .A(n_145), .B(n_147), .Y(n_144) );
INVx1_ASAP7_75t_L g453 ( .A(n_145), .Y(n_453) );
INVx1_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx2_ASAP7_75t_L g154 ( .A(n_146), .Y(n_154) );
INVx1_ASAP7_75t_L g235 ( .A(n_146), .Y(n_235) );
INVx1_ASAP7_75t_L g155 ( .A(n_147), .Y(n_155) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_147), .Y(n_158) );
INVx3_ASAP7_75t_L g175 ( .A(n_147), .Y(n_175) );
INVx1_ASAP7_75t_L g177 ( .A(n_147), .Y(n_177) );
BUFx6f_ASAP7_75t_L g192 ( .A(n_147), .Y(n_192) );
INVx4_ASAP7_75t_SL g163 ( .A(n_148), .Y(n_163) );
BUFx3_ASAP7_75t_L g454 ( .A(n_148), .Y(n_454) );
O2A1O1Ixp33_ASAP7_75t_L g150 ( .A1(n_151), .A2(n_152), .B(n_156), .C(n_163), .Y(n_150) );
O2A1O1Ixp33_ASAP7_75t_L g222 ( .A1(n_152), .A2(n_163), .B(n_223), .C(n_224), .Y(n_222) );
O2A1O1Ixp33_ASAP7_75t_L g245 ( .A1(n_152), .A2(n_163), .B(n_246), .C(n_247), .Y(n_245) );
O2A1O1Ixp33_ASAP7_75t_L g460 ( .A1(n_152), .A2(n_163), .B(n_461), .C(n_462), .Y(n_460) );
O2A1O1Ixp33_ASAP7_75t_SL g471 ( .A1(n_152), .A2(n_163), .B(n_472), .C(n_473), .Y(n_471) );
O2A1O1Ixp33_ASAP7_75t_SL g511 ( .A1(n_152), .A2(n_163), .B(n_512), .C(n_513), .Y(n_511) );
O2A1O1Ixp33_ASAP7_75t_SL g519 ( .A1(n_152), .A2(n_163), .B(n_520), .C(n_521), .Y(n_519) );
O2A1O1Ixp33_ASAP7_75t_SL g550 ( .A1(n_152), .A2(n_163), .B(n_551), .C(n_552), .Y(n_550) );
INVx5_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
AND2x6_ASAP7_75t_L g153 ( .A(n_154), .B(n_155), .Y(n_153) );
BUFx3_ASAP7_75t_L g162 ( .A(n_154), .Y(n_162) );
BUFx6f_ASAP7_75t_L g210 ( .A(n_154), .Y(n_210) );
NOR2xp33_ASAP7_75t_L g159 ( .A(n_157), .B(n_160), .Y(n_159) );
OAI22xp33_ASAP7_75t_L g474 ( .A1(n_157), .A2(n_174), .B1(n_475), .B2(n_476), .Y(n_474) );
NOR2xp33_ASAP7_75t_L g514 ( .A(n_157), .B(n_515), .Y(n_514) );
NOR2xp33_ASAP7_75t_L g522 ( .A(n_157), .B(n_523), .Y(n_522) );
INVx4_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
OAI22xp5_ASAP7_75t_SL g236 ( .A1(n_158), .A2(n_237), .B1(n_238), .B2(n_239), .Y(n_236) );
INVx2_ASAP7_75t_L g238 ( .A(n_158), .Y(n_238) );
INVx1_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
INVx2_ASAP7_75t_L g179 ( .A(n_162), .Y(n_179) );
OAI22xp33_ASAP7_75t_L g232 ( .A1(n_163), .A2(n_188), .B1(n_233), .B2(n_240), .Y(n_232) );
INVx1_ASAP7_75t_L g488 ( .A(n_163), .Y(n_488) );
INVx4_ASAP7_75t_L g184 ( .A(n_165), .Y(n_184) );
OA21x2_ASAP7_75t_L g243 ( .A1(n_165), .A2(n_244), .B(n_250), .Y(n_243) );
HB1xp67_ASAP7_75t_L g458 ( .A(n_165), .Y(n_458) );
BUFx6f_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
INVx1_ASAP7_75t_L g181 ( .A(n_166), .Y(n_181) );
INVx4_ASAP7_75t_L g272 ( .A(n_167), .Y(n_272) );
OAI21xp5_ASAP7_75t_L g327 ( .A1(n_167), .A2(n_328), .B(n_330), .Y(n_327) );
AND2x2_ASAP7_75t_L g408 ( .A(n_167), .B(n_409), .Y(n_408) );
AND2x2_ASAP7_75t_L g167 ( .A(n_168), .B(n_185), .Y(n_167) );
INVx1_ASAP7_75t_L g215 ( .A(n_168), .Y(n_215) );
AND2x2_ASAP7_75t_L g277 ( .A(n_168), .B(n_217), .Y(n_277) );
OR2x2_ASAP7_75t_L g306 ( .A(n_168), .B(n_307), .Y(n_306) );
INVx2_ASAP7_75t_L g320 ( .A(n_168), .Y(n_320) );
INVx3_ASAP7_75t_L g329 ( .A(n_168), .Y(n_329) );
AND2x2_ASAP7_75t_L g339 ( .A(n_168), .B(n_340), .Y(n_339) );
AND2x2_ASAP7_75t_L g372 ( .A(n_168), .B(n_278), .Y(n_372) );
AND2x2_ASAP7_75t_L g396 ( .A(n_168), .B(n_352), .Y(n_396) );
OR2x6_ASAP7_75t_L g168 ( .A(n_169), .B(n_182), .Y(n_168) );
AOI21xp5_ASAP7_75t_SL g169 ( .A1(n_170), .A2(n_171), .B(n_180), .Y(n_169) );
AOI21xp5_ASAP7_75t_L g172 ( .A1(n_173), .A2(n_176), .B(n_178), .Y(n_172) );
O2A1O1Ixp33_ASAP7_75t_L g259 ( .A1(n_174), .A2(n_260), .B(n_261), .C(n_262), .Y(n_259) );
O2A1O1Ixp33_ASAP7_75t_L g449 ( .A1(n_174), .A2(n_450), .B(n_451), .C(n_452), .Y(n_449) );
INVx5_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
NOR2xp33_ASAP7_75t_L g226 ( .A(n_175), .B(n_227), .Y(n_226) );
NOR2xp33_ASAP7_75t_L g248 ( .A(n_175), .B(n_249), .Y(n_248) );
NOR2xp33_ASAP7_75t_L g553 ( .A(n_175), .B(n_554), .Y(n_553) );
AOI21xp5_ASAP7_75t_L g190 ( .A1(n_178), .A2(n_191), .B(n_193), .Y(n_190) );
O2A1O1Ixp33_ASAP7_75t_L g484 ( .A1(n_178), .A2(n_485), .B(n_486), .C(n_487), .Y(n_484) );
O2A1O1Ixp5_ASAP7_75t_L g503 ( .A1(n_178), .A2(n_486), .B(n_504), .C(n_505), .Y(n_503) );
INVx2_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
INVx1_ASAP7_75t_L g194 ( .A(n_180), .Y(n_194) );
INVx2_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
AO21x2_ASAP7_75t_L g231 ( .A1(n_181), .A2(n_232), .B(n_241), .Y(n_231) );
NOR2xp33_ASAP7_75t_L g241 ( .A(n_181), .B(n_242), .Y(n_241) );
AO21x2_ASAP7_75t_L g255 ( .A1(n_181), .A2(n_256), .B(n_263), .Y(n_255) );
NOR2xp33_ASAP7_75t_SL g182 ( .A(n_183), .B(n_184), .Y(n_182) );
INVx3_ASAP7_75t_L g220 ( .A(n_184), .Y(n_220) );
NOR2xp33_ASAP7_75t_L g455 ( .A(n_184), .B(n_456), .Y(n_455) );
AO21x2_ASAP7_75t_L g480 ( .A1(n_184), .A2(n_481), .B(n_489), .Y(n_480) );
NOR2xp33_ASAP7_75t_L g506 ( .A(n_184), .B(n_507), .Y(n_506) );
INVx2_ASAP7_75t_L g217 ( .A(n_185), .Y(n_217) );
AND2x2_ASAP7_75t_L g432 ( .A(n_185), .B(n_274), .Y(n_432) );
AO21x2_ASAP7_75t_L g185 ( .A1(n_186), .A2(n_194), .B(n_195), .Y(n_185) );
OAI21xp5_ASAP7_75t_L g186 ( .A1(n_187), .A2(n_188), .B(n_189), .Y(n_186) );
OAI21xp5_ASAP7_75t_L g256 ( .A1(n_188), .A2(n_257), .B(n_258), .Y(n_256) );
OAI21xp5_ASAP7_75t_L g481 ( .A1(n_188), .A2(n_482), .B(n_483), .Y(n_481) );
OAI21xp5_ASAP7_75t_L g500 ( .A1(n_188), .A2(n_501), .B(n_502), .Y(n_500) );
INVx4_ASAP7_75t_L g208 ( .A(n_192), .Y(n_208) );
INVx2_ASAP7_75t_L g225 ( .A(n_192), .Y(n_225) );
INVx1_ASAP7_75t_L g469 ( .A(n_194), .Y(n_469) );
AO21x2_ASAP7_75t_L g493 ( .A1(n_194), .A2(n_494), .B(n_495), .Y(n_493) );
NOR2xp33_ASAP7_75t_L g195 ( .A(n_196), .B(n_197), .Y(n_195) );
NOR2xp33_ASAP7_75t_L g212 ( .A(n_197), .B(n_213), .Y(n_212) );
NOR2xp33_ASAP7_75t_L g263 ( .A(n_197), .B(n_264), .Y(n_263) );
AO21x2_ASAP7_75t_L g499 ( .A1(n_197), .A2(n_500), .B(n_506), .Y(n_499) );
AND2x2_ASAP7_75t_L g198 ( .A(n_199), .B(n_214), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
NOR2xp33_ASAP7_75t_L g328 ( .A(n_200), .B(n_329), .Y(n_328) );
AND2x2_ASAP7_75t_L g352 ( .A(n_200), .B(n_340), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_200), .B(n_329), .Y(n_414) );
INVx1_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
INVx2_ASAP7_75t_L g274 ( .A(n_201), .Y(n_274) );
AND2x2_ASAP7_75t_L g278 ( .A(n_201), .B(n_279), .Y(n_278) );
AND2x2_ASAP7_75t_L g319 ( .A(n_201), .B(n_320), .Y(n_319) );
AO21x2_ASAP7_75t_L g201 ( .A1(n_202), .A2(n_203), .B(n_212), .Y(n_201) );
INVx1_ASAP7_75t_L g478 ( .A(n_202), .Y(n_478) );
NOR2xp33_ASAP7_75t_L g489 ( .A(n_202), .B(n_490), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_204), .B(n_211), .Y(n_203) );
AOI21xp5_ASAP7_75t_L g205 ( .A1(n_206), .A2(n_207), .B(n_209), .Y(n_205) );
NOR2xp33_ASAP7_75t_L g463 ( .A(n_208), .B(n_464), .Y(n_463) );
HB1xp67_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
INVx3_ASAP7_75t_L g228 ( .A(n_210), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_214), .B(n_315), .Y(n_337) );
INVx1_ASAP7_75t_L g376 ( .A(n_214), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_214), .B(n_303), .Y(n_420) );
AND2x2_ASAP7_75t_L g214 ( .A(n_215), .B(n_216), .Y(n_214) );
AND2x2_ASAP7_75t_L g283 ( .A(n_215), .B(n_278), .Y(n_283) );
INVx2_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_217), .B(n_274), .Y(n_307) );
INVx1_ASAP7_75t_L g386 ( .A(n_217), .Y(n_386) );
AOI322xp5_ASAP7_75t_L g410 ( .A1(n_218), .A2(n_325), .A3(n_385), .B1(n_411), .B2(n_413), .C1(n_415), .C2(n_417), .Y(n_410) );
AND2x2_ASAP7_75t_SL g218 ( .A(n_219), .B(n_230), .Y(n_218) );
AND2x2_ASAP7_75t_L g265 ( .A(n_219), .B(n_243), .Y(n_265) );
INVx1_ASAP7_75t_SL g268 ( .A(n_219), .Y(n_268) );
AND2x2_ASAP7_75t_L g270 ( .A(n_219), .B(n_231), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_219), .B(n_287), .Y(n_293) );
INVx2_ASAP7_75t_L g312 ( .A(n_219), .Y(n_312) );
AND2x2_ASAP7_75t_L g325 ( .A(n_219), .B(n_326), .Y(n_325) );
OR2x2_ASAP7_75t_L g363 ( .A(n_219), .B(n_287), .Y(n_363) );
BUFx2_ASAP7_75t_L g380 ( .A(n_219), .Y(n_380) );
AND2x2_ASAP7_75t_L g394 ( .A(n_219), .B(n_254), .Y(n_394) );
OA21x2_ASAP7_75t_L g219 ( .A1(n_220), .A2(n_221), .B(n_229), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_230), .B(n_282), .Y(n_309) );
AND2x2_ASAP7_75t_L g436 ( .A(n_230), .B(n_312), .Y(n_436) );
AND2x2_ASAP7_75t_L g230 ( .A(n_231), .B(n_243), .Y(n_230) );
OR2x2_ASAP7_75t_L g281 ( .A(n_231), .B(n_282), .Y(n_281) );
INVx3_ASAP7_75t_L g287 ( .A(n_231), .Y(n_287) );
AND2x2_ASAP7_75t_L g332 ( .A(n_231), .B(n_255), .Y(n_332) );
NOR2xp33_ASAP7_75t_L g379 ( .A(n_231), .B(n_380), .Y(n_379) );
HB1xp67_ASAP7_75t_L g416 ( .A(n_231), .Y(n_416) );
INVx2_ASAP7_75t_L g262 ( .A(n_234), .Y(n_262) );
INVx3_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
INVx2_ASAP7_75t_L g486 ( .A(n_238), .Y(n_486) );
AND2x2_ASAP7_75t_L g267 ( .A(n_243), .B(n_268), .Y(n_267) );
INVx1_ASAP7_75t_L g289 ( .A(n_243), .Y(n_289) );
BUFx2_ASAP7_75t_L g295 ( .A(n_243), .Y(n_295) );
AND2x2_ASAP7_75t_L g314 ( .A(n_243), .B(n_287), .Y(n_314) );
INVx3_ASAP7_75t_L g326 ( .A(n_243), .Y(n_326) );
OR2x2_ASAP7_75t_L g336 ( .A(n_243), .B(n_287), .Y(n_336) );
AOI31xp33_ASAP7_75t_SL g251 ( .A1(n_252), .A2(n_266), .A3(n_269), .B(n_271), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_253), .B(n_265), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_253), .B(n_288), .Y(n_299) );
OR2x2_ASAP7_75t_L g323 ( .A(n_253), .B(n_293), .Y(n_323) );
INVx1_ASAP7_75t_SL g253 ( .A(n_254), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_254), .B(n_267), .Y(n_266) );
OR2x2_ASAP7_75t_L g344 ( .A(n_254), .B(n_336), .Y(n_344) );
NOR2xp33_ASAP7_75t_L g354 ( .A(n_254), .B(n_326), .Y(n_354) );
AND2x2_ASAP7_75t_L g361 ( .A(n_254), .B(n_362), .Y(n_361) );
NAND2x1_ASAP7_75t_L g389 ( .A(n_254), .B(n_325), .Y(n_389) );
NOR2xp33_ASAP7_75t_L g390 ( .A(n_254), .B(n_380), .Y(n_390) );
AND2x2_ASAP7_75t_L g402 ( .A(n_254), .B(n_287), .Y(n_402) );
INVx3_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
INVx3_ASAP7_75t_L g282 ( .A(n_255), .Y(n_282) );
INVx1_ASAP7_75t_L g348 ( .A(n_265), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_265), .B(n_402), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_267), .B(n_343), .Y(n_377) );
AND2x4_ASAP7_75t_L g288 ( .A(n_268), .B(n_289), .Y(n_288) );
CKINVDCx16_ASAP7_75t_R g269 ( .A(n_270), .Y(n_269) );
OR2x2_ASAP7_75t_L g271 ( .A(n_272), .B(n_273), .Y(n_271) );
INVx2_ASAP7_75t_L g367 ( .A(n_273), .Y(n_367) );
NOR2xp33_ASAP7_75t_L g384 ( .A(n_273), .B(n_385), .Y(n_384) );
AND2x2_ASAP7_75t_L g315 ( .A(n_274), .B(n_305), .Y(n_315) );
AND2x2_ASAP7_75t_L g409 ( .A(n_274), .B(n_279), .Y(n_409) );
INVx1_ASAP7_75t_L g434 ( .A(n_274), .Y(n_434) );
AOI221xp5_ASAP7_75t_L g275 ( .A1(n_276), .A2(n_280), .B1(n_283), .B2(n_284), .C(n_290), .Y(n_275) );
CKINVDCx14_ASAP7_75t_R g296 ( .A(n_276), .Y(n_296) );
AND2x2_ASAP7_75t_L g276 ( .A(n_277), .B(n_278), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_277), .B(n_298), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_280), .B(n_331), .Y(n_350) );
INVx3_ASAP7_75t_SL g280 ( .A(n_281), .Y(n_280) );
OR2x2_ASAP7_75t_L g399 ( .A(n_281), .B(n_295), .Y(n_399) );
AND2x2_ASAP7_75t_L g313 ( .A(n_282), .B(n_314), .Y(n_313) );
INVx1_ASAP7_75t_L g343 ( .A(n_282), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_282), .B(n_326), .Y(n_371) );
NOR3xp33_ASAP7_75t_L g413 ( .A(n_282), .B(n_383), .C(n_414), .Y(n_413) );
AOI211xp5_ASAP7_75t_SL g346 ( .A1(n_283), .A2(n_347), .B(n_349), .C(n_357), .Y(n_346) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
OAI22xp33_ASAP7_75t_L g335 ( .A1(n_285), .A2(n_336), .B1(n_337), .B2(n_338), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_286), .B(n_288), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_286), .B(n_325), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_286), .B(n_370), .Y(n_369) );
BUFx2_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
AND2x2_ASAP7_75t_L g428 ( .A(n_288), .B(n_402), .Y(n_428) );
OAI22xp5_ASAP7_75t_L g290 ( .A1(n_291), .A2(n_296), .B1(n_297), .B2(n_299), .Y(n_290) );
NOR2xp33_ASAP7_75t_SL g291 ( .A(n_292), .B(n_294), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_294), .B(n_343), .Y(n_374) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
OAI22xp5_ASAP7_75t_L g426 ( .A1(n_297), .A2(n_389), .B1(n_420), .B2(n_427), .Y(n_426) );
AOI221xp5_ASAP7_75t_L g300 ( .A1(n_301), .A2(n_308), .B1(n_310), .B2(n_315), .C(n_316), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
OR2x2_ASAP7_75t_L g302 ( .A(n_303), .B(n_306), .Y(n_302) );
HB1xp67_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
INVxp67_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
OAI221xp5_ASAP7_75t_L g316 ( .A1(n_306), .A2(n_317), .B1(n_323), .B2(n_324), .C(n_327), .Y(n_316) );
INVx1_ASAP7_75t_L g359 ( .A(n_307), .Y(n_359) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_312), .B(n_313), .Y(n_311) );
INVx1_ASAP7_75t_SL g331 ( .A(n_312), .Y(n_331) );
OR2x2_ASAP7_75t_L g404 ( .A(n_312), .B(n_336), .Y(n_404) );
AND2x2_ASAP7_75t_L g406 ( .A(n_312), .B(n_314), .Y(n_406) );
INVx1_ASAP7_75t_L g345 ( .A(n_315), .Y(n_345) );
OR2x2_ASAP7_75t_L g317 ( .A(n_318), .B(n_321), .Y(n_317) );
AOI21xp33_ASAP7_75t_SL g375 ( .A1(n_318), .A2(n_376), .B(n_377), .Y(n_375) );
OR2x2_ASAP7_75t_L g382 ( .A(n_318), .B(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
AND2x2_ASAP7_75t_L g356 ( .A(n_319), .B(n_340), .Y(n_356) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
NAND2xp33_ASAP7_75t_SL g373 ( .A(n_324), .B(n_374), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_325), .B(n_343), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_326), .B(n_362), .Y(n_425) );
O2A1O1Ixp33_ASAP7_75t_L g341 ( .A1(n_329), .A2(n_342), .B(n_344), .C(n_345), .Y(n_341) );
NAND2x1_ASAP7_75t_SL g366 ( .A(n_329), .B(n_367), .Y(n_366) );
AOI22xp5_ASAP7_75t_L g378 ( .A1(n_330), .A2(n_379), .B1(n_381), .B2(n_384), .Y(n_378) );
AND2x2_ASAP7_75t_L g330 ( .A(n_331), .B(n_332), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_332), .B(n_422), .Y(n_421) );
NAND5xp2_ASAP7_75t_L g333 ( .A(n_334), .B(n_346), .C(n_364), .D(n_378), .E(n_387), .Y(n_333) );
NOR2xp33_ASAP7_75t_L g334 ( .A(n_335), .B(n_341), .Y(n_334) );
INVx1_ASAP7_75t_L g391 ( .A(n_337), .Y(n_391) );
INVx1_ASAP7_75t_SL g338 ( .A(n_339), .Y(n_338) );
AOI221xp5_ASAP7_75t_L g397 ( .A1(n_339), .A2(n_358), .B1(n_398), .B2(n_400), .C(n_403), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_340), .B(n_434), .Y(n_433) );
NOR2xp33_ASAP7_75t_L g347 ( .A(n_343), .B(n_348), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_343), .B(n_409), .Y(n_412) );
OAI22xp5_ASAP7_75t_L g349 ( .A1(n_350), .A2(n_351), .B1(n_353), .B2(n_355), .Y(n_349) );
INVx1_ASAP7_75t_SL g351 ( .A(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
AND2x2_ASAP7_75t_L g357 ( .A(n_358), .B(n_361), .Y(n_357) );
AND2x2_ASAP7_75t_L g358 ( .A(n_359), .B(n_360), .Y(n_358) );
AND2x2_ASAP7_75t_L g431 ( .A(n_360), .B(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
AOI221xp5_ASAP7_75t_L g364 ( .A1(n_365), .A2(n_368), .B1(n_372), .B2(n_373), .C(n_375), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
AND2x2_ASAP7_75t_L g415 ( .A(n_370), .B(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVx1_ASAP7_75t_SL g422 ( .A(n_380), .Y(n_422) );
INVx1_ASAP7_75t_SL g381 ( .A(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
OAI21xp5_ASAP7_75t_SL g387 ( .A1(n_388), .A2(n_390), .B(n_391), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
OAI211xp5_ASAP7_75t_SL g392 ( .A1(n_393), .A2(n_395), .B(n_397), .C(n_410), .Y(n_392) );
INVx1_ASAP7_75t_SL g393 ( .A(n_394), .Y(n_393) );
A2O1A1Ixp33_ASAP7_75t_L g419 ( .A1(n_395), .A2(n_420), .B(n_421), .C(n_423), .Y(n_419) );
INVx1_ASAP7_75t_SL g395 ( .A(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
NAND2xp5_ASAP7_75t_SL g400 ( .A(n_399), .B(n_401), .Y(n_400) );
AOI21xp33_ASAP7_75t_L g403 ( .A1(n_404), .A2(n_405), .B(n_407), .Y(n_403) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx2_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
AOI21xp33_ASAP7_75t_L g429 ( .A1(n_430), .A2(n_433), .B(n_435), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx2_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g706 ( .A(n_437), .Y(n_706) );
INVx1_ASAP7_75t_L g707 ( .A(n_438), .Y(n_707) );
OR3x1_ASAP7_75t_L g438 ( .A(n_439), .B(n_612), .C(n_659), .Y(n_438) );
NAND3xp33_ASAP7_75t_SL g439 ( .A(n_440), .B(n_558), .C(n_583), .Y(n_439) );
AOI221xp5_ASAP7_75t_L g440 ( .A1(n_441), .A2(n_498), .B1(n_525), .B2(n_528), .C(n_536), .Y(n_440) );
OAI21xp5_ASAP7_75t_L g441 ( .A1(n_442), .A2(n_466), .B(n_491), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_443), .B(n_538), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_443), .B(n_541), .Y(n_656) );
AND2x2_ASAP7_75t_L g443 ( .A(n_444), .B(n_457), .Y(n_443) );
AND2x2_ASAP7_75t_L g527 ( .A(n_444), .B(n_497), .Y(n_527) );
AND2x2_ASAP7_75t_L g576 ( .A(n_444), .B(n_496), .Y(n_576) );
AND2x2_ASAP7_75t_L g597 ( .A(n_444), .B(n_598), .Y(n_597) );
AND2x2_ASAP7_75t_L g602 ( .A(n_444), .B(n_569), .Y(n_602) );
OR2x2_ASAP7_75t_L g610 ( .A(n_444), .B(n_611), .Y(n_610) );
AND2x2_ASAP7_75t_L g682 ( .A(n_444), .B(n_479), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_444), .B(n_631), .Y(n_696) );
INVx3_ASAP7_75t_SL g444 ( .A(n_445), .Y(n_444) );
AND2x2_ASAP7_75t_L g542 ( .A(n_445), .B(n_457), .Y(n_542) );
OR2x2_ASAP7_75t_L g543 ( .A(n_445), .B(n_479), .Y(n_543) );
AND2x4_ASAP7_75t_L g564 ( .A(n_445), .B(n_497), .Y(n_564) );
AND2x2_ASAP7_75t_L g594 ( .A(n_445), .B(n_468), .Y(n_594) );
AND2x2_ASAP7_75t_L g603 ( .A(n_445), .B(n_593), .Y(n_603) );
AND2x2_ASAP7_75t_L g619 ( .A(n_445), .B(n_480), .Y(n_619) );
OR2x2_ASAP7_75t_L g628 ( .A(n_445), .B(n_611), .Y(n_628) );
AND2x2_ASAP7_75t_L g634 ( .A(n_445), .B(n_569), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_445), .B(n_640), .Y(n_639) );
OR2x2_ASAP7_75t_L g648 ( .A(n_445), .B(n_493), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_445), .B(n_538), .Y(n_658) );
NAND2xp5_ASAP7_75t_SL g687 ( .A(n_445), .B(n_598), .Y(n_687) );
OR2x6_ASAP7_75t_L g445 ( .A(n_446), .B(n_455), .Y(n_445) );
INVx2_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
NAND2xp5_ASAP7_75t_SL g473 ( .A(n_453), .B(n_474), .Y(n_473) );
INVx2_ASAP7_75t_L g497 ( .A(n_457), .Y(n_497) );
AND2x2_ASAP7_75t_L g593 ( .A(n_457), .B(n_479), .Y(n_593) );
AND2x2_ASAP7_75t_L g598 ( .A(n_457), .B(n_480), .Y(n_598) );
INVx1_ASAP7_75t_L g654 ( .A(n_457), .Y(n_654) );
OA21x2_ASAP7_75t_L g457 ( .A1(n_458), .A2(n_459), .B(n_465), .Y(n_457) );
OA21x2_ASAP7_75t_L g509 ( .A1(n_458), .A2(n_510), .B(n_516), .Y(n_509) );
OA21x2_ASAP7_75t_L g517 ( .A1(n_458), .A2(n_518), .B(n_524), .Y(n_517) );
INVx1_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
AND2x2_ASAP7_75t_L g563 ( .A(n_467), .B(n_564), .Y(n_563) );
AND2x2_ASAP7_75t_L g467 ( .A(n_468), .B(n_479), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_468), .B(n_527), .Y(n_526) );
BUFx3_ASAP7_75t_L g541 ( .A(n_468), .Y(n_541) );
OR2x2_ASAP7_75t_L g611 ( .A(n_468), .B(n_479), .Y(n_611) );
OR2x2_ASAP7_75t_L g672 ( .A(n_468), .B(n_579), .Y(n_672) );
OA21x2_ASAP7_75t_L g468 ( .A1(n_469), .A2(n_470), .B(n_477), .Y(n_468) );
INVx1_ASAP7_75t_L g494 ( .A(n_470), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_477), .Y(n_495) );
AND2x2_ASAP7_75t_L g496 ( .A(n_479), .B(n_497), .Y(n_496) );
AND2x2_ASAP7_75t_L g631 ( .A(n_479), .B(n_493), .Y(n_631) );
INVx2_ASAP7_75t_SL g479 ( .A(n_480), .Y(n_479) );
BUFx2_ASAP7_75t_L g570 ( .A(n_480), .Y(n_570) );
INVx1_ASAP7_75t_SL g491 ( .A(n_492), .Y(n_491) );
AOI221xp5_ASAP7_75t_L g675 ( .A1(n_492), .A2(n_676), .B1(n_680), .B2(n_683), .C(n_684), .Y(n_675) );
AND2x2_ASAP7_75t_L g492 ( .A(n_493), .B(n_496), .Y(n_492) );
INVx1_ASAP7_75t_SL g539 ( .A(n_493), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_493), .B(n_654), .Y(n_653) );
AND2x2_ASAP7_75t_L g670 ( .A(n_493), .B(n_527), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_496), .B(n_541), .Y(n_662) );
AND2x2_ASAP7_75t_L g569 ( .A(n_497), .B(n_570), .Y(n_569) );
INVx1_ASAP7_75t_SL g573 ( .A(n_498), .Y(n_573) );
NAND2xp5_ASAP7_75t_SL g609 ( .A(n_498), .B(n_579), .Y(n_609) );
AND2x2_ASAP7_75t_L g498 ( .A(n_499), .B(n_508), .Y(n_498) );
AND2x2_ASAP7_75t_L g535 ( .A(n_499), .B(n_509), .Y(n_535) );
INVx4_ASAP7_75t_L g547 ( .A(n_499), .Y(n_547) );
BUFx3_ASAP7_75t_L g589 ( .A(n_499), .Y(n_589) );
AND3x2_ASAP7_75t_L g604 ( .A(n_499), .B(n_605), .C(n_606), .Y(n_604) );
AND2x2_ASAP7_75t_L g686 ( .A(n_508), .B(n_600), .Y(n_686) );
AND2x2_ASAP7_75t_L g694 ( .A(n_508), .B(n_579), .Y(n_694) );
INVx1_ASAP7_75t_SL g699 ( .A(n_508), .Y(n_699) );
AND2x2_ASAP7_75t_L g508 ( .A(n_509), .B(n_517), .Y(n_508) );
INVx1_ASAP7_75t_SL g557 ( .A(n_509), .Y(n_557) );
AND2x2_ASAP7_75t_L g580 ( .A(n_509), .B(n_547), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_509), .B(n_531), .Y(n_582) );
HB1xp67_ASAP7_75t_L g622 ( .A(n_509), .Y(n_622) );
OR2x2_ASAP7_75t_L g627 ( .A(n_509), .B(n_547), .Y(n_627) );
INVx2_ASAP7_75t_L g533 ( .A(n_517), .Y(n_533) );
AND2x2_ASAP7_75t_L g567 ( .A(n_517), .B(n_548), .Y(n_567) );
OR2x2_ASAP7_75t_L g587 ( .A(n_517), .B(n_548), .Y(n_587) );
HB1xp67_ASAP7_75t_L g607 ( .A(n_517), .Y(n_607) );
INVx1_ASAP7_75t_SL g525 ( .A(n_526), .Y(n_525) );
AOI21xp33_ASAP7_75t_L g657 ( .A1(n_526), .A2(n_566), .B(n_658), .Y(n_657) );
AOI322xp5_ASAP7_75t_L g693 ( .A1(n_528), .A2(n_538), .A3(n_564), .B1(n_694), .B2(n_695), .C1(n_697), .C2(n_700), .Y(n_693) );
INVx1_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
OR2x2_ASAP7_75t_L g529 ( .A(n_530), .B(n_534), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_530), .B(n_637), .Y(n_636) );
INVx1_ASAP7_75t_SL g530 ( .A(n_531), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_531), .B(n_561), .Y(n_560) );
INVx2_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
AND2x2_ASAP7_75t_L g556 ( .A(n_532), .B(n_557), .Y(n_556) );
INVx2_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
AND2x2_ASAP7_75t_L g624 ( .A(n_533), .B(n_547), .Y(n_624) );
AND2x2_ASAP7_75t_L g691 ( .A(n_533), .B(n_548), .Y(n_691) );
INVx1_ASAP7_75t_SL g534 ( .A(n_535), .Y(n_534) );
AND2x2_ASAP7_75t_L g632 ( .A(n_535), .B(n_586), .Y(n_632) );
AOI31xp33_ASAP7_75t_L g536 ( .A1(n_537), .A2(n_540), .A3(n_543), .B(n_544), .Y(n_536) );
AND2x2_ASAP7_75t_L g591 ( .A(n_538), .B(n_569), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_538), .B(n_561), .Y(n_673) );
AND2x2_ASAP7_75t_L g692 ( .A(n_538), .B(n_597), .Y(n_692) );
INVx2_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_541), .B(n_542), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_541), .B(n_569), .Y(n_581) );
NAND2x1p5_ASAP7_75t_L g615 ( .A(n_541), .B(n_598), .Y(n_615) );
NAND2xp5_ASAP7_75t_SL g618 ( .A(n_541), .B(n_619), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_541), .B(n_682), .Y(n_681) );
NOR2xp33_ASAP7_75t_L g630 ( .A(n_542), .B(n_598), .Y(n_630) );
INVx1_ASAP7_75t_L g674 ( .A(n_542), .Y(n_674) );
INVx1_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
AND2x2_ASAP7_75t_L g545 ( .A(n_546), .B(n_556), .Y(n_545) );
INVxp67_ASAP7_75t_L g626 ( .A(n_546), .Y(n_626) );
NOR2xp33_ASAP7_75t_L g546 ( .A(n_547), .B(n_548), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_547), .B(n_557), .Y(n_562) );
INVx1_ASAP7_75t_L g668 ( .A(n_547), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_547), .B(n_645), .Y(n_679) );
BUFx3_ASAP7_75t_L g579 ( .A(n_548), .Y(n_579) );
AND2x2_ASAP7_75t_L g605 ( .A(n_548), .B(n_557), .Y(n_605) );
INVx2_ASAP7_75t_L g645 ( .A(n_548), .Y(n_645) );
NAND2xp5_ASAP7_75t_SL g677 ( .A(n_556), .B(n_678), .Y(n_677) );
AOI211xp5_ASAP7_75t_L g558 ( .A1(n_559), .A2(n_563), .B(n_565), .C(n_574), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
AOI21xp33_ASAP7_75t_L g608 ( .A1(n_560), .A2(n_609), .B(n_610), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_561), .B(n_567), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_561), .B(n_600), .Y(n_599) );
INVx1_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
OR2x2_ASAP7_75t_L g641 ( .A(n_562), .B(n_587), .Y(n_641) );
INVx3_ASAP7_75t_L g572 ( .A(n_564), .Y(n_572) );
OAI22xp5_ASAP7_75t_SL g565 ( .A1(n_566), .A2(n_568), .B1(n_571), .B2(n_573), .Y(n_565) );
OAI21xp5_ASAP7_75t_SL g590 ( .A1(n_567), .A2(n_591), .B(n_592), .Y(n_590) );
AND2x2_ASAP7_75t_L g616 ( .A(n_567), .B(n_580), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_567), .B(n_668), .Y(n_667) );
INVxp67_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
OR2x2_ASAP7_75t_L g571 ( .A(n_570), .B(n_572), .Y(n_571) );
INVx1_ASAP7_75t_L g640 ( .A(n_570), .Y(n_640) );
OAI21xp5_ASAP7_75t_SL g584 ( .A1(n_571), .A2(n_585), .B(n_590), .Y(n_584) );
OAI22xp33_ASAP7_75t_SL g574 ( .A1(n_575), .A2(n_577), .B1(n_581), .B2(n_582), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
NOR2xp33_ASAP7_75t_L g651 ( .A(n_576), .B(n_652), .Y(n_651) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
AND2x2_ASAP7_75t_L g578 ( .A(n_579), .B(n_580), .Y(n_578) );
INVx1_ASAP7_75t_L g600 ( .A(n_579), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_579), .B(n_622), .Y(n_621) );
NOR3xp33_ASAP7_75t_L g583 ( .A(n_584), .B(n_595), .C(n_608), .Y(n_583) );
OAI22xp5_ASAP7_75t_SL g650 ( .A1(n_585), .A2(n_651), .B1(n_655), .B2(n_656), .Y(n_650) );
NAND2xp5_ASAP7_75t_SL g585 ( .A(n_586), .B(n_588), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
OR2x2_ASAP7_75t_L g655 ( .A(n_587), .B(n_588), .Y(n_655) );
AND2x2_ASAP7_75t_L g663 ( .A(n_588), .B(n_644), .Y(n_663) );
CKINVDCx16_ASAP7_75t_R g588 ( .A(n_589), .Y(n_588) );
O2A1O1Ixp33_ASAP7_75t_SL g671 ( .A1(n_589), .A2(n_672), .B(n_673), .C(n_674), .Y(n_671) );
OR2x2_ASAP7_75t_L g698 ( .A(n_589), .B(n_699), .Y(n_698) );
AND2x2_ASAP7_75t_L g592 ( .A(n_593), .B(n_594), .Y(n_592) );
OAI21xp33_ASAP7_75t_L g595 ( .A1(n_596), .A2(n_599), .B(n_601), .Y(n_595) );
INVx1_ASAP7_75t_SL g596 ( .A(n_597), .Y(n_596) );
O2A1O1Ixp33_ASAP7_75t_L g633 ( .A1(n_597), .A2(n_634), .B(n_635), .C(n_638), .Y(n_633) );
OAI21xp33_ASAP7_75t_SL g601 ( .A1(n_602), .A2(n_603), .B(n_604), .Y(n_601) );
AND2x2_ASAP7_75t_L g666 ( .A(n_605), .B(n_624), .Y(n_666) );
INVxp67_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
AND2x2_ASAP7_75t_L g644 ( .A(n_607), .B(n_645), .Y(n_644) );
INVx1_ASAP7_75t_L g649 ( .A(n_609), .Y(n_649) );
NAND3xp33_ASAP7_75t_SL g612 ( .A(n_613), .B(n_633), .C(n_646), .Y(n_612) );
AOI211xp5_ASAP7_75t_L g613 ( .A1(n_614), .A2(n_616), .B(n_617), .C(n_625), .Y(n_613) );
INVx1_ASAP7_75t_SL g614 ( .A(n_615), .Y(n_614) );
NOR2xp33_ASAP7_75t_L g617 ( .A(n_618), .B(n_620), .Y(n_617) );
INVx1_ASAP7_75t_L g683 ( .A(n_620), .Y(n_683) );
OR2x2_ASAP7_75t_L g620 ( .A(n_621), .B(n_623), .Y(n_620) );
INVx1_ASAP7_75t_L g643 ( .A(n_622), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_622), .B(n_691), .Y(n_690) );
INVxp67_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
A2O1A1Ixp33_ASAP7_75t_L g625 ( .A1(n_626), .A2(n_627), .B(n_628), .C(n_629), .Y(n_625) );
INVx2_ASAP7_75t_SL g637 ( .A(n_627), .Y(n_637) );
OAI22xp5_ASAP7_75t_L g638 ( .A1(n_628), .A2(n_639), .B1(n_641), .B2(n_642), .Y(n_638) );
OAI21xp33_ASAP7_75t_SL g629 ( .A1(n_630), .A2(n_631), .B(n_632), .Y(n_629) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_643), .B(n_644), .Y(n_642) );
AOI211xp5_ASAP7_75t_L g646 ( .A1(n_647), .A2(n_649), .B(n_650), .C(n_657), .Y(n_646) );
INVx1_ASAP7_75t_SL g647 ( .A(n_648), .Y(n_647) );
INVxp33_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
INVx1_ASAP7_75t_L g700 ( .A(n_654), .Y(n_700) );
NAND4xp25_ASAP7_75t_L g659 ( .A(n_660), .B(n_675), .C(n_688), .D(n_693), .Y(n_659) );
AOI211xp5_ASAP7_75t_L g660 ( .A1(n_661), .A2(n_663), .B(n_664), .C(n_671), .Y(n_660) );
INVx1_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
AOI21xp5_ASAP7_75t_L g664 ( .A1(n_665), .A2(n_667), .B(n_669), .Y(n_664) );
AOI21xp33_ASAP7_75t_L g684 ( .A1(n_665), .A2(n_685), .B(n_687), .Y(n_684) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
NOR2xp33_ASAP7_75t_L g697 ( .A(n_672), .B(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_689), .B(n_692), .Y(n_688) );
INVxp67_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
INVx1_ASAP7_75t_L g709 ( .A(n_701), .Y(n_709) );
OAI22xp5_ASAP7_75t_SL g703 ( .A1(n_704), .A2(n_705), .B1(n_707), .B2(n_708), .Y(n_703) );
INVx2_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVx2_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
INVx1_ASAP7_75t_SL g710 ( .A(n_711), .Y(n_710) );
INVx3_ASAP7_75t_SL g711 ( .A(n_712), .Y(n_711) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
endmodule