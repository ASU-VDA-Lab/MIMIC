module fake_jpeg_21104_n_39 (n_3, n_2, n_1, n_0, n_4, n_5, n_39);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_39;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

CKINVDCx20_ASAP7_75t_R g6 ( 
.A(n_2),
.Y(n_6)
);

BUFx12f_ASAP7_75t_L g7 ( 
.A(n_5),
.Y(n_7)
);

INVx3_ASAP7_75t_L g8 ( 
.A(n_0),
.Y(n_8)
);

INVx6_ASAP7_75t_L g9 ( 
.A(n_1),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_1),
.Y(n_10)
);

INVx1_ASAP7_75t_SL g11 ( 
.A(n_4),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_7),
.Y(n_12)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx6_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_13),
.B(n_14),
.Y(n_19)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

AOI22xp5_ASAP7_75t_L g15 ( 
.A1(n_9),
.A2(n_8),
.B1(n_11),
.B2(n_10),
.Y(n_15)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_15),
.A2(n_11),
.B(n_6),
.Y(n_20)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_16),
.Y(n_22)
);

HB1xp67_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_17),
.Y(n_18)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_20),
.A2(n_9),
.B1(n_8),
.B2(n_3),
.Y(n_24)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_19),
.Y(n_23)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_24),
.B(n_25),
.Y(n_29)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_21),
.Y(n_25)
);

NOR3xp33_ASAP7_75t_SL g26 ( 
.A(n_18),
.B(n_17),
.C(n_12),
.Y(n_26)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_26),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_26),
.B(n_22),
.Y(n_28)
);

XNOR2xp5_ASAP7_75t_L g32 ( 
.A(n_28),
.B(n_29),
.Y(n_32)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_30),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_31),
.B(n_32),
.Y(n_34)
);

HB1xp67_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

AOI21xp33_ASAP7_75t_SL g35 ( 
.A1(n_33),
.A2(n_27),
.B(n_2),
.Y(n_35)
);

OAI21xp5_ASAP7_75t_L g37 ( 
.A1(n_35),
.A2(n_36),
.B(n_27),
.Y(n_37)
);

AO21x1_ASAP7_75t_L g36 ( 
.A1(n_33),
.A2(n_27),
.B(n_18),
.Y(n_36)
);

XOR2xp5_ASAP7_75t_L g39 ( 
.A(n_37),
.B(n_38),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_34),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_38)
);


endmodule