module fake_jpeg_27793_n_415 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_415);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_415;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx5p33_ASAP7_75t_R g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVxp67_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx4f_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_10),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_15),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_6),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g126 ( 
.A(n_45),
.Y(n_126)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_46),
.Y(n_98)
);

INVx3_ASAP7_75t_SL g47 ( 
.A(n_20),
.Y(n_47)
);

INVx5_ASAP7_75t_SL g127 ( 
.A(n_47),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_48),
.Y(n_95)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_49),
.Y(n_92)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_50),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_27),
.B(n_14),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_51),
.B(n_53),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_19),
.Y(n_52)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_52),
.Y(n_105)
);

INVx1_ASAP7_75t_SL g53 ( 
.A(n_23),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_23),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_54),
.B(n_58),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_55),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_56),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_57),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_33),
.B(n_7),
.Y(n_58)
);

BUFx10_ASAP7_75t_L g59 ( 
.A(n_30),
.Y(n_59)
);

INVx8_ASAP7_75t_L g133 ( 
.A(n_59),
.Y(n_133)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_28),
.Y(n_60)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_60),
.Y(n_116)
);

HB1xp67_ASAP7_75t_L g61 ( 
.A(n_30),
.Y(n_61)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_61),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

BUFx2_ASAP7_75t_L g104 ( 
.A(n_62),
.Y(n_104)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g131 ( 
.A(n_63),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_28),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_64),
.Y(n_93)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_28),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_65),
.Y(n_99)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_34),
.Y(n_66)
);

BUFx2_ASAP7_75t_L g124 ( 
.A(n_66),
.Y(n_124)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_67),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_68),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_69),
.Y(n_114)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_29),
.Y(n_70)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_70),
.Y(n_110)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_71),
.Y(n_103)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_72),
.Y(n_109)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_30),
.Y(n_73)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_73),
.Y(n_94)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_41),
.Y(n_74)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_74),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_30),
.Y(n_75)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_75),
.Y(n_108)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_29),
.Y(n_76)
);

INVx11_ASAP7_75t_L g112 ( 
.A(n_76),
.Y(n_112)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_41),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_77),
.B(n_78),
.Y(n_90)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_42),
.Y(n_78)
);

HB1xp67_ASAP7_75t_L g79 ( 
.A(n_20),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_79),
.Y(n_88)
);

INVx11_ASAP7_75t_L g80 ( 
.A(n_29),
.Y(n_80)
);

INVx11_ASAP7_75t_L g113 ( 
.A(n_80),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_33),
.B(n_7),
.Y(n_81)
);

OR2x2_ASAP7_75t_L g115 ( 
.A(n_81),
.B(n_83),
.Y(n_115)
);

BUFx5_ASAP7_75t_L g82 ( 
.A(n_24),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_82),
.Y(n_102)
);

NOR2xp67_ASAP7_75t_L g83 ( 
.A(n_42),
.B(n_44),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_40),
.B(n_7),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_84),
.B(n_18),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_44),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_85),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_40),
.B(n_6),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_86),
.B(n_11),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_86),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_91),
.B(n_24),
.Y(n_135)
);

INVx13_ASAP7_75t_L g96 ( 
.A(n_47),
.Y(n_96)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_96),
.Y(n_138)
);

BUFx12_ASAP7_75t_L g97 ( 
.A(n_62),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g142 ( 
.A(n_97),
.Y(n_142)
);

BUFx12_ASAP7_75t_L g106 ( 
.A(n_67),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g156 ( 
.A(n_106),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_48),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_117),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_118),
.A2(n_130),
.B(n_26),
.Y(n_157)
);

AND2x2_ASAP7_75t_SL g119 ( 
.A(n_68),
.B(n_42),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_119),
.B(n_121),
.C(n_89),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_53),
.B(n_18),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_70),
.A2(n_32),
.B1(n_21),
.B2(n_36),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_122),
.A2(n_16),
.B1(n_35),
.B2(n_31),
.Y(n_144)
);

INVx2_ASAP7_75t_R g129 ( 
.A(n_63),
.Y(n_129)
);

INVx1_ASAP7_75t_SL g159 ( 
.A(n_129),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_135),
.B(n_157),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_115),
.A2(n_76),
.B1(n_80),
.B2(n_17),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_136),
.A2(n_39),
.B1(n_169),
.B2(n_166),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_95),
.A2(n_45),
.B1(n_17),
.B2(n_71),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_137),
.A2(n_145),
.B1(n_96),
.B2(n_108),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_129),
.Y(n_139)
);

INVx13_ASAP7_75t_L g198 ( 
.A(n_139),
.Y(n_198)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_98),
.Y(n_140)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_140),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g190 ( 
.A(n_141),
.B(n_144),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_123),
.B(n_26),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_143),
.B(n_150),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_95),
.A2(n_65),
.B1(n_60),
.B2(n_22),
.Y(n_145)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_100),
.Y(n_146)
);

INVx6_ASAP7_75t_L g185 ( 
.A(n_146),
.Y(n_185)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_125),
.Y(n_147)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_147),
.Y(n_200)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_100),
.Y(n_148)
);

INVx1_ASAP7_75t_SL g197 ( 
.A(n_148),
.Y(n_197)
);

INVx8_ASAP7_75t_L g149 ( 
.A(n_92),
.Y(n_149)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_149),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_88),
.B(n_36),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_115),
.B(n_25),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_151),
.B(n_152),
.Y(n_179)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_90),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_91),
.B(n_25),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_153),
.B(n_155),
.Y(n_182)
);

INVx6_ASAP7_75t_L g154 ( 
.A(n_110),
.Y(n_154)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_154),
.Y(n_209)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_87),
.Y(n_155)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_87),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_158),
.B(n_161),
.Y(n_186)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_131),
.Y(n_160)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_160),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_119),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_101),
.B(n_35),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_162),
.B(n_165),
.Y(n_195)
);

BUFx3_ASAP7_75t_L g163 ( 
.A(n_97),
.Y(n_163)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_163),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_112),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_164),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_127),
.B(n_21),
.Y(n_165)
);

INVx6_ASAP7_75t_L g166 ( 
.A(n_93),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_166),
.B(n_167),
.Y(n_204)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_132),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_127),
.B(n_31),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_168),
.B(n_169),
.Y(n_208)
);

INVx6_ASAP7_75t_L g169 ( 
.A(n_93),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_92),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_170),
.B(n_146),
.Y(n_203)
);

INVx8_ASAP7_75t_L g171 ( 
.A(n_113),
.Y(n_171)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_171),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_113),
.Y(n_172)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_172),
.Y(n_191)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_105),
.Y(n_173)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_173),
.Y(n_196)
);

INVx4_ASAP7_75t_L g174 ( 
.A(n_131),
.Y(n_174)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_174),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_120),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g205 ( 
.A(n_175),
.B(n_164),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_134),
.B(n_107),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_176),
.B(n_187),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_145),
.A2(n_108),
.B1(n_128),
.B2(n_109),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_177),
.A2(n_207),
.B1(n_212),
.B2(n_158),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_139),
.B(n_16),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_159),
.B(n_103),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_188),
.B(n_69),
.C(n_56),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_159),
.B(n_75),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_192),
.B(n_193),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_175),
.B(n_59),
.Y(n_193)
);

AND2x2_ASAP7_75t_SL g194 ( 
.A(n_149),
.B(n_133),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g238 ( 
.A(n_194),
.B(n_126),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_155),
.B(n_59),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_201),
.B(n_203),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_202),
.A2(n_138),
.B1(n_38),
.B2(n_99),
.Y(n_235)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_205),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_137),
.A2(n_73),
.B1(n_94),
.B2(n_133),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_154),
.A2(n_39),
.B(n_22),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_210),
.A2(n_102),
.B(n_124),
.Y(n_246)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_206),
.Y(n_213)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_213),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_L g251 ( 
.A1(n_214),
.A2(n_209),
.B1(n_177),
.B2(n_185),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_215),
.B(n_207),
.Y(n_247)
);

INVx13_ASAP7_75t_L g216 ( 
.A(n_211),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_216),
.B(n_222),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_202),
.A2(n_148),
.B1(n_94),
.B2(n_116),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_218),
.A2(n_235),
.B1(n_197),
.B2(n_198),
.Y(n_272)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_206),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_198),
.A2(n_171),
.B1(n_174),
.B2(n_160),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g265 ( 
.A(n_223),
.Y(n_265)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_176),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_224),
.B(n_229),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_208),
.B(n_156),
.Y(n_225)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_225),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_178),
.B(n_156),
.Y(n_226)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_226),
.Y(n_259)
);

BUFx24_ASAP7_75t_L g227 ( 
.A(n_211),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_227),
.B(n_230),
.Y(n_270)
);

A2O1A1Ixp33_ASAP7_75t_L g228 ( 
.A1(n_190),
.A2(n_38),
.B(n_10),
.C(n_12),
.Y(n_228)
);

A2O1A1Ixp33_ASAP7_75t_L g266 ( 
.A1(n_228),
.A2(n_210),
.B(n_187),
.C(n_205),
.Y(n_266)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_193),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_180),
.Y(n_230)
);

BUFx4f_ASAP7_75t_SL g231 ( 
.A(n_209),
.Y(n_231)
);

INVx3_ASAP7_75t_L g250 ( 
.A(n_231),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_201),
.A2(n_49),
.B1(n_85),
.B2(n_99),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_232),
.A2(n_240),
.B1(n_197),
.B2(n_184),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_204),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_233),
.B(n_234),
.Y(n_271)
);

NOR3xp33_ASAP7_75t_L g234 ( 
.A(n_179),
.B(n_126),
.C(n_131),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_198),
.A2(n_138),
.B1(n_102),
.B2(n_124),
.Y(n_236)
);

CKINVDCx14_ASAP7_75t_R g274 ( 
.A(n_236),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_195),
.B(n_163),
.Y(n_237)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_237),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_L g252 ( 
.A1(n_238),
.A2(n_242),
.B(n_246),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_203),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_239),
.B(n_243),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_189),
.A2(n_44),
.B1(n_114),
.B2(n_111),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_182),
.B(n_142),
.Y(n_241)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_241),
.Y(n_261)
);

O2A1O1Ixp33_ASAP7_75t_L g242 ( 
.A1(n_192),
.A2(n_64),
.B(n_55),
.C(n_52),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_180),
.Y(n_243)
);

BUFx12f_ASAP7_75t_L g244 ( 
.A(n_199),
.Y(n_244)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_244),
.Y(n_262)
);

INVx3_ASAP7_75t_L g245 ( 
.A(n_185),
.Y(n_245)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_245),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_247),
.B(n_248),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_215),
.B(n_188),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_224),
.B(n_186),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_249),
.B(n_254),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_251),
.A2(n_268),
.B1(n_233),
.B2(n_245),
.Y(n_279)
);

OA22x2_ASAP7_75t_L g253 ( 
.A1(n_214),
.A2(n_194),
.B1(n_205),
.B2(n_212),
.Y(n_253)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_253),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_229),
.B(n_190),
.C(n_189),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_217),
.B(n_190),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_256),
.B(n_257),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_238),
.B(n_194),
.C(n_181),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_239),
.B(n_194),
.Y(n_263)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_263),
.Y(n_304)
);

AO21x1_ASAP7_75t_L g300 ( 
.A1(n_266),
.A2(n_231),
.B(n_9),
.Y(n_300)
);

AOI22xp33_ASAP7_75t_L g293 ( 
.A1(n_272),
.A2(n_200),
.B1(n_216),
.B2(n_230),
.Y(n_293)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_220),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_273),
.B(n_199),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_235),
.A2(n_181),
.B1(n_196),
.B2(n_183),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_276),
.A2(n_222),
.B1(n_213),
.B2(n_243),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_219),
.B(n_196),
.Y(n_277)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_277),
.Y(n_287)
);

OAI22x1_ASAP7_75t_L g278 ( 
.A1(n_265),
.A2(n_246),
.B1(n_238),
.B2(n_218),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_278),
.A2(n_301),
.B1(n_302),
.B2(n_274),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_279),
.A2(n_280),
.B1(n_281),
.B2(n_290),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_268),
.A2(n_221),
.B1(n_219),
.B2(n_242),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_253),
.A2(n_232),
.B1(n_183),
.B2(n_228),
.Y(n_281)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_270),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_283),
.B(n_291),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_275),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_284),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_255),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_285),
.Y(n_327)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_277),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_288),
.B(n_295),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_253),
.A2(n_191),
.B1(n_200),
.B2(n_184),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_267),
.Y(n_291)
);

CKINVDCx14_ASAP7_75t_R g322 ( 
.A(n_293),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_250),
.B(n_227),
.Y(n_294)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_294),
.Y(n_308)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_271),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_250),
.B(n_227),
.Y(n_296)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_296),
.Y(n_310)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_263),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_297),
.B(n_299),
.Y(n_314)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_298),
.Y(n_318)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_276),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_300),
.B(n_266),
.Y(n_319)
);

OAI22x1_ASAP7_75t_L g302 ( 
.A1(n_265),
.A2(n_231),
.B1(n_244),
.B2(n_142),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_253),
.A2(n_191),
.B1(n_244),
.B2(n_114),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_303),
.A2(n_272),
.B1(n_262),
.B2(n_264),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_289),
.B(n_248),
.C(n_247),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_305),
.B(n_313),
.C(n_328),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_289),
.B(n_254),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g342 ( 
.A(n_307),
.B(n_315),
.Y(n_342)
);

BUFx2_ASAP7_75t_L g311 ( 
.A(n_302),
.Y(n_311)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_311),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_312),
.A2(n_269),
.B1(n_111),
.B2(n_172),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_282),
.B(n_256),
.C(n_257),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_282),
.B(n_249),
.Y(n_315)
);

HB1xp67_ASAP7_75t_L g316 ( 
.A(n_292),
.Y(n_316)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_316),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_319),
.B(n_324),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_L g321 ( 
.A1(n_286),
.A2(n_252),
.B(n_258),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_L g334 ( 
.A1(n_321),
.A2(n_300),
.B(n_278),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_287),
.B(n_261),
.Y(n_323)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_323),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_287),
.B(n_260),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_325),
.A2(n_286),
.B1(n_299),
.B2(n_301),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_292),
.B(n_252),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g348 ( 
.A(n_326),
.B(n_57),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_288),
.B(n_259),
.C(n_244),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_305),
.B(n_290),
.C(n_304),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_330),
.B(n_332),
.C(n_313),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_307),
.B(n_304),
.C(n_297),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_333),
.A2(n_340),
.B1(n_343),
.B2(n_322),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_334),
.B(n_348),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_306),
.B(n_280),
.Y(n_336)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_336),
.Y(n_356)
);

INVxp67_ASAP7_75t_L g337 ( 
.A(n_317),
.Y(n_337)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_337),
.Y(n_358)
);

INVxp67_ASAP7_75t_L g338 ( 
.A(n_328),
.Y(n_338)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_338),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_320),
.A2(n_303),
.B1(n_281),
.B2(n_269),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_341),
.A2(n_310),
.B1(n_308),
.B2(n_309),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_320),
.A2(n_104),
.B1(n_1),
.B2(n_2),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_SL g344 ( 
.A1(n_311),
.A2(n_106),
.B(n_1),
.Y(n_344)
);

CKINVDCx16_ASAP7_75t_R g357 ( 
.A(n_344),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_306),
.B(n_0),
.Y(n_346)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_346),
.Y(n_363)
);

AOI21xp5_ASAP7_75t_L g347 ( 
.A1(n_321),
.A2(n_0),
.B(n_1),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_347),
.B(n_319),
.Y(n_355)
);

XOR2xp5_ASAP7_75t_L g365 ( 
.A(n_349),
.B(n_359),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_350),
.A2(n_352),
.B1(n_360),
.B2(n_341),
.Y(n_374)
);

XOR2xp5_ASAP7_75t_SL g351 ( 
.A(n_334),
.B(n_326),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_SL g375 ( 
.A(n_351),
.B(n_348),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_340),
.A2(n_312),
.B1(n_325),
.B2(n_314),
.Y(n_352)
);

INVx2_ASAP7_75t_SL g353 ( 
.A(n_339),
.Y(n_353)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_353),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_330),
.B(n_315),
.C(n_324),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_354),
.B(n_359),
.Y(n_371)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_355),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_329),
.B(n_323),
.C(n_314),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_346),
.B(n_327),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_SL g368 ( 
.A(n_362),
.B(n_318),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_365),
.B(n_332),
.C(n_361),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_L g366 ( 
.A(n_349),
.B(n_329),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_366),
.B(n_373),
.Y(n_385)
);

HB1xp67_ASAP7_75t_L g367 ( 
.A(n_354),
.Y(n_367)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_367),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_368),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_L g369 ( 
.A1(n_357),
.A2(n_336),
.B1(n_331),
.B2(n_345),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_369),
.B(n_370),
.Y(n_386)
);

INVx1_ASAP7_75t_SL g370 ( 
.A(n_353),
.Y(n_370)
);

HB1xp67_ASAP7_75t_L g373 ( 
.A(n_351),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_374),
.B(n_376),
.Y(n_382)
);

XNOR2x1_ASAP7_75t_L g380 ( 
.A(n_375),
.B(n_364),
.Y(n_380)
);

INVx13_ASAP7_75t_L g376 ( 
.A(n_358),
.Y(n_376)
);

OAI21xp5_ASAP7_75t_SL g379 ( 
.A1(n_371),
.A2(n_338),
.B(n_337),
.Y(n_379)
);

AOI21xp5_ASAP7_75t_SL g390 ( 
.A1(n_379),
.A2(n_372),
.B(n_347),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g394 ( 
.A(n_380),
.B(n_333),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_381),
.B(n_383),
.C(n_366),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_365),
.B(n_342),
.C(n_364),
.Y(n_383)
);

FAx1_ASAP7_75t_SL g384 ( 
.A(n_375),
.B(n_335),
.CI(n_352),
.CON(n_384),
.SN(n_384)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_384),
.B(n_342),
.Y(n_392)
);

OAI21xp5_ASAP7_75t_L g388 ( 
.A1(n_377),
.A2(n_356),
.B(n_335),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_SL g396 ( 
.A(n_388),
.B(n_376),
.Y(n_396)
);

XOR2xp5_ASAP7_75t_L g402 ( 
.A(n_389),
.B(n_394),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_390),
.B(n_386),
.Y(n_400)
);

AND2x2_ASAP7_75t_L g391 ( 
.A(n_381),
.B(n_360),
.Y(n_391)
);

AOI21xp5_ASAP7_75t_L g398 ( 
.A1(n_391),
.A2(n_393),
.B(n_380),
.Y(n_398)
);

OR2x2_ASAP7_75t_L g401 ( 
.A(n_392),
.B(n_395),
.Y(n_401)
);

AND2x2_ASAP7_75t_L g393 ( 
.A(n_385),
.B(n_370),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_385),
.B(n_350),
.C(n_363),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_SL g399 ( 
.A(n_396),
.B(n_397),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_SL g397 ( 
.A1(n_382),
.A2(n_343),
.B1(n_344),
.B2(n_12),
.Y(n_397)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_398),
.Y(n_405)
);

AOI21xp5_ASAP7_75t_L g404 ( 
.A1(n_400),
.A2(n_378),
.B(n_396),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_392),
.B(n_387),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_403),
.B(n_388),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_404),
.B(n_399),
.C(n_384),
.Y(n_409)
);

AOI21xp5_ASAP7_75t_L g408 ( 
.A1(n_406),
.A2(n_407),
.B(n_401),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_L g407 ( 
.A(n_402),
.B(n_383),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_408),
.Y(n_410)
);

A2O1A1Ixp33_ASAP7_75t_L g411 ( 
.A1(n_410),
.A2(n_409),
.B(n_399),
.C(n_405),
.Y(n_411)
);

AOI322xp5_ASAP7_75t_L g412 ( 
.A1(n_411),
.A2(n_384),
.A3(n_104),
.B1(n_126),
.B2(n_9),
.C1(n_5),
.C2(n_2),
.Y(n_412)
);

AOI221xp5_ASAP7_75t_L g413 ( 
.A1(n_412),
.A2(n_9),
.B1(n_1),
.B2(n_2),
.C(n_5),
.Y(n_413)
);

XOR2xp5_ASAP7_75t_L g414 ( 
.A(n_413),
.B(n_0),
.Y(n_414)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_414),
.B(n_5),
.Y(n_415)
);


endmodule