module fake_jpeg_25506_n_335 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_335);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_335;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_260;
wire n_199;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_8),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_6),
.B(n_12),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_14),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_14),
.Y(n_27)
);

INVx1_ASAP7_75t_SL g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

INVx1_ASAP7_75t_SL g34 ( 
.A(n_0),
.Y(n_34)
);

AND2x2_ASAP7_75t_SL g35 ( 
.A(n_30),
.B(n_0),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_35),
.B(n_39),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

INVx2_ASAP7_75t_SL g39 ( 
.A(n_30),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_41),
.B(n_43),
.Y(n_64)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_45),
.Y(n_51)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_46),
.Y(n_101)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_47),
.B(n_49),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_35),
.B(n_21),
.Y(n_49)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_52),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_41),
.A2(n_21),
.B1(n_20),
.B2(n_24),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_54),
.A2(n_56),
.B1(n_61),
.B2(n_34),
.Y(n_81)
);

OAI22xp33_ASAP7_75t_L g56 ( 
.A1(n_37),
.A2(n_25),
.B1(n_24),
.B2(n_42),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_57),
.Y(n_80)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_58),
.Y(n_87)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_59),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_43),
.A2(n_21),
.B1(n_24),
.B2(n_25),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_41),
.B(n_18),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_62),
.B(n_28),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_49),
.A2(n_44),
.B1(n_25),
.B2(n_37),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_66),
.A2(n_75),
.B1(n_40),
.B2(n_38),
.Y(n_118)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_55),
.Y(n_67)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_67),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_61),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_68),
.B(n_77),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_60),
.Y(n_69)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_69),
.Y(n_114)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_65),
.Y(n_70)
);

INVx1_ASAP7_75t_SL g130 ( 
.A(n_70),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_60),
.Y(n_72)
);

INVx2_ASAP7_75t_SL g119 ( 
.A(n_72),
.Y(n_119)
);

BUFx2_ASAP7_75t_L g73 ( 
.A(n_65),
.Y(n_73)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_73),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_50),
.A2(n_27),
.B1(n_23),
.B2(n_22),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_74),
.A2(n_99),
.B1(n_26),
.B2(n_17),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_64),
.A2(n_44),
.B1(n_37),
.B2(n_42),
.Y(n_75)
);

AO22x1_ASAP7_75t_L g76 ( 
.A1(n_46),
.A2(n_35),
.B1(n_43),
.B2(n_36),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_76),
.A2(n_40),
.B(n_38),
.Y(n_113)
);

OR2x2_ASAP7_75t_L g77 ( 
.A(n_64),
.B(n_27),
.Y(n_77)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_65),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_78),
.B(n_83),
.Y(n_121)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_55),
.Y(n_79)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_79),
.Y(n_104)
);

OAI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_81),
.A2(n_93),
.B1(n_96),
.B2(n_63),
.Y(n_115)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_55),
.Y(n_82)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_82),
.Y(n_111)
);

BUFx12f_ASAP7_75t_L g84 ( 
.A(n_51),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_84),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_48),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_85),
.B(n_97),
.Y(n_125)
);

BUFx2_ASAP7_75t_L g86 ( 
.A(n_48),
.Y(n_86)
);

INVxp33_ASAP7_75t_L g102 ( 
.A(n_86),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_47),
.A2(n_28),
.B1(n_34),
.B2(n_23),
.Y(n_88)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_88),
.Y(n_122)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_51),
.Y(n_89)
);

HB1xp67_ASAP7_75t_L g123 ( 
.A(n_89),
.Y(n_123)
);

OAI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_51),
.A2(n_35),
.B1(n_16),
.B2(n_22),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g116 ( 
.A1(n_92),
.A2(n_63),
.B1(n_29),
.B2(n_33),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_62),
.A2(n_35),
.B1(n_16),
.B2(n_34),
.Y(n_93)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_50),
.Y(n_94)
);

INVx2_ASAP7_75t_SL g105 ( 
.A(n_94),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_53),
.B(n_28),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_95),
.A2(n_83),
.B(n_77),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_53),
.A2(n_26),
.B1(n_17),
.B2(n_32),
.Y(n_96)
);

HB1xp67_ASAP7_75t_L g97 ( 
.A(n_50),
.Y(n_97)
);

INVx11_ASAP7_75t_L g98 ( 
.A(n_46),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_98),
.B(n_100),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_63),
.A2(n_26),
.B1(n_17),
.B2(n_13),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_52),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_91),
.B(n_59),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_106),
.B(n_110),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_91),
.B(n_58),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_107),
.B(n_112),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_109),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_95),
.B(n_57),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_113),
.A2(n_90),
.B(n_87),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_115),
.A2(n_118),
.B1(n_129),
.B2(n_80),
.Y(n_139)
);

OAI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_116),
.A2(n_98),
.B1(n_101),
.B2(n_70),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_95),
.B(n_36),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_117),
.B(n_124),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_76),
.B(n_40),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_83),
.B(n_38),
.C(n_32),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_126),
.B(n_84),
.C(n_72),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_76),
.B(n_33),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_128),
.B(n_88),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_68),
.A2(n_32),
.B1(n_30),
.B2(n_33),
.Y(n_129)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_103),
.Y(n_133)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_133),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_102),
.B(n_71),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_134),
.B(n_138),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_135),
.B(n_126),
.Y(n_168)
);

AND2x2_ASAP7_75t_L g191 ( 
.A(n_136),
.B(n_0),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_137),
.A2(n_149),
.B1(n_151),
.B2(n_156),
.Y(n_163)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_125),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_139),
.A2(n_121),
.B1(n_116),
.B2(n_129),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_123),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_140),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_107),
.B(n_100),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_141),
.B(n_157),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_122),
.A2(n_71),
.B(n_80),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_144),
.A2(n_152),
.B(n_131),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_125),
.B(n_82),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_145),
.B(n_19),
.Y(n_188)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_123),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_146),
.B(n_147),
.Y(n_183)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_127),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_127),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_148),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_124),
.A2(n_90),
.B1(n_87),
.B2(n_101),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_150),
.A2(n_161),
.B(n_0),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_122),
.A2(n_89),
.B1(n_94),
.B2(n_67),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_128),
.A2(n_29),
.B(n_86),
.Y(n_152)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_103),
.Y(n_154)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_154),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_108),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_155),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_113),
.A2(n_78),
.B1(n_79),
.B2(n_69),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_105),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_112),
.B(n_19),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_SL g185 ( 
.A(n_158),
.B(n_29),
.Y(n_185)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_105),
.Y(n_159)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_159),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_106),
.A2(n_73),
.B1(n_32),
.B2(n_30),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_160),
.A2(n_119),
.B1(n_114),
.B2(n_130),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_114),
.A2(n_15),
.B1(n_14),
.B2(n_13),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_120),
.B(n_84),
.Y(n_162)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_162),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_143),
.B(n_117),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_SL g208 ( 
.A(n_165),
.B(n_182),
.Y(n_208)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_155),
.Y(n_167)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_167),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_168),
.B(n_181),
.C(n_189),
.Y(n_212)
);

OAI32xp33_ASAP7_75t_L g169 ( 
.A1(n_132),
.A2(n_110),
.A3(n_121),
.B1(n_120),
.B2(n_118),
.Y(n_169)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_169),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_171),
.A2(n_172),
.B1(n_177),
.B2(n_179),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_139),
.A2(n_114),
.B1(n_119),
.B2(n_131),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_174),
.A2(n_180),
.B(n_190),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_L g215 ( 
.A1(n_176),
.A2(n_140),
.B1(n_157),
.B2(n_172),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_142),
.A2(n_119),
.B1(n_130),
.B2(n_105),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_150),
.A2(n_119),
.B1(n_130),
.B2(n_111),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_143),
.B(n_111),
.C(n_104),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_158),
.B(n_104),
.Y(n_182)
);

OA21x2_ASAP7_75t_L g184 ( 
.A1(n_144),
.A2(n_162),
.B(n_147),
.Y(n_184)
);

OA21x2_ASAP7_75t_L g205 ( 
.A1(n_184),
.A2(n_146),
.B(n_159),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_SL g224 ( 
.A(n_185),
.B(n_4),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_156),
.A2(n_108),
.B1(n_84),
.B2(n_19),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_187),
.A2(n_194),
.B1(n_152),
.B2(n_132),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_188),
.B(n_192),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_141),
.B(n_15),
.C(n_13),
.Y(n_189)
);

XNOR2x1_ASAP7_75t_SL g190 ( 
.A(n_153),
.B(n_12),
.Y(n_190)
);

INVx1_ASAP7_75t_SL g216 ( 
.A(n_191),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_138),
.B(n_12),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_149),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_151),
.Y(n_195)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_195),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_166),
.B(n_170),
.Y(n_197)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_197),
.Y(n_231)
);

OAI22x1_ASAP7_75t_L g198 ( 
.A1(n_180),
.A2(n_152),
.B1(n_136),
.B2(n_148),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_198),
.A2(n_215),
.B1(n_218),
.B2(n_223),
.Y(n_229)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_183),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_200),
.B(n_206),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_165),
.B(n_135),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_201),
.B(n_220),
.Y(n_236)
);

CKINVDCx14_ASAP7_75t_R g242 ( 
.A(n_203),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_SL g234 ( 
.A1(n_205),
.A2(n_213),
.B(n_221),
.Y(n_234)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_186),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_164),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_209),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_167),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_211),
.B(n_175),
.Y(n_243)
);

AND2x4_ASAP7_75t_SL g213 ( 
.A(n_174),
.B(n_160),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_179),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_214),
.B(n_219),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_166),
.B(n_153),
.Y(n_217)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_217),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_171),
.A2(n_154),
.B1(n_133),
.B2(n_3),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_176),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_168),
.B(n_1),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_184),
.A2(n_1),
.B(n_2),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_177),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_222),
.B(n_226),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_193),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_SL g232 ( 
.A(n_224),
.B(n_189),
.Y(n_232)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_184),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_203),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_227),
.B(n_238),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_201),
.B(n_181),
.C(n_182),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_228),
.B(n_230),
.C(n_212),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_212),
.B(n_185),
.C(n_178),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_SL g261 ( 
.A(n_232),
.B(n_241),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_217),
.B(n_190),
.Y(n_237)
);

CKINVDCx14_ASAP7_75t_R g271 ( 
.A(n_237),
.Y(n_271)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_197),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_210),
.A2(n_163),
.B1(n_196),
.B2(n_169),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_240),
.A2(n_248),
.B1(n_202),
.B2(n_213),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_SL g241 ( 
.A(n_208),
.B(n_191),
.Y(n_241)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_243),
.Y(n_257)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_218),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_244),
.B(n_246),
.Y(n_269)
);

BUFx2_ASAP7_75t_L g245 ( 
.A(n_207),
.Y(n_245)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_245),
.Y(n_258)
);

INVx1_ASAP7_75t_SL g246 ( 
.A(n_205),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_210),
.A2(n_163),
.B1(n_196),
.B2(n_191),
.Y(n_248)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_205),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_250),
.B(n_221),
.Y(n_262)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_245),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_251),
.B(n_254),
.Y(n_273)
);

XNOR2x1_ASAP7_75t_L g252 ( 
.A(n_241),
.B(n_198),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_252),
.A2(n_255),
.B1(n_216),
.B2(n_204),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_228),
.B(n_208),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_253),
.B(n_232),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_235),
.B(n_225),
.Y(n_254)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_235),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_256),
.B(n_267),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_259),
.B(n_236),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_230),
.B(n_236),
.C(n_220),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_260),
.B(n_224),
.C(n_204),
.Y(n_287)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_262),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_227),
.A2(n_242),
.B1(n_240),
.B2(n_246),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_264),
.A2(n_255),
.B1(n_229),
.B2(n_250),
.Y(n_275)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_239),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_265),
.B(n_266),
.Y(n_279)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_239),
.Y(n_266)
);

HB1xp67_ASAP7_75t_L g267 ( 
.A(n_247),
.Y(n_267)
);

BUFx5_ASAP7_75t_L g268 ( 
.A(n_248),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_268),
.B(n_270),
.Y(n_285)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_249),
.Y(n_270)
);

A2O1A1Ixp33_ASAP7_75t_L g272 ( 
.A1(n_263),
.A2(n_233),
.B(n_234),
.C(n_249),
.Y(n_272)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_272),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_275),
.A2(n_276),
.B1(n_283),
.B2(n_288),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_264),
.A2(n_244),
.B1(n_213),
.B2(n_238),
.Y(n_276)
);

AND2x2_ASAP7_75t_L g277 ( 
.A(n_263),
.B(n_237),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_SL g298 ( 
.A1(n_277),
.A2(n_256),
.B(n_187),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_269),
.A2(n_247),
.B1(n_202),
.B2(n_231),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_278),
.A2(n_252),
.B1(n_269),
.B2(n_251),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_271),
.A2(n_233),
.B1(n_199),
.B2(n_231),
.Y(n_281)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_281),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_282),
.B(n_260),
.C(n_253),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_268),
.A2(n_234),
.B1(n_207),
.B2(n_216),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_257),
.B(n_223),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_284),
.B(n_5),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_286),
.B(n_287),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_289),
.B(n_298),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_282),
.B(n_259),
.C(n_266),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_290),
.B(n_299),
.Y(n_304)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_291),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_283),
.B(n_261),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_296),
.B(n_297),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_279),
.B(n_261),
.Y(n_297)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_274),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_277),
.A2(n_258),
.B1(n_173),
.B2(n_194),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_300),
.B(n_302),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_SL g301 ( 
.A1(n_273),
.A2(n_280),
.B(n_285),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_SL g307 ( 
.A1(n_301),
.A2(n_288),
.B(n_287),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_275),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_303),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_294),
.A2(n_278),
.B1(n_272),
.B2(n_276),
.Y(n_305)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_305),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_307),
.B(n_310),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_290),
.B(n_286),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_309),
.B(n_314),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_293),
.A2(n_7),
.B(n_8),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_292),
.B(n_8),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_313),
.B(n_298),
.C(n_291),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_306),
.A2(n_295),
.B1(n_294),
.B2(n_303),
.Y(n_316)
);

OR2x2_ASAP7_75t_L g325 ( 
.A(n_316),
.B(n_318),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_SL g318 ( 
.A(n_312),
.B(n_296),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_SL g319 ( 
.A(n_304),
.B(n_297),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_319),
.B(n_321),
.Y(n_327)
);

AND2x2_ASAP7_75t_L g323 ( 
.A(n_320),
.B(n_311),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_312),
.B(n_313),
.C(n_289),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_323),
.A2(n_324),
.B(n_326),
.Y(n_328)
);

A2O1A1Ixp33_ASAP7_75t_SL g324 ( 
.A1(n_315),
.A2(n_308),
.B(n_300),
.C(n_305),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_L g326 ( 
.A1(n_321),
.A2(n_311),
.B(n_292),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_L g329 ( 
.A1(n_327),
.A2(n_322),
.B(n_325),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_SL g330 ( 
.A1(n_329),
.A2(n_317),
.B(n_318),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_330),
.B(n_328),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_331),
.B(n_9),
.C(n_10),
.Y(n_332)
);

OAI211xp5_ASAP7_75t_L g333 ( 
.A1(n_332),
.A2(n_11),
.B(n_9),
.C(n_10),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_333),
.B(n_10),
.Y(n_334)
);

AOI21xp5_ASAP7_75t_L g335 ( 
.A1(n_334),
.A2(n_11),
.B(n_235),
.Y(n_335)
);


endmodule