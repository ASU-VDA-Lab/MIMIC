module real_jpeg_29911_n_18 (n_17, n_8, n_0, n_2, n_10, n_9, n_330, n_12, n_6, n_11, n_14, n_7, n_329, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_330;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_329;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

OAI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_0),
.A2(n_29),
.B1(n_34),
.B2(n_35),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_0),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_0),
.A2(n_35),
.B1(n_45),
.B2(n_46),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_0),
.A2(n_35),
.B1(n_63),
.B2(n_64),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_0),
.A2(n_35),
.B1(n_57),
.B2(n_58),
.Y(n_297)
);

HB1xp67_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

INVx5_ASAP7_75t_L g221 ( 
.A(n_1),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_2),
.A2(n_63),
.B1(n_64),
.B2(n_77),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_2),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_2),
.A2(n_57),
.B1(n_58),
.B2(n_77),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_2),
.A2(n_45),
.B1(n_46),
.B2(n_77),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_2),
.A2(n_29),
.B1(n_34),
.B2(n_77),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_3),
.Y(n_90)
);

AOI21xp33_ASAP7_75t_SL g91 ( 
.A1(n_3),
.A2(n_60),
.B(n_64),
.Y(n_91)
);

OAI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_3),
.A2(n_57),
.B1(n_58),
.B2(n_90),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_3),
.B(n_62),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_3),
.A2(n_46),
.B(n_190),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_3),
.B(n_46),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_3),
.B(n_79),
.Y(n_199)
);

OAI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_3),
.A2(n_27),
.B1(n_217),
.B2(n_221),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_3),
.A2(n_63),
.B(n_233),
.Y(n_232)
);

BUFx12_ASAP7_75t_L g60 ( 
.A(n_4),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_5),
.A2(n_57),
.B1(n_58),
.B2(n_85),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_5),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g166 ( 
.A1(n_5),
.A2(n_63),
.B1(n_64),
.B2(n_85),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_5),
.A2(n_45),
.B1(n_46),
.B2(n_85),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_5),
.A2(n_29),
.B1(n_34),
.B2(n_85),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_6),
.A2(n_45),
.B1(n_46),
.B2(n_52),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_6),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_6),
.A2(n_29),
.B1(n_34),
.B2(n_52),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_6),
.A2(n_52),
.B1(n_63),
.B2(n_64),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g282 ( 
.A1(n_6),
.A2(n_52),
.B1(n_57),
.B2(n_58),
.Y(n_282)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_8),
.A2(n_29),
.B1(n_34),
.B2(n_101),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_8),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_8),
.A2(n_45),
.B1(n_46),
.B2(n_101),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g300 ( 
.A1(n_8),
.A2(n_63),
.B1(n_64),
.B2(n_101),
.Y(n_300)
);

BUFx10_ASAP7_75t_L g57 ( 
.A(n_9),
.Y(n_57)
);

OAI22xp33_ASAP7_75t_L g43 ( 
.A1(n_10),
.A2(n_44),
.B1(n_45),
.B2(n_46),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_10),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_10),
.A2(n_44),
.B1(n_63),
.B2(n_64),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_10),
.A2(n_44),
.B1(n_57),
.B2(n_58),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_10),
.A2(n_29),
.B1(n_34),
.B2(n_44),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_11),
.A2(n_29),
.B1(n_34),
.B2(n_49),
.Y(n_48)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_11),
.Y(n_49)
);

OAI22xp33_ASAP7_75t_L g50 ( 
.A1(n_11),
.A2(n_45),
.B1(n_46),
.B2(n_49),
.Y(n_50)
);

OAI32xp33_ASAP7_75t_L g193 ( 
.A1(n_11),
.A2(n_34),
.A3(n_46),
.B1(n_194),
.B2(n_195),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_12),
.A2(n_57),
.B1(n_58),
.B2(n_68),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_12),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_12),
.A2(n_63),
.B1(n_64),
.B2(n_68),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g204 ( 
.A1(n_12),
.A2(n_29),
.B1(n_34),
.B2(n_68),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_12),
.A2(n_45),
.B1(n_46),
.B2(n_68),
.Y(n_237)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_13),
.Y(n_65)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_14),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_14),
.B(n_63),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_14),
.A2(n_45),
.B1(n_46),
.B2(n_73),
.Y(n_75)
);

INVx4_ASAP7_75t_L g243 ( 
.A(n_14),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_L g39 ( 
.A1(n_15),
.A2(n_29),
.B1(n_34),
.B2(n_40),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_15),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_15),
.A2(n_40),
.B1(n_45),
.B2(n_46),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_15),
.A2(n_40),
.B1(n_63),
.B2(n_64),
.Y(n_286)
);

AOI22xp33_ASAP7_75t_SL g321 ( 
.A1(n_15),
.A2(n_40),
.B1(n_57),
.B2(n_58),
.Y(n_321)
);

INVx11_ASAP7_75t_SL g30 ( 
.A(n_16),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_17),
.A2(n_56),
.B1(n_57),
.B2(n_58),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_17),
.Y(n_56)
);

OAI22xp33_ASAP7_75t_L g154 ( 
.A1(n_17),
.A2(n_56),
.B1(n_63),
.B2(n_64),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_17),
.A2(n_45),
.B1(n_46),
.B2(n_56),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_17),
.A2(n_29),
.B1(n_34),
.B2(n_56),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_309),
.Y(n_18)
);

OAI321xp33_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_277),
.A3(n_304),
.B1(n_307),
.B2(n_308),
.C(n_329),
.Y(n_19)
);

AOI321xp33_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_123),
.A3(n_146),
.B1(n_271),
.B2(n_276),
.C(n_330),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

OAI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_22),
.A2(n_272),
.B(n_275),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_104),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_23),
.B(n_104),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_80),
.C(n_98),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_24),
.B(n_98),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_SL g24 ( 
.A(n_25),
.B(n_53),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_25),
.B(n_54),
.C(n_69),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_41),
.Y(n_25)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_26),
.B(n_41),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_32),
.B1(n_36),
.B2(n_39),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_27),
.A2(n_38),
.B1(n_39),
.B2(n_100),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_27),
.A2(n_36),
.B(n_100),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_27),
.A2(n_204),
.B1(n_205),
.B2(n_206),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_27),
.A2(n_38),
.B1(n_211),
.B2(n_217),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_27),
.A2(n_205),
.B1(n_206),
.B2(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_28),
.A2(n_33),
.B1(n_93),
.B2(n_94),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_28),
.A2(n_37),
.B1(n_93),
.B2(n_168),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_28),
.A2(n_37),
.B1(n_210),
.B2(n_212),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_31),
.Y(n_28)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_29),
.B(n_49),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_29),
.B(n_223),
.Y(n_222)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_33),
.Y(n_32)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_36),
.Y(n_94)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx5_ASAP7_75t_SL g206 ( 
.A(n_37),
.Y(n_206)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_47),
.B1(n_48),
.B2(n_51),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_43),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_43),
.A2(n_110),
.B1(n_113),
.B2(n_157),
.Y(n_156)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_45),
.Y(n_46)
);

OAI32xp33_ASAP7_75t_L g241 ( 
.A1(n_45),
.A2(n_63),
.A3(n_234),
.B1(n_242),
.B2(n_244),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_46),
.B(n_245),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_47),
.A2(n_48),
.B1(n_51),
.B2(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_47),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_47),
.A2(n_48),
.B1(n_112),
.B2(n_133),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_47),
.A2(n_48),
.B1(n_189),
.B2(n_191),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_47),
.A2(n_48),
.B1(n_191),
.B2(n_202),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_47),
.A2(n_48),
.B1(n_158),
.B2(n_261),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_47),
.A2(n_48),
.B(n_133),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_48),
.B(n_50),
.Y(n_47)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_48),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_48),
.B(n_90),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_69),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_59),
.B1(n_62),
.B2(n_67),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_55),
.Y(n_87)
);

INVx13_ASAP7_75t_L g58 ( 
.A(n_57),
.Y(n_58)
);

A2O1A1Ixp33_ASAP7_75t_L g89 ( 
.A1(n_57),
.A2(n_66),
.B(n_90),
.C(n_91),
.Y(n_89)
);

O2A1O1Ixp33_ASAP7_75t_L g59 ( 
.A1(n_58),
.A2(n_60),
.B(n_61),
.C(n_62),
.Y(n_59)
);

NAND2xp33_ASAP7_75t_SL g61 ( 
.A(n_58),
.B(n_60),
.Y(n_61)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_59),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_59),
.A2(n_62),
.B1(n_67),
.B2(n_118),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_59),
.A2(n_62),
.B1(n_84),
.B2(n_160),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_59),
.A2(n_62),
.B1(n_296),
.B2(n_297),
.Y(n_295)
);

AO22x1_ASAP7_75t_L g62 ( 
.A1(n_60),
.A2(n_63),
.B1(n_64),
.B2(n_66),
.Y(n_62)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_60),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_62),
.Y(n_86)
);

A2O1A1Ixp33_ASAP7_75t_L g71 ( 
.A1(n_63),
.A2(n_72),
.B(n_74),
.C(n_75),
.Y(n_71)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_64),
.B(n_90),
.Y(n_234)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_70),
.A2(n_76),
.B1(n_78),
.B2(n_79),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_70),
.A2(n_78),
.B1(n_79),
.B2(n_120),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_70),
.A2(n_79),
.B1(n_154),
.B2(n_165),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_70),
.A2(n_79),
.B1(n_285),
.B2(n_286),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_70),
.A2(n_79),
.B1(n_286),
.B2(n_300),
.Y(n_299)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_71),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_71),
.A2(n_75),
.B1(n_96),
.B2(n_97),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_71),
.A2(n_75),
.B1(n_130),
.B2(n_131),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_71),
.A2(n_75),
.B1(n_96),
.B2(n_153),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_71),
.A2(n_75),
.B1(n_166),
.B2(n_232),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g316 ( 
.A1(n_71),
.A2(n_75),
.B(n_317),
.Y(n_316)
);

INVx1_ASAP7_75t_SL g72 ( 
.A(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_75),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_76),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_80),
.B(n_180),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_88),
.C(n_95),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_81),
.B(n_95),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_82),
.A2(n_83),
.B1(n_86),
.B2(n_87),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_82),
.A2(n_86),
.B1(n_139),
.B2(n_140),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_82),
.A2(n_86),
.B1(n_140),
.B2(n_282),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_82),
.A2(n_86),
.B1(n_320),
.B2(n_321),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_84),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_SL g174 ( 
.A(n_88),
.B(n_175),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_92),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_89),
.B(n_92),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_90),
.B(n_221),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_102),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_99),
.B(n_102),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_103),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_122),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_116),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_106),
.B(n_116),
.C(n_122),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_107),
.A2(n_108),
.B1(n_114),
.B2(n_115),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_107),
.B(n_115),
.Y(n_142)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_109),
.A2(n_110),
.B1(n_111),
.B2(n_113),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_110),
.A2(n_113),
.B1(n_236),
.B2(n_237),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_112),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_114),
.A2(n_115),
.B1(n_137),
.B2(n_138),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g291 ( 
.A1(n_114),
.A2(n_138),
.B(n_141),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_115),
.Y(n_114)
);

BUFx24_ASAP7_75t_SL g327 ( 
.A(n_116),
.Y(n_327)
);

FAx1_ASAP7_75t_SL g116 ( 
.A(n_117),
.B(n_119),
.CI(n_121),
.CON(n_116),
.SN(n_116)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_117),
.B(n_119),
.C(n_121),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_118),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_120),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_125),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_124),
.B(n_125),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_126),
.A2(n_127),
.B1(n_144),
.B2(n_145),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_135),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_128),
.B(n_135),
.C(n_145),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_132),
.B(n_134),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_129),
.B(n_132),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_131),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_134),
.B(n_279),
.C(n_291),
.Y(n_278)
);

FAx1_ASAP7_75t_SL g306 ( 
.A(n_134),
.B(n_279),
.CI(n_291),
.CON(n_306),
.SN(n_306)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_141),
.B1(n_142),
.B2(n_143),
.Y(n_135)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_136),
.Y(n_143)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_144),
.Y(n_145)
);

NOR3xp33_ASAP7_75t_SL g146 ( 
.A(n_147),
.B(n_176),
.C(n_181),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_170),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g273 ( 
.A(n_148),
.B(n_170),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_161),
.C(n_162),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_149),
.B(n_268),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_159),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_152),
.B1(n_155),
.B2(n_156),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_151),
.B(n_156),
.C(n_159),
.Y(n_173)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_158),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_161),
.A2(n_162),
.B1(n_163),
.B2(n_269),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_161),
.Y(n_269)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_167),
.C(n_169),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_164),
.B(n_256),
.Y(n_255)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_167),
.B(n_169),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_168),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_174),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_173),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_172),
.B(n_173),
.C(n_174),
.Y(n_178)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

AOI21xp33_ASAP7_75t_L g272 ( 
.A1(n_177),
.A2(n_273),
.B(n_274),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_179),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_178),
.B(n_179),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_182),
.A2(n_265),
.B(n_270),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_183),
.A2(n_251),
.B(n_264),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_227),
.B(n_250),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_185),
.A2(n_207),
.B(n_226),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_196),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_186),
.B(n_196),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_187),
.B(n_192),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_187),
.A2(n_188),
.B1(n_192),
.B2(n_193),
.Y(n_213)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_190),
.Y(n_194)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_203),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_198),
.A2(n_199),
.B1(n_200),
.B2(n_201),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_198),
.B(n_201),
.C(n_203),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_199),
.Y(n_198)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_202),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_204),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_208),
.A2(n_214),
.B(n_225),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_213),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_209),
.B(n_213),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_211),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_215),
.A2(n_219),
.B(n_224),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_218),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_216),
.B(n_218),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_220),
.B(n_222),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_229),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_228),
.B(n_229),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_230),
.A2(n_240),
.B1(n_248),
.B2(n_249),
.Y(n_229)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_230),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_231),
.A2(n_235),
.B1(n_238),
.B2(n_239),
.Y(n_230)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_231),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_235),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_235),
.B(n_239),
.C(n_249),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_237),
.Y(n_261)
);

CKINVDCx16_ASAP7_75t_R g249 ( 
.A(n_240),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_246),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_241),
.B(n_246),
.Y(n_259)
);

INVx6_ASAP7_75t_L g245 ( 
.A(n_242),
.Y(n_245)
);

INVx8_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_253),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_252),
.B(n_253),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_254),
.A2(n_255),
.B1(n_257),
.B2(n_258),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_254),
.B(n_260),
.C(n_262),
.Y(n_266)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_259),
.A2(n_260),
.B1(n_262),
.B2(n_263),
.Y(n_258)
);

CKINVDCx16_ASAP7_75t_R g262 ( 
.A(n_259),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_260),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_267),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_266),
.B(n_267),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_292),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_278),
.B(n_292),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_280),
.A2(n_281),
.B1(n_283),
.B2(n_290),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_280),
.A2(n_281),
.B1(n_294),
.B2(n_302),
.Y(n_293)
);

CKINVDCx14_ASAP7_75t_R g280 ( 
.A(n_281),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_281),
.B(n_284),
.C(n_289),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_281),
.B(n_302),
.C(n_303),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_282),
.Y(n_296)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_283),
.Y(n_290)
);

AOI22xp33_ASAP7_75t_L g283 ( 
.A1(n_284),
.A2(n_287),
.B1(n_288),
.B2(n_289),
.Y(n_283)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_284),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_287),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_287),
.A2(n_289),
.B1(n_299),
.B2(n_301),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_287),
.B(n_295),
.C(n_299),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_303),
.Y(n_292)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_294),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_SL g294 ( 
.A(n_295),
.B(n_298),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_297),
.Y(n_320)
);

CKINVDCx16_ASAP7_75t_R g301 ( 
.A(n_299),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g317 ( 
.A(n_300),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_306),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_305),
.B(n_306),
.Y(n_307)
);

BUFx24_ASAP7_75t_SL g326 ( 
.A(n_306),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_324),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_311),
.B(n_312),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_311),
.B(n_312),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_313),
.A2(n_314),
.B1(n_322),
.B2(n_323),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_315),
.A2(n_316),
.B1(n_318),
.B2(n_319),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_316),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_319),
.Y(n_318)
);

CKINVDCx16_ASAP7_75t_R g322 ( 
.A(n_323),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);


endmodule