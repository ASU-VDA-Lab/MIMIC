module fake_jpeg_16859_n_290 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_290);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_290;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx11_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_3),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx16f_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx2_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_6),
.Y(n_29)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_27),
.Y(n_30)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_31),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_22),
.B(n_13),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_32),
.B(n_36),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx3_ASAP7_75t_SL g55 ( 
.A(n_33),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_20),
.B(n_0),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_20),
.B(n_0),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_26),
.Y(n_50)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_31),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_41),
.B(n_49),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g43 ( 
.A1(n_35),
.A2(n_14),
.B1(n_29),
.B2(n_27),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_43),
.A2(n_35),
.B1(n_14),
.B2(n_26),
.Y(n_63)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_31),
.Y(n_49)
);

CKINVDCx14_ASAP7_75t_R g76 ( 
.A(n_50),
.Y(n_76)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_31),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_51),
.A2(n_30),
.B1(n_35),
.B2(n_14),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_33),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_53),
.B(n_40),
.Y(n_69)
);

BUFx4f_ASAP7_75t_SL g56 ( 
.A(n_33),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_56),
.Y(n_61)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_57),
.Y(n_67)
);

AND2x4_ASAP7_75t_L g59 ( 
.A(n_50),
.B(n_27),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_59),
.B(n_0),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_60),
.A2(n_48),
.B1(n_46),
.B2(n_45),
.Y(n_106)
);

INVx1_ASAP7_75t_SL g62 ( 
.A(n_58),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_62),
.B(n_65),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_63),
.A2(n_46),
.B1(n_57),
.B2(n_45),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_42),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_52),
.Y(n_66)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_66),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_44),
.A2(n_37),
.B1(n_36),
.B2(n_38),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_68),
.A2(n_76),
.B1(n_59),
.B2(n_82),
.Y(n_90)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_69),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_51),
.A2(n_15),
.B1(n_21),
.B2(n_27),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_70),
.A2(n_73),
.B(n_74),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_42),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_72),
.B(n_75),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_51),
.A2(n_15),
.B1(n_21),
.B2(n_27),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_48),
.A2(n_15),
.B1(n_21),
.B2(n_30),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_56),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_44),
.B(n_37),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_77),
.B(n_79),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_56),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_78),
.B(n_48),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_41),
.B(n_36),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_52),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_80),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g81 ( 
.A1(n_49),
.A2(n_32),
.B(n_26),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_81),
.A2(n_82),
.B(n_23),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_54),
.A2(n_20),
.B(n_1),
.Y(n_82)
);

AO22x1_ASAP7_75t_SL g83 ( 
.A1(n_55),
.A2(n_40),
.B1(n_39),
.B2(n_33),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_83),
.A2(n_58),
.B1(n_38),
.B2(n_30),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_85),
.A2(n_107),
.B(n_19),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_71),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_86),
.B(n_90),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_63),
.A2(n_55),
.B1(n_47),
.B2(n_54),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_88),
.A2(n_102),
.B1(n_106),
.B2(n_74),
.Y(n_115)
);

OAI32xp33_ASAP7_75t_L g89 ( 
.A1(n_68),
.A2(n_59),
.A3(n_77),
.B1(n_79),
.B2(n_81),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_89),
.A2(n_97),
.B1(n_109),
.B2(n_61),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_71),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_91),
.B(n_59),
.Y(n_112)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_65),
.Y(n_92)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_92),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_93),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_76),
.B(n_53),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_96),
.B(n_19),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_60),
.A2(n_55),
.B1(n_57),
.B2(n_46),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_69),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_98),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_59),
.B(n_34),
.C(n_56),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_100),
.B(n_61),
.C(n_78),
.Y(n_113)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_83),
.Y(n_101)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_101),
.Y(n_119)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_83),
.Y(n_103)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_103),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_59),
.B(n_58),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_108),
.B(n_39),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_SL g138 ( 
.A(n_112),
.B(n_129),
.C(n_132),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_113),
.B(n_134),
.C(n_87),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_92),
.B(n_72),
.Y(n_114)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_114),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_115),
.A2(n_117),
.B1(n_120),
.B2(n_107),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_87),
.B(n_75),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_116),
.B(n_105),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_101),
.A2(n_73),
.B1(n_70),
.B2(n_83),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_93),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_118),
.B(n_104),
.Y(n_150)
);

OR2x2_ASAP7_75t_L g121 ( 
.A(n_86),
.B(n_28),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_121),
.A2(n_96),
.B(n_91),
.Y(n_146)
);

AO21x1_ASAP7_75t_L g142 ( 
.A1(n_123),
.A2(n_127),
.B(n_130),
.Y(n_142)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_84),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_124),
.B(n_128),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_103),
.A2(n_64),
.B1(n_67),
.B2(n_62),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_125),
.A2(n_97),
.B1(n_104),
.B2(n_98),
.Y(n_149)
);

OA21x2_ASAP7_75t_L g127 ( 
.A1(n_95),
.A2(n_28),
.B(n_40),
.Y(n_127)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_99),
.Y(n_128)
);

MAJx2_ASAP7_75t_L g129 ( 
.A(n_89),
.B(n_28),
.C(n_34),
.Y(n_129)
);

AO22x1_ASAP7_75t_L g131 ( 
.A1(n_109),
.A2(n_62),
.B1(n_40),
.B2(n_39),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_131),
.B(n_106),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_94),
.B(n_34),
.C(n_67),
.Y(n_134)
);

INVx13_ASAP7_75t_L g135 ( 
.A(n_128),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_135),
.B(n_143),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_110),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_136),
.B(n_140),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_111),
.B(n_108),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_137),
.A2(n_145),
.B1(n_148),
.B2(n_153),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_133),
.B(n_90),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_139),
.B(n_154),
.C(n_159),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_110),
.Y(n_140)
);

AND2x6_ASAP7_75t_L g141 ( 
.A(n_129),
.B(n_85),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_141),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_113),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_111),
.B(n_100),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_146),
.B(n_121),
.Y(n_161)
);

INVx13_ASAP7_75t_L g147 ( 
.A(n_118),
.Y(n_147)
);

CKINVDCx14_ASAP7_75t_R g177 ( 
.A(n_147),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_125),
.B(n_84),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_149),
.A2(n_151),
.B1(n_152),
.B2(n_155),
.Y(n_182)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_150),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_119),
.A2(n_107),
.B1(n_95),
.B2(n_94),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_119),
.A2(n_107),
.B1(n_88),
.B2(n_64),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_122),
.B(n_105),
.Y(n_157)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_157),
.Y(n_167)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_158),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_134),
.B(n_99),
.C(n_39),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_120),
.A2(n_38),
.B1(n_29),
.B2(n_23),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_160),
.A2(n_24),
.B1(n_25),
.B2(n_23),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_161),
.A2(n_152),
.B(n_142),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_157),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_165),
.B(n_166),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_156),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_144),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_168),
.B(n_175),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_154),
.B(n_123),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_170),
.B(n_185),
.C(n_155),
.Y(n_189)
);

XNOR2x1_ASAP7_75t_SL g173 ( 
.A(n_138),
.B(n_124),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_173),
.A2(n_145),
.B1(n_143),
.B2(n_147),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_146),
.B(n_122),
.Y(n_174)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_174),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_148),
.Y(n_175)
);

AND2x2_ASAP7_75t_SL g178 ( 
.A(n_151),
.B(n_132),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_178),
.A2(n_183),
.B(n_171),
.Y(n_191)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_149),
.Y(n_179)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_179),
.Y(n_201)
);

CKINVDCx14_ASAP7_75t_R g205 ( 
.A(n_180),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_148),
.A2(n_126),
.B1(n_117),
.B2(n_127),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_181),
.A2(n_131),
.B1(n_28),
.B2(n_18),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_137),
.B(n_126),
.Y(n_183)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_183),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_137),
.B(n_130),
.Y(n_184)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_184),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_139),
.B(n_115),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_172),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_186),
.B(n_194),
.Y(n_215)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_187),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_176),
.B(n_159),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_188),
.B(n_189),
.C(n_200),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_165),
.B(n_142),
.Y(n_190)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_190),
.Y(n_219)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_191),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_193),
.B(n_171),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_168),
.B(n_135),
.Y(n_194)
);

O2A1O1Ixp33_ASAP7_75t_L g195 ( 
.A1(n_175),
.A2(n_127),
.B(n_138),
.C(n_141),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_195),
.B(n_204),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_161),
.A2(n_174),
.B(n_173),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_197),
.A2(n_203),
.B1(n_181),
.B2(n_184),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_169),
.B(n_145),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_199),
.B(n_206),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_176),
.B(n_131),
.Y(n_200)
);

INVx1_ASAP7_75t_SL g204 ( 
.A(n_178),
.Y(n_204)
);

HB1xp67_ASAP7_75t_L g206 ( 
.A(n_179),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_209),
.B(n_220),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_211),
.A2(n_212),
.B1(n_218),
.B2(n_9),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_204),
.A2(n_163),
.B1(n_169),
.B2(n_164),
.Y(n_212)
);

INVx1_ASAP7_75t_SL g213 ( 
.A(n_198),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_213),
.B(n_217),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_201),
.A2(n_178),
.B1(n_182),
.B2(n_192),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_214),
.A2(n_223),
.B1(n_19),
.B2(n_18),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_188),
.B(n_162),
.C(n_170),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_216),
.B(n_200),
.C(n_193),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_196),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_191),
.A2(n_163),
.B1(n_164),
.B2(n_166),
.Y(n_218)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_202),
.B(n_185),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_220),
.A2(n_197),
.B(n_187),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_192),
.B(n_167),
.Y(n_222)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_222),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_202),
.A2(n_207),
.B1(n_190),
.B2(n_189),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_226),
.B(n_235),
.C(n_237),
.Y(n_251)
);

A2O1A1Ixp33_ASAP7_75t_SL g227 ( 
.A1(n_225),
.A2(n_207),
.B(n_167),
.C(n_195),
.Y(n_227)
);

NOR3xp33_ASAP7_75t_L g252 ( 
.A(n_227),
.B(n_1),
.C(n_2),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_228),
.B(n_239),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_208),
.A2(n_205),
.B1(n_203),
.B2(n_177),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_229),
.B(n_234),
.Y(n_242)
);

OR2x2_ASAP7_75t_L g230 ( 
.A(n_219),
.B(n_180),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_230),
.B(n_240),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_213),
.A2(n_25),
.B(n_24),
.Y(n_231)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_231),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_233),
.A2(n_220),
.B1(n_222),
.B2(n_3),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_210),
.B(n_17),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_210),
.B(n_216),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_209),
.B(n_17),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_238),
.B(n_221),
.C(n_223),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_224),
.B(n_17),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_241),
.B(n_248),
.C(n_227),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_230),
.B(n_214),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_244),
.B(n_246),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_236),
.B(n_215),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_235),
.B(n_221),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_249),
.B(n_2),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_232),
.B(n_238),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_250),
.B(n_10),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_252),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_253)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_253),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_243),
.A2(n_245),
.B(n_239),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_254),
.B(n_258),
.Y(n_266)
);

AND2x2_ASAP7_75t_L g255 ( 
.A(n_243),
.B(n_226),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_255),
.B(n_262),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_242),
.A2(n_227),
.B1(n_10),
.B2(n_6),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_256),
.B(n_263),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_259),
.B(n_7),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_251),
.B(n_227),
.C(n_18),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_260),
.B(n_261),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_241),
.B(n_11),
.Y(n_262)
);

AND2x2_ASAP7_75t_L g263 ( 
.A(n_247),
.B(n_11),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_257),
.B(n_252),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_267),
.B(n_270),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_269),
.B(n_260),
.C(n_20),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_262),
.B(n_7),
.Y(n_270)
);

NOR2x1_ASAP7_75t_L g272 ( 
.A(n_263),
.B(n_8),
.Y(n_272)
);

NAND3xp33_ASAP7_75t_SL g274 ( 
.A(n_272),
.B(n_9),
.C(n_12),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_273),
.B(n_274),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_265),
.A2(n_255),
.B(n_9),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_276),
.B(n_272),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_266),
.B(n_12),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_277),
.B(n_279),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_268),
.A2(n_12),
.B1(n_13),
.B2(n_4),
.Y(n_278)
);

INVxp33_ASAP7_75t_L g280 ( 
.A(n_278),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_264),
.B(n_13),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_282),
.A2(n_284),
.B(n_283),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_275),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_SL g285 ( 
.A1(n_281),
.A2(n_279),
.B(n_265),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_285),
.B(n_286),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_280),
.B(n_271),
.C(n_4),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_288),
.B(n_287),
.C(n_4),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_SL g290 ( 
.A(n_289),
.B(n_4),
.Y(n_290)
);


endmodule