module fake_jpeg_2315_n_161 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_161);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_161;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_39),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_4),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_15),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_21),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_32),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_4),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_17),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_30),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_10),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_29),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_20),
.Y(n_55)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_8),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_9),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_11),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_15),
.Y(n_61)
);

BUFx8_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_10),
.Y(n_63)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_62),
.Y(n_64)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_64),
.Y(n_78)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_62),
.Y(n_65)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_65),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_66),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_L g67 ( 
.A1(n_53),
.A2(n_62),
.B(n_58),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_67),
.B(n_69),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_68),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_53),
.B(n_41),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_51),
.B(n_19),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_70),
.B(n_71),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_51),
.B(n_52),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_59),
.B(n_61),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_72),
.A2(n_52),
.B1(n_63),
.B2(n_46),
.Y(n_85)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_66),
.Y(n_76)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_76),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_65),
.Y(n_77)
);

BUFx2_ASAP7_75t_L g99 ( 
.A(n_77),
.Y(n_99)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_65),
.Y(n_79)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_79),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_66),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_81),
.Y(n_97)
);

BUFx2_ASAP7_75t_L g82 ( 
.A(n_64),
.Y(n_82)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_82),
.Y(n_91)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_68),
.Y(n_84)
);

BUFx5_ASAP7_75t_L g98 ( 
.A(n_84),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_85),
.B(n_67),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_68),
.A2(n_60),
.B1(n_63),
.B2(n_46),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_86),
.A2(n_60),
.B1(n_56),
.B2(n_44),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_87),
.B(n_96),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_75),
.B(n_72),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_89),
.B(n_90),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_83),
.B(n_69),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_73),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_92),
.B(n_101),
.Y(n_108)
);

O2A1O1Ixp33_ASAP7_75t_SL g93 ( 
.A1(n_86),
.A2(n_71),
.B(n_50),
.C(n_43),
.Y(n_93)
);

A2O1A1Ixp33_ASAP7_75t_L g120 ( 
.A1(n_93),
.A2(n_0),
.B(n_1),
.C(n_2),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_83),
.B(n_70),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_94),
.B(n_95),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_73),
.A2(n_81),
.B1(n_80),
.B2(n_85),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_74),
.A2(n_57),
.B1(n_45),
.B2(n_49),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_100),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_78),
.B(n_48),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_82),
.B(n_47),
.Y(n_103)
);

NAND3xp33_ASAP7_75t_L g121 ( 
.A(n_103),
.B(n_95),
.C(n_97),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_103),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_104),
.B(n_116),
.Y(n_126)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_98),
.Y(n_105)
);

INVx2_ASAP7_75t_SL g124 ( 
.A(n_105),
.Y(n_124)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_102),
.Y(n_106)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_106),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_90),
.A2(n_54),
.B(n_55),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_110),
.A2(n_12),
.B(n_13),
.Y(n_135)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_88),
.Y(n_112)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_112),
.Y(n_133)
);

INVx1_ASAP7_75t_SL g114 ( 
.A(n_99),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_114),
.B(n_117),
.Y(n_122)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_91),
.Y(n_115)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_115),
.Y(n_137)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_98),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_99),
.Y(n_117)
);

INVxp33_ASAP7_75t_L g118 ( 
.A(n_97),
.Y(n_118)
);

FAx1_ASAP7_75t_SL g119 ( 
.A(n_93),
.B(n_0),
.CI(n_1),
.CON(n_119),
.SN(n_119)
);

NOR4xp25_ASAP7_75t_L g125 ( 
.A(n_119),
.B(n_2),
.C(n_3),
.D(n_5),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_125),
.B(n_135),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_111),
.B(n_113),
.C(n_109),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_127),
.B(n_129),
.C(n_24),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_108),
.B(n_3),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_128),
.B(n_134),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_109),
.B(n_107),
.C(n_118),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_121),
.B(n_37),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_120),
.A2(n_5),
.B(n_6),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_131),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_107),
.A2(n_7),
.B(n_9),
.Y(n_132)
);

A2O1A1O1Ixp25_ASAP7_75t_L g141 ( 
.A1(n_132),
.A2(n_12),
.B(n_13),
.C(n_14),
.D(n_16),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_105),
.B(n_11),
.Y(n_134)
);

AOI21xp33_ASAP7_75t_SL g136 ( 
.A1(n_104),
.A2(n_22),
.B(n_33),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_136),
.B(n_25),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_122),
.Y(n_138)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_138),
.Y(n_147)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_123),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_139),
.B(n_146),
.Y(n_150)
);

MAJx2_ASAP7_75t_L g149 ( 
.A(n_144),
.B(n_135),
.C(n_136),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_126),
.B(n_14),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_144),
.B(n_130),
.C(n_133),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_148),
.B(n_145),
.C(n_137),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_149),
.B(n_142),
.C(n_140),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_147),
.B(n_143),
.Y(n_151)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_151),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_152),
.B(n_153),
.C(n_150),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_155),
.A2(n_152),
.B1(n_141),
.B2(n_124),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_156),
.A2(n_154),
.B1(n_26),
.B2(n_27),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_157),
.B(n_23),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_158),
.B(n_28),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_159),
.B(n_31),
.Y(n_160)
);

HB1xp67_ASAP7_75t_L g161 ( 
.A(n_160),
.Y(n_161)
);


endmodule