module real_aes_11139_n_16 (n_13, n_4, n_0, n_3, n_5, n_2, n_15, n_7, n_8, n_6, n_9, n_12, n_1, n_14, n_10, n_11, n_16);
input n_13;
input n_4;
input n_0;
input n_3;
input n_5;
input n_2;
input n_15;
input n_7;
input n_8;
input n_6;
input n_9;
input n_12;
input n_1;
input n_14;
input n_10;
input n_11;
output n_16;
wire n_28;
wire n_17;
wire n_22;
wire n_24;
wire n_34;
wire n_19;
wire n_25;
wire n_32;
wire n_30;
wire n_37;
wire n_35;
wire n_39;
wire n_27;
wire n_23;
wire n_38;
wire n_29;
wire n_20;
wire n_26;
wire n_18;
wire n_21;
wire n_31;
wire n_33;
wire n_36;
NOR2xp33_ASAP7_75t_R g26 ( .A(n_0), .B(n_5), .Y(n_26) );
NOR3xp33_ASAP7_75t_SL g24 ( .A(n_1), .B(n_8), .C(n_25), .Y(n_24) );
NAND2xp33_ASAP7_75t_R g25 ( .A(n_2), .B(n_26), .Y(n_25) );
OAI22xp33_ASAP7_75t_SL g17 ( .A1(n_3), .A2(n_15), .B1(n_18), .B2(n_20), .Y(n_17) );
CKINVDCx5p33_ASAP7_75t_R g27 ( .A(n_4), .Y(n_27) );
NOR4xp25_ASAP7_75t_SL g22 ( .A(n_6), .B(n_23), .C(n_27), .D(n_28), .Y(n_22) );
CKINVDCx5p33_ASAP7_75t_R g39 ( .A(n_6), .Y(n_39) );
NOR2xp33_ASAP7_75t_R g19 ( .A(n_7), .B(n_12), .Y(n_19) );
NAND2xp33_ASAP7_75t_R g20 ( .A(n_7), .B(n_12), .Y(n_20) );
NAND2xp33_ASAP7_75t_SL g30 ( .A(n_7), .B(n_31), .Y(n_30) );
NOR2xp33_ASAP7_75t_R g33 ( .A(n_7), .B(n_31), .Y(n_33) );
INVx1_ASAP7_75t_L g36 ( .A(n_9), .Y(n_36) );
OAI22xp33_ASAP7_75t_SL g29 ( .A1(n_10), .A2(n_13), .B1(n_30), .B2(n_32), .Y(n_29) );
OAI33xp33_ASAP7_75t_R g16 ( .A1(n_11), .A2(n_17), .A3(n_21), .B1(n_29), .B2(n_34), .B3(n_39), .Y(n_16) );
CKINVDCx5p33_ASAP7_75t_R g28 ( .A(n_11), .Y(n_28) );
CKINVDCx5p33_ASAP7_75t_R g31 ( .A(n_12), .Y(n_31) );
A2O1A1Ixp33_ASAP7_75t_R g34 ( .A1(n_14), .A2(n_33), .B(n_35), .C(n_37), .Y(n_34) );
NOR2xp33_ASAP7_75t_R g35 ( .A(n_18), .B(n_36), .Y(n_35) );
CKINVDCx5p33_ASAP7_75t_R g18 ( .A(n_19), .Y(n_18) );
CKINVDCx5p33_ASAP7_75t_R g21 ( .A(n_22), .Y(n_21) );
CKINVDCx5p33_ASAP7_75t_R g23 ( .A(n_24), .Y(n_23) );
NAND2xp33_ASAP7_75t_R g38 ( .A(n_24), .B(n_27), .Y(n_38) );
CKINVDCx5p33_ASAP7_75t_R g32 ( .A(n_33), .Y(n_32) );
CKINVDCx5p33_ASAP7_75t_R g37 ( .A(n_38), .Y(n_37) );
endmodule