module real_aes_4150_n_407 (n_76, n_113, n_187, n_90, n_257, n_390, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_357, n_386, n_64, n_254, n_207, n_10, n_83, n_181, n_362, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_355, n_239, n_100, n_54, n_112, n_319, n_364, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_376, n_308, n_172, n_341, n_232, n_6, n_401, n_69, n_317, n_353, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_379, n_374, n_26, n_235, n_399, n_378, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_388, n_395, n_332, n_292, n_400, n_116, n_94, n_289, n_280, n_333, n_213, n_356, n_184, n_28, n_372, n_202, n_56, n_370, n_34, n_98, n_384, n_121, n_352, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_369, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_383, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_381, n_311, n_324, n_25, n_278, n_236, n_367, n_267, n_218, n_48, n_204, n_339, n_398, n_89, n_277, n_331, n_93, n_182, n_363, n_323, n_199, n_350, n_142, n_223, n_67, n_405, n_368, n_250, n_85, n_406, n_45, n_5, n_244, n_118, n_139, n_402, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_391, n_360, n_58, n_165, n_361, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_387, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_351, n_126, n_200, n_115, n_96, n_110, n_392, n_150, n_147, n_288, n_404, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_366, n_346, n_193, n_397, n_293, n_162, n_358, n_385, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_377, n_273, n_114, n_276, n_295, n_382, n_265, n_354, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_373, n_60, n_233, n_290, n_365, n_155, n_243, n_268, n_136, n_157, n_282, n_389, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_359, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_371, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_375, n_340, n_13, n_380, n_394, n_168, n_175, n_241, n_105, n_84, n_294, n_393, n_258, n_206, n_307, n_396, n_342, n_348, n_14, n_403, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_407);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_390;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_357;
input n_386;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_362;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_355;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_364;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_376;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_401;
input n_69;
input n_317;
input n_353;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_379;
input n_374;
input n_26;
input n_235;
input n_399;
input n_378;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_388;
input n_395;
input n_332;
input n_292;
input n_400;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_356;
input n_184;
input n_28;
input n_372;
input n_202;
input n_56;
input n_370;
input n_34;
input n_98;
input n_384;
input n_121;
input n_352;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_369;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_383;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_381;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_367;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_398;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_363;
input n_323;
input n_199;
input n_350;
input n_142;
input n_223;
input n_67;
input n_405;
input n_368;
input n_250;
input n_85;
input n_406;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_402;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_391;
input n_360;
input n_58;
input n_165;
input n_361;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_387;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_351;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_392;
input n_150;
input n_147;
input n_288;
input n_404;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_366;
input n_346;
input n_193;
input n_397;
input n_293;
input n_162;
input n_358;
input n_385;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_377;
input n_273;
input n_114;
input n_276;
input n_295;
input n_382;
input n_265;
input n_354;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_373;
input n_60;
input n_233;
input n_290;
input n_365;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_389;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_359;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_371;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_375;
input n_340;
input n_13;
input n_380;
input n_394;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_393;
input n_258;
input n_206;
input n_307;
input n_396;
input n_342;
input n_348;
input n_14;
input n_403;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_407;
wire n_476;
wire n_599;
wire n_887;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_761;
wire n_421;
wire n_919;
wire n_1217;
wire n_571;
wire n_549;
wire n_1034;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_870;
wire n_1248;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_786;
wire n_512;
wire n_795;
wire n_1379;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_553;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1225;
wire n_1382;
wire n_875;
wire n_951;
wire n_1199;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_595;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_796;
wire n_874;
wire n_1126;
wire n_455;
wire n_682;
wire n_812;
wire n_817;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_1317;
wire n_417;
wire n_690;
wire n_499;
wire n_1142;
wire n_947;
wire n_970;
wire n_1149;
wire n_527;
wire n_1342;
wire n_552;
wire n_1346;
wire n_1383;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_805;
wire n_619;
wire n_1095;
wire n_1250;
wire n_1284;
wire n_859;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_501;
wire n_488;
wire n_1380;
wire n_954;
wire n_702;
wire n_1007;
wire n_898;
wire n_562;
wire n_1022;
wire n_1073;
wire n_728;
wire n_1301;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_1003;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_648;
wire n_939;
wire n_928;
wire n_1384;
wire n_789;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_712;
wire n_422;
wire n_861;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_829;
wire n_1030;
wire n_1348;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_652;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_480;
wire n_684;
wire n_1178;
wire n_821;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_635;
wire n_792;
wire n_1392;
wire n_665;
wire n_667;
wire n_991;
wire n_580;
wire n_1004;
wire n_1370;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_1260;
wire n_1129;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_461;
wire n_1047;
wire n_1016;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_538;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_704;
wire n_453;
wire n_647;
wire n_948;
wire n_700;
wire n_677;
wire n_1269;
wire n_591;
wire n_1366;
wire n_678;
wire n_415;
wire n_564;
wire n_638;
wire n_1361;
wire n_510;
wire n_1358;
wire n_550;
wire n_966;
wire n_1368;
wire n_994;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_535;
wire n_882;
wire n_1210;
wire n_746;
wire n_656;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_651;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_428;
wire n_783;
wire n_1107;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1386;
wire n_617;
wire n_602;
wire n_733;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_807;
wire n_1011;
wire n_416;
wire n_895;
wire n_799;
wire n_490;
wire n_695;
wire n_1181;
wire n_881;
wire n_645;
wire n_1145;
wire n_557;
wire n_777;
wire n_985;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_1347;
wire n_1163;
wire n_1278;
wire n_734;
wire n_735;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_649;
wire n_1234;
wire n_622;
wire n_1353;
wire n_1002;
wire n_1165;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_720;
wire n_1026;
wire n_492;
wire n_419;
wire n_1023;
wire n_730;
wire n_643;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_526;
wire n_1194;
wire n_701;
wire n_809;
wire n_679;
wire n_520;
wire n_926;
wire n_942;
wire n_1374;
wire n_1120;
wire n_689;
wire n_946;
wire n_753;
wire n_1188;
wire n_623;
wire n_1032;
wire n_721;
wire n_1133;
wire n_739;
wire n_1322;
wire n_1162;
wire n_762;
wire n_1298;
wire n_442;
wire n_740;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_459;
wire n_1172;
wire n_998;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_473;
wire n_967;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_1377;
wire n_800;
wire n_778;
wire n_1170;
wire n_1175;
wire n_522;
wire n_977;
wire n_943;
wire n_905;
wire n_878;
wire n_1333;
wire n_577;
wire n_759;
wire n_1235;
wire n_900;
wire n_841;
wire n_1218;
wire n_736;
wire n_766;
wire n_852;
wire n_1113;
wire n_1268;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_773;
wire n_865;
wire n_594;
wire n_856;
wire n_1146;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_519;
wire n_1116;
wire n_709;
wire n_816;
wire n_625;
wire n_953;
wire n_1373;
wire n_716;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_935;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_1168;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1263;
wire n_1115;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_1303;
wire n_443;
wire n_1029;
wire n_1207;
wire n_664;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_561;
wire n_437;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_502;
wire n_769;
wire n_434;
wire n_1212;
wire n_1054;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1134;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1060;
wire n_1154;
wire n_632;
wire n_1344;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_912;
wire n_464;
wire n_1227;
wire n_945;
wire n_563;
wire n_891;
wire n_568;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1028;
wire n_1083;
wire n_727;
wire n_1056;
wire n_663;
wire n_588;
wire n_707;
wire n_915;
wire n_1001;
wire n_711;
wire n_864;
wire n_1169;
wire n_1139;
wire n_1038;
wire n_1085;
wire n_845;
wire n_1127;
wire n_484;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_697;
wire n_978;
wire n_847;
wire n_826;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1051;
wire n_1355;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_1378;
wire n_524;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_525;
wire n_1226;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_929;
wire n_1143;
wire n_1190;
wire n_543;
wire n_585;
wire n_465;
wire n_719;
wire n_1343;
wire n_1156;
wire n_988;
wire n_921;
wire n_640;
wire n_1176;
wire n_1151;
wire n_1254;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_1096;
wire n_1316;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1240;
wire n_987;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_460;
wire n_666;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_489;
wire n_1381;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_408;
wire n_578;
wire n_892;
wire n_938;
wire n_774;
wire n_559;
wire n_466;
wire n_1049;
wire n_1277;
wire n_984;
wire n_726;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_532;
wire n_1025;
wire n_924;
wire n_1264;
wire n_1245;
wire n_1152;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1318;
wire n_1290;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_1100;
wire n_425;
wire n_879;
wire n_449;
wire n_1340;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_655;
wire n_654;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1334;
wire n_1291;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1356;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1077;
wire n_1111;
wire n_1249;
wire n_1239;
wire n_969;
wire n_1009;
wire n_1202;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_1252;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_536;
wire n_851;
wire n_470;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_1296;
wire n_1043;
wire n_435;
wire n_511;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1087;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1273;
wire n_959;
wire n_1130;
wire n_794;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1253;
wire n_1183;
wire n_516;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_1372;
wire n_698;
wire n_1345;
wire n_587;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_793;
wire n_1390;
wire n_757;
wire n_803;
wire n_514;
wire n_507;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1388;
wire n_483;
wire n_1352;
wire n_729;
wire n_1280;
wire n_1323;
wire n_703;
wire n_1097;
wire n_1369;
wire n_601;
wire n_463;
wire n_1236;
wire n_603;
wire n_1288;
wire n_868;
wire n_1024;
wire n_1144;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_429;
INVx1_ASAP7_75t_L g656 ( .A(n_0), .Y(n_656) );
AOI22xp33_ASAP7_75t_L g1171 ( .A1(n_1), .A2(n_396), .B1(n_556), .B2(n_602), .Y(n_1171) );
AOI22xp33_ASAP7_75t_L g1124 ( .A1(n_2), .A2(n_246), .B1(n_505), .B2(n_709), .Y(n_1124) );
AOI22xp33_ASAP7_75t_L g736 ( .A1(n_3), .A2(n_329), .B1(n_582), .B2(n_737), .Y(n_736) );
AOI22xp33_ASAP7_75t_L g1288 ( .A1(n_4), .A2(n_305), .B1(n_553), .B2(n_745), .Y(n_1288) );
AOI21xp33_ASAP7_75t_SL g1165 ( .A1(n_5), .A2(n_1166), .B(n_1167), .Y(n_1165) );
AOI22xp33_ASAP7_75t_L g1191 ( .A1(n_6), .A2(n_394), .B1(n_623), .B2(n_629), .Y(n_1191) );
AO22x1_ASAP7_75t_L g1201 ( .A1(n_7), .A2(n_252), .B1(n_639), .B2(n_640), .Y(n_1201) );
AOI22xp33_ASAP7_75t_L g694 ( .A1(n_8), .A2(n_298), .B1(n_654), .B2(n_695), .Y(n_694) );
INVx1_ASAP7_75t_L g1295 ( .A(n_9), .Y(n_1295) );
AOI22xp5_ASAP7_75t_L g673 ( .A1(n_10), .A2(n_335), .B1(n_555), .B2(n_556), .Y(n_673) );
AOI22xp5_ASAP7_75t_L g627 ( .A1(n_11), .A2(n_215), .B1(n_628), .B2(n_629), .Y(n_627) );
AOI22xp5_ASAP7_75t_L g1255 ( .A1(n_12), .A2(n_181), .B1(n_518), .B2(n_525), .Y(n_1255) );
AOI22xp33_ASAP7_75t_L g1333 ( .A1(n_13), .A2(n_137), .B1(n_621), .B2(n_645), .Y(n_1333) );
AOI22xp33_ASAP7_75t_L g1181 ( .A1(n_14), .A2(n_374), .B1(n_703), .B2(n_1182), .Y(n_1181) );
AOI21xp33_ASAP7_75t_SL g590 ( .A1(n_15), .A2(n_564), .B(n_591), .Y(n_590) );
AOI22xp33_ASAP7_75t_L g767 ( .A1(n_16), .A2(n_223), .B1(n_768), .B2(n_769), .Y(n_767) );
AOI22xp5_ASAP7_75t_L g1214 ( .A1(n_17), .A2(n_235), .B1(n_513), .B2(n_632), .Y(n_1214) );
NAND2xp5_ASAP7_75t_SL g445 ( .A(n_18), .B(n_434), .Y(n_445) );
AOI22xp33_ASAP7_75t_L g1376 ( .A1(n_19), .A2(n_189), .B1(n_568), .B2(n_598), .Y(n_1376) );
AOI22xp33_ASAP7_75t_L g1148 ( .A1(n_20), .A2(n_337), .B1(n_1149), .B2(n_1150), .Y(n_1148) );
AOI22xp33_ASAP7_75t_L g732 ( .A1(n_21), .A2(n_200), .B1(n_654), .B2(n_665), .Y(n_732) );
AOI22xp33_ASAP7_75t_L g1334 ( .A1(n_22), .A2(n_132), .B1(n_626), .B2(n_628), .Y(n_1334) );
AOI22xp5_ASAP7_75t_L g875 ( .A1(n_23), .A2(n_363), .B1(n_836), .B2(n_844), .Y(n_875) );
OAI22x1_ASAP7_75t_L g1054 ( .A1(n_23), .A2(n_1055), .B1(n_1080), .B2(n_1081), .Y(n_1054) );
INVx1_ASAP7_75t_L g1081 ( .A(n_23), .Y(n_1081) );
AOI22xp33_ASAP7_75t_L g1086 ( .A1(n_23), .A2(n_1087), .B1(n_1090), .B2(n_1092), .Y(n_1086) );
AOI21xp33_ASAP7_75t_L g1222 ( .A1(n_24), .A2(n_662), .B(n_1223), .Y(n_1222) );
AOI22xp5_ASAP7_75t_L g1285 ( .A1(n_25), .A2(n_390), .B1(n_518), .B2(n_1070), .Y(n_1285) );
AOI22xp33_ASAP7_75t_L g708 ( .A1(n_26), .A2(n_369), .B1(n_506), .B2(n_709), .Y(n_708) );
AOI22xp33_ASAP7_75t_L g1357 ( .A1(n_27), .A2(n_72), .B1(n_633), .B2(n_643), .Y(n_1357) );
AOI22xp5_ASAP7_75t_L g1381 ( .A1(n_28), .A2(n_323), .B1(n_555), .B2(n_556), .Y(n_1381) );
AOI221xp5_ASAP7_75t_L g1372 ( .A1(n_29), .A2(n_313), .B1(n_1312), .B2(n_1373), .C(n_1374), .Y(n_1372) );
BUFx6f_ASAP7_75t_L g434 ( .A(n_30), .Y(n_434) );
INVx1_ASAP7_75t_L g647 ( .A(n_31), .Y(n_647) );
AOI22xp5_ASAP7_75t_L g1104 ( .A1(n_32), .A2(n_75), .B1(n_1105), .B2(n_1106), .Y(n_1104) );
NAND2xp5_ASAP7_75t_L g1276 ( .A(n_33), .B(n_775), .Y(n_1276) );
AOI22xp5_ASAP7_75t_L g1229 ( .A1(n_34), .A2(n_96), .B1(n_632), .B2(n_1230), .Y(n_1229) );
AOI22xp5_ASAP7_75t_L g805 ( .A1(n_35), .A2(n_395), .B1(n_513), .B2(n_552), .Y(n_805) );
AOI22xp33_ASAP7_75t_L g1072 ( .A1(n_36), .A2(n_128), .B1(n_1073), .B2(n_1074), .Y(n_1072) );
AO22x1_ASAP7_75t_L g1139 ( .A1(n_37), .A2(n_166), .B1(n_775), .B2(n_781), .Y(n_1139) );
AOI22xp33_ASAP7_75t_L g604 ( .A1(n_38), .A2(n_41), .B1(n_558), .B2(n_605), .Y(n_604) );
INVx1_ASAP7_75t_L g1224 ( .A(n_39), .Y(n_1224) );
AOI22xp33_ASAP7_75t_L g711 ( .A1(n_40), .A2(n_159), .B1(n_519), .B2(n_712), .Y(n_711) );
AOI22xp33_ASAP7_75t_L g746 ( .A1(n_42), .A2(n_94), .B1(n_550), .B2(n_747), .Y(n_746) );
OA21x2_ASAP7_75t_L g1345 ( .A1(n_43), .A2(n_1346), .B(n_1361), .Y(n_1345) );
INVx1_ASAP7_75t_L g1364 ( .A(n_43), .Y(n_1364) );
INVx1_ASAP7_75t_L g815 ( .A(n_44), .Y(n_815) );
AOI22xp33_ASAP7_75t_L g770 ( .A1(n_45), .A2(n_229), .B1(n_771), .B2(n_772), .Y(n_770) );
AOI22xp33_ASAP7_75t_L g674 ( .A1(n_46), .A2(n_224), .B1(n_553), .B2(n_675), .Y(n_674) );
AOI22xp5_ASAP7_75t_L g1382 ( .A1(n_47), .A2(n_392), .B1(n_675), .B2(n_1383), .Y(n_1382) );
AOI21xp5_ASAP7_75t_L g1135 ( .A1(n_48), .A2(n_1136), .B(n_1139), .Y(n_1135) );
AOI22xp33_ASAP7_75t_L g1147 ( .A1(n_49), .A2(n_265), .B1(n_555), .B2(n_793), .Y(n_1147) );
AOI21xp33_ASAP7_75t_SL g1266 ( .A1(n_50), .A2(n_564), .B(n_1267), .Y(n_1266) );
AOI22x1_ASAP7_75t_L g1280 ( .A1(n_51), .A2(n_1281), .B1(n_1282), .B2(n_1296), .Y(n_1280) );
INVx1_ASAP7_75t_L g1296 ( .A(n_51), .Y(n_1296) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_52), .B(n_481), .Y(n_589) );
INVx1_ASAP7_75t_L g1353 ( .A(n_53), .Y(n_1353) );
AOI22xp33_ASAP7_75t_L g725 ( .A1(n_54), .A2(n_350), .B1(n_506), .B2(n_707), .Y(n_725) );
INVx1_ASAP7_75t_L g427 ( .A(n_55), .Y(n_427) );
AOI22xp33_ASAP7_75t_SL g1141 ( .A1(n_56), .A2(n_69), .B1(n_1059), .B2(n_1142), .Y(n_1141) );
AOI22xp33_ASAP7_75t_L g1349 ( .A1(n_57), .A2(n_195), .B1(n_623), .B2(n_1350), .Y(n_1349) );
OA22x2_ASAP7_75t_L g432 ( .A1(n_58), .A2(n_169), .B1(n_433), .B2(n_434), .Y(n_432) );
INVx1_ASAP7_75t_L g475 ( .A(n_58), .Y(n_475) );
AOI22xp5_ASAP7_75t_L g1217 ( .A1(n_59), .A2(n_118), .B1(n_529), .B2(n_714), .Y(n_1217) );
AOI22xp5_ASAP7_75t_L g727 ( .A1(n_60), .A2(n_238), .B1(n_555), .B2(n_556), .Y(n_727) );
AOI22xp33_ASAP7_75t_L g794 ( .A1(n_61), .A2(n_151), .B1(n_540), .B2(n_795), .Y(n_794) );
AOI22xp33_ASAP7_75t_L g548 ( .A1(n_62), .A2(n_406), .B1(n_549), .B2(n_550), .Y(n_548) );
AOI22xp33_ASAP7_75t_L g965 ( .A1(n_63), .A2(n_217), .B1(n_843), .B2(n_870), .Y(n_965) );
INVx1_ASAP7_75t_L g1259 ( .A(n_64), .Y(n_1259) );
AOI22xp33_ASAP7_75t_L g730 ( .A1(n_65), .A2(n_77), .B1(n_703), .B2(n_731), .Y(n_730) );
AOI22xp5_ASAP7_75t_L g1380 ( .A1(n_66), .A2(n_110), .B1(n_549), .B2(n_787), .Y(n_1380) );
AOI22xp33_ASAP7_75t_L g1144 ( .A1(n_67), .A2(n_180), .B1(n_786), .B2(n_788), .Y(n_1144) );
AOI22xp33_ASAP7_75t_L g860 ( .A1(n_68), .A2(n_194), .B1(n_828), .B2(n_849), .Y(n_860) );
AOI22xp33_ASAP7_75t_L g557 ( .A1(n_70), .A2(n_142), .B1(n_558), .B2(n_559), .Y(n_557) );
INVx1_ASAP7_75t_L g592 ( .A(n_71), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g1354 ( .A(n_73), .B(n_1355), .Y(n_1354) );
AOI22xp5_ASAP7_75t_L g638 ( .A1(n_74), .A2(n_388), .B1(n_639), .B2(n_640), .Y(n_638) );
AOI22xp33_ASAP7_75t_L g1384 ( .A1(n_76), .A2(n_201), .B1(n_541), .B2(n_558), .Y(n_1384) );
AOI22xp33_ASAP7_75t_L g757 ( .A1(n_78), .A2(n_254), .B1(n_758), .B2(n_759), .Y(n_757) );
AOI22xp5_ASAP7_75t_L g1338 ( .A1(n_79), .A2(n_247), .B1(n_633), .B2(n_643), .Y(n_1338) );
AOI22xp5_ASAP7_75t_L g1220 ( .A1(n_80), .A2(n_144), .B1(n_665), .B2(n_669), .Y(n_1220) );
INVx1_ASAP7_75t_SL g1274 ( .A(n_81), .Y(n_1274) );
INVx1_ASAP7_75t_L g1113 ( .A(n_82), .Y(n_1113) );
AOI22xp5_ASAP7_75t_L g641 ( .A1(n_83), .A2(n_404), .B1(n_642), .B2(n_643), .Y(n_641) );
AOI22xp33_ASAP7_75t_L g726 ( .A1(n_84), .A2(n_327), .B1(n_549), .B2(n_706), .Y(n_726) );
INVx1_ASAP7_75t_SL g1323 ( .A(n_85), .Y(n_1323) );
NOR2xp33_ASAP7_75t_L g417 ( .A(n_86), .B(n_187), .Y(n_417) );
INVx1_ASAP7_75t_L g440 ( .A(n_86), .Y(n_440) );
OAI21xp33_ASAP7_75t_L g476 ( .A1(n_86), .A2(n_169), .B(n_477), .Y(n_476) );
AO221x2_ASAP7_75t_L g841 ( .A1(n_87), .A2(n_367), .B1(n_828), .B2(n_833), .C(n_842), .Y(n_841) );
AOI22xp33_ASAP7_75t_L g1340 ( .A1(n_88), .A2(n_248), .B1(n_636), .B2(n_642), .Y(n_1340) );
AOI22xp33_ASAP7_75t_L g1284 ( .A1(n_89), .A2(n_343), .B1(n_532), .B2(n_1105), .Y(n_1284) );
AOI22xp5_ASAP7_75t_L g803 ( .A1(n_90), .A2(n_266), .B1(n_558), .B2(n_559), .Y(n_803) );
AOI22xp5_ASAP7_75t_L g809 ( .A1(n_91), .A2(n_393), .B1(n_665), .B2(n_669), .Y(n_809) );
AOI21xp5_ASAP7_75t_L g751 ( .A1(n_92), .A2(n_481), .B(n_752), .Y(n_751) );
AOI22xp5_ASAP7_75t_L g846 ( .A1(n_93), .A2(n_351), .B1(n_847), .B2(n_849), .Y(n_846) );
AOI22xp33_ASAP7_75t_L g1076 ( .A1(n_95), .A2(n_271), .B1(n_709), .B2(n_1077), .Y(n_1076) );
XNOR2x1_ASAP7_75t_L g423 ( .A(n_97), .B(n_424), .Y(n_423) );
AOI22xp33_ASAP7_75t_L g869 ( .A1(n_97), .A2(n_377), .B1(n_836), .B2(n_870), .Y(n_869) );
AOI22xp5_ASAP7_75t_L g1339 ( .A1(n_98), .A2(n_239), .B1(n_632), .B2(n_635), .Y(n_1339) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_99), .B(n_734), .Y(n_733) );
INVx1_ASAP7_75t_L g832 ( .A(n_100), .Y(n_832) );
AND2x4_ASAP7_75t_L g837 ( .A(n_100), .B(n_299), .Y(n_837) );
INVx1_ASAP7_75t_L g1066 ( .A(n_101), .Y(n_1066) );
INVx1_ASAP7_75t_L g690 ( .A(n_102), .Y(n_690) );
AO22x1_ASAP7_75t_L g842 ( .A1(n_103), .A2(n_193), .B1(n_843), .B2(n_844), .Y(n_842) );
AOI22xp33_ASAP7_75t_L g1240 ( .A1(n_104), .A2(n_230), .B1(n_635), .B2(n_636), .Y(n_1240) );
AOI22xp5_ASAP7_75t_L g1198 ( .A1(n_105), .A2(n_359), .B1(n_632), .B2(n_633), .Y(n_1198) );
AOI22xp33_ASAP7_75t_L g1192 ( .A1(n_106), .A2(n_292), .B1(n_626), .B2(n_628), .Y(n_1192) );
AOI22xp5_ASAP7_75t_L g607 ( .A1(n_107), .A2(n_306), .B1(n_526), .B2(n_608), .Y(n_607) );
INVx1_ASAP7_75t_L g616 ( .A(n_108), .Y(n_616) );
AOI22xp5_ASAP7_75t_L g850 ( .A1(n_108), .A2(n_145), .B1(n_838), .B2(n_851), .Y(n_850) );
AOI22xp33_ASAP7_75t_L g1219 ( .A1(n_109), .A2(n_354), .B1(n_429), .B2(n_581), .Y(n_1219) );
AOI22xp33_ASAP7_75t_L g504 ( .A1(n_111), .A2(n_231), .B1(n_505), .B2(n_511), .Y(n_504) );
INVx1_ASAP7_75t_L g1319 ( .A(n_112), .Y(n_1319) );
AOI22xp33_ASAP7_75t_L g808 ( .A1(n_113), .A2(n_274), .B1(n_429), .B2(n_731), .Y(n_808) );
AOI221xp5_ASAP7_75t_L g1232 ( .A1(n_114), .A2(n_321), .B1(n_621), .B2(n_645), .C(n_1233), .Y(n_1232) );
AOI22xp33_ASAP7_75t_L g789 ( .A1(n_115), .A2(n_260), .B1(n_505), .B2(n_709), .Y(n_789) );
AOI22xp33_ASAP7_75t_L g1287 ( .A1(n_116), .A2(n_183), .B1(n_538), .B2(n_541), .Y(n_1287) );
INVx1_ASAP7_75t_SL g1270 ( .A(n_117), .Y(n_1270) );
AOI22xp33_ASAP7_75t_L g1360 ( .A1(n_119), .A2(n_178), .B1(n_639), .B2(n_640), .Y(n_1360) );
NAND2xp5_ASAP7_75t_L g1190 ( .A(n_120), .B(n_621), .Y(n_1190) );
AOI22xp33_ASAP7_75t_L g597 ( .A1(n_121), .A2(n_172), .B1(n_568), .B2(n_598), .Y(n_597) );
INVx1_ASAP7_75t_L g830 ( .A(n_122), .Y(n_830) );
AND2x4_ASAP7_75t_L g834 ( .A(n_122), .B(n_413), .Y(n_834) );
INVx1_ASAP7_75t_SL g848 ( .A(n_122), .Y(n_848) );
NAND2xp5_ASAP7_75t_L g1310 ( .A(n_123), .B(n_1138), .Y(n_1310) );
AOI22xp33_ASAP7_75t_L g1145 ( .A1(n_124), .A2(n_300), .B1(n_505), .B2(n_1146), .Y(n_1145) );
AOI22xp5_ASAP7_75t_L g677 ( .A1(n_125), .A2(n_346), .B1(n_519), .B2(n_550), .Y(n_677) );
AOI22xp5_ASAP7_75t_L g1239 ( .A1(n_126), .A2(n_158), .B1(n_519), .B2(n_706), .Y(n_1239) );
AOI22xp5_ASAP7_75t_L g622 ( .A1(n_127), .A2(n_272), .B1(n_623), .B2(n_624), .Y(n_622) );
AOI22xp5_ASAP7_75t_L g1176 ( .A1(n_129), .A2(n_339), .B1(n_558), .B2(n_605), .Y(n_1176) );
AOI22xp33_ASAP7_75t_L g1236 ( .A1(n_130), .A2(n_370), .B1(n_623), .B2(n_629), .Y(n_1236) );
AOI22xp33_ASAP7_75t_L g1291 ( .A1(n_131), .A2(n_133), .B1(n_462), .B2(n_469), .Y(n_1291) );
AOI22xp33_ASAP7_75t_L g859 ( .A1(n_134), .A2(n_165), .B1(n_836), .B2(n_844), .Y(n_859) );
OAI22x1_ASAP7_75t_L g1101 ( .A1(n_134), .A2(n_1102), .B1(n_1117), .B2(n_1127), .Y(n_1101) );
NAND3xp33_ASAP7_75t_L g1102 ( .A(n_134), .B(n_1103), .C(n_1109), .Y(n_1102) );
INVx1_ASAP7_75t_L g1234 ( .A(n_135), .Y(n_1234) );
AOI22xp33_ASAP7_75t_L g1140 ( .A1(n_136), .A2(n_176), .B1(n_759), .B2(n_771), .Y(n_1140) );
INVx1_ASAP7_75t_L g460 ( .A(n_138), .Y(n_460) );
XOR2x2_ASAP7_75t_L g1132 ( .A(n_139), .B(n_1133), .Y(n_1132) );
AOI22xp33_ASAP7_75t_L g748 ( .A1(n_140), .A2(n_196), .B1(n_608), .B2(n_749), .Y(n_748) );
AOI221xp5_ASAP7_75t_L g774 ( .A1(n_141), .A2(n_152), .B1(n_775), .B2(n_776), .C(n_778), .Y(n_774) );
AOI221xp5_ASAP7_75t_L g797 ( .A1(n_141), .A2(n_152), .B1(n_775), .B2(n_776), .C(n_778), .Y(n_797) );
AOI22xp33_ASAP7_75t_L g1172 ( .A1(n_143), .A2(n_341), .B1(n_552), .B2(n_553), .Y(n_1172) );
XNOR2x1_ASAP7_75t_L g799 ( .A(n_146), .B(n_800), .Y(n_799) );
AOI22xp33_ASAP7_75t_L g537 ( .A1(n_147), .A2(n_202), .B1(n_538), .B2(n_540), .Y(n_537) );
INVx1_ASAP7_75t_L g573 ( .A(n_148), .Y(n_573) );
INVx1_ASAP7_75t_L g1253 ( .A(n_149), .Y(n_1253) );
AOI22xp33_ASAP7_75t_L g678 ( .A1(n_150), .A2(n_276), .B1(n_558), .B2(n_679), .Y(n_678) );
AO22x1_ASAP7_75t_L g1199 ( .A1(n_153), .A2(n_309), .B1(n_635), .B2(n_636), .Y(n_1199) );
INVx1_ASAP7_75t_L g738 ( .A(n_154), .Y(n_738) );
AOI22xp33_ASAP7_75t_L g1216 ( .A1(n_155), .A2(n_385), .B1(n_635), .B2(n_636), .Y(n_1216) );
AOI22xp33_ASAP7_75t_L g1107 ( .A1(n_156), .A2(n_357), .B1(n_608), .B2(n_1108), .Y(n_1107) );
AOI22xp33_ASAP7_75t_L g1079 ( .A1(n_157), .A2(n_317), .B1(n_505), .B2(n_788), .Y(n_1079) );
XNOR2xp5_ASAP7_75t_L g1088 ( .A(n_160), .B(n_1089), .Y(n_1088) );
AOI22xp33_ASAP7_75t_L g713 ( .A1(n_161), .A2(n_342), .B1(n_555), .B2(n_714), .Y(n_713) );
AOI22xp33_ASAP7_75t_L g517 ( .A1(n_162), .A2(n_378), .B1(n_518), .B2(n_525), .Y(n_517) );
AOI22xp33_ASAP7_75t_L g1228 ( .A1(n_163), .A2(n_209), .B1(n_714), .B2(n_792), .Y(n_1228) );
AOI22xp33_ASAP7_75t_L g791 ( .A1(n_164), .A2(n_288), .B1(n_792), .B2(n_793), .Y(n_791) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_167), .B(n_658), .Y(n_657) );
INVx1_ASAP7_75t_L g451 ( .A(n_168), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_168), .B(n_227), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_168), .B(n_473), .Y(n_502) );
NOR2xp33_ASAP7_75t_L g416 ( .A(n_169), .B(n_308), .Y(n_416) );
AOI22xp33_ASAP7_75t_L g962 ( .A1(n_170), .A2(n_241), .B1(n_867), .B2(n_963), .Y(n_962) );
AOI22xp33_ASAP7_75t_L g1341 ( .A1(n_171), .A2(n_216), .B1(n_639), .B2(n_640), .Y(n_1341) );
AOI221xp5_ASAP7_75t_L g810 ( .A1(n_173), .A2(n_365), .B1(n_811), .B2(n_812), .C(n_814), .Y(n_810) );
AOI22xp33_ASAP7_75t_L g705 ( .A1(n_174), .A2(n_331), .B1(n_706), .B2(n_707), .Y(n_705) );
INVx1_ASAP7_75t_L g660 ( .A(n_175), .Y(n_660) );
AOI22xp33_ASAP7_75t_L g580 ( .A1(n_177), .A2(n_368), .B1(n_581), .B2(n_582), .Y(n_580) );
INVx1_ASAP7_75t_SL g1258 ( .A(n_179), .Y(n_1258) );
INVx1_ASAP7_75t_L g1211 ( .A(n_182), .Y(n_1211) );
NAND2xp5_ASAP7_75t_L g755 ( .A(n_184), .B(n_756), .Y(n_755) );
AOI22xp33_ASAP7_75t_L g1058 ( .A1(n_185), .A2(n_213), .B1(n_769), .B2(n_1059), .Y(n_1058) );
AOI21xp33_ASAP7_75t_L g1311 ( .A1(n_186), .A2(n_1312), .B(n_1313), .Y(n_1311) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_187), .B(n_444), .Y(n_443) );
AO22x1_ASAP7_75t_L g1200 ( .A1(n_188), .A2(n_344), .B1(n_642), .B2(n_643), .Y(n_1200) );
AOI22xp33_ASAP7_75t_L g1305 ( .A1(n_190), .A2(n_208), .B1(n_608), .B2(n_787), .Y(n_1305) );
NAND2xp5_ASAP7_75t_L g1164 ( .A(n_191), .B(n_1138), .Y(n_1164) );
AOI22xp33_ASAP7_75t_L g551 ( .A1(n_192), .A2(n_282), .B1(n_552), .B2(n_553), .Y(n_551) );
XOR2x2_ASAP7_75t_L g545 ( .A(n_193), .B(n_546), .Y(n_545) );
XNOR2xp5_ASAP7_75t_L g611 ( .A(n_193), .B(n_546), .Y(n_611) );
AOI22xp33_ASAP7_75t_L g485 ( .A1(n_197), .A2(n_236), .B1(n_486), .B2(n_496), .Y(n_485) );
AOI21xp33_ASAP7_75t_SL g696 ( .A1(n_198), .A2(n_697), .B(n_698), .Y(n_696) );
INVx1_ASAP7_75t_L g562 ( .A(n_199), .Y(n_562) );
AOI21xp5_ASAP7_75t_L g1193 ( .A1(n_203), .A2(n_645), .B(n_1194), .Y(n_1193) );
AOI22xp33_ASAP7_75t_L g1256 ( .A1(n_204), .A2(n_322), .B1(n_538), .B2(n_1108), .Y(n_1256) );
AOI22xp33_ASAP7_75t_L g1122 ( .A1(n_205), .A2(n_400), .B1(n_462), .B2(n_469), .Y(n_1122) );
NAND2xp5_ASAP7_75t_SL g700 ( .A(n_206), .B(n_701), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g1221 ( .A(n_207), .B(n_658), .Y(n_1221) );
AOI22xp33_ASAP7_75t_L g702 ( .A1(n_210), .A2(n_383), .B1(n_665), .B2(n_703), .Y(n_702) );
NAND2xp33_ASAP7_75t_L g619 ( .A(n_211), .B(n_620), .Y(n_619) );
AOI22xp33_ASAP7_75t_L g1215 ( .A1(n_212), .A2(n_302), .B1(n_519), .B2(n_526), .Y(n_1215) );
INVx1_ASAP7_75t_L g1318 ( .A(n_214), .Y(n_1318) );
AOI22xp33_ASAP7_75t_L g742 ( .A1(n_218), .A2(n_255), .B1(n_602), .B2(n_743), .Y(n_742) );
AOI22xp33_ASAP7_75t_L g1060 ( .A1(n_219), .A2(n_301), .B1(n_1061), .B2(n_1062), .Y(n_1060) );
XOR2x2_ASAP7_75t_L g1244 ( .A(n_220), .B(n_1245), .Y(n_1244) );
AOI22xp33_ASAP7_75t_SL g1335 ( .A1(n_221), .A2(n_253), .B1(n_623), .B2(n_629), .Y(n_1335) );
AOI221xp5_ASAP7_75t_L g1292 ( .A1(n_222), .A2(n_381), .B1(n_429), .B2(n_1293), .C(n_1294), .Y(n_1292) );
AOI22xp5_ASAP7_75t_L g827 ( .A1(n_225), .A2(n_258), .B1(n_828), .B2(n_833), .Y(n_827) );
AOI22xp33_ASAP7_75t_L g785 ( .A1(n_226), .A2(n_228), .B1(n_786), .B2(n_788), .Y(n_785) );
INVx1_ASAP7_75t_L g438 ( .A(n_227), .Y(n_438) );
AOI22xp33_ASAP7_75t_L g1069 ( .A1(n_232), .A2(n_293), .B1(n_795), .B2(n_1070), .Y(n_1069) );
AOI22xp33_ASAP7_75t_L g864 ( .A1(n_233), .A2(n_338), .B1(n_828), .B2(n_849), .Y(n_864) );
AOI22xp33_ASAP7_75t_L g554 ( .A1(n_234), .A2(n_376), .B1(n_555), .B2(n_556), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g1322 ( .A(n_237), .B(n_731), .Y(n_1322) );
INVx1_ASAP7_75t_L g699 ( .A(n_240), .Y(n_699) );
AOI22xp33_ASAP7_75t_L g1175 ( .A1(n_242), .A2(n_311), .B1(n_519), .B2(n_787), .Y(n_1175) );
AOI22xp5_ASAP7_75t_L g876 ( .A1(n_243), .A2(n_295), .B1(n_828), .B2(n_849), .Y(n_876) );
AOI22xp33_ASAP7_75t_L g601 ( .A1(n_244), .A2(n_250), .B1(n_602), .B2(n_603), .Y(n_601) );
AOI22xp33_ASAP7_75t_L g528 ( .A1(n_245), .A2(n_373), .B1(n_529), .B2(n_532), .Y(n_528) );
AOI22xp33_ASAP7_75t_L g802 ( .A1(n_249), .A2(n_281), .B1(n_549), .B2(n_787), .Y(n_802) );
AOI22xp33_ASAP7_75t_L g599 ( .A1(n_251), .A2(n_347), .B1(n_462), .B2(n_469), .Y(n_599) );
CKINVDCx14_ASAP7_75t_R g1329 ( .A(n_256), .Y(n_1329) );
AOI22xp5_ASAP7_75t_L g1119 ( .A1(n_257), .A2(n_277), .B1(n_1120), .B2(n_1121), .Y(n_1119) );
AOI22xp33_ASAP7_75t_L g1306 ( .A1(n_259), .A2(n_264), .B1(n_556), .B2(n_602), .Y(n_1306) );
XNOR2x2_ASAP7_75t_L g1187 ( .A(n_261), .B(n_1188), .Y(n_1187) );
AOI22xp33_ASAP7_75t_L g866 ( .A1(n_262), .A2(n_334), .B1(n_828), .B2(n_867), .Y(n_866) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_263), .B(n_581), .Y(n_670) );
AOI22xp33_ASAP7_75t_L g863 ( .A1(n_267), .A2(n_330), .B1(n_843), .B2(n_844), .Y(n_863) );
AOI22xp33_ASAP7_75t_L g1358 ( .A1(n_268), .A2(n_340), .B1(n_632), .B2(n_635), .Y(n_1358) );
INVx1_ASAP7_75t_L g570 ( .A(n_269), .Y(n_570) );
AOI22xp33_ASAP7_75t_L g1237 ( .A1(n_270), .A2(n_324), .B1(n_626), .B2(n_628), .Y(n_1237) );
AOI22xp33_ASAP7_75t_L g1307 ( .A1(n_273), .A2(n_356), .B1(n_558), .B2(n_1108), .Y(n_1307) );
INVx1_ASAP7_75t_L g1321 ( .A(n_275), .Y(n_1321) );
AOI22xp5_ASAP7_75t_L g806 ( .A1(n_278), .A2(n_303), .B1(n_555), .B2(n_714), .Y(n_806) );
INVx1_ASAP7_75t_L g586 ( .A(n_279), .Y(n_586) );
AOI22xp5_ASAP7_75t_L g835 ( .A1(n_279), .A2(n_358), .B1(n_836), .B2(n_838), .Y(n_835) );
INVx1_ASAP7_75t_L g1314 ( .A(n_280), .Y(n_1314) );
INVx1_ASAP7_75t_L g467 ( .A(n_283), .Y(n_467) );
AOI221xp5_ASAP7_75t_L g1063 ( .A1(n_284), .A2(n_402), .B1(n_486), .B2(n_1064), .C(n_1065), .Y(n_1063) );
AOI22xp33_ASAP7_75t_L g1125 ( .A1(n_285), .A2(n_291), .B1(n_550), .B2(n_1126), .Y(n_1125) );
CKINVDCx5p33_ASAP7_75t_R g1168 ( .A(n_286), .Y(n_1168) );
AOI22xp33_ASAP7_75t_L g1377 ( .A1(n_287), .A2(n_314), .B1(n_572), .B2(n_1378), .Y(n_1377) );
AOI22xp5_ASAP7_75t_L g728 ( .A1(n_289), .A2(n_401), .B1(n_541), .B2(n_558), .Y(n_728) );
INVx1_ASAP7_75t_L g754 ( .A(n_290), .Y(n_754) );
INVx1_ASAP7_75t_L g779 ( .A(n_294), .Y(n_779) );
AOI22xp33_ASAP7_75t_L g760 ( .A1(n_296), .A2(n_371), .B1(n_454), .B2(n_564), .Y(n_760) );
INVx1_ASAP7_75t_L g566 ( .A(n_297), .Y(n_566) );
HB1xp67_ASAP7_75t_L g418 ( .A(n_299), .Y(n_418) );
AND2x4_ASAP7_75t_L g831 ( .A(n_299), .B(n_832), .Y(n_831) );
AOI22xp33_ASAP7_75t_L g1290 ( .A1(n_304), .A2(n_349), .B1(n_486), .B2(n_1121), .Y(n_1290) );
INVx1_ASAP7_75t_L g576 ( .A(n_307), .Y(n_576) );
INVx1_ASAP7_75t_L g449 ( .A(n_308), .Y(n_449) );
INVxp67_ASAP7_75t_L g495 ( .A(n_308), .Y(n_495) );
AOI22xp33_ASAP7_75t_L g1348 ( .A1(n_310), .A2(n_386), .B1(n_626), .B2(n_662), .Y(n_1348) );
OAI21x1_ASAP7_75t_L g1225 ( .A1(n_312), .A2(n_1226), .B(n_1241), .Y(n_1225) );
NAND4xp25_ASAP7_75t_L g1241 ( .A(n_312), .B(n_1227), .C(n_1231), .D(n_1238), .Y(n_1241) );
INVxp67_ASAP7_75t_R g1160 ( .A(n_315), .Y(n_1160) );
INVx1_ASAP7_75t_L g1185 ( .A(n_315), .Y(n_1185) );
INVx1_ASAP7_75t_L g1272 ( .A(n_316), .Y(n_1272) );
INVx2_ASAP7_75t_L g413 ( .A(n_318), .Y(n_413) );
INVx1_ASAP7_75t_L g452 ( .A(n_319), .Y(n_452) );
XOR2x2_ASAP7_75t_L g739 ( .A(n_320), .B(n_740), .Y(n_739) );
INVx1_ASAP7_75t_L g667 ( .A(n_325), .Y(n_667) );
INVx1_ASAP7_75t_L g1268 ( .A(n_326), .Y(n_1268) );
INVx1_ASAP7_75t_L g1115 ( .A(n_328), .Y(n_1115) );
XNOR2x1_ASAP7_75t_L g649 ( .A(n_330), .B(n_650), .Y(n_649) );
AOI22xp33_ASAP7_75t_L g1359 ( .A1(n_332), .A2(n_366), .B1(n_636), .B2(n_642), .Y(n_1359) );
AOI22xp33_ASAP7_75t_L g1304 ( .A1(n_333), .A2(n_389), .B1(n_553), .B2(n_675), .Y(n_1304) );
INVx1_ASAP7_75t_L g1195 ( .A(n_336), .Y(n_1195) );
AOI22xp5_ASAP7_75t_L g634 ( .A1(n_345), .A2(n_382), .B1(n_635), .B2(n_636), .Y(n_634) );
INVx1_ASAP7_75t_L g1250 ( .A(n_348), .Y(n_1250) );
AOI22xp5_ASAP7_75t_L g631 ( .A1(n_352), .A2(n_361), .B1(n_632), .B2(n_633), .Y(n_631) );
AOI22xp33_ASAP7_75t_L g744 ( .A1(n_353), .A2(n_362), .B1(n_538), .B2(n_745), .Y(n_744) );
INVx1_ASAP7_75t_L g479 ( .A(n_355), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g1336 ( .A(n_360), .B(n_781), .Y(n_1336) );
AOI21xp33_ASAP7_75t_L g653 ( .A1(n_364), .A2(n_654), .B(n_655), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g1263 ( .A(n_372), .B(n_1264), .Y(n_1263) );
INVx1_ASAP7_75t_L g663 ( .A(n_375), .Y(n_663) );
AOI22xp33_ASAP7_75t_L g609 ( .A1(n_379), .A2(n_391), .B1(n_553), .B2(n_610), .Y(n_609) );
AOI21xp5_ASAP7_75t_L g1109 ( .A1(n_380), .A2(n_1110), .B(n_1112), .Y(n_1109) );
CKINVDCx5p33_ASAP7_75t_R g1369 ( .A(n_384), .Y(n_1369) );
INVxp67_ASAP7_75t_SL g782 ( .A(n_387), .Y(n_782) );
AOI21xp33_ASAP7_75t_L g1351 ( .A1(n_397), .A2(n_628), .B(n_1352), .Y(n_1351) );
AOI21xp33_ASAP7_75t_SL g644 ( .A1(n_398), .A2(n_645), .B(n_646), .Y(n_644) );
AOI22xp33_ASAP7_75t_L g1179 ( .A1(n_399), .A2(n_405), .B1(n_697), .B2(n_1180), .Y(n_1179) );
CKINVDCx20_ASAP7_75t_R g1375 ( .A(n_403), .Y(n_1375) );
OAI21xp5_ASAP7_75t_L g407 ( .A1(n_408), .A2(n_1095), .B(n_1392), .Y(n_407) );
OAI21xp33_ASAP7_75t_L g408 ( .A1(n_409), .A2(n_419), .B(n_819), .Y(n_408) );
INVx2_ASAP7_75t_R g1391 ( .A(n_409), .Y(n_1391) );
BUFx4_ASAP7_75t_SL g409 ( .A(n_410), .Y(n_409) );
NAND3xp33_ASAP7_75t_L g410 ( .A(n_411), .B(n_414), .C(n_418), .Y(n_410) );
AND2x2_ASAP7_75t_L g1083 ( .A(n_411), .B(n_1084), .Y(n_1083) );
AND2x2_ASAP7_75t_L g1091 ( .A(n_411), .B(n_1085), .Y(n_1091) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
OA21x2_ASAP7_75t_L g1093 ( .A1(n_412), .A2(n_848), .B(n_1094), .Y(n_1093) );
HB1xp67_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
AND2x2_ASAP7_75t_L g829 ( .A(n_413), .B(n_830), .Y(n_829) );
AND3x4_ASAP7_75t_L g847 ( .A(n_413), .B(n_831), .C(n_848), .Y(n_847) );
NOR2xp33_ASAP7_75t_L g1084 ( .A(n_414), .B(n_1085), .Y(n_1084) );
HB1xp67_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
AO21x2_ASAP7_75t_L g499 ( .A1(n_415), .A2(n_500), .B(n_501), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_416), .B(n_417), .Y(n_415) );
INVx1_ASAP7_75t_L g1085 ( .A(n_418), .Y(n_1085) );
INVx2_ASAP7_75t_L g1393 ( .A(n_419), .Y(n_1393) );
XNOR2xp5_ASAP7_75t_L g419 ( .A(n_420), .B(n_682), .Y(n_419) );
XOR2xp5_ASAP7_75t_L g420 ( .A(n_421), .B(n_612), .Y(n_420) );
XOR2x2_ASAP7_75t_L g421 ( .A(n_422), .B(n_544), .Y(n_421) );
INVx1_ASAP7_75t_SL g422 ( .A(n_423), .Y(n_422) );
AND2x4_ASAP7_75t_L g424 ( .A(n_425), .B(n_503), .Y(n_424) );
NOR3xp33_ASAP7_75t_L g425 ( .A(n_426), .B(n_459), .C(n_478), .Y(n_425) );
OAI22xp5_ASAP7_75t_L g426 ( .A1(n_427), .A2(n_428), .B1(n_452), .B2(n_453), .Y(n_426) );
INVx2_ASAP7_75t_L g768 ( .A(n_428), .Y(n_768) );
INVx2_ASAP7_75t_L g1120 ( .A(n_428), .Y(n_1120) );
INVx2_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
BUFx3_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g565 ( .A(n_430), .Y(n_565) );
BUFx3_ASAP7_75t_L g654 ( .A(n_430), .Y(n_654) );
BUFx6f_ASAP7_75t_L g1312 ( .A(n_430), .Y(n_1312) );
AND2x4_ASAP7_75t_L g430 ( .A(n_431), .B(n_441), .Y(n_430) );
AND2x4_ASAP7_75t_L g464 ( .A(n_431), .B(n_465), .Y(n_464) );
AND2x4_ASAP7_75t_L g628 ( .A(n_431), .B(n_441), .Y(n_628) );
AND2x2_ASAP7_75t_L g645 ( .A(n_431), .B(n_465), .Y(n_645) );
AND2x2_ASAP7_75t_L g431 ( .A(n_432), .B(n_435), .Y(n_431) );
AND2x2_ASAP7_75t_L g458 ( .A(n_432), .B(n_436), .Y(n_458) );
AND2x2_ASAP7_75t_L g493 ( .A(n_432), .B(n_494), .Y(n_493) );
INVx1_ASAP7_75t_L g522 ( .A(n_432), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_433), .B(n_440), .Y(n_439) );
INVx2_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
NAND2xp33_ASAP7_75t_L g437 ( .A(n_434), .B(n_438), .Y(n_437) );
INVx3_ASAP7_75t_L g444 ( .A(n_434), .Y(n_444) );
NAND2xp33_ASAP7_75t_L g450 ( .A(n_434), .B(n_451), .Y(n_450) );
INVx1_ASAP7_75t_L g477 ( .A(n_434), .Y(n_477) );
HB1xp67_ASAP7_75t_L g491 ( .A(n_434), .Y(n_491) );
AND2x4_ASAP7_75t_L g521 ( .A(n_435), .B(n_522), .Y(n_521) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_437), .B(n_439), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_438), .B(n_475), .Y(n_474) );
OAI21xp5_ASAP7_75t_L g494 ( .A1(n_440), .A2(n_477), .B(n_495), .Y(n_494) );
AND2x2_ASAP7_75t_L g457 ( .A(n_441), .B(n_458), .Y(n_457) );
AND2x4_ASAP7_75t_L g531 ( .A(n_441), .B(n_521), .Y(n_531) );
AND2x4_ASAP7_75t_L g623 ( .A(n_441), .B(n_458), .Y(n_623) );
AND2x4_ASAP7_75t_L g639 ( .A(n_441), .B(n_521), .Y(n_639) );
AND2x4_ASAP7_75t_L g441 ( .A(n_442), .B(n_446), .Y(n_441) );
INVx2_ASAP7_75t_L g466 ( .A(n_442), .Y(n_466) );
AND2x2_ASAP7_75t_L g489 ( .A(n_442), .B(n_490), .Y(n_489) );
OR2x2_ASAP7_75t_L g509 ( .A(n_442), .B(n_510), .Y(n_509) );
AND2x4_ASAP7_75t_L g523 ( .A(n_442), .B(n_524), .Y(n_523) );
AND2x4_ASAP7_75t_L g442 ( .A(n_443), .B(n_445), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_444), .B(n_449), .Y(n_448) );
INVxp67_ASAP7_75t_L g473 ( .A(n_444), .Y(n_473) );
NAND3xp33_ASAP7_75t_L g501 ( .A(n_445), .B(n_472), .C(n_502), .Y(n_501) );
AND2x4_ASAP7_75t_L g465 ( .A(n_446), .B(n_466), .Y(n_465) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx1_ASAP7_75t_L g510 ( .A(n_447), .Y(n_510) );
AND2x2_ASAP7_75t_L g447 ( .A(n_448), .B(n_450), .Y(n_447) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx2_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx2_ASAP7_75t_L g1121 ( .A(n_455), .Y(n_1121) );
BUFx6f_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVx2_ASAP7_75t_L g669 ( .A(n_456), .Y(n_669) );
INVx2_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
BUFx3_ASAP7_75t_L g568 ( .A(n_457), .Y(n_568) );
BUFx6f_ASAP7_75t_L g703 ( .A(n_457), .Y(n_703) );
AND2x2_ASAP7_75t_L g484 ( .A(n_458), .B(n_465), .Y(n_484) );
AND2x4_ASAP7_75t_L g507 ( .A(n_458), .B(n_508), .Y(n_507) );
AND2x2_ASAP7_75t_L g539 ( .A(n_458), .B(n_523), .Y(n_539) );
AND2x2_ASAP7_75t_L g621 ( .A(n_458), .B(n_465), .Y(n_621) );
AND2x4_ASAP7_75t_L g632 ( .A(n_458), .B(n_516), .Y(n_632) );
AND2x4_ASAP7_75t_L g635 ( .A(n_458), .B(n_523), .Y(n_635) );
AND2x2_ASAP7_75t_L g710 ( .A(n_458), .B(n_523), .Y(n_710) );
OAI22xp5_ASAP7_75t_L g459 ( .A1(n_460), .A2(n_461), .B1(n_467), .B2(n_468), .Y(n_459) );
OAI22xp5_ASAP7_75t_L g1317 ( .A1(n_461), .A2(n_468), .B1(n_1318), .B2(n_1319), .Y(n_1317) );
INVx2_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx2_ASAP7_75t_SL g462 ( .A(n_463), .Y(n_462) );
INVx2_ASAP7_75t_SL g811 ( .A(n_463), .Y(n_811) );
INVx2_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
BUFx3_ASAP7_75t_L g572 ( .A(n_464), .Y(n_572) );
BUFx6f_ASAP7_75t_L g662 ( .A(n_464), .Y(n_662) );
BUFx6f_ASAP7_75t_L g697 ( .A(n_464), .Y(n_697) );
INVx2_ASAP7_75t_L g735 ( .A(n_464), .Y(n_735) );
BUFx8_ASAP7_75t_SL g758 ( .A(n_464), .Y(n_758) );
AND2x4_ASAP7_75t_L g470 ( .A(n_465), .B(n_471), .Y(n_470) );
AND2x2_ASAP7_75t_L g536 ( .A(n_465), .B(n_521), .Y(n_536) );
AND2x4_ASAP7_75t_L g626 ( .A(n_465), .B(n_471), .Y(n_626) );
AND2x4_ASAP7_75t_L g640 ( .A(n_465), .B(n_521), .Y(n_640) );
INVx4_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
BUFx3_ASAP7_75t_L g759 ( .A(n_469), .Y(n_759) );
BUFx6f_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
INVx3_ASAP7_75t_L g574 ( .A(n_470), .Y(n_574) );
BUFx6f_ASAP7_75t_L g665 ( .A(n_470), .Y(n_665) );
AND2x4_ASAP7_75t_L g515 ( .A(n_471), .B(n_516), .Y(n_515) );
AND2x4_ASAP7_75t_L g543 ( .A(n_471), .B(n_523), .Y(n_543) );
AND2x4_ASAP7_75t_L g633 ( .A(n_471), .B(n_516), .Y(n_633) );
AND2x4_ASAP7_75t_L g636 ( .A(n_471), .B(n_523), .Y(n_636) );
AND2x2_ASAP7_75t_L g471 ( .A(n_472), .B(n_476), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_473), .B(n_474), .Y(n_472) );
OAI21xp33_ASAP7_75t_L g478 ( .A1(n_479), .A2(n_480), .B(n_485), .Y(n_478) );
INVx1_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
INVx2_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx1_ASAP7_75t_L g701 ( .A(n_482), .Y(n_701) );
INVx2_ASAP7_75t_L g1138 ( .A(n_482), .Y(n_1138) );
BUFx6f_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
INVx2_ASAP7_75t_L g1265 ( .A(n_483), .Y(n_1265) );
INVx2_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
INVx3_ASAP7_75t_L g579 ( .A(n_484), .Y(n_579) );
BUFx3_ASAP7_75t_L g737 ( .A(n_484), .Y(n_737) );
INVx1_ASAP7_75t_L g1114 ( .A(n_486), .Y(n_1114) );
INVx3_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
INVx2_ASAP7_75t_L g598 ( .A(n_487), .Y(n_598) );
INVx4_ASAP7_75t_L g731 ( .A(n_487), .Y(n_731) );
INVx2_ASAP7_75t_L g775 ( .A(n_487), .Y(n_775) );
INVx2_ASAP7_75t_L g1182 ( .A(n_487), .Y(n_1182) );
INVx5_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
BUFx4f_ASAP7_75t_L g581 ( .A(n_488), .Y(n_581) );
BUFx2_ASAP7_75t_L g695 ( .A(n_488), .Y(n_695) );
AND2x4_ASAP7_75t_L g488 ( .A(n_489), .B(n_493), .Y(n_488) );
AND2x4_ASAP7_75t_L g629 ( .A(n_489), .B(n_493), .Y(n_629) );
AND2x2_ASAP7_75t_L g1350 ( .A(n_489), .B(n_493), .Y(n_1350) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_491), .B(n_492), .Y(n_490) );
INVx1_ASAP7_75t_L g500 ( .A(n_491), .Y(n_500) );
INVx4_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
NOR2xp33_ASAP7_75t_L g1065 ( .A(n_497), .B(n_1066), .Y(n_1065) );
NOR2xp33_ASAP7_75t_L g1223 ( .A(n_497), .B(n_1224), .Y(n_1223) );
NOR2xp33_ASAP7_75t_L g1233 ( .A(n_497), .B(n_1234), .Y(n_1233) );
NOR2xp33_ASAP7_75t_L g1294 ( .A(n_497), .B(n_1295), .Y(n_1294) );
INVx3_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
INVx4_ASAP7_75t_L g583 ( .A(n_498), .Y(n_583) );
INVx3_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
BUFx6f_ASAP7_75t_L g595 ( .A(n_499), .Y(n_595) );
AND4x1_ASAP7_75t_L g503 ( .A(n_504), .B(n_517), .C(n_528), .D(n_537), .Y(n_503) );
BUFx3_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
BUFx12f_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
BUFx6f_ASAP7_75t_L g552 ( .A(n_507), .Y(n_552) );
BUFx6f_ASAP7_75t_L g610 ( .A(n_507), .Y(n_610) );
BUFx6f_ASAP7_75t_L g675 ( .A(n_507), .Y(n_675) );
BUFx3_ASAP7_75t_L g745 ( .A(n_507), .Y(n_745) );
AND2x4_ASAP7_75t_L g643 ( .A(n_508), .B(n_521), .Y(n_643) );
INVx2_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
INVx2_ASAP7_75t_L g516 ( .A(n_509), .Y(n_516) );
INVx1_ASAP7_75t_L g524 ( .A(n_510), .Y(n_524) );
INVx1_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
INVx1_ASAP7_75t_L g1252 ( .A(n_512), .Y(n_1252) );
INVx1_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
INVx2_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
INVx5_ASAP7_75t_L g707 ( .A(n_514), .Y(n_707) );
INVx1_ASAP7_75t_L g747 ( .A(n_514), .Y(n_747) );
INVx1_ASAP7_75t_L g1126 ( .A(n_514), .Y(n_1126) );
INVx3_ASAP7_75t_L g1230 ( .A(n_514), .Y(n_1230) );
INVx2_ASAP7_75t_L g1383 ( .A(n_514), .Y(n_1383) );
INVx6_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
BUFx12f_ASAP7_75t_L g553 ( .A(n_515), .Y(n_553) );
AND2x4_ASAP7_75t_L g527 ( .A(n_516), .B(n_521), .Y(n_527) );
BUFx12f_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
BUFx6f_ASAP7_75t_L g795 ( .A(n_519), .Y(n_795) );
BUFx12f_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
BUFx6f_ASAP7_75t_L g549 ( .A(n_520), .Y(n_549) );
BUFx6f_ASAP7_75t_L g608 ( .A(n_520), .Y(n_608) );
AND2x4_ASAP7_75t_L g520 ( .A(n_521), .B(n_523), .Y(n_520) );
AND2x4_ASAP7_75t_L g642 ( .A(n_521), .B(n_523), .Y(n_642) );
BUFx3_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
INVx1_ASAP7_75t_L g1071 ( .A(n_526), .Y(n_1071) );
BUFx6f_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
BUFx6f_ASAP7_75t_L g550 ( .A(n_527), .Y(n_550) );
BUFx6f_ASAP7_75t_L g706 ( .A(n_527), .Y(n_706) );
BUFx6f_ASAP7_75t_L g787 ( .A(n_527), .Y(n_787) );
BUFx4f_ASAP7_75t_L g1105 ( .A(n_529), .Y(n_1105) );
INVx2_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
INVx1_ASAP7_75t_L g792 ( .A(n_530), .Y(n_792) );
INVx1_ASAP7_75t_L g1073 ( .A(n_530), .Y(n_1073) );
OAI22xp5_ASAP7_75t_L g1257 ( .A1(n_530), .A2(n_1258), .B1(n_1259), .B2(n_1260), .Y(n_1257) );
INVx3_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
BUFx12f_ASAP7_75t_L g555 ( .A(n_531), .Y(n_555) );
BUFx6f_ASAP7_75t_L g602 ( .A(n_531), .Y(n_602) );
INVx1_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
INVx1_ASAP7_75t_L g743 ( .A(n_533), .Y(n_743) );
INVx1_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
BUFx6f_ASAP7_75t_L g1106 ( .A(n_534), .Y(n_1106) );
INVx2_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
BUFx6f_ASAP7_75t_L g556 ( .A(n_536), .Y(n_556) );
BUFx5_ASAP7_75t_L g603 ( .A(n_536), .Y(n_603) );
BUFx3_ASAP7_75t_L g714 ( .A(n_536), .Y(n_714) );
BUFx8_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
BUFx6f_ASAP7_75t_L g558 ( .A(n_539), .Y(n_558) );
BUFx2_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
INVx4_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
INVx4_ASAP7_75t_L g559 ( .A(n_542), .Y(n_559) );
INVx2_ASAP7_75t_L g605 ( .A(n_542), .Y(n_605) );
INVx2_ASAP7_75t_SL g679 ( .A(n_542), .Y(n_679) );
INVx1_ASAP7_75t_L g712 ( .A(n_542), .Y(n_712) );
INVx1_ASAP7_75t_L g749 ( .A(n_542), .Y(n_749) );
INVx1_ASAP7_75t_L g1078 ( .A(n_542), .Y(n_1078) );
INVx4_ASAP7_75t_L g1108 ( .A(n_542), .Y(n_1108) );
INVx2_ASAP7_75t_L g1151 ( .A(n_542), .Y(n_1151) );
INVx8_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
AOI22x1_ASAP7_75t_L g544 ( .A1(n_545), .A2(n_584), .B1(n_585), .B2(n_611), .Y(n_544) );
AO22x2_ASAP7_75t_L g613 ( .A1(n_545), .A2(n_614), .B1(n_680), .B2(n_681), .Y(n_613) );
INVx1_ASAP7_75t_L g680 ( .A(n_545), .Y(n_680) );
AND2x4_ASAP7_75t_L g546 ( .A(n_547), .B(n_560), .Y(n_546) );
AND4x1_ASAP7_75t_L g547 ( .A(n_548), .B(n_551), .C(n_554), .D(n_557), .Y(n_547) );
BUFx2_ASAP7_75t_SL g1149 ( .A(n_549), .Y(n_1149) );
BUFx3_ASAP7_75t_L g1249 ( .A(n_552), .Y(n_1249) );
BUFx3_ASAP7_75t_L g788 ( .A(n_553), .Y(n_788) );
BUFx2_ASAP7_75t_SL g1074 ( .A(n_556), .Y(n_1074) );
INVx1_ASAP7_75t_L g1260 ( .A(n_556), .Y(n_1260) );
BUFx3_ASAP7_75t_L g1146 ( .A(n_558), .Y(n_1146) );
NOR3xp33_ASAP7_75t_L g560 ( .A(n_561), .B(n_569), .C(n_575), .Y(n_560) );
OAI22xp5_ASAP7_75t_L g561 ( .A1(n_562), .A2(n_563), .B1(n_566), .B2(n_567), .Y(n_561) );
INVx2_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
INVx2_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
INVx2_ASAP7_75t_L g1166 ( .A(n_565), .Y(n_1166) );
INVx2_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
BUFx2_ASAP7_75t_L g1142 ( .A(n_568), .Y(n_1142) );
OAI22xp5_ASAP7_75t_L g569 ( .A1(n_570), .A2(n_571), .B1(n_573), .B2(n_574), .Y(n_569) );
INVx2_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
INVx2_ASAP7_75t_L g1062 ( .A(n_574), .Y(n_1062) );
INVx3_ASAP7_75t_L g1180 ( .A(n_574), .Y(n_1180) );
INVx2_ASAP7_75t_L g1378 ( .A(n_574), .Y(n_1378) );
OAI21xp33_ASAP7_75t_L g575 ( .A1(n_576), .A2(n_577), .B(n_580), .Y(n_575) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
INVx1_ASAP7_75t_L g1111 ( .A(n_578), .Y(n_1111) );
INVx2_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
INVx2_ASAP7_75t_L g658 ( .A(n_579), .Y(n_658) );
INVx2_ASAP7_75t_L g777 ( .A(n_579), .Y(n_777) );
INVx2_ASAP7_75t_L g1355 ( .A(n_579), .Y(n_1355) );
INVx2_ASAP7_75t_L g1373 ( .A(n_579), .Y(n_1373) );
INVx2_ASAP7_75t_L g1116 ( .A(n_582), .Y(n_1116) );
INVx4_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
NOR2xp33_ASAP7_75t_L g1194 ( .A(n_583), .B(n_1195), .Y(n_1194) );
NOR2xp33_ASAP7_75t_L g1352 ( .A(n_583), .B(n_1353), .Y(n_1352) );
INVx2_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
XNOR2x1_ASAP7_75t_L g585 ( .A(n_586), .B(n_587), .Y(n_585) );
NOR4xp75_ASAP7_75t_L g587 ( .A(n_588), .B(n_596), .C(n_600), .D(n_606), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_589), .B(n_590), .Y(n_588) );
NOR2xp33_ASAP7_75t_L g591 ( .A(n_592), .B(n_593), .Y(n_591) );
NOR2xp33_ASAP7_75t_L g655 ( .A(n_593), .B(n_656), .Y(n_655) );
NOR2xp33_ASAP7_75t_L g1167 ( .A(n_593), .B(n_1168), .Y(n_1167) );
INVx3_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
INVx2_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
BUFx6f_ASAP7_75t_L g648 ( .A(n_595), .Y(n_648) );
INVx2_ASAP7_75t_SL g781 ( .A(n_595), .Y(n_781) );
INVx1_ASAP7_75t_L g1316 ( .A(n_595), .Y(n_1316) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_597), .B(n_599), .Y(n_596) );
NAND2xp5_ASAP7_75t_SL g600 ( .A(n_601), .B(n_604), .Y(n_600) );
BUFx3_ASAP7_75t_L g793 ( .A(n_603), .Y(n_793) );
NAND2xp5_ASAP7_75t_SL g606 ( .A(n_607), .B(n_609), .Y(n_606) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
INVx1_ASAP7_75t_L g681 ( .A(n_614), .Y(n_681) );
XNOR2xp5_ASAP7_75t_L g614 ( .A(n_615), .B(n_649), .Y(n_614) );
INVx3_ASAP7_75t_SL g1129 ( .A(n_615), .Y(n_1129) );
XNOR2x1_ASAP7_75t_L g615 ( .A(n_616), .B(n_617), .Y(n_615) );
NOR2x1_ASAP7_75t_L g617 ( .A(n_618), .B(n_630), .Y(n_617) );
NAND3xp33_ASAP7_75t_L g618 ( .A(n_619), .B(n_622), .C(n_627), .Y(n_618) );
HB1xp67_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
INVx2_ASAP7_75t_L g813 ( .A(n_621), .Y(n_813) );
INVxp67_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
INVx2_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
INVx4_ASAP7_75t_L g753 ( .A(n_629), .Y(n_753) );
NAND4xp25_ASAP7_75t_SL g630 ( .A(n_631), .B(n_634), .C(n_637), .D(n_644), .Y(n_630) );
AND2x2_ASAP7_75t_L g637 ( .A(n_638), .B(n_641), .Y(n_637) );
NOR2xp33_ASAP7_75t_L g646 ( .A(n_647), .B(n_648), .Y(n_646) );
NOR2xp33_ASAP7_75t_L g698 ( .A(n_648), .B(n_699), .Y(n_698) );
INVx1_ASAP7_75t_L g756 ( .A(n_648), .Y(n_756) );
NOR2xp33_ASAP7_75t_L g1374 ( .A(n_648), .B(n_1375), .Y(n_1374) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_651), .B(n_671), .Y(n_650) );
NOR3xp33_ASAP7_75t_L g651 ( .A(n_652), .B(n_659), .C(n_666), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_653), .B(n_657), .Y(n_652) );
BUFx2_ASAP7_75t_L g1059 ( .A(n_654), .Y(n_1059) );
OAI22xp5_ASAP7_75t_L g659 ( .A1(n_660), .A2(n_661), .B1(n_663), .B2(n_664), .Y(n_659) );
INVx1_ASAP7_75t_L g1061 ( .A(n_661), .Y(n_1061) );
INVx2_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
OAI22xp5_ASAP7_75t_L g1269 ( .A1(n_664), .A2(n_1270), .B1(n_1271), .B2(n_1272), .Y(n_1269) );
INVx3_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
BUFx3_ASAP7_75t_L g772 ( .A(n_665), .Y(n_772) );
OAI21xp33_ASAP7_75t_L g666 ( .A1(n_667), .A2(n_668), .B(n_670), .Y(n_666) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
NOR2xp33_ASAP7_75t_SL g671 ( .A(n_672), .B(n_676), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_673), .B(n_674), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_677), .B(n_678), .Y(n_676) );
OAI22xp5_ASAP7_75t_L g682 ( .A1(n_683), .A2(n_684), .B1(n_761), .B2(n_818), .Y(n_682) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
XOR2x1_ASAP7_75t_L g685 ( .A(n_686), .B(n_739), .Y(n_685) );
XNOR2x1_ASAP7_75t_L g686 ( .A(n_687), .B(n_721), .Y(n_686) );
INVx2_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
XNOR2x2_ASAP7_75t_L g798 ( .A(n_688), .B(n_799), .Y(n_798) );
OAI21x1_ASAP7_75t_L g688 ( .A1(n_689), .A2(n_691), .B(n_715), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_689), .B(n_702), .Y(n_718) );
CKINVDCx5p33_ASAP7_75t_R g689 ( .A(n_690), .Y(n_689) );
NOR2xp67_ASAP7_75t_L g691 ( .A(n_692), .B(n_704), .Y(n_691) );
NAND3xp33_ASAP7_75t_L g692 ( .A(n_693), .B(n_700), .C(n_702), .Y(n_692) );
INVx1_ASAP7_75t_L g719 ( .A(n_693), .Y(n_719) );
AND2x2_ASAP7_75t_L g693 ( .A(n_694), .B(n_696), .Y(n_693) );
BUFx3_ASAP7_75t_L g771 ( .A(n_697), .Y(n_771) );
INVxp67_ASAP7_75t_L g717 ( .A(n_700), .Y(n_717) );
HB1xp67_ASAP7_75t_L g1064 ( .A(n_701), .Y(n_1064) );
BUFx3_ASAP7_75t_L g769 ( .A(n_703), .Y(n_769) );
INVx3_ASAP7_75t_L g1275 ( .A(n_703), .Y(n_1275) );
INVx1_ASAP7_75t_L g720 ( .A(n_704), .Y(n_720) );
NAND4xp25_ASAP7_75t_L g704 ( .A(n_705), .B(n_708), .C(n_711), .D(n_713), .Y(n_704) );
BUFx6f_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_716), .B(n_720), .Y(n_715) );
NOR3xp33_ASAP7_75t_L g716 ( .A(n_717), .B(n_718), .C(n_719), .Y(n_716) );
INVx2_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
XOR2x2_ASAP7_75t_L g722 ( .A(n_723), .B(n_738), .Y(n_722) );
NOR2x1_ASAP7_75t_L g723 ( .A(n_724), .B(n_729), .Y(n_723) );
NAND4xp25_ASAP7_75t_L g724 ( .A(n_725), .B(n_726), .C(n_727), .D(n_728), .Y(n_724) );
NAND4xp25_ASAP7_75t_L g729 ( .A(n_730), .B(n_732), .C(n_733), .D(n_736), .Y(n_729) );
INVx2_ASAP7_75t_L g1271 ( .A(n_734), .Y(n_1271) );
INVx3_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
BUFx3_ASAP7_75t_L g1293 ( .A(n_737), .Y(n_1293) );
NOR2x1_ASAP7_75t_L g740 ( .A(n_741), .B(n_750), .Y(n_740) );
NAND4xp25_ASAP7_75t_L g741 ( .A(n_742), .B(n_744), .C(n_746), .D(n_748), .Y(n_741) );
NAND3xp33_ASAP7_75t_L g750 ( .A(n_751), .B(n_757), .C(n_760), .Y(n_750) );
OAI21xp5_ASAP7_75t_L g752 ( .A1(n_753), .A2(n_754), .B(n_755), .Y(n_752) );
INVxp67_ASAP7_75t_SL g818 ( .A(n_761), .Y(n_818) );
INVx2_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
OAI22x1_ASAP7_75t_L g762 ( .A1(n_763), .A2(n_798), .B1(n_816), .B2(n_817), .Y(n_762) );
INVx1_ASAP7_75t_L g817 ( .A(n_763), .Y(n_817) );
AO22x2_ASAP7_75t_SL g763 ( .A1(n_764), .A2(n_782), .B1(n_783), .B2(n_796), .Y(n_763) );
NOR3xp33_ASAP7_75t_L g764 ( .A(n_765), .B(n_773), .C(n_782), .Y(n_764) );
INVxp67_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
NAND4xp75_ASAP7_75t_SL g796 ( .A(n_766), .B(n_784), .C(n_790), .D(n_797), .Y(n_796) );
AND2x2_ASAP7_75t_L g766 ( .A(n_767), .B(n_770), .Y(n_766) );
INVx1_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
HB1xp67_ASAP7_75t_L g776 ( .A(n_777), .Y(n_776) );
NOR2xp33_ASAP7_75t_R g778 ( .A(n_779), .B(n_780), .Y(n_778) );
NOR2xp33_ASAP7_75t_L g814 ( .A(n_780), .B(n_815), .Y(n_814) );
INVx2_ASAP7_75t_SL g780 ( .A(n_781), .Y(n_780) );
AND2x2_ASAP7_75t_L g783 ( .A(n_784), .B(n_790), .Y(n_783) );
AND2x2_ASAP7_75t_L g784 ( .A(n_785), .B(n_789), .Y(n_784) );
BUFx3_ASAP7_75t_L g786 ( .A(n_787), .Y(n_786) );
AND2x2_ASAP7_75t_L g790 ( .A(n_791), .B(n_794), .Y(n_790) );
INVx3_ASAP7_75t_L g816 ( .A(n_798), .Y(n_816) );
NAND4xp75_ASAP7_75t_L g800 ( .A(n_801), .B(n_804), .C(n_807), .D(n_810), .Y(n_800) );
AND2x2_ASAP7_75t_L g801 ( .A(n_802), .B(n_803), .Y(n_801) );
AND2x2_ASAP7_75t_L g804 ( .A(n_805), .B(n_806), .Y(n_804) );
AND2x2_ASAP7_75t_L g807 ( .A(n_808), .B(n_809), .Y(n_807) );
INVx2_ASAP7_75t_L g812 ( .A(n_813), .Y(n_812) );
NAND3xp33_ASAP7_75t_L g1392 ( .A(n_819), .B(n_1097), .C(n_1393), .Y(n_1392) );
INVx1_ASAP7_75t_L g819 ( .A(n_820), .Y(n_819) );
OAI221xp5_ASAP7_75t_L g820 ( .A1(n_821), .A2(n_1051), .B1(n_1053), .B2(n_1082), .C(n_1086), .Y(n_820) );
AND5x1_ASAP7_75t_L g821 ( .A(n_822), .B(n_1013), .C(n_1022), .D(n_1037), .E(n_1047), .Y(n_821) );
OAI33xp33_ASAP7_75t_L g822 ( .A1(n_823), .A2(n_916), .A3(n_942), .B1(n_966), .B2(n_981), .B3(n_990), .Y(n_822) );
NAND3xp33_ASAP7_75t_L g823 ( .A(n_824), .B(n_890), .C(n_901), .Y(n_823) );
AOI221xp5_ASAP7_75t_L g824 ( .A1(n_825), .A2(n_852), .B1(n_871), .B2(n_877), .C(n_880), .Y(n_824) );
INVx1_ASAP7_75t_L g1006 ( .A(n_825), .Y(n_1006) );
AND2x2_ASAP7_75t_L g825 ( .A(n_826), .B(n_839), .Y(n_825) );
AND2x2_ASAP7_75t_L g887 ( .A(n_826), .B(n_872), .Y(n_887) );
CKINVDCx6p67_ASAP7_75t_R g900 ( .A(n_826), .Y(n_900) );
AND2x2_ASAP7_75t_L g913 ( .A(n_826), .B(n_885), .Y(n_913) );
AND2x2_ASAP7_75t_L g922 ( .A(n_826), .B(n_895), .Y(n_922) );
AND2x2_ASAP7_75t_L g932 ( .A(n_826), .B(n_845), .Y(n_932) );
AND2x2_ASAP7_75t_L g954 ( .A(n_826), .B(n_926), .Y(n_954) );
AND2x2_ASAP7_75t_L g985 ( .A(n_826), .B(n_894), .Y(n_985) );
AND2x2_ASAP7_75t_L g993 ( .A(n_826), .B(n_946), .Y(n_993) );
NAND2xp5_ASAP7_75t_L g996 ( .A(n_826), .B(n_904), .Y(n_996) );
OAI332xp33_ASAP7_75t_L g998 ( .A1(n_826), .A2(n_879), .A3(n_900), .B1(n_999), .B2(n_1000), .B3(n_1001), .C1(n_1003), .C2(n_1004), .Y(n_998) );
AND2x2_ASAP7_75t_L g826 ( .A(n_827), .B(n_835), .Y(n_826) );
INVx3_ASAP7_75t_L g964 ( .A(n_828), .Y(n_964) );
AND2x4_ASAP7_75t_L g828 ( .A(n_829), .B(n_831), .Y(n_828) );
AND2x2_ASAP7_75t_L g836 ( .A(n_829), .B(n_837), .Y(n_836) );
AND2x4_ASAP7_75t_L g843 ( .A(n_829), .B(n_837), .Y(n_843) );
AND2x2_ASAP7_75t_L g851 ( .A(n_829), .B(n_837), .Y(n_851) );
AND2x4_ASAP7_75t_L g833 ( .A(n_831), .B(n_834), .Y(n_833) );
AND2x4_ASAP7_75t_L g849 ( .A(n_831), .B(n_834), .Y(n_849) );
AND2x2_ASAP7_75t_L g838 ( .A(n_834), .B(n_837), .Y(n_838) );
AND2x2_ASAP7_75t_L g844 ( .A(n_834), .B(n_837), .Y(n_844) );
AND2x4_ASAP7_75t_L g870 ( .A(n_834), .B(n_837), .Y(n_870) );
CKINVDCx5p33_ASAP7_75t_R g1094 ( .A(n_837), .Y(n_1094) );
NAND2xp5_ASAP7_75t_L g940 ( .A(n_839), .B(n_905), .Y(n_940) );
AND2x2_ASAP7_75t_L g959 ( .A(n_839), .B(n_899), .Y(n_959) );
NAND3xp33_ASAP7_75t_L g978 ( .A(n_839), .B(n_957), .C(n_979), .Y(n_978) );
AND2x2_ASAP7_75t_L g1030 ( .A(n_839), .B(n_887), .Y(n_1030) );
AND2x2_ASAP7_75t_L g1039 ( .A(n_839), .B(n_900), .Y(n_1039) );
INVx1_ASAP7_75t_L g839 ( .A(n_840), .Y(n_839) );
NOR2x1_ASAP7_75t_L g871 ( .A(n_840), .B(n_872), .Y(n_871) );
NOR2xp33_ASAP7_75t_L g1008 ( .A(n_840), .B(n_952), .Y(n_1008) );
OR2x2_ASAP7_75t_L g840 ( .A(n_841), .B(n_845), .Y(n_840) );
AND2x2_ASAP7_75t_L g885 ( .A(n_841), .B(n_845), .Y(n_885) );
AND2x2_ASAP7_75t_L g894 ( .A(n_841), .B(n_895), .Y(n_894) );
INVx1_ASAP7_75t_L g904 ( .A(n_841), .Y(n_904) );
AND2x2_ASAP7_75t_L g1036 ( .A(n_841), .B(n_900), .Y(n_1036) );
INVx1_ASAP7_75t_L g895 ( .A(n_845), .Y(n_895) );
AND2x2_ASAP7_75t_L g926 ( .A(n_845), .B(n_904), .Y(n_926) );
AND2x2_ASAP7_75t_L g845 ( .A(n_846), .B(n_850), .Y(n_845) );
INVx2_ASAP7_75t_SL g868 ( .A(n_849), .Y(n_868) );
NOR2xp33_ASAP7_75t_L g852 ( .A(n_853), .B(n_861), .Y(n_852) );
NAND2xp5_ASAP7_75t_L g892 ( .A(n_853), .B(n_893), .Y(n_892) );
INVx1_ASAP7_75t_L g853 ( .A(n_854), .Y(n_853) );
INVx1_ASAP7_75t_L g854 ( .A(n_855), .Y(n_854) );
HB1xp67_ASAP7_75t_L g937 ( .A(n_855), .Y(n_937) );
NOR2xp33_ASAP7_75t_L g1046 ( .A(n_855), .B(n_952), .Y(n_1046) );
INVx1_ASAP7_75t_L g855 ( .A(n_856), .Y(n_855) );
INVx1_ASAP7_75t_L g911 ( .A(n_856), .Y(n_911) );
INVx1_ASAP7_75t_L g856 ( .A(n_857), .Y(n_856) );
INVx2_ASAP7_75t_L g878 ( .A(n_857), .Y(n_878) );
OR2x2_ASAP7_75t_L g935 ( .A(n_857), .B(n_889), .Y(n_935) );
INVx4_ASAP7_75t_L g857 ( .A(n_858), .Y(n_857) );
OR2x2_ASAP7_75t_L g907 ( .A(n_858), .B(n_889), .Y(n_907) );
AND2x2_ASAP7_75t_L g944 ( .A(n_858), .B(n_889), .Y(n_944) );
NAND2xp5_ASAP7_75t_L g951 ( .A(n_858), .B(n_952), .Y(n_951) );
OR2x2_ASAP7_75t_L g973 ( .A(n_858), .B(n_862), .Y(n_973) );
NOR2xp33_ASAP7_75t_L g979 ( .A(n_858), .B(n_952), .Y(n_979) );
AND2x2_ASAP7_75t_L g858 ( .A(n_859), .B(n_860), .Y(n_858) );
AOI222xp33_ASAP7_75t_L g927 ( .A1(n_861), .A2(n_928), .B1(n_933), .B2(n_936), .C1(n_937), .C2(n_938), .Y(n_927) );
AOI211xp5_ASAP7_75t_L g976 ( .A1(n_861), .A2(n_920), .B(n_977), .C(n_980), .Y(n_976) );
AND2x2_ASAP7_75t_L g997 ( .A(n_861), .B(n_937), .Y(n_997) );
AND2x2_ASAP7_75t_L g861 ( .A(n_862), .B(n_865), .Y(n_861) );
INVx2_ASAP7_75t_L g889 ( .A(n_862), .Y(n_889) );
NAND2xp5_ASAP7_75t_L g862 ( .A(n_863), .B(n_864), .Y(n_862) );
INVx4_ASAP7_75t_L g879 ( .A(n_865), .Y(n_879) );
INVx1_ASAP7_75t_L g915 ( .A(n_865), .Y(n_915) );
AND2x2_ASAP7_75t_L g958 ( .A(n_865), .B(n_934), .Y(n_958) );
AND2x2_ASAP7_75t_L g986 ( .A(n_865), .B(n_878), .Y(n_986) );
NAND2xp5_ASAP7_75t_L g1009 ( .A(n_865), .B(n_911), .Y(n_1009) );
AND2x2_ASAP7_75t_L g865 ( .A(n_866), .B(n_869), .Y(n_865) );
INVx2_ASAP7_75t_L g867 ( .A(n_868), .Y(n_867) );
BUFx2_ASAP7_75t_L g1052 ( .A(n_870), .Y(n_1052) );
NAND2xp5_ASAP7_75t_L g975 ( .A(n_871), .B(n_900), .Y(n_975) );
AND2x2_ASAP7_75t_L g923 ( .A(n_872), .B(n_924), .Y(n_923) );
NAND2xp5_ASAP7_75t_L g999 ( .A(n_872), .B(n_906), .Y(n_999) );
NAND2xp5_ASAP7_75t_L g1004 ( .A(n_872), .B(n_926), .Y(n_1004) );
INVx3_ASAP7_75t_L g872 ( .A(n_873), .Y(n_872) );
AND2x2_ASAP7_75t_L g905 ( .A(n_873), .B(n_906), .Y(n_905) );
AND2x2_ASAP7_75t_L g946 ( .A(n_873), .B(n_885), .Y(n_946) );
INVx3_ASAP7_75t_L g873 ( .A(n_874), .Y(n_873) );
INVx2_ASAP7_75t_L g883 ( .A(n_874), .Y(n_883) );
AND2x2_ASAP7_75t_L g899 ( .A(n_874), .B(n_900), .Y(n_899) );
NOR2xp33_ASAP7_75t_L g938 ( .A(n_874), .B(n_939), .Y(n_938) );
INVx2_ASAP7_75t_L g952 ( .A(n_874), .Y(n_952) );
NAND2xp5_ASAP7_75t_L g1000 ( .A(n_874), .B(n_879), .Y(n_1000) );
NAND2xp5_ASAP7_75t_L g1012 ( .A(n_874), .B(n_944), .Y(n_1012) );
NAND2xp5_ASAP7_75t_L g1028 ( .A(n_874), .B(n_922), .Y(n_1028) );
AND2x2_ASAP7_75t_L g874 ( .A(n_875), .B(n_876), .Y(n_874) );
INVx1_ASAP7_75t_L g1003 ( .A(n_877), .Y(n_1003) );
AND2x2_ASAP7_75t_L g877 ( .A(n_878), .B(n_879), .Y(n_877) );
O2A1O1Ixp33_ASAP7_75t_L g880 ( .A1(n_878), .A2(n_881), .B(n_886), .C(n_888), .Y(n_880) );
AND2x2_ASAP7_75t_L g893 ( .A(n_879), .B(n_889), .Y(n_893) );
NAND2xp5_ASAP7_75t_L g897 ( .A(n_879), .B(n_898), .Y(n_897) );
OR2x2_ASAP7_75t_L g956 ( .A(n_879), .B(n_957), .Y(n_956) );
NAND2xp5_ASAP7_75t_L g967 ( .A(n_879), .B(n_906), .Y(n_967) );
A2O1A1Ixp33_ASAP7_75t_L g1025 ( .A1(n_879), .A2(n_1026), .B(n_1029), .C(n_1031), .Y(n_1025) );
NOR2xp33_ASAP7_75t_L g1034 ( .A(n_879), .B(n_973), .Y(n_1034) );
A2O1A1Ixp33_ASAP7_75t_L g1047 ( .A1(n_879), .A2(n_932), .B(n_1048), .C(n_1049), .Y(n_1047) );
INVx1_ASAP7_75t_L g881 ( .A(n_882), .Y(n_881) );
NAND2xp5_ASAP7_75t_L g909 ( .A(n_882), .B(n_910), .Y(n_909) );
NOR2xp33_ASAP7_75t_L g882 ( .A(n_883), .B(n_884), .Y(n_882) );
A2O1A1Ixp33_ASAP7_75t_L g917 ( .A1(n_883), .A2(n_893), .B(n_918), .C(n_923), .Y(n_917) );
AND2x2_ASAP7_75t_L g933 ( .A(n_883), .B(n_934), .Y(n_933) );
NAND2xp5_ASAP7_75t_L g968 ( .A(n_883), .B(n_969), .Y(n_968) );
AND2x2_ASAP7_75t_L g984 ( .A(n_883), .B(n_985), .Y(n_984) );
NOR2xp33_ASAP7_75t_L g1016 ( .A(n_883), .B(n_1017), .Y(n_1016) );
O2A1O1Ixp33_ASAP7_75t_SL g1020 ( .A1(n_883), .A2(n_892), .B(n_939), .C(n_1021), .Y(n_1020) );
INVx1_ASAP7_75t_L g884 ( .A(n_885), .Y(n_884) );
NAND2xp5_ASAP7_75t_L g886 ( .A(n_885), .B(n_887), .Y(n_886) );
AND2x2_ASAP7_75t_L g920 ( .A(n_885), .B(n_900), .Y(n_920) );
NAND2xp5_ASAP7_75t_L g1042 ( .A(n_885), .B(n_899), .Y(n_1042) );
INVx1_ASAP7_75t_L g936 ( .A(n_886), .Y(n_936) );
INVx3_ASAP7_75t_SL g914 ( .A(n_888), .Y(n_914) );
INVx2_ASAP7_75t_L g888 ( .A(n_889), .Y(n_888) );
INVxp67_ASAP7_75t_L g957 ( .A(n_889), .Y(n_957) );
AOI21xp5_ASAP7_75t_L g890 ( .A1(n_891), .A2(n_894), .B(n_896), .Y(n_890) );
INVx1_ASAP7_75t_L g891 ( .A(n_892), .Y(n_891) );
INVx1_ASAP7_75t_L g982 ( .A(n_893), .Y(n_982) );
AND2x2_ASAP7_75t_L g898 ( .A(n_894), .B(n_899), .Y(n_898) );
AND2x2_ASAP7_75t_L g930 ( .A(n_894), .B(n_900), .Y(n_930) );
INVx1_ASAP7_75t_L g939 ( .A(n_894), .Y(n_939) );
NAND2xp5_ASAP7_75t_L g970 ( .A(n_895), .B(n_900), .Y(n_970) );
AOI211xp5_ASAP7_75t_L g1013 ( .A1(n_896), .A2(n_934), .B(n_1014), .C(n_1020), .Y(n_1013) );
INVx1_ASAP7_75t_L g896 ( .A(n_897), .Y(n_896) );
NAND2xp5_ASAP7_75t_L g903 ( .A(n_900), .B(n_904), .Y(n_903) );
NAND2xp5_ASAP7_75t_L g925 ( .A(n_900), .B(n_926), .Y(n_925) );
NAND2xp5_ASAP7_75t_L g945 ( .A(n_900), .B(n_946), .Y(n_945) );
NAND2xp5_ASAP7_75t_L g1033 ( .A(n_900), .B(n_952), .Y(n_1033) );
A2O1A1Ixp33_ASAP7_75t_L g901 ( .A1(n_902), .A2(n_905), .B(n_908), .C(n_915), .Y(n_901) );
INVx1_ASAP7_75t_L g902 ( .A(n_903), .Y(n_902) );
NOR2xp33_ASAP7_75t_L g1011 ( .A(n_903), .B(n_1012), .Y(n_1011) );
OAI22xp33_ASAP7_75t_L g1040 ( .A1(n_903), .A2(n_1041), .B1(n_1042), .B2(n_1043), .Y(n_1040) );
NAND2xp5_ASAP7_75t_L g941 ( .A(n_905), .B(n_922), .Y(n_941) );
INVx1_ASAP7_75t_L g906 ( .A(n_907), .Y(n_906) );
AOI21xp33_ASAP7_75t_L g908 ( .A1(n_909), .A2(n_912), .B(n_914), .Y(n_908) );
INVxp67_ASAP7_75t_SL g1023 ( .A(n_909), .Y(n_1023) );
INVx2_ASAP7_75t_L g910 ( .A(n_911), .Y(n_910) );
INVx1_ASAP7_75t_L g912 ( .A(n_913), .Y(n_912) );
NAND2xp5_ASAP7_75t_L g1050 ( .A(n_913), .B(n_934), .Y(n_1050) );
INVx1_ASAP7_75t_L g991 ( .A(n_914), .Y(n_991) );
NAND2xp5_ASAP7_75t_L g1026 ( .A(n_914), .B(n_1027), .Y(n_1026) );
NOR2xp33_ASAP7_75t_L g948 ( .A(n_915), .B(n_949), .Y(n_948) );
NAND4xp25_ASAP7_75t_SL g916 ( .A(n_917), .B(n_927), .C(n_940), .D(n_941), .Y(n_916) );
NAND2xp5_ASAP7_75t_SL g918 ( .A(n_919), .B(n_921), .Y(n_918) );
INVx1_ASAP7_75t_L g919 ( .A(n_920), .Y(n_919) );
INVx1_ASAP7_75t_L g921 ( .A(n_922), .Y(n_921) );
AOI221xp5_ASAP7_75t_L g1037 ( .A1(n_923), .A2(n_944), .B1(n_1038), .B2(n_1039), .C(n_1040), .Y(n_1037) );
INVx1_ASAP7_75t_L g924 ( .A(n_925), .Y(n_924) );
NOR2xp33_ASAP7_75t_L g988 ( .A(n_925), .B(n_989), .Y(n_988) );
INVx1_ASAP7_75t_L g1002 ( .A(n_926), .Y(n_1002) );
NAND2xp5_ASAP7_75t_SL g928 ( .A(n_929), .B(n_931), .Y(n_928) );
INVx1_ASAP7_75t_L g929 ( .A(n_930), .Y(n_929) );
NAND2xp5_ASAP7_75t_L g949 ( .A(n_930), .B(n_950), .Y(n_949) );
INVx1_ASAP7_75t_L g931 ( .A(n_932), .Y(n_931) );
INVx1_ASAP7_75t_L g989 ( .A(n_933), .Y(n_989) );
INVx1_ASAP7_75t_L g934 ( .A(n_935), .Y(n_934) );
NAND2xp5_ASAP7_75t_L g1029 ( .A(n_937), .B(n_1030), .Y(n_1029) );
INVx1_ASAP7_75t_L g1018 ( .A(n_938), .Y(n_1018) );
AND2x2_ASAP7_75t_L g1001 ( .A(n_939), .B(n_1002), .Y(n_1001) );
OAI211xp5_ASAP7_75t_L g942 ( .A1(n_943), .A2(n_945), .B(n_947), .C(n_953), .Y(n_942) );
INVx1_ASAP7_75t_L g943 ( .A(n_944), .Y(n_943) );
OAI211xp5_ASAP7_75t_L g1031 ( .A1(n_946), .A2(n_1032), .B(n_1034), .C(n_1035), .Y(n_1031) );
INVx1_ASAP7_75t_L g947 ( .A(n_948), .Y(n_947) );
OAI211xp5_ASAP7_75t_L g981 ( .A1(n_949), .A2(n_982), .B(n_983), .C(n_987), .Y(n_981) );
INVx1_ASAP7_75t_L g950 ( .A(n_951), .Y(n_950) );
NAND2xp33_ASAP7_75t_L g955 ( .A(n_951), .B(n_956), .Y(n_955) );
AOI221xp5_ASAP7_75t_L g953 ( .A1(n_954), .A2(n_955), .B1(n_958), .B2(n_959), .C(n_960), .Y(n_953) );
INVx1_ASAP7_75t_L g1017 ( .A(n_954), .Y(n_1017) );
INVx1_ASAP7_75t_L g1024 ( .A(n_956), .Y(n_1024) );
INVx1_ASAP7_75t_L g1019 ( .A(n_958), .Y(n_1019) );
INVx2_ASAP7_75t_L g980 ( .A(n_960), .Y(n_980) );
CKINVDCx5p33_ASAP7_75t_R g960 ( .A(n_961), .Y(n_960) );
AND2x2_ASAP7_75t_L g961 ( .A(n_962), .B(n_965), .Y(n_961) );
INVx1_ASAP7_75t_L g963 ( .A(n_964), .Y(n_963) );
OAI211xp5_ASAP7_75t_L g966 ( .A1(n_967), .A2(n_968), .B(n_971), .C(n_976), .Y(n_966) );
INVx1_ASAP7_75t_L g1038 ( .A(n_967), .Y(n_1038) );
INVx1_ASAP7_75t_L g969 ( .A(n_970), .Y(n_969) );
NAND2xp5_ASAP7_75t_L g971 ( .A(n_972), .B(n_974), .Y(n_971) );
INVx1_ASAP7_75t_L g972 ( .A(n_973), .Y(n_972) );
OAI21xp5_ASAP7_75t_SL g983 ( .A1(n_974), .A2(n_984), .B(n_986), .Y(n_983) );
O2A1O1Ixp33_ASAP7_75t_L g1022 ( .A1(n_974), .A2(n_1023), .B(n_1024), .C(n_1025), .Y(n_1022) );
INVx1_ASAP7_75t_L g974 ( .A(n_975), .Y(n_974) );
INVxp67_ASAP7_75t_L g977 ( .A(n_978), .Y(n_977) );
NOR2xp33_ASAP7_75t_L g1044 ( .A(n_982), .B(n_1045), .Y(n_1044) );
INVx1_ASAP7_75t_L g1021 ( .A(n_985), .Y(n_1021) );
INVxp67_ASAP7_75t_SL g987 ( .A(n_988), .Y(n_987) );
OAI211xp5_ASAP7_75t_L g990 ( .A1(n_991), .A2(n_992), .B(n_994), .C(n_1010), .Y(n_990) );
INVx1_ASAP7_75t_L g992 ( .A(n_993), .Y(n_992) );
AOI211xp5_ASAP7_75t_SL g994 ( .A1(n_995), .A2(n_997), .B(n_998), .C(n_1005), .Y(n_994) );
INVx1_ASAP7_75t_L g995 ( .A(n_996), .Y(n_995) );
INVx1_ASAP7_75t_L g1041 ( .A(n_997), .Y(n_1041) );
INVx1_ASAP7_75t_L g1048 ( .A(n_999), .Y(n_1048) );
AOI21xp33_ASAP7_75t_SL g1005 ( .A1(n_1006), .A2(n_1007), .B(n_1009), .Y(n_1005) );
INVxp33_ASAP7_75t_SL g1007 ( .A(n_1008), .Y(n_1007) );
INVxp67_ASAP7_75t_SL g1010 ( .A(n_1011), .Y(n_1010) );
AOI21xp33_ASAP7_75t_L g1014 ( .A1(n_1015), .A2(n_1018), .B(n_1019), .Y(n_1014) );
INVxp33_ASAP7_75t_L g1015 ( .A(n_1016), .Y(n_1015) );
INVxp67_ASAP7_75t_SL g1027 ( .A(n_1028), .Y(n_1027) );
INVxp67_ASAP7_75t_SL g1032 ( .A(n_1033), .Y(n_1032) );
INVx1_ASAP7_75t_L g1035 ( .A(n_1036), .Y(n_1035) );
INVxp33_ASAP7_75t_L g1043 ( .A(n_1044), .Y(n_1043) );
INVxp33_ASAP7_75t_L g1045 ( .A(n_1046), .Y(n_1045) );
INVxp67_ASAP7_75t_SL g1049 ( .A(n_1050), .Y(n_1049) );
CKINVDCx5p33_ASAP7_75t_R g1051 ( .A(n_1052), .Y(n_1051) );
BUFx3_ASAP7_75t_L g1053 ( .A(n_1054), .Y(n_1053) );
BUFx2_ASAP7_75t_L g1089 ( .A(n_1055), .Y(n_1089) );
OR2x2_ASAP7_75t_L g1055 ( .A(n_1056), .B(n_1067), .Y(n_1055) );
NOR2xp33_ASAP7_75t_L g1080 ( .A(n_1056), .B(n_1067), .Y(n_1080) );
NAND2xp5_ASAP7_75t_L g1056 ( .A(n_1057), .B(n_1063), .Y(n_1056) );
AND2x2_ASAP7_75t_L g1057 ( .A(n_1058), .B(n_1060), .Y(n_1057) );
NAND2x1p5_ASAP7_75t_L g1067 ( .A(n_1068), .B(n_1075), .Y(n_1067) );
AND2x2_ASAP7_75t_L g1068 ( .A(n_1069), .B(n_1072), .Y(n_1068) );
INVx1_ASAP7_75t_L g1070 ( .A(n_1071), .Y(n_1070) );
AND2x2_ASAP7_75t_L g1075 ( .A(n_1076), .B(n_1079), .Y(n_1075) );
BUFx2_ASAP7_75t_L g1077 ( .A(n_1078), .Y(n_1077) );
CKINVDCx20_ASAP7_75t_R g1082 ( .A(n_1083), .Y(n_1082) );
INVx1_ASAP7_75t_L g1087 ( .A(n_1088), .Y(n_1087) );
BUFx3_ASAP7_75t_L g1090 ( .A(n_1091), .Y(n_1090) );
BUFx2_ASAP7_75t_L g1092 ( .A(n_1093), .Y(n_1092) );
INVx1_ASAP7_75t_L g1095 ( .A(n_1096), .Y(n_1095) );
NAND2xp5_ASAP7_75t_L g1096 ( .A(n_1097), .B(n_1391), .Y(n_1096) );
XNOR2xp5_ASAP7_75t_L g1097 ( .A(n_1098), .B(n_1203), .Y(n_1097) );
AOI22xp5_ASAP7_75t_L g1098 ( .A1(n_1099), .A2(n_1154), .B1(n_1155), .B2(n_1202), .Y(n_1098) );
INVx1_ASAP7_75t_L g1202 ( .A(n_1099), .Y(n_1202) );
AOI22xp5_ASAP7_75t_L g1099 ( .A1(n_1100), .A2(n_1131), .B1(n_1152), .B2(n_1153), .Y(n_1099) );
INVx2_ASAP7_75t_SL g1153 ( .A(n_1100), .Y(n_1153) );
OA22x2_ASAP7_75t_L g1100 ( .A1(n_1101), .A2(n_1128), .B1(n_1129), .B2(n_1130), .Y(n_1100) );
INVx2_ASAP7_75t_L g1130 ( .A(n_1101), .Y(n_1130) );
AND4x1_ASAP7_75t_L g1127 ( .A(n_1103), .B(n_1109), .C(n_1118), .D(n_1123), .Y(n_1127) );
AND2x2_ASAP7_75t_L g1103 ( .A(n_1104), .B(n_1107), .Y(n_1103) );
INVx1_ASAP7_75t_L g1110 ( .A(n_1111), .Y(n_1110) );
OAI22xp5_ASAP7_75t_L g1112 ( .A1(n_1113), .A2(n_1114), .B1(n_1115), .B2(n_1116), .Y(n_1112) );
NOR2xp33_ASAP7_75t_L g1267 ( .A(n_1116), .B(n_1268), .Y(n_1267) );
NAND2xp5_ASAP7_75t_L g1117 ( .A(n_1118), .B(n_1123), .Y(n_1117) );
AND2x2_ASAP7_75t_L g1118 ( .A(n_1119), .B(n_1122), .Y(n_1118) );
AND2x2_ASAP7_75t_L g1123 ( .A(n_1124), .B(n_1125), .Y(n_1123) );
INVx2_ASAP7_75t_SL g1128 ( .A(n_1129), .Y(n_1128) );
INVx2_ASAP7_75t_L g1131 ( .A(n_1132), .Y(n_1131) );
BUFx2_ASAP7_75t_SL g1152 ( .A(n_1132), .Y(n_1152) );
NOR2x1_ASAP7_75t_L g1133 ( .A(n_1134), .B(n_1143), .Y(n_1133) );
NAND3xp33_ASAP7_75t_L g1134 ( .A(n_1135), .B(n_1140), .C(n_1141), .Y(n_1134) );
INVx2_ASAP7_75t_SL g1136 ( .A(n_1137), .Y(n_1136) );
INVx2_ASAP7_75t_L g1137 ( .A(n_1138), .Y(n_1137) );
NAND4xp25_ASAP7_75t_SL g1143 ( .A(n_1144), .B(n_1145), .C(n_1147), .D(n_1148), .Y(n_1143) );
BUFx2_ASAP7_75t_SL g1150 ( .A(n_1151), .Y(n_1150) );
INVx1_ASAP7_75t_L g1154 ( .A(n_1155), .Y(n_1154) );
BUFx2_ASAP7_75t_L g1155 ( .A(n_1156), .Y(n_1155) );
INVx1_ASAP7_75t_L g1156 ( .A(n_1157), .Y(n_1156) );
OA22x2_ASAP7_75t_L g1157 ( .A1(n_1158), .A2(n_1159), .B1(n_1186), .B2(n_1187), .Y(n_1157) );
INVx2_ASAP7_75t_L g1158 ( .A(n_1159), .Y(n_1158) );
OAI21x1_ASAP7_75t_L g1159 ( .A1(n_1160), .A2(n_1161), .B(n_1183), .Y(n_1159) );
NOR4xp75_ASAP7_75t_L g1161 ( .A(n_1162), .B(n_1169), .C(n_1173), .D(n_1177), .Y(n_1161) );
INVx3_ASAP7_75t_L g1162 ( .A(n_1163), .Y(n_1162) );
NAND4xp75_ASAP7_75t_L g1183 ( .A(n_1163), .B(n_1170), .C(n_1174), .D(n_1184), .Y(n_1183) );
AND2x2_ASAP7_75t_L g1163 ( .A(n_1164), .B(n_1165), .Y(n_1163) );
INVx2_ASAP7_75t_L g1169 ( .A(n_1170), .Y(n_1169) );
AND2x2_ASAP7_75t_L g1170 ( .A(n_1171), .B(n_1172), .Y(n_1170) );
INVx2_ASAP7_75t_SL g1173 ( .A(n_1174), .Y(n_1173) );
AND2x2_ASAP7_75t_L g1174 ( .A(n_1175), .B(n_1176), .Y(n_1174) );
INVx1_ASAP7_75t_L g1177 ( .A(n_1178), .Y(n_1177) );
AND2x2_ASAP7_75t_L g1184 ( .A(n_1178), .B(n_1185), .Y(n_1184) );
AND2x2_ASAP7_75t_L g1178 ( .A(n_1179), .B(n_1181), .Y(n_1178) );
INVx1_ASAP7_75t_L g1186 ( .A(n_1187), .Y(n_1186) );
NAND2xp5_ASAP7_75t_L g1188 ( .A(n_1189), .B(n_1196), .Y(n_1188) );
AND4x1_ASAP7_75t_L g1189 ( .A(n_1190), .B(n_1191), .C(n_1192), .D(n_1193), .Y(n_1189) );
NOR4xp25_ASAP7_75t_L g1196 ( .A(n_1197), .B(n_1199), .C(n_1200), .D(n_1201), .Y(n_1196) );
INVx1_ASAP7_75t_L g1197 ( .A(n_1198), .Y(n_1197) );
AOI22xp5_ASAP7_75t_L g1203 ( .A1(n_1204), .A2(n_1298), .B1(n_1299), .B2(n_1390), .Y(n_1203) );
INVx2_ASAP7_75t_L g1390 ( .A(n_1204), .Y(n_1390) );
AOI22xp5_ASAP7_75t_L g1204 ( .A1(n_1205), .A2(n_1206), .B1(n_1277), .B2(n_1297), .Y(n_1204) );
INVx2_ASAP7_75t_SL g1205 ( .A(n_1206), .Y(n_1205) );
AOI22x1_ASAP7_75t_L g1206 ( .A1(n_1207), .A2(n_1208), .B1(n_1243), .B2(n_1244), .Y(n_1206) );
INVx2_ASAP7_75t_L g1207 ( .A(n_1208), .Y(n_1207) );
AO22x2_ASAP7_75t_L g1208 ( .A1(n_1209), .A2(n_1210), .B1(n_1225), .B2(n_1242), .Y(n_1208) );
INVx2_ASAP7_75t_L g1209 ( .A(n_1210), .Y(n_1209) );
XNOR2x1_ASAP7_75t_L g1210 ( .A(n_1211), .B(n_1212), .Y(n_1210) );
NOR2x1_ASAP7_75t_L g1212 ( .A(n_1213), .B(n_1218), .Y(n_1212) );
NAND4xp25_ASAP7_75t_L g1213 ( .A(n_1214), .B(n_1215), .C(n_1216), .D(n_1217), .Y(n_1213) );
NAND4xp25_ASAP7_75t_L g1218 ( .A(n_1219), .B(n_1220), .C(n_1221), .D(n_1222), .Y(n_1218) );
INVx2_ASAP7_75t_L g1242 ( .A(n_1225), .Y(n_1242) );
AND3x1_ASAP7_75t_L g1226 ( .A(n_1227), .B(n_1231), .C(n_1238), .Y(n_1226) );
AND2x2_ASAP7_75t_L g1227 ( .A(n_1228), .B(n_1229), .Y(n_1227) );
AND2x2_ASAP7_75t_L g1231 ( .A(n_1232), .B(n_1235), .Y(n_1231) );
AND2x2_ASAP7_75t_L g1235 ( .A(n_1236), .B(n_1237), .Y(n_1235) );
AND2x2_ASAP7_75t_L g1238 ( .A(n_1239), .B(n_1240), .Y(n_1238) );
INVx1_ASAP7_75t_L g1243 ( .A(n_1244), .Y(n_1243) );
NAND2xp5_ASAP7_75t_L g1245 ( .A(n_1246), .B(n_1261), .Y(n_1245) );
NOR3xp33_ASAP7_75t_L g1246 ( .A(n_1247), .B(n_1254), .C(n_1257), .Y(n_1246) );
OAI22xp5_ASAP7_75t_L g1247 ( .A1(n_1248), .A2(n_1250), .B1(n_1251), .B2(n_1253), .Y(n_1247) );
INVx1_ASAP7_75t_L g1248 ( .A(n_1249), .Y(n_1248) );
INVx1_ASAP7_75t_L g1251 ( .A(n_1252), .Y(n_1251) );
NAND2xp5_ASAP7_75t_SL g1254 ( .A(n_1255), .B(n_1256), .Y(n_1254) );
NOR3xp33_ASAP7_75t_L g1261 ( .A(n_1262), .B(n_1269), .C(n_1273), .Y(n_1261) );
NAND2xp5_ASAP7_75t_SL g1262 ( .A(n_1263), .B(n_1266), .Y(n_1262) );
BUFx3_ASAP7_75t_L g1264 ( .A(n_1265), .Y(n_1264) );
OAI21xp5_ASAP7_75t_L g1273 ( .A1(n_1274), .A2(n_1275), .B(n_1276), .Y(n_1273) );
OAI21xp33_ASAP7_75t_L g1320 ( .A1(n_1275), .A2(n_1321), .B(n_1322), .Y(n_1320) );
INVx1_ASAP7_75t_L g1297 ( .A(n_1277), .Y(n_1297) );
BUFx2_ASAP7_75t_SL g1277 ( .A(n_1278), .Y(n_1277) );
INVx1_ASAP7_75t_L g1278 ( .A(n_1279), .Y(n_1278) );
INVx2_ASAP7_75t_L g1279 ( .A(n_1280), .Y(n_1279) );
INVx2_ASAP7_75t_L g1281 ( .A(n_1282), .Y(n_1281) );
NAND4xp75_ASAP7_75t_L g1282 ( .A(n_1283), .B(n_1286), .C(n_1289), .D(n_1292), .Y(n_1282) );
AND2x2_ASAP7_75t_L g1283 ( .A(n_1284), .B(n_1285), .Y(n_1283) );
AND2x2_ASAP7_75t_L g1286 ( .A(n_1287), .B(n_1288), .Y(n_1286) );
AND2x2_ASAP7_75t_L g1289 ( .A(n_1290), .B(n_1291), .Y(n_1289) );
INVx1_ASAP7_75t_L g1298 ( .A(n_1299), .Y(n_1298) );
AO22x2_ASAP7_75t_L g1299 ( .A1(n_1300), .A2(n_1324), .B1(n_1387), .B2(n_1389), .Y(n_1299) );
INVx1_ASAP7_75t_L g1300 ( .A(n_1301), .Y(n_1300) );
INVx2_ASAP7_75t_L g1388 ( .A(n_1301), .Y(n_1388) );
XOR2x1_ASAP7_75t_L g1301 ( .A(n_1302), .B(n_1323), .Y(n_1301) );
AND2x2_ASAP7_75t_L g1302 ( .A(n_1303), .B(n_1308), .Y(n_1302) );
AND4x1_ASAP7_75t_L g1303 ( .A(n_1304), .B(n_1305), .C(n_1306), .D(n_1307), .Y(n_1303) );
NOR3xp33_ASAP7_75t_L g1308 ( .A(n_1309), .B(n_1317), .C(n_1320), .Y(n_1308) );
NAND2xp5_ASAP7_75t_SL g1309 ( .A(n_1310), .B(n_1311), .Y(n_1309) );
NOR2xp33_ASAP7_75t_L g1313 ( .A(n_1314), .B(n_1315), .Y(n_1313) );
INVx1_ASAP7_75t_L g1315 ( .A(n_1316), .Y(n_1315) );
INVx2_ASAP7_75t_L g1389 ( .A(n_1324), .Y(n_1389) );
AO22x2_ASAP7_75t_L g1324 ( .A1(n_1325), .A2(n_1326), .B1(n_1367), .B2(n_1385), .Y(n_1324) );
INVx1_ASAP7_75t_L g1325 ( .A(n_1326), .Y(n_1325) );
OAI21xp5_ASAP7_75t_L g1326 ( .A1(n_1327), .A2(n_1345), .B(n_1365), .Y(n_1326) );
INVxp67_ASAP7_75t_L g1327 ( .A(n_1328), .Y(n_1327) );
INVx1_ASAP7_75t_L g1366 ( .A(n_1328), .Y(n_1366) );
OAI21x1_ASAP7_75t_L g1328 ( .A1(n_1329), .A2(n_1330), .B(n_1342), .Y(n_1328) );
NAND3xp33_ASAP7_75t_SL g1342 ( .A(n_1329), .B(n_1343), .C(n_1344), .Y(n_1342) );
INVx1_ASAP7_75t_L g1330 ( .A(n_1331), .Y(n_1330) );
OR2x2_ASAP7_75t_L g1331 ( .A(n_1332), .B(n_1337), .Y(n_1331) );
INVx1_ASAP7_75t_L g1344 ( .A(n_1332), .Y(n_1344) );
NAND4xp25_ASAP7_75t_L g1332 ( .A(n_1333), .B(n_1334), .C(n_1335), .D(n_1336), .Y(n_1332) );
INVxp67_ASAP7_75t_L g1343 ( .A(n_1337), .Y(n_1343) );
NAND4xp25_ASAP7_75t_L g1337 ( .A(n_1338), .B(n_1339), .C(n_1340), .D(n_1341), .Y(n_1337) );
NAND2xp5_ASAP7_75t_L g1365 ( .A(n_1345), .B(n_1366), .Y(n_1365) );
NOR2xp33_ASAP7_75t_L g1346 ( .A(n_1347), .B(n_1356), .Y(n_1346) );
INVxp67_ASAP7_75t_L g1362 ( .A(n_1347), .Y(n_1362) );
NAND4xp25_ASAP7_75t_L g1347 ( .A(n_1348), .B(n_1349), .C(n_1351), .D(n_1354), .Y(n_1347) );
NOR2xp33_ASAP7_75t_L g1363 ( .A(n_1356), .B(n_1364), .Y(n_1363) );
NAND4xp25_ASAP7_75t_L g1356 ( .A(n_1357), .B(n_1358), .C(n_1359), .D(n_1360), .Y(n_1356) );
NAND2xp5_ASAP7_75t_L g1361 ( .A(n_1362), .B(n_1363), .Y(n_1361) );
INVxp67_ASAP7_75t_SL g1367 ( .A(n_1368), .Y(n_1367) );
INVx1_ASAP7_75t_L g1386 ( .A(n_1368), .Y(n_1386) );
XNOR2x1_ASAP7_75t_L g1368 ( .A(n_1369), .B(n_1370), .Y(n_1368) );
OR2x2_ASAP7_75t_L g1370 ( .A(n_1371), .B(n_1379), .Y(n_1370) );
NAND3xp33_ASAP7_75t_L g1371 ( .A(n_1372), .B(n_1376), .C(n_1377), .Y(n_1371) );
NAND4xp25_ASAP7_75t_SL g1379 ( .A(n_1380), .B(n_1381), .C(n_1382), .D(n_1384), .Y(n_1379) );
INVx1_ASAP7_75t_L g1385 ( .A(n_1386), .Y(n_1385) );
INVx1_ASAP7_75t_L g1387 ( .A(n_1388), .Y(n_1387) );
endmodule