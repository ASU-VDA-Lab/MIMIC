module fake_aes_2930_n_19 (n_3, n_1, n_2, n_0, n_19);
input n_3;
input n_1;
input n_2;
input n_0;
output n_19;
wire n_5;
wire n_8;
wire n_11;
wire n_16;
wire n_13;
wire n_18;
wire n_12;
wire n_9;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_6;
wire n_4;
wire n_7;
INVx3_ASAP7_75t_L g4 ( .A(n_1), .Y(n_4) );
INVx1_ASAP7_75t_L g5 ( .A(n_2), .Y(n_5) );
BUFx3_ASAP7_75t_L g6 ( .A(n_4), .Y(n_6) );
INVx2_ASAP7_75t_L g7 ( .A(n_4), .Y(n_7) );
NAND2x1p5_ASAP7_75t_L g8 ( .A(n_6), .B(n_5), .Y(n_8) );
AND2x2_ASAP7_75t_L g9 ( .A(n_7), .B(n_4), .Y(n_9) );
INVx1_ASAP7_75t_L g10 ( .A(n_9), .Y(n_10) );
INVx1_ASAP7_75t_L g11 ( .A(n_10), .Y(n_11) );
INVx1_ASAP7_75t_SL g12 ( .A(n_11), .Y(n_12) );
AND2x2_ASAP7_75t_L g13 ( .A(n_11), .B(n_8), .Y(n_13) );
CKINVDCx16_ASAP7_75t_R g14 ( .A(n_13), .Y(n_14) );
INVx1_ASAP7_75t_L g15 ( .A(n_12), .Y(n_15) );
OR2x2_ASAP7_75t_L g16 ( .A(n_14), .B(n_12), .Y(n_16) );
INVx2_ASAP7_75t_L g17 ( .A(n_15), .Y(n_17) );
INVx1_ASAP7_75t_L g18 ( .A(n_17), .Y(n_18) );
AOI22xp5_ASAP7_75t_SL g19 ( .A1(n_18), .A2(n_16), .B1(n_0), .B2(n_3), .Y(n_19) );
endmodule