module fake_ibex_516_n_630 (n_85, n_84, n_64, n_3, n_73, n_65, n_95, n_55, n_63, n_98, n_29, n_2, n_76, n_8, n_67, n_9, n_38, n_37, n_47, n_10, n_82, n_21, n_27, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_48, n_57, n_59, n_28, n_39, n_5, n_62, n_71, n_93, n_13, n_61, n_14, n_0, n_94, n_12, n_42, n_77, n_88, n_44, n_51, n_46, n_80, n_49, n_40, n_66, n_17, n_74, n_90, n_58, n_43, n_22, n_4, n_33, n_30, n_6, n_72, n_26, n_34, n_97, n_15, n_24, n_52, n_1, n_25, n_36, n_41, n_45, n_18, n_89, n_83, n_32, n_53, n_50, n_11, n_92, n_96, n_68, n_79, n_81, n_35, n_31, n_56, n_23, n_91, n_54, n_19, n_630);

input n_85;
input n_84;
input n_64;
input n_3;
input n_73;
input n_65;
input n_95;
input n_55;
input n_63;
input n_98;
input n_29;
input n_2;
input n_76;
input n_8;
input n_67;
input n_9;
input n_38;
input n_37;
input n_47;
input n_10;
input n_82;
input n_21;
input n_27;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_48;
input n_57;
input n_59;
input n_28;
input n_39;
input n_5;
input n_62;
input n_71;
input n_93;
input n_13;
input n_61;
input n_14;
input n_0;
input n_94;
input n_12;
input n_42;
input n_77;
input n_88;
input n_44;
input n_51;
input n_46;
input n_80;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_58;
input n_43;
input n_22;
input n_4;
input n_33;
input n_30;
input n_6;
input n_72;
input n_26;
input n_34;
input n_97;
input n_15;
input n_24;
input n_52;
input n_1;
input n_25;
input n_36;
input n_41;
input n_45;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_50;
input n_11;
input n_92;
input n_96;
input n_68;
input n_79;
input n_81;
input n_35;
input n_31;
input n_56;
input n_23;
input n_91;
input n_54;
input n_19;

output n_630;

wire n_151;
wire n_599;
wire n_507;
wire n_540;
wire n_395;
wire n_171;
wire n_103;
wire n_529;
wire n_389;
wire n_204;
wire n_626;
wire n_274;
wire n_387;
wire n_130;
wire n_177;
wire n_273;
wire n_330;
wire n_309;
wire n_328;
wire n_293;
wire n_341;
wire n_372;
wire n_124;
wire n_256;
wire n_418;
wire n_193;
wire n_510;
wire n_446;
wire n_108;
wire n_350;
wire n_601;
wire n_621;
wire n_610;
wire n_165;
wire n_452;
wire n_255;
wire n_175;
wire n_586;
wire n_398;
wire n_125;
wire n_304;
wire n_191;
wire n_593;
wire n_153;
wire n_545;
wire n_583;
wire n_194;
wire n_249;
wire n_334;
wire n_312;
wire n_622;
wire n_578;
wire n_478;
wire n_239;
wire n_134;
wire n_432;
wire n_371;
wire n_403;
wire n_423;
wire n_608;
wire n_357;
wire n_412;
wire n_457;
wire n_494;
wire n_142;
wire n_226;
wire n_336;
wire n_258;
wire n_449;
wire n_547;
wire n_176;
wire n_216;
wire n_421;
wire n_475;
wire n_166;
wire n_163;
wire n_500;
wire n_542;
wire n_114;
wire n_236;
wire n_376;
wire n_377;
wire n_584;
wire n_531;
wire n_556;
wire n_189;
wire n_498;
wire n_280;
wire n_317;
wire n_340;
wire n_375;
wire n_105;
wire n_187;
wire n_154;
wire n_182;
wire n_196;
wire n_327;
wire n_326;
wire n_144;
wire n_170;
wire n_270;
wire n_383;
wire n_346;
wire n_113;
wire n_561;
wire n_117;
wire n_417;
wire n_471;
wire n_265;
wire n_504;
wire n_158;
wire n_259;
wire n_339;
wire n_276;
wire n_470;
wire n_210;
wire n_348;
wire n_220;
wire n_481;
wire n_287;
wire n_243;
wire n_497;
wire n_228;
wire n_147;
wire n_552;
wire n_251;
wire n_384;
wire n_373;
wire n_458;
wire n_244;
wire n_343;
wire n_310;
wire n_426;
wire n_323;
wire n_469;
wire n_598;
wire n_143;
wire n_106;
wire n_386;
wire n_549;
wire n_224;
wire n_183;
wire n_533;
wire n_508;
wire n_453;
wire n_591;
wire n_333;
wire n_110;
wire n_400;
wire n_306;
wire n_550;
wire n_169;
wire n_242;
wire n_278;
wire n_316;
wire n_404;
wire n_557;
wire n_109;
wire n_127;
wire n_121;
wire n_527;
wire n_590;
wire n_465;
wire n_325;
wire n_301;
wire n_496;
wire n_617;
wire n_434;
wire n_296;
wire n_120;
wire n_168;
wire n_526;
wire n_155;
wire n_315;
wire n_441;
wire n_604;
wire n_122;
wire n_523;
wire n_116;
wire n_614;
wire n_370;
wire n_431;
wire n_574;
wire n_289;
wire n_515;
wire n_150;
wire n_286;
wire n_321;
wire n_133;
wire n_569;
wire n_600;
wire n_215;
wire n_279;
wire n_374;
wire n_235;
wire n_464;
wire n_538;
wire n_136;
wire n_261;
wire n_521;
wire n_459;
wire n_518;
wire n_367;
wire n_221;
wire n_437;
wire n_602;
wire n_355;
wire n_474;
wire n_594;
wire n_407;
wire n_102;
wire n_490;
wire n_568;
wire n_448;
wire n_595;
wire n_99;
wire n_466;
wire n_269;
wire n_156;
wire n_570;
wire n_126;
wire n_623;
wire n_585;
wire n_530;
wire n_356;
wire n_104;
wire n_420;
wire n_483;
wire n_543;
wire n_580;
wire n_141;
wire n_487;
wire n_222;
wire n_186;
wire n_524;
wire n_349;
wire n_454;
wire n_295;
wire n_331;
wire n_576;
wire n_230;
wire n_185;
wire n_388;
wire n_625;
wire n_619;
wire n_536;
wire n_611;
wire n_352;
wire n_290;
wire n_558;
wire n_174;
wire n_467;
wire n_427;
wire n_607;
wire n_157;
wire n_219;
wire n_246;
wire n_442;
wire n_146;
wire n_207;
wire n_438;
wire n_167;
wire n_128;
wire n_253;
wire n_208;
wire n_234;
wire n_152;
wire n_300;
wire n_145;
wire n_358;
wire n_205;
wire n_618;
wire n_488;
wire n_139;
wire n_514;
wire n_429;
wire n_560;
wire n_275;
wire n_541;
wire n_129;
wire n_613;
wire n_267;
wire n_245;
wire n_589;
wire n_571;
wire n_229;
wire n_209;
wire n_472;
wire n_347;
wire n_473;
wire n_445;
wire n_629;
wire n_335;
wire n_413;
wire n_263;
wire n_573;
wire n_353;
wire n_359;
wire n_299;
wire n_262;
wire n_433;
wire n_439;
wire n_137;
wire n_338;
wire n_173;
wire n_477;
wire n_363;
wire n_402;
wire n_180;
wire n_369;
wire n_596;
wire n_201;
wire n_351;
wire n_368;
wire n_456;
wire n_257;
wire n_401;
wire n_554;
wire n_553;
wire n_305;
wire n_307;
wire n_192;
wire n_140;
wire n_484;
wire n_566;
wire n_480;
wire n_416;
wire n_581;
wire n_365;
wire n_605;
wire n_539;
wire n_100;
wire n_179;
wire n_354;
wire n_206;
wire n_392;
wire n_516;
wire n_567;
wire n_548;
wire n_329;
wire n_447;
wire n_188;
wire n_200;
wire n_444;
wire n_506;
wire n_562;
wire n_564;
wire n_546;
wire n_199;
wire n_592;
wire n_495;
wire n_410;
wire n_308;
wire n_463;
wire n_624;
wire n_411;
wire n_135;
wire n_520;
wire n_512;
wire n_615;
wire n_283;
wire n_397;
wire n_366;
wire n_111;
wire n_627;
wire n_322;
wire n_227;
wire n_499;
wire n_115;
wire n_248;
wire n_451;
wire n_101;
wire n_190;
wire n_138;
wire n_409;
wire n_582;
wire n_238;
wire n_214;
wire n_579;
wire n_332;
wire n_517;
wire n_211;
wire n_218;
wire n_314;
wire n_563;
wire n_132;
wire n_277;
wire n_555;
wire n_337;
wire n_522;
wire n_479;
wire n_534;
wire n_225;
wire n_360;
wire n_272;
wire n_511;
wire n_468;
wire n_223;
wire n_381;
wire n_525;
wire n_535;
wire n_382;
wire n_502;
wire n_532;
wire n_405;
wire n_415;
wire n_597;
wire n_320;
wire n_285;
wire n_247;
wire n_288;
wire n_379;
wire n_551;
wire n_612;
wire n_291;
wire n_318;
wire n_161;
wire n_237;
wire n_203;
wire n_268;
wire n_440;
wire n_148;
wire n_385;
wire n_233;
wire n_342;
wire n_414;
wire n_430;
wire n_118;
wire n_603;
wire n_378;
wire n_486;
wire n_422;
wire n_164;
wire n_198;
wire n_264;
wire n_616;
wire n_217;
wire n_324;
wire n_391;
wire n_537;
wire n_390;
wire n_544;
wire n_178;
wire n_509;
wire n_303;
wire n_362;
wire n_505;
wire n_162;
wire n_482;
wire n_240;
wire n_282;
wire n_501;
wire n_266;
wire n_294;
wire n_112;
wire n_485;
wire n_284;
wire n_172;
wire n_250;
wire n_493;
wire n_460;
wire n_609;
wire n_476;
wire n_461;
wire n_575;
wire n_313;
wire n_519;
wire n_345;
wire n_408;
wire n_119;
wire n_361;
wire n_455;
wire n_419;
wire n_319;
wire n_195;
wire n_513;
wire n_212;
wire n_588;
wire n_311;
wire n_406;
wire n_606;
wire n_197;
wire n_528;
wire n_181;
wire n_131;
wire n_123;
wire n_260;
wire n_620;
wire n_462;
wire n_302;
wire n_450;
wire n_443;
wire n_572;
wire n_577;
wire n_344;
wire n_393;
wire n_436;
wire n_428;
wire n_491;
wire n_297;
wire n_435;
wire n_628;
wire n_252;
wire n_396;
wire n_107;
wire n_149;
wire n_489;
wire n_399;
wire n_254;
wire n_213;
wire n_424;
wire n_565;
wire n_271;
wire n_241;
wire n_503;
wire n_292;
wire n_394;
wire n_364;
wire n_159;
wire n_202;
wire n_231;
wire n_298;
wire n_587;
wire n_160;
wire n_184;
wire n_492;
wire n_232;
wire n_380;
wire n_281;
wire n_559;
wire n_425;

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_10),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_65),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_75),
.Y(n_101)
);

INVx1_ASAP7_75t_SL g102 ( 
.A(n_87),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_1),
.Y(n_103)
);

CKINVDCx14_ASAP7_75t_R g104 ( 
.A(n_3),
.Y(n_104)
);

CKINVDCx5p33_ASAP7_75t_R g105 ( 
.A(n_34),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_11),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_46),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_1),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_57),
.Y(n_109)
);

CKINVDCx5p33_ASAP7_75t_R g110 ( 
.A(n_33),
.Y(n_110)
);

CKINVDCx5p33_ASAP7_75t_R g111 ( 
.A(n_94),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_53),
.Y(n_112)
);

HB1xp67_ASAP7_75t_L g113 ( 
.A(n_45),
.Y(n_113)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_50),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_98),
.Y(n_115)
);

CKINVDCx5p33_ASAP7_75t_R g116 ( 
.A(n_48),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_59),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_8),
.Y(n_118)
);

CKINVDCx5p33_ASAP7_75t_R g119 ( 
.A(n_97),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_26),
.Y(n_120)
);

INVx1_ASAP7_75t_SL g121 ( 
.A(n_43),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_17),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_40),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_86),
.Y(n_124)
);

NOR2xp67_ASAP7_75t_L g125 ( 
.A(n_10),
.B(n_39),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_25),
.Y(n_126)
);

CKINVDCx5p33_ASAP7_75t_R g127 ( 
.A(n_5),
.Y(n_127)
);

CKINVDCx5p33_ASAP7_75t_R g128 ( 
.A(n_16),
.Y(n_128)
);

CKINVDCx5p33_ASAP7_75t_R g129 ( 
.A(n_13),
.Y(n_129)
);

INVxp33_ASAP7_75t_L g130 ( 
.A(n_56),
.Y(n_130)
);

BUFx2_ASAP7_75t_L g131 ( 
.A(n_49),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_91),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_44),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_62),
.Y(n_134)
);

INVx2_ASAP7_75t_SL g135 ( 
.A(n_22),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_35),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g137 ( 
.A(n_29),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_21),
.Y(n_138)
);

CKINVDCx5p33_ASAP7_75t_R g139 ( 
.A(n_19),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_60),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_68),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_9),
.Y(n_142)
);

CKINVDCx5p33_ASAP7_75t_R g143 ( 
.A(n_38),
.Y(n_143)
);

INVx2_ASAP7_75t_SL g144 ( 
.A(n_2),
.Y(n_144)
);

BUFx3_ASAP7_75t_L g145 ( 
.A(n_51),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_42),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_63),
.Y(n_147)
);

CKINVDCx5p33_ASAP7_75t_R g148 ( 
.A(n_3),
.Y(n_148)
);

CKINVDCx5p33_ASAP7_75t_R g149 ( 
.A(n_58),
.Y(n_149)
);

BUFx2_ASAP7_75t_SL g150 ( 
.A(n_90),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_20),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_80),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_30),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_7),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_18),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_55),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_23),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_84),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_21),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_85),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_12),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_37),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_66),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_77),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_16),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_32),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_61),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_31),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_78),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_67),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_28),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_22),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_6),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_93),
.Y(n_174)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_27),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_17),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_47),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_131),
.B(n_0),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_156),
.Y(n_179)
);

BUFx12f_ASAP7_75t_L g180 ( 
.A(n_131),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_114),
.Y(n_181)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_114),
.Y(n_182)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_167),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_167),
.Y(n_184)
);

HB1xp67_ASAP7_75t_L g185 ( 
.A(n_104),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_137),
.Y(n_186)
);

AND2x6_ASAP7_75t_L g187 ( 
.A(n_137),
.B(n_41),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_173),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_145),
.Y(n_189)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_173),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_145),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_113),
.B(n_0),
.Y(n_192)
);

AND2x4_ASAP7_75t_L g193 ( 
.A(n_175),
.B(n_2),
.Y(n_193)
);

AND2x4_ASAP7_75t_L g194 ( 
.A(n_175),
.B(n_135),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g195 ( 
.A(n_99),
.B(n_4),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_135),
.B(n_4),
.Y(n_196)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_118),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_156),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_100),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_156),
.Y(n_200)
);

AND2x4_ASAP7_75t_L g201 ( 
.A(n_144),
.B(n_5),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_101),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_156),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_107),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_115),
.B(n_54),
.Y(n_205)
);

OA21x2_ASAP7_75t_L g206 ( 
.A1(n_109),
.A2(n_177),
.B(n_174),
.Y(n_206)
);

OAI21x1_ASAP7_75t_L g207 ( 
.A1(n_112),
.A2(n_52),
.B(n_95),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_117),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_123),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_118),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_124),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_144),
.B(n_9),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_132),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_120),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_156),
.Y(n_215)
);

AND2x4_ASAP7_75t_L g216 ( 
.A(n_120),
.B(n_103),
.Y(n_216)
);

INVx2_ASAP7_75t_SL g217 ( 
.A(n_133),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_127),
.A2(n_14),
.B1(n_15),
.B2(n_18),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_134),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_136),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_141),
.Y(n_221)
);

OAI22x1_ASAP7_75t_L g222 ( 
.A1(n_127),
.A2(n_14),
.B1(n_15),
.B2(n_19),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_146),
.Y(n_223)
);

AND2x4_ASAP7_75t_L g224 ( 
.A(n_106),
.B(n_20),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_152),
.Y(n_225)
);

AND2x6_ASAP7_75t_L g226 ( 
.A(n_153),
.B(n_72),
.Y(n_226)
);

OR2x2_ASAP7_75t_L g227 ( 
.A(n_108),
.B(n_23),
.Y(n_227)
);

INVx5_ASAP7_75t_L g228 ( 
.A(n_140),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_160),
.Y(n_229)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_122),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_162),
.Y(n_231)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_163),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_170),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_147),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_138),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_142),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_128),
.B(n_24),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_151),
.Y(n_238)
);

BUFx2_ASAP7_75t_L g239 ( 
.A(n_128),
.Y(n_239)
);

AND2x6_ASAP7_75t_L g240 ( 
.A(n_102),
.B(n_73),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_155),
.Y(n_241)
);

INVx3_ASAP7_75t_L g242 ( 
.A(n_159),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_129),
.B(n_24),
.Y(n_243)
);

OAI21x1_ASAP7_75t_L g244 ( 
.A1(n_125),
.A2(n_74),
.B(n_92),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_161),
.Y(n_245)
);

AND2x4_ASAP7_75t_L g246 ( 
.A(n_172),
.B(n_25),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_150),
.Y(n_247)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_105),
.Y(n_248)
);

CKINVDCx6p67_ASAP7_75t_R g249 ( 
.A(n_150),
.Y(n_249)
);

AND2x4_ASAP7_75t_L g250 ( 
.A(n_171),
.B(n_26),
.Y(n_250)
);

BUFx2_ASAP7_75t_L g251 ( 
.A(n_239),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_245),
.Y(n_252)
);

OR2x6_ASAP7_75t_L g253 ( 
.A(n_180),
.B(n_176),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_179),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_184),
.B(n_169),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_245),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_247),
.B(n_130),
.Y(n_257)
);

NOR2x1p5_ASAP7_75t_L g258 ( 
.A(n_180),
.B(n_165),
.Y(n_258)
);

BUFx10_ASAP7_75t_L g259 ( 
.A(n_185),
.Y(n_259)
);

INVx2_ASAP7_75t_SL g260 ( 
.A(n_228),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_247),
.B(n_105),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_184),
.B(n_169),
.Y(n_262)
);

AND2x2_ASAP7_75t_L g263 ( 
.A(n_239),
.B(n_139),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_217),
.B(n_194),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_201),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_201),
.Y(n_266)
);

NAND2xp33_ASAP7_75t_R g267 ( 
.A(n_234),
.B(n_195),
.Y(n_267)
);

BUFx3_ASAP7_75t_L g268 ( 
.A(n_248),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_201),
.Y(n_269)
);

BUFx3_ASAP7_75t_L g270 ( 
.A(n_248),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_193),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_193),
.Y(n_272)
);

HB1xp67_ASAP7_75t_L g273 ( 
.A(n_234),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_199),
.B(n_168),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_245),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_245),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g277 ( 
.A(n_179),
.Y(n_277)
);

NAND3xp33_ASAP7_75t_L g278 ( 
.A(n_178),
.B(n_139),
.C(n_148),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_228),
.B(n_148),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_193),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_195),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_193),
.Y(n_282)
);

INVxp67_ASAP7_75t_SL g283 ( 
.A(n_237),
.Y(n_283)
);

INVx5_ASAP7_75t_L g284 ( 
.A(n_187),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_224),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_224),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_228),
.B(n_154),
.Y(n_287)
);

INVx2_ASAP7_75t_SL g288 ( 
.A(n_228),
.Y(n_288)
);

NAND2xp33_ASAP7_75t_L g289 ( 
.A(n_187),
.B(n_168),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_224),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_249),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_245),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_205),
.B(n_187),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_194),
.B(n_166),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_199),
.B(n_166),
.Y(n_295)
);

OAI22xp33_ASAP7_75t_L g296 ( 
.A1(n_218),
.A2(n_126),
.B1(n_157),
.B2(n_158),
.Y(n_296)
);

NOR2x1p5_ASAP7_75t_L g297 ( 
.A(n_249),
.B(n_164),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_202),
.B(n_164),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_250),
.A2(n_158),
.B1(n_149),
.B2(n_143),
.Y(n_299)
);

NOR3xp33_ASAP7_75t_L g300 ( 
.A(n_210),
.B(n_121),
.C(n_149),
.Y(n_300)
);

INVx4_ASAP7_75t_SL g301 ( 
.A(n_187),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_202),
.B(n_143),
.Y(n_302)
);

INVx3_ASAP7_75t_L g303 ( 
.A(n_194),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_224),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_246),
.Y(n_305)
);

BUFx3_ASAP7_75t_L g306 ( 
.A(n_248),
.Y(n_306)
);

BUFx10_ASAP7_75t_L g307 ( 
.A(n_250),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_246),
.Y(n_308)
);

BUFx3_ASAP7_75t_L g309 ( 
.A(n_248),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_250),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_194),
.B(n_119),
.Y(n_311)
);

INVx4_ASAP7_75t_L g312 ( 
.A(n_187),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_208),
.B(n_119),
.Y(n_313)
);

AND2x2_ASAP7_75t_L g314 ( 
.A(n_216),
.B(n_116),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_246),
.Y(n_315)
);

INVx4_ASAP7_75t_SL g316 ( 
.A(n_187),
.Y(n_316)
);

NAND3xp33_ASAP7_75t_L g317 ( 
.A(n_206),
.B(n_116),
.C(n_111),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_179),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_246),
.Y(n_319)
);

AND2x2_ASAP7_75t_L g320 ( 
.A(n_216),
.B(n_110),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_208),
.B(n_111),
.Y(n_321)
);

BUFx3_ASAP7_75t_L g322 ( 
.A(n_226),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_250),
.A2(n_110),
.B1(n_27),
.B2(n_36),
.Y(n_323)
);

INVx3_ASAP7_75t_L g324 ( 
.A(n_197),
.Y(n_324)
);

INVx3_ASAP7_75t_L g325 ( 
.A(n_197),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_179),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_197),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_179),
.Y(n_328)
);

NAND2xp33_ASAP7_75t_L g329 ( 
.A(n_187),
.B(n_64),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_209),
.B(n_69),
.Y(n_330)
);

INVx5_ASAP7_75t_L g331 ( 
.A(n_226),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_196),
.Y(n_332)
);

INVx1_ASAP7_75t_SL g333 ( 
.A(n_243),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_212),
.Y(n_334)
);

INVx4_ASAP7_75t_L g335 ( 
.A(n_226),
.Y(n_335)
);

OR2x2_ASAP7_75t_L g336 ( 
.A(n_238),
.B(n_70),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_198),
.Y(n_337)
);

AND2x4_ASAP7_75t_L g338 ( 
.A(n_216),
.B(n_71),
.Y(n_338)
);

BUFx10_ASAP7_75t_L g339 ( 
.A(n_216),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_332),
.B(n_209),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_334),
.B(n_229),
.Y(n_341)
);

A2O1A1Ixp33_ASAP7_75t_L g342 ( 
.A1(n_265),
.A2(n_211),
.B(n_229),
.C(n_223),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_257),
.B(n_220),
.Y(n_343)
);

OR2x6_ASAP7_75t_L g344 ( 
.A(n_253),
.B(n_222),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_283),
.B(n_225),
.Y(n_345)
);

AOI22xp33_ASAP7_75t_L g346 ( 
.A1(n_271),
.A2(n_206),
.B1(n_183),
.B2(n_225),
.Y(n_346)
);

AND2x4_ASAP7_75t_L g347 ( 
.A(n_297),
.B(n_227),
.Y(n_347)
);

OR2x2_ASAP7_75t_L g348 ( 
.A(n_251),
.B(n_227),
.Y(n_348)
);

INVx2_ASAP7_75t_SL g349 ( 
.A(n_259),
.Y(n_349)
);

INVx4_ASAP7_75t_L g350 ( 
.A(n_339),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_321),
.B(n_211),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_339),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_321),
.B(n_220),
.Y(n_353)
);

INVx4_ASAP7_75t_L g354 ( 
.A(n_339),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_SL g355 ( 
.A(n_312),
.B(n_231),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_314),
.B(n_241),
.Y(n_356)
);

AOI21xp5_ASAP7_75t_L g357 ( 
.A1(n_289),
.A2(n_206),
.B(n_244),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_320),
.B(n_241),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_295),
.B(n_238),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_257),
.B(n_230),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_294),
.B(n_242),
.Y(n_361)
);

BUFx3_ASAP7_75t_L g362 ( 
.A(n_268),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_SL g363 ( 
.A(n_312),
.B(n_335),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_294),
.B(n_242),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_303),
.Y(n_365)
);

AOI22x1_ASAP7_75t_L g366 ( 
.A1(n_335),
.A2(n_189),
.B1(n_186),
.B2(n_191),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_252),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_311),
.B(n_242),
.Y(n_368)
);

AND2x2_ASAP7_75t_L g369 ( 
.A(n_263),
.B(n_192),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_311),
.B(n_213),
.Y(n_370)
);

NAND3xp33_ASAP7_75t_L g371 ( 
.A(n_299),
.B(n_206),
.C(n_218),
.Y(n_371)
);

AND2x2_ASAP7_75t_L g372 ( 
.A(n_333),
.B(n_235),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_261),
.B(n_204),
.Y(n_373)
);

INVx4_ASAP7_75t_L g374 ( 
.A(n_338),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_261),
.B(n_204),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_252),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_264),
.B(n_219),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_264),
.B(n_219),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_SL g379 ( 
.A(n_293),
.B(n_231),
.Y(n_379)
);

O2A1O1Ixp33_ASAP7_75t_L g380 ( 
.A1(n_272),
.A2(n_282),
.B(n_280),
.C(n_266),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_310),
.B(n_221),
.Y(n_381)
);

INVxp33_ASAP7_75t_L g382 ( 
.A(n_273),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_324),
.B(n_221),
.Y(n_383)
);

AND2x4_ASAP7_75t_L g384 ( 
.A(n_278),
.B(n_236),
.Y(n_384)
);

INVxp67_ASAP7_75t_L g385 ( 
.A(n_259),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_324),
.B(n_233),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_325),
.B(n_233),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_325),
.B(n_232),
.Y(n_388)
);

INVx2_ASAP7_75t_SL g389 ( 
.A(n_307),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_255),
.B(n_232),
.Y(n_390)
);

NAND2xp33_ASAP7_75t_SL g391 ( 
.A(n_291),
.B(n_222),
.Y(n_391)
);

AOI22xp33_ASAP7_75t_L g392 ( 
.A1(n_269),
.A2(n_183),
.B1(n_226),
.B2(n_181),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_255),
.B(n_235),
.Y(n_393)
);

HB1xp67_ASAP7_75t_L g394 ( 
.A(n_267),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_262),
.B(n_236),
.Y(n_395)
);

BUFx3_ASAP7_75t_L g396 ( 
.A(n_268),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_262),
.B(n_226),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_327),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_274),
.B(n_226),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_274),
.B(n_226),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_298),
.B(n_190),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_298),
.B(n_186),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_L g403 ( 
.A1(n_300),
.A2(n_214),
.B1(n_191),
.B2(n_189),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_L g404 ( 
.A1(n_285),
.A2(n_181),
.B1(n_182),
.B2(n_188),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_302),
.B(n_190),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_L g406 ( 
.A1(n_286),
.A2(n_182),
.B1(n_188),
.B2(n_231),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_290),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_313),
.B(n_231),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_313),
.B(n_240),
.Y(n_409)
);

OR2x2_ASAP7_75t_L g410 ( 
.A(n_253),
.B(n_244),
.Y(n_410)
);

OAI22xp33_ASAP7_75t_L g411 ( 
.A1(n_281),
.A2(n_215),
.B1(n_203),
.B2(n_200),
.Y(n_411)
);

OAI221xp5_ASAP7_75t_L g412 ( 
.A1(n_323),
.A2(n_215),
.B1(n_203),
.B2(n_200),
.C(n_198),
.Y(n_412)
);

AOI22xp33_ASAP7_75t_L g413 ( 
.A1(n_304),
.A2(n_240),
.B1(n_207),
.B2(n_215),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_SL g414 ( 
.A(n_284),
.B(n_207),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_279),
.B(n_240),
.Y(n_415)
);

OR2x2_ASAP7_75t_L g416 ( 
.A(n_253),
.B(n_296),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_287),
.B(n_240),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_L g418 ( 
.A1(n_374),
.A2(n_319),
.B1(n_305),
.B2(n_308),
.Y(n_418)
);

AO22x1_ASAP7_75t_L g419 ( 
.A1(n_382),
.A2(n_338),
.B1(n_267),
.B2(n_315),
.Y(n_419)
);

BUFx3_ASAP7_75t_L g420 ( 
.A(n_349),
.Y(n_420)
);

AOI22xp33_ASAP7_75t_SL g421 ( 
.A1(n_344),
.A2(n_281),
.B1(n_338),
.B2(n_289),
.Y(n_421)
);

AOI21xp5_ASAP7_75t_L g422 ( 
.A1(n_397),
.A2(n_322),
.B(n_284),
.Y(n_422)
);

OR2x2_ASAP7_75t_L g423 ( 
.A(n_348),
.B(n_258),
.Y(n_423)
);

AOI21xp5_ASAP7_75t_L g424 ( 
.A1(n_399),
.A2(n_322),
.B(n_331),
.Y(n_424)
);

AOI21xp5_ASAP7_75t_L g425 ( 
.A1(n_400),
.A2(n_331),
.B(n_329),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_L g426 ( 
.A1(n_374),
.A2(n_336),
.B1(n_317),
.B2(n_330),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_340),
.B(n_288),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_347),
.B(n_260),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_340),
.B(n_270),
.Y(n_429)
);

BUFx2_ASAP7_75t_L g430 ( 
.A(n_385),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_365),
.Y(n_431)
);

A2O1A1Ixp33_ASAP7_75t_L g432 ( 
.A1(n_343),
.A2(n_329),
.B(n_330),
.C(n_270),
.Y(n_432)
);

A2O1A1Ixp33_ASAP7_75t_L g433 ( 
.A1(n_343),
.A2(n_306),
.B(n_309),
.C(n_331),
.Y(n_433)
);

BUFx6f_ASAP7_75t_L g434 ( 
.A(n_350),
.Y(n_434)
);

BUFx6f_ASAP7_75t_L g435 ( 
.A(n_350),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_SL g436 ( 
.A(n_354),
.B(n_301),
.Y(n_436)
);

INVx3_ASAP7_75t_L g437 ( 
.A(n_354),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_345),
.B(n_316),
.Y(n_438)
);

INVx5_ASAP7_75t_L g439 ( 
.A(n_389),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_341),
.B(n_240),
.Y(n_440)
);

INVx1_ASAP7_75t_SL g441 ( 
.A(n_362),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_360),
.B(n_240),
.Y(n_442)
);

BUFx2_ASAP7_75t_L g443 ( 
.A(n_394),
.Y(n_443)
);

OAI21xp33_ASAP7_75t_SL g444 ( 
.A1(n_360),
.A2(n_256),
.B(n_275),
.Y(n_444)
);

A2O1A1Ixp33_ASAP7_75t_L g445 ( 
.A1(n_380),
.A2(n_276),
.B(n_292),
.C(n_198),
.Y(n_445)
);

INVxp33_ASAP7_75t_SL g446 ( 
.A(n_416),
.Y(n_446)
);

OAI22x1_ASAP7_75t_L g447 ( 
.A1(n_371),
.A2(n_276),
.B1(n_292),
.B2(n_81),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_369),
.B(n_76),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_359),
.B(n_203),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_356),
.B(n_203),
.Y(n_450)
);

O2A1O1Ixp33_ASAP7_75t_L g451 ( 
.A1(n_342),
.A2(n_358),
.B(n_353),
.C(n_351),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_362),
.Y(n_452)
);

BUFx6f_ASAP7_75t_L g453 ( 
.A(n_396),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_381),
.B(n_79),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_L g455 ( 
.A1(n_407),
.A2(n_203),
.B1(n_215),
.B2(n_200),
.Y(n_455)
);

INVx3_ASAP7_75t_L g456 ( 
.A(n_396),
.Y(n_456)
);

A2O1A1Ixp33_ASAP7_75t_L g457 ( 
.A1(n_375),
.A2(n_215),
.B(n_200),
.C(n_337),
.Y(n_457)
);

AOI21xp5_ASAP7_75t_L g458 ( 
.A1(n_363),
.A2(n_357),
.B(n_414),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g459 ( 
.A(n_352),
.B(n_200),
.Y(n_459)
);

A2O1A1Ixp33_ASAP7_75t_L g460 ( 
.A1(n_375),
.A2(n_326),
.B(n_318),
.C(n_328),
.Y(n_460)
);

AOI22xp33_ASAP7_75t_L g461 ( 
.A1(n_384),
.A2(n_326),
.B1(n_318),
.B2(n_277),
.Y(n_461)
);

INVx4_ASAP7_75t_L g462 ( 
.A(n_344),
.Y(n_462)
);

AOI22xp33_ASAP7_75t_L g463 ( 
.A1(n_384),
.A2(n_277),
.B1(n_254),
.B2(n_83),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_SL g464 ( 
.A(n_410),
.B(n_277),
.Y(n_464)
);

HB1xp67_ASAP7_75t_L g465 ( 
.A(n_383),
.Y(n_465)
);

OR2x6_ASAP7_75t_L g466 ( 
.A(n_405),
.B(n_254),
.Y(n_466)
);

INVx6_ASAP7_75t_L g467 ( 
.A(n_403),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_L g468 ( 
.A1(n_346),
.A2(n_254),
.B1(n_82),
.B2(n_88),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_L g469 ( 
.A1(n_373),
.A2(n_89),
.B1(n_96),
.B2(n_378),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_370),
.B(n_361),
.Y(n_470)
);

AOI21xp5_ASAP7_75t_L g471 ( 
.A1(n_355),
.A2(n_409),
.B(n_379),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_364),
.B(n_368),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_398),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_401),
.B(n_377),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_SL g475 ( 
.A(n_411),
.B(n_392),
.Y(n_475)
);

OA22x2_ASAP7_75t_L g476 ( 
.A1(n_390),
.A2(n_395),
.B1(n_393),
.B2(n_404),
.Y(n_476)
);

BUFx2_ASAP7_75t_L g477 ( 
.A(n_386),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_401),
.B(n_387),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_402),
.Y(n_479)
);

AOI21xp5_ASAP7_75t_L g480 ( 
.A1(n_355),
.A2(n_417),
.B(n_415),
.Y(n_480)
);

NOR2xp67_ASAP7_75t_L g481 ( 
.A(n_412),
.B(n_408),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_388),
.B(n_392),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_406),
.B(n_417),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_366),
.Y(n_484)
);

AOI222xp33_ASAP7_75t_SL g485 ( 
.A1(n_430),
.A2(n_367),
.B1(n_376),
.B2(n_413),
.C1(n_443),
.C2(n_423),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_467),
.B(n_465),
.Y(n_486)
);

O2A1O1Ixp33_ASAP7_75t_SL g487 ( 
.A1(n_432),
.A2(n_445),
.B(n_433),
.C(n_457),
.Y(n_487)
);

AOI21xp5_ASAP7_75t_L g488 ( 
.A1(n_425),
.A2(n_480),
.B(n_471),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_470),
.B(n_477),
.Y(n_489)
);

AOI21xp5_ASAP7_75t_L g490 ( 
.A1(n_442),
.A2(n_424),
.B(n_422),
.Y(n_490)
);

NOR4xp25_ASAP7_75t_L g491 ( 
.A(n_444),
.B(n_469),
.C(n_448),
.D(n_418),
.Y(n_491)
);

BUFx2_ASAP7_75t_L g492 ( 
.A(n_434),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_472),
.B(n_479),
.Y(n_493)
);

AOI21xp5_ASAP7_75t_L g494 ( 
.A1(n_438),
.A2(n_440),
.B(n_474),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_428),
.B(n_420),
.Y(n_495)
);

AO31x2_ASAP7_75t_L g496 ( 
.A1(n_460),
.A2(n_426),
.A3(n_482),
.B(n_483),
.Y(n_496)
);

A2O1A1Ixp33_ASAP7_75t_L g497 ( 
.A1(n_454),
.A2(n_478),
.B(n_427),
.C(n_481),
.Y(n_497)
);

AND2x4_ASAP7_75t_L g498 ( 
.A(n_437),
.B(n_434),
.Y(n_498)
);

AOI21xp5_ASAP7_75t_L g499 ( 
.A1(n_464),
.A2(n_449),
.B(n_450),
.Y(n_499)
);

BUFx6f_ASAP7_75t_L g500 ( 
.A(n_435),
.Y(n_500)
);

AO31x2_ASAP7_75t_L g501 ( 
.A1(n_455),
.A2(n_429),
.A3(n_476),
.B(n_431),
.Y(n_501)
);

O2A1O1Ixp33_ASAP7_75t_SL g502 ( 
.A1(n_475),
.A2(n_436),
.B(n_459),
.C(n_441),
.Y(n_502)
);

BUFx3_ASAP7_75t_L g503 ( 
.A(n_439),
.Y(n_503)
);

AOI21xp5_ASAP7_75t_L g504 ( 
.A1(n_466),
.A2(n_452),
.B(n_461),
.Y(n_504)
);

O2A1O1Ixp33_ASAP7_75t_SL g505 ( 
.A1(n_456),
.A2(n_466),
.B(n_463),
.C(n_453),
.Y(n_505)
);

AOI21xp5_ASAP7_75t_L g506 ( 
.A1(n_453),
.A2(n_458),
.B(n_425),
.Y(n_506)
);

BUFx6f_ASAP7_75t_L g507 ( 
.A(n_434),
.Y(n_507)
);

OAI22xp5_ASAP7_75t_L g508 ( 
.A1(n_467),
.A2(n_421),
.B1(n_374),
.B2(n_470),
.Y(n_508)
);

AOI21xp5_ASAP7_75t_L g509 ( 
.A1(n_458),
.A2(n_425),
.B(n_312),
.Y(n_509)
);

O2A1O1Ixp33_ASAP7_75t_SL g510 ( 
.A1(n_432),
.A2(n_445),
.B(n_433),
.C(n_457),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_467),
.B(n_372),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_467),
.B(n_372),
.Y(n_512)
);

OAI22xp5_ASAP7_75t_L g513 ( 
.A1(n_467),
.A2(n_421),
.B1(n_374),
.B2(n_470),
.Y(n_513)
);

OA21x2_ASAP7_75t_L g514 ( 
.A1(n_458),
.A2(n_357),
.B(n_484),
.Y(n_514)
);

INVx3_ASAP7_75t_SL g515 ( 
.A(n_462),
.Y(n_515)
);

AOI21xp5_ASAP7_75t_L g516 ( 
.A1(n_458),
.A2(n_425),
.B(n_312),
.Y(n_516)
);

INVx8_ASAP7_75t_L g517 ( 
.A(n_434),
.Y(n_517)
);

AO31x2_ASAP7_75t_L g518 ( 
.A1(n_447),
.A2(n_432),
.A3(n_468),
.B(n_458),
.Y(n_518)
);

AOI22xp5_ASAP7_75t_L g519 ( 
.A1(n_467),
.A2(n_470),
.B1(n_371),
.B2(n_391),
.Y(n_519)
);

AOI211x1_ASAP7_75t_L g520 ( 
.A1(n_419),
.A2(n_371),
.B(n_474),
.C(n_412),
.Y(n_520)
);

NAND3xp33_ASAP7_75t_L g521 ( 
.A(n_469),
.B(n_448),
.C(n_432),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_473),
.Y(n_522)
);

AO31x2_ASAP7_75t_L g523 ( 
.A1(n_447),
.A2(n_432),
.A3(n_468),
.B(n_458),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_446),
.B(n_382),
.Y(n_524)
);

INVx3_ASAP7_75t_L g525 ( 
.A(n_434),
.Y(n_525)
);

AOI21xp5_ASAP7_75t_L g526 ( 
.A1(n_458),
.A2(n_425),
.B(n_312),
.Y(n_526)
);

INVxp67_ASAP7_75t_SL g527 ( 
.A(n_465),
.Y(n_527)
);

AO31x2_ASAP7_75t_L g528 ( 
.A1(n_447),
.A2(n_432),
.A3(n_468),
.B(n_458),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_446),
.B(n_382),
.Y(n_529)
);

AOI21xp5_ASAP7_75t_L g530 ( 
.A1(n_458),
.A2(n_425),
.B(n_312),
.Y(n_530)
);

CKINVDCx16_ASAP7_75t_R g531 ( 
.A(n_420),
.Y(n_531)
);

AO32x2_ASAP7_75t_L g532 ( 
.A1(n_469),
.A2(n_468),
.A3(n_426),
.B1(n_404),
.B2(n_406),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_SL g533 ( 
.A(n_434),
.B(n_349),
.Y(n_533)
);

AOI21xp5_ASAP7_75t_L g534 ( 
.A1(n_458),
.A2(n_425),
.B(n_312),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_467),
.B(n_372),
.Y(n_535)
);

A2O1A1Ixp33_ASAP7_75t_L g536 ( 
.A1(n_451),
.A2(n_470),
.B(n_343),
.C(n_360),
.Y(n_536)
);

AOI21xp5_ASAP7_75t_L g537 ( 
.A1(n_458),
.A2(n_425),
.B(n_312),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_467),
.B(n_372),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_467),
.B(n_372),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_467),
.B(n_372),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_430),
.Y(n_541)
);

INVxp67_ASAP7_75t_L g542 ( 
.A(n_430),
.Y(n_542)
);

BUFx6f_ASAP7_75t_SL g543 ( 
.A(n_503),
.Y(n_543)
);

AOI21xp5_ASAP7_75t_L g544 ( 
.A1(n_497),
.A2(n_521),
.B(n_510),
.Y(n_544)
);

AOI21xp5_ASAP7_75t_L g545 ( 
.A1(n_487),
.A2(n_536),
.B(n_488),
.Y(n_545)
);

INVx4_ASAP7_75t_L g546 ( 
.A(n_517),
.Y(n_546)
);

AND2x2_ASAP7_75t_L g547 ( 
.A(n_489),
.B(n_493),
.Y(n_547)
);

AND2x2_ASAP7_75t_L g548 ( 
.A(n_522),
.B(n_527),
.Y(n_548)
);

CKINVDCx20_ASAP7_75t_R g549 ( 
.A(n_531),
.Y(n_549)
);

A2O1A1Ixp33_ASAP7_75t_L g550 ( 
.A1(n_519),
.A2(n_512),
.B(n_540),
.C(n_539),
.Y(n_550)
);

AO31x2_ASAP7_75t_L g551 ( 
.A1(n_506),
.A2(n_490),
.A3(n_494),
.B(n_526),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_514),
.Y(n_552)
);

AO21x2_ASAP7_75t_L g553 ( 
.A1(n_491),
.A2(n_509),
.B(n_537),
.Y(n_553)
);

AO21x1_ASAP7_75t_L g554 ( 
.A1(n_516),
.A2(n_534),
.B(n_530),
.Y(n_554)
);

AOI22xp5_ASAP7_75t_L g555 ( 
.A1(n_524),
.A2(n_529),
.B1(n_508),
.B2(n_513),
.Y(n_555)
);

OAI221xp5_ASAP7_75t_L g556 ( 
.A1(n_519),
.A2(n_511),
.B1(n_538),
.B2(n_535),
.C(n_486),
.Y(n_556)
);

AND2x4_ASAP7_75t_L g557 ( 
.A(n_498),
.B(n_500),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_542),
.B(n_495),
.Y(n_558)
);

NAND3xp33_ASAP7_75t_L g559 ( 
.A(n_485),
.B(n_520),
.C(n_504),
.Y(n_559)
);

NAND2x1p5_ASAP7_75t_L g560 ( 
.A(n_500),
.B(n_507),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_492),
.Y(n_561)
);

OA21x2_ASAP7_75t_L g562 ( 
.A1(n_499),
.A2(n_518),
.B(n_523),
.Y(n_562)
);

BUFx2_ASAP7_75t_L g563 ( 
.A(n_517),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_515),
.B(n_498),
.Y(n_564)
);

OAI21x1_ASAP7_75t_L g565 ( 
.A1(n_525),
.A2(n_518),
.B(n_528),
.Y(n_565)
);

INVx5_ASAP7_75t_SL g566 ( 
.A(n_500),
.Y(n_566)
);

AOI21xp5_ASAP7_75t_L g567 ( 
.A1(n_502),
.A2(n_505),
.B(n_533),
.Y(n_567)
);

OAI21x1_ASAP7_75t_L g568 ( 
.A1(n_523),
.A2(n_528),
.B(n_496),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_501),
.Y(n_569)
);

BUFx6f_ASAP7_75t_L g570 ( 
.A(n_532),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_520),
.B(n_501),
.Y(n_571)
);

AOI22xp33_ASAP7_75t_L g572 ( 
.A1(n_508),
.A2(n_467),
.B1(n_446),
.B2(n_513),
.Y(n_572)
);

BUFx12f_ASAP7_75t_L g573 ( 
.A(n_541),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_514),
.Y(n_574)
);

CKINVDCx6p67_ASAP7_75t_R g575 ( 
.A(n_543),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_569),
.Y(n_576)
);

INVx3_ASAP7_75t_L g577 ( 
.A(n_560),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_552),
.Y(n_578)
);

AO21x2_ASAP7_75t_L g579 ( 
.A1(n_545),
.A2(n_544),
.B(n_550),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_574),
.Y(n_580)
);

AO21x2_ASAP7_75t_L g581 ( 
.A1(n_571),
.A2(n_554),
.B(n_559),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_573),
.Y(n_582)
);

AOI22xp5_ASAP7_75t_L g583 ( 
.A1(n_572),
.A2(n_556),
.B1(n_555),
.B2(n_547),
.Y(n_583)
);

INVx3_ASAP7_75t_L g584 ( 
.A(n_566),
.Y(n_584)
);

AND2x2_ASAP7_75t_L g585 ( 
.A(n_570),
.B(n_568),
.Y(n_585)
);

AND2x4_ASAP7_75t_L g586 ( 
.A(n_565),
.B(n_551),
.Y(n_586)
);

AND2x4_ASAP7_75t_L g587 ( 
.A(n_551),
.B(n_553),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_576),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_576),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_576),
.Y(n_590)
);

INVx3_ASAP7_75t_L g591 ( 
.A(n_586),
.Y(n_591)
);

INVx4_ASAP7_75t_L g592 ( 
.A(n_577),
.Y(n_592)
);

INVxp67_ASAP7_75t_SL g593 ( 
.A(n_578),
.Y(n_593)
);

BUFx2_ASAP7_75t_L g594 ( 
.A(n_580),
.Y(n_594)
);

AND2x2_ASAP7_75t_L g595 ( 
.A(n_587),
.B(n_562),
.Y(n_595)
);

INVxp67_ASAP7_75t_SL g596 ( 
.A(n_580),
.Y(n_596)
);

AND2x2_ASAP7_75t_L g597 ( 
.A(n_587),
.B(n_562),
.Y(n_597)
);

OR2x2_ASAP7_75t_L g598 ( 
.A(n_594),
.B(n_581),
.Y(n_598)
);

OR2x2_ASAP7_75t_L g599 ( 
.A(n_594),
.B(n_581),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_588),
.Y(n_600)
);

AND2x2_ASAP7_75t_L g601 ( 
.A(n_595),
.B(n_585),
.Y(n_601)
);

AND2x2_ASAP7_75t_L g602 ( 
.A(n_595),
.B(n_585),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_589),
.Y(n_603)
);

AND2x2_ASAP7_75t_L g604 ( 
.A(n_595),
.B(n_585),
.Y(n_604)
);

BUFx2_ASAP7_75t_SL g605 ( 
.A(n_592),
.Y(n_605)
);

AND2x4_ASAP7_75t_L g606 ( 
.A(n_601),
.B(n_591),
.Y(n_606)
);

AND2x2_ASAP7_75t_L g607 ( 
.A(n_601),
.B(n_597),
.Y(n_607)
);

INVx1_ASAP7_75t_SL g608 ( 
.A(n_605),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_603),
.Y(n_609)
);

AND2x2_ASAP7_75t_L g610 ( 
.A(n_602),
.B(n_597),
.Y(n_610)
);

OR2x2_ASAP7_75t_L g611 ( 
.A(n_602),
.B(n_594),
.Y(n_611)
);

INVxp67_ASAP7_75t_SL g612 ( 
.A(n_611),
.Y(n_612)
);

CKINVDCx14_ASAP7_75t_R g613 ( 
.A(n_607),
.Y(n_613)
);

OAI33xp33_ASAP7_75t_L g614 ( 
.A1(n_609),
.A2(n_600),
.A3(n_599),
.B1(n_598),
.B2(n_590),
.B3(n_558),
.Y(n_614)
);

OR2x2_ASAP7_75t_L g615 ( 
.A(n_607),
.B(n_604),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_SL g616 ( 
.A(n_612),
.B(n_608),
.Y(n_616)
);

OA22x2_ASAP7_75t_L g617 ( 
.A1(n_613),
.A2(n_606),
.B1(n_610),
.B2(n_582),
.Y(n_617)
);

AOI21xp5_ASAP7_75t_L g618 ( 
.A1(n_614),
.A2(n_593),
.B(n_596),
.Y(n_618)
);

OAI22xp5_ASAP7_75t_L g619 ( 
.A1(n_617),
.A2(n_615),
.B1(n_575),
.B2(n_583),
.Y(n_619)
);

AOI21xp5_ASAP7_75t_L g620 ( 
.A1(n_619),
.A2(n_616),
.B(n_618),
.Y(n_620)
);

AND2x4_ASAP7_75t_L g621 ( 
.A(n_620),
.B(n_549),
.Y(n_621)
);

NAND5xp2_ASAP7_75t_L g622 ( 
.A(n_621),
.B(n_575),
.C(n_563),
.D(n_567),
.E(n_564),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_622),
.Y(n_623)
);

XNOR2x1_ASAP7_75t_L g624 ( 
.A(n_623),
.B(n_575),
.Y(n_624)
);

AOI22xp5_ASAP7_75t_L g625 ( 
.A1(n_624),
.A2(n_543),
.B1(n_587),
.B2(n_546),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_625),
.Y(n_626)
);

OAI21xp33_ASAP7_75t_L g627 ( 
.A1(n_626),
.A2(n_584),
.B(n_561),
.Y(n_627)
);

OAI21xp33_ASAP7_75t_L g628 ( 
.A1(n_627),
.A2(n_584),
.B(n_548),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_628),
.Y(n_629)
);

AOI22xp5_ASAP7_75t_L g630 ( 
.A1(n_629),
.A2(n_566),
.B1(n_557),
.B2(n_579),
.Y(n_630)
);


endmodule