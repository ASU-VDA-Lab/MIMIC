module fake_jpeg_17067_n_137 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_137);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_137;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_4),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_7),
.Y(n_44)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_8),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_8),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_17),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_28),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_42),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_10),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_36),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_21),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_2),
.Y(n_55)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_2),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_0),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_40),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_54),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_60),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_54),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_61),
.Y(n_75)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_55),
.Y(n_62)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_62),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_46),
.B(n_0),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_63),
.B(n_43),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_50),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_64),
.B(n_62),
.Y(n_69)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_58),
.Y(n_65)
);

HAxp5_ASAP7_75t_SL g71 ( 
.A(n_65),
.B(n_48),
.CON(n_71),
.SN(n_71)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_58),
.Y(n_66)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_66),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_57),
.Y(n_67)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_67),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_65),
.A2(n_45),
.B1(n_46),
.B2(n_56),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_68),
.A2(n_74),
.B1(n_57),
.B2(n_59),
.Y(n_93)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_69),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_70),
.B(n_80),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_71),
.A2(n_61),
.B(n_48),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_66),
.A2(n_45),
.B1(n_56),
.B2(n_49),
.Y(n_74)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_67),
.Y(n_77)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_77),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_63),
.B(n_44),
.Y(n_78)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_78),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_64),
.B(n_47),
.Y(n_80)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_60),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_81),
.B(n_61),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_60),
.A2(n_49),
.B1(n_53),
.B2(n_52),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_82),
.A2(n_51),
.B1(n_3),
.B2(n_4),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_72),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_83),
.B(n_87),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g104 ( 
.A1(n_85),
.A2(n_93),
.B(n_94),
.Y(n_104)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_86),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_73),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_73),
.B(n_1),
.Y(n_88)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_88),
.Y(n_100)
);

INVxp67_ASAP7_75t_SL g90 ( 
.A(n_76),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_90),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_75),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_91),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_75),
.Y(n_92)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_92),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_74),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_97),
.A2(n_98),
.B1(n_3),
.B2(n_5),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_71),
.B(n_1),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_93),
.A2(n_68),
.B(n_23),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_105),
.A2(n_104),
.B(n_103),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_106),
.B(n_107),
.Y(n_114)
);

AO22x1_ASAP7_75t_SL g107 ( 
.A1(n_97),
.A2(n_79),
.B1(n_6),
.B2(n_7),
.Y(n_107)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_109),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_102),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_110),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_100),
.B(n_89),
.C(n_96),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_111),
.A2(n_108),
.B1(n_103),
.B2(n_95),
.Y(n_118)
);

OR2x2_ASAP7_75t_L g112 ( 
.A(n_99),
.B(n_84),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_112),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_107),
.B(n_84),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_113),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_118),
.B(n_114),
.Y(n_123)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_116),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_120),
.A2(n_121),
.B1(n_122),
.B2(n_117),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_115),
.B(n_114),
.Y(n_121)
);

INVx1_ASAP7_75t_SL g122 ( 
.A(n_118),
.Y(n_122)
);

AOI21xp33_ASAP7_75t_L g126 ( 
.A1(n_123),
.A2(n_101),
.B(n_90),
.Y(n_126)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_124),
.Y(n_128)
);

OAI322xp33_ASAP7_75t_L g125 ( 
.A1(n_122),
.A2(n_119),
.A3(n_101),
.B1(n_9),
.B2(n_11),
.C1(n_12),
.C2(n_13),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_125),
.A2(n_126),
.B1(n_25),
.B2(n_38),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_127),
.B(n_24),
.C(n_35),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_129),
.B(n_26),
.Y(n_130)
);

AOI21xp33_ASAP7_75t_L g131 ( 
.A1(n_130),
.A2(n_22),
.B(n_41),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_131),
.B(n_20),
.Y(n_132)
);

AOI322xp5_ASAP7_75t_L g133 ( 
.A1(n_132),
.A2(n_128),
.A3(n_27),
.B1(n_14),
.B2(n_15),
.C1(n_16),
.C2(n_18),
.Y(n_133)
);

AOI322xp5_ASAP7_75t_L g134 ( 
.A1(n_133),
.A2(n_30),
.A3(n_32),
.B1(n_19),
.B2(n_29),
.C1(n_33),
.C2(n_31),
.Y(n_134)
);

BUFx24_ASAP7_75t_SL g135 ( 
.A(n_134),
.Y(n_135)
);

XNOR2x2_ASAP7_75t_SL g136 ( 
.A(n_135),
.B(n_5),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_136),
.B(n_6),
.Y(n_137)
);


endmodule