module fake_jpeg_25408_n_199 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_199);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_199;

wire n_159;
wire n_117;
wire n_144;
wire n_10;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_2),
.Y(n_10)
);

INVx11_ASAP7_75t_L g11 ( 
.A(n_5),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_9),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

BUFx5_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

INVx4_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx12_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

INVx13_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_27),
.B(n_28),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_14),
.B(n_5),
.Y(n_28)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx8_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_30),
.A2(n_15),
.B1(n_16),
.B2(n_14),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_20),
.B(n_6),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_31),
.B(n_32),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

OAI22xp33_ASAP7_75t_L g33 ( 
.A1(n_23),
.A2(n_15),
.B1(n_10),
.B2(n_17),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_33),
.A2(n_40),
.B1(n_43),
.B2(n_23),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_23),
.A2(n_15),
.B1(n_19),
.B2(n_22),
.Y(n_40)
);

OA22x2_ASAP7_75t_L g56 ( 
.A1(n_42),
.A2(n_29),
.B1(n_24),
.B2(n_30),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_27),
.B(n_10),
.C(n_18),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_44),
.Y(n_80)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

A2O1A1Ixp33_ASAP7_75t_L g46 ( 
.A1(n_39),
.A2(n_28),
.B(n_31),
.C(n_27),
.Y(n_46)
);

NAND3xp33_ASAP7_75t_L g69 ( 
.A(n_46),
.B(n_30),
.C(n_1),
.Y(n_69)
);

NOR2x1_ASAP7_75t_L g47 ( 
.A(n_39),
.B(n_20),
.Y(n_47)
);

OR2x2_ASAP7_75t_L g62 ( 
.A(n_47),
.B(n_53),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_40),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_48),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_49),
.A2(n_58),
.B1(n_25),
.B2(n_37),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_28),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_50),
.B(n_17),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_35),
.B(n_19),
.Y(n_51)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_51),
.Y(n_67)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_52),
.B(n_54),
.Y(n_74)
);

OR2x2_ASAP7_75t_L g53 ( 
.A(n_35),
.B(n_21),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_34),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_55),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_56),
.A2(n_42),
.B(n_0),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_57),
.B(n_61),
.Y(n_76)
);

OAI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_43),
.A2(n_30),
.B1(n_29),
.B2(n_24),
.Y(n_58)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

INVx2_ASAP7_75t_SL g68 ( 
.A(n_59),
.Y(n_68)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_60),
.Y(n_78)
);

BUFx2_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

AND2x6_ASAP7_75t_L g64 ( 
.A(n_55),
.B(n_6),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_64),
.B(n_69),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_66),
.A2(n_65),
.B1(n_37),
.B2(n_60),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_70),
.B(n_73),
.Y(n_90)
);

BUFx24_ASAP7_75t_SL g71 ( 
.A(n_50),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_71),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_49),
.B(n_34),
.C(n_38),
.Y(n_72)
);

XOR2xp5_ASAP7_75t_L g85 ( 
.A(n_72),
.B(n_56),
.Y(n_85)
);

AND2x6_ASAP7_75t_L g73 ( 
.A(n_47),
.B(n_1),
.Y(n_73)
);

OR2x2_ASAP7_75t_L g75 ( 
.A(n_53),
.B(n_20),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_75),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_79),
.A2(n_0),
.B(n_1),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_74),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_82),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_80),
.Y(n_83)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_83),
.Y(n_107)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_76),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_84),
.B(n_86),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_85),
.B(n_25),
.Y(n_116)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_63),
.Y(n_86)
);

AOI22x1_ASAP7_75t_SL g87 ( 
.A1(n_79),
.A2(n_56),
.B1(n_46),
.B2(n_48),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_87),
.A2(n_89),
.B(n_95),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_88),
.A2(n_89),
.B1(n_87),
.B2(n_68),
.Y(n_105)
);

AND2x4_ASAP7_75t_L g89 ( 
.A(n_66),
.B(n_56),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_70),
.B(n_77),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_91),
.B(n_93),
.Y(n_111)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_80),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_92),
.B(n_94),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_77),
.B(n_54),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_62),
.Y(n_94)
);

NAND2xp33_ASAP7_75t_SL g95 ( 
.A(n_72),
.B(n_16),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_68),
.Y(n_96)
);

INVxp33_ASAP7_75t_L g103 ( 
.A(n_96),
.Y(n_103)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_62),
.Y(n_97)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_97),
.Y(n_119)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_75),
.Y(n_98)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_98),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_101),
.A2(n_13),
.B(n_12),
.Y(n_112)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_78),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_102),
.B(n_45),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_88),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_104),
.B(n_121),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_105),
.A2(n_101),
.B1(n_96),
.B2(n_99),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_89),
.A2(n_64),
.B(n_73),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_108),
.A2(n_112),
.B(n_100),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_85),
.B(n_91),
.C(n_93),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_113),
.B(n_114),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_95),
.B(n_67),
.C(n_38),
.Y(n_114)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_83),
.Y(n_115)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_115),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_116),
.B(n_120),
.Y(n_139)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_118),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_90),
.B(n_44),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_90),
.B(n_34),
.C(n_32),
.Y(n_121)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_102),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_123),
.B(n_124),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_89),
.B(n_25),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_125),
.A2(n_137),
.B1(n_140),
.B2(n_142),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_109),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_126),
.B(n_131),
.Y(n_149)
);

INVx6_ASAP7_75t_SL g129 ( 
.A(n_103),
.Y(n_129)
);

CKINVDCx14_ASAP7_75t_R g154 ( 
.A(n_129),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_110),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_117),
.B(n_68),
.Y(n_133)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_133),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_134),
.A2(n_135),
.B(n_13),
.Y(n_155)
);

OAI21x1_ASAP7_75t_L g135 ( 
.A1(n_106),
.A2(n_108),
.B(n_112),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_118),
.Y(n_136)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_136),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_120),
.A2(n_52),
.B1(n_59),
.B2(n_21),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_111),
.Y(n_138)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_138),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_122),
.B(n_10),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_111),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_106),
.A2(n_37),
.B1(n_29),
.B2(n_24),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_143),
.A2(n_115),
.B1(n_107),
.B2(n_114),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_141),
.B(n_116),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_145),
.B(n_147),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_141),
.B(n_113),
.Y(n_147)
);

OAI21xp33_ASAP7_75t_R g150 ( 
.A1(n_125),
.A2(n_121),
.B(n_124),
.Y(n_150)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_150),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_151),
.A2(n_152),
.B1(n_157),
.B2(n_128),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_127),
.A2(n_119),
.B1(n_107),
.B2(n_103),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_139),
.B(n_81),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_153),
.B(n_134),
.C(n_132),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_155),
.A2(n_21),
.B(n_22),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_139),
.A2(n_13),
.B1(n_22),
.B2(n_12),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_158),
.B(n_166),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_147),
.B(n_136),
.C(n_130),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_159),
.B(n_160),
.C(n_167),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_145),
.B(n_130),
.C(n_138),
.Y(n_160)
);

AOI31xp33_ASAP7_75t_L g162 ( 
.A1(n_150),
.A2(n_143),
.A3(n_129),
.B(n_16),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_162),
.B(n_163),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_153),
.B(n_128),
.C(n_32),
.Y(n_163)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_164),
.Y(n_169)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_149),
.Y(n_166)
);

MAJx2_ASAP7_75t_L g167 ( 
.A(n_155),
.B(n_17),
.C(n_18),
.Y(n_167)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_168),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_161),
.A2(n_148),
.B1(n_144),
.B2(n_154),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_170),
.B(n_173),
.Y(n_180)
);

OAI22xp33_ASAP7_75t_L g171 ( 
.A1(n_167),
.A2(n_146),
.B1(n_156),
.B2(n_152),
.Y(n_171)
);

AOI21x1_ASAP7_75t_SL g178 ( 
.A1(n_171),
.A2(n_57),
.B(n_37),
.Y(n_178)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_159),
.Y(n_173)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_160),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_176),
.B(n_8),
.Y(n_184)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_178),
.Y(n_188)
);

A2O1A1O1Ixp25_ASAP7_75t_L g179 ( 
.A1(n_172),
.A2(n_165),
.B(n_3),
.C(n_4),
.D(n_7),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_179),
.B(n_181),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_177),
.B(n_32),
.C(n_12),
.Y(n_181)
);

XNOR2x1_ASAP7_75t_L g182 ( 
.A(n_177),
.B(n_3),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_182),
.B(n_174),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_175),
.B(n_26),
.C(n_3),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_183),
.B(n_184),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_185),
.B(n_186),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_180),
.B(n_169),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_189),
.B(n_8),
.Y(n_191)
);

OAI21x1_ASAP7_75t_L g190 ( 
.A1(n_185),
.A2(n_184),
.B(n_171),
.Y(n_190)
);

AOI322xp5_ASAP7_75t_L g195 ( 
.A1(n_190),
.A2(n_0),
.A3(n_26),
.B1(n_41),
.B2(n_61),
.C1(n_188),
.C2(n_162),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_191),
.B(n_192),
.C(n_193),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_187),
.A2(n_61),
.B(n_9),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_195),
.A2(n_41),
.B(n_26),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_196),
.Y(n_197)
);

HB1xp67_ASAP7_75t_L g198 ( 
.A(n_197),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_198),
.B(n_194),
.Y(n_199)
);


endmodule