module fake_jpeg_9027_n_340 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_340);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_340;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_SL g17 ( 
.A(n_10),
.Y(n_17)
);

BUFx12_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

INVx2_ASAP7_75t_SL g19 ( 
.A(n_13),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_0),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_5),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_38),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_39),
.Y(n_55)
);

INVx4_ASAP7_75t_SL g40 ( 
.A(n_26),
.Y(n_40)
);

INVx3_ASAP7_75t_SL g49 ( 
.A(n_40),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_19),
.B(n_16),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_41),
.B(n_42),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_19),
.B(n_16),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

INVx4_ASAP7_75t_SL g62 ( 
.A(n_43),
.Y(n_62)
);

BUFx12_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

INVx13_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_22),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_45),
.A2(n_19),
.B1(n_22),
.B2(n_32),
.Y(n_53)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_46),
.B(n_47),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_24),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_26),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_48),
.B(n_22),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_41),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_50),
.B(n_60),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_51),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_42),
.B(n_29),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_52),
.B(n_29),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_SL g71 ( 
.A1(n_53),
.A2(n_32),
.B(n_29),
.Y(n_71)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_57),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_44),
.B(n_25),
.Y(n_58)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_58),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_44),
.B(n_25),
.Y(n_59)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_59),
.Y(n_95)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_48),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_48),
.A2(n_32),
.B1(n_34),
.B2(n_23),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_61),
.A2(n_40),
.B1(n_19),
.B2(n_25),
.Y(n_79)
);

INVx2_ASAP7_75t_SL g63 ( 
.A(n_39),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_63),
.B(n_67),
.Y(n_84)
);

INVx6_ASAP7_75t_SL g65 ( 
.A(n_47),
.Y(n_65)
);

BUFx4f_ASAP7_75t_SL g82 ( 
.A(n_65),
.Y(n_82)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

CKINVDCx5p33_ASAP7_75t_R g68 ( 
.A(n_40),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_68),
.B(n_38),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_57),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_70),
.B(n_74),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_71),
.A2(n_20),
.B1(n_23),
.B2(n_66),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_52),
.B(n_43),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_73),
.B(n_75),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_50),
.B(n_30),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_65),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_76),
.B(n_88),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_77),
.B(n_78),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_58),
.B(n_59),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_79),
.A2(n_81),
.B1(n_67),
.B2(n_38),
.Y(n_119)
);

AO22x1_ASAP7_75t_SL g81 ( 
.A1(n_49),
.A2(n_65),
.B1(n_37),
.B2(n_38),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_49),
.B(n_20),
.Y(n_83)
);

NAND3xp33_ASAP7_75t_L g111 ( 
.A(n_83),
.B(n_78),
.C(n_77),
.Y(n_111)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_49),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_86),
.A2(n_63),
.B1(n_55),
.B2(n_66),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_60),
.A2(n_46),
.B1(n_40),
.B2(n_45),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_87),
.A2(n_62),
.B1(n_55),
.B2(n_63),
.Y(n_114)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_49),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_51),
.Y(n_89)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_89),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_56),
.B(n_39),
.C(n_44),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_90),
.B(n_55),
.C(n_39),
.Y(n_104)
);

HB1xp67_ASAP7_75t_L g91 ( 
.A(n_51),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_91),
.B(n_92),
.Y(n_110)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_61),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_61),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_93),
.B(n_96),
.Y(n_116)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_67),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_56),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_97),
.B(n_98),
.Y(n_127)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_62),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_72),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_99),
.B(n_102),
.Y(n_136)
);

NOR2x1_ASAP7_75t_L g100 ( 
.A(n_81),
.B(n_68),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_100),
.A2(n_82),
.B(n_31),
.Y(n_146)
);

FAx1_ASAP7_75t_SL g101 ( 
.A(n_73),
.B(n_68),
.CI(n_54),
.CON(n_101),
.SN(n_101)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_101),
.B(n_122),
.Y(n_132)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_84),
.Y(n_102)
);

OR2x2_ASAP7_75t_L g103 ( 
.A(n_97),
.B(n_54),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_103),
.B(n_128),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_104),
.B(n_128),
.C(n_126),
.Y(n_138)
);

OAI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_92),
.A2(n_53),
.B1(n_45),
.B2(n_60),
.Y(n_105)
);

OAI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_105),
.A2(n_108),
.B1(n_118),
.B2(n_119),
.Y(n_141)
);

NAND3xp33_ASAP7_75t_L g137 ( 
.A(n_111),
.B(n_83),
.C(n_82),
.Y(n_137)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_79),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_112),
.B(n_115),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_L g139 ( 
.A1(n_114),
.A2(n_123),
.B1(n_96),
.B2(n_80),
.Y(n_139)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_89),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_93),
.A2(n_66),
.B1(n_63),
.B2(n_62),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_90),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_120),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_121),
.A2(n_18),
.B(n_35),
.Y(n_150)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_75),
.Y(n_122)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_81),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_74),
.Y(n_124)
);

OAI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_124),
.A2(n_126),
.B1(n_21),
.B2(n_27),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_70),
.A2(n_62),
.B1(n_66),
.B2(n_37),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_125),
.A2(n_80),
.B1(n_69),
.B2(n_64),
.Y(n_143)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_83),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_77),
.B(n_37),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_112),
.A2(n_85),
.B1(n_71),
.B2(n_95),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_129),
.A2(n_134),
.B1(n_135),
.B2(n_153),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_104),
.B(n_85),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_130),
.A2(n_140),
.B(n_150),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_107),
.B(n_95),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_131),
.B(n_138),
.C(n_148),
.Y(n_164)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_116),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_133),
.B(n_142),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_123),
.A2(n_94),
.B1(n_86),
.B2(n_98),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_123),
.A2(n_76),
.B1(n_88),
.B2(n_94),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_137),
.A2(n_146),
.B(n_156),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_L g173 ( 
.A1(n_139),
.A2(n_143),
.B1(n_109),
.B2(n_127),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_110),
.A2(n_82),
.B(n_39),
.Y(n_140)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_116),
.Y(n_142)
);

OAI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_147),
.A2(n_27),
.B1(n_35),
.B2(n_33),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_SL g148 ( 
.A(n_107),
.B(n_82),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_110),
.A2(n_69),
.B1(n_64),
.B2(n_31),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_149),
.A2(n_106),
.B1(n_99),
.B2(n_127),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_122),
.B(n_117),
.C(n_124),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_152),
.B(n_44),
.C(n_36),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_119),
.A2(n_69),
.B1(n_64),
.B2(n_21),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_109),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_154),
.B(n_30),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_100),
.A2(n_69),
.B1(n_64),
.B2(n_34),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_155),
.A2(n_125),
.B1(n_106),
.B2(n_102),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_117),
.B(n_0),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_145),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_157),
.B(n_158),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_136),
.Y(n_158)
);

INVx2_ASAP7_75t_SL g159 ( 
.A(n_154),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_159),
.B(n_171),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_132),
.B(n_103),
.Y(n_160)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_160),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_144),
.A2(n_113),
.B1(n_115),
.B2(n_100),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_161),
.A2(n_173),
.B1(n_176),
.B2(n_181),
.Y(n_204)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_145),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_163),
.B(n_167),
.Y(n_188)
);

OA21x2_ASAP7_75t_L g165 ( 
.A1(n_133),
.A2(n_121),
.B(n_101),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_165),
.A2(n_151),
.B(n_156),
.Y(n_195)
);

MAJx2_ASAP7_75t_L g166 ( 
.A(n_132),
.B(n_111),
.C(n_101),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_166),
.B(n_182),
.C(n_148),
.Y(n_197)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_136),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_135),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_168),
.B(n_177),
.Y(n_192)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_143),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_172),
.A2(n_179),
.B1(n_183),
.B2(n_171),
.Y(n_208)
);

INVx1_ASAP7_75t_SL g174 ( 
.A(n_151),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_174),
.B(n_187),
.Y(n_214)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_134),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_131),
.B(n_103),
.Y(n_178)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_178),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_144),
.A2(n_101),
.B1(n_114),
.B2(n_113),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_149),
.B(n_36),
.Y(n_180)
);

CKINVDCx14_ASAP7_75t_R g194 ( 
.A(n_180),
.Y(n_194)
);

OAI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_142),
.A2(n_33),
.B1(n_26),
.B2(n_34),
.Y(n_183)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_184),
.Y(n_198)
);

A2O1A1O1Ixp25_ASAP7_75t_L g185 ( 
.A1(n_137),
.A2(n_36),
.B(n_30),
.C(n_28),
.D(n_24),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_185),
.B(n_153),
.Y(n_209)
);

BUFx16f_ASAP7_75t_L g186 ( 
.A(n_140),
.Y(n_186)
);

INVx4_ASAP7_75t_L g191 ( 
.A(n_186),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_129),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_168),
.A2(n_141),
.B1(n_150),
.B2(n_146),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_190),
.A2(n_195),
.B(n_212),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_174),
.B(n_152),
.Y(n_196)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_196),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_197),
.B(n_202),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_169),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_199),
.B(n_209),
.Y(n_235)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_169),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_200),
.B(n_213),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_160),
.B(n_156),
.Y(n_201)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_201),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_164),
.B(n_138),
.C(n_148),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_187),
.A2(n_130),
.B1(n_155),
.B2(n_146),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_205),
.A2(n_179),
.B1(n_172),
.B2(n_186),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_164),
.B(n_130),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_206),
.B(n_207),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_182),
.B(n_130),
.C(n_156),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_208),
.A2(n_28),
.B1(n_18),
.B2(n_16),
.Y(n_237)
);

A2O1A1O1Ixp25_ASAP7_75t_L g211 ( 
.A1(n_166),
.A2(n_36),
.B(n_30),
.C(n_28),
.D(n_24),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_211),
.B(n_185),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_170),
.A2(n_36),
.B(n_30),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_178),
.B(n_36),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_170),
.A2(n_24),
.B(n_28),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_215),
.A2(n_18),
.B(n_28),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_158),
.B(n_18),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_216),
.B(n_0),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_162),
.B(n_30),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_217),
.B(n_184),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_219),
.B(n_223),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_192),
.A2(n_177),
.B1(n_175),
.B2(n_176),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_220),
.A2(n_222),
.B1(n_225),
.B2(n_232),
.Y(n_246)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_221),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_205),
.A2(n_186),
.B1(n_157),
.B2(n_163),
.Y(n_222)
);

INVxp33_ASAP7_75t_L g223 ( 
.A(n_203),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_214),
.A2(n_165),
.B1(n_175),
.B2(n_162),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_200),
.B(n_167),
.Y(n_226)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_226),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_189),
.B(n_165),
.Y(n_229)
);

CKINVDCx14_ASAP7_75t_R g262 ( 
.A(n_229),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_230),
.B(n_206),
.Y(n_253)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_210),
.Y(n_231)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_231),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_189),
.A2(n_159),
.B1(n_34),
.B2(n_33),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_188),
.B(n_198),
.Y(n_233)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_233),
.Y(n_247)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_188),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_234),
.B(n_239),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_192),
.A2(n_159),
.B1(n_33),
.B2(n_2),
.Y(n_236)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_236),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_237),
.A2(n_241),
.B1(n_194),
.B2(n_191),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_208),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g265 ( 
.A1(n_240),
.A2(n_215),
.B(n_212),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_191),
.A2(n_28),
.B1(n_1),
.B2(n_2),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_243),
.B(n_244),
.Y(n_254)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_201),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_236),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_248),
.B(n_259),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_252),
.A2(n_241),
.B1(n_240),
.B2(n_211),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_253),
.B(n_230),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_225),
.B(n_202),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_255),
.B(n_260),
.C(n_266),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_234),
.B(n_198),
.Y(n_256)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_256),
.Y(n_272)
);

HB1xp67_ASAP7_75t_L g258 ( 
.A(n_231),
.Y(n_258)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_258),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_232),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_228),
.B(n_227),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_239),
.A2(n_190),
.B1(n_193),
.B2(n_204),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_261),
.A2(n_222),
.B1(n_221),
.B2(n_242),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_218),
.B(n_193),
.Y(n_264)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_264),
.Y(n_281)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_265),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_227),
.B(n_197),
.C(n_207),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_267),
.A2(n_268),
.B1(n_257),
.B2(n_263),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_246),
.A2(n_242),
.B1(n_224),
.B2(n_244),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_245),
.A2(n_220),
.B1(n_262),
.B2(n_218),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_269),
.A2(n_280),
.B1(n_265),
.B2(n_257),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_254),
.B(n_224),
.Y(n_271)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_271),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_260),
.B(n_238),
.C(n_228),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_275),
.B(n_278),
.C(n_253),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_250),
.B(n_229),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_276),
.B(n_282),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_SL g277 ( 
.A(n_255),
.B(n_195),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_277),
.B(n_279),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_266),
.B(n_238),
.C(n_196),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_249),
.A2(n_235),
.B(n_217),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g282 ( 
.A(n_249),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_284),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_286),
.B(n_287),
.C(n_288),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_270),
.B(n_256),
.C(n_264),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_270),
.B(n_246),
.C(n_247),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_289),
.A2(n_298),
.B1(n_281),
.B2(n_274),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_278),
.B(n_247),
.C(n_261),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_290),
.B(n_292),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_291),
.B(n_1),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_275),
.B(n_251),
.C(n_252),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_269),
.B(n_254),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_293),
.B(n_295),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_277),
.B(n_279),
.C(n_280),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_267),
.A2(n_209),
.B1(n_213),
.B2(n_15),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_283),
.B(n_15),
.C(n_14),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_299),
.B(n_12),
.C(n_11),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_296),
.A2(n_268),
.B1(n_282),
.B2(n_272),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_301),
.B(n_308),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_287),
.B(n_273),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_302),
.B(n_303),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_286),
.B(n_271),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_304),
.A2(n_311),
.B1(n_294),
.B2(n_4),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_306),
.B(n_310),
.Y(n_313)
);

MAJx2_ASAP7_75t_L g307 ( 
.A(n_285),
.B(n_14),
.C(n_13),
.Y(n_307)
);

OAI21x1_ASAP7_75t_L g321 ( 
.A1(n_307),
.A2(n_4),
.B(n_5),
.Y(n_321)
);

XNOR2x1_ASAP7_75t_L g310 ( 
.A(n_296),
.B(n_1),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_288),
.A2(n_12),
.B1(n_11),
.B2(n_3),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_297),
.B(n_1),
.C(n_2),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_L g316 ( 
.A1(n_312),
.A2(n_3),
.B(n_4),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_314),
.B(n_319),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_316),
.B(n_320),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_300),
.B(n_285),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_318),
.B(n_300),
.C(n_305),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_312),
.B(n_18),
.Y(n_319)
);

OR2x2_ASAP7_75t_L g320 ( 
.A(n_310),
.B(n_3),
.Y(n_320)
);

INVxp33_ASAP7_75t_SL g325 ( 
.A(n_321),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_306),
.B(n_4),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_322),
.B(n_308),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_315),
.B(n_309),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_323),
.B(n_326),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_SL g330 ( 
.A(n_328),
.B(n_329),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_317),
.B(n_307),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_325),
.A2(n_313),
.B1(n_318),
.B2(n_320),
.Y(n_331)
);

AOI21xp5_ASAP7_75t_L g335 ( 
.A1(n_331),
.A2(n_332),
.B(n_5),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_SL g332 ( 
.A(n_324),
.B(n_313),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_SL g334 ( 
.A1(n_333),
.A2(n_327),
.B(n_6),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_334),
.B(n_335),
.Y(n_336)
);

OAI321xp33_ASAP7_75t_L g337 ( 
.A1(n_336),
.A2(n_7),
.A3(n_8),
.B1(n_9),
.B2(n_330),
.C(n_335),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_337),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_338)
);

AOI21xp5_ASAP7_75t_L g339 ( 
.A1(n_338),
.A2(n_9),
.B(n_7),
.Y(n_339)
);

AOI21xp5_ASAP7_75t_L g340 ( 
.A1(n_339),
.A2(n_8),
.B(n_9),
.Y(n_340)
);


endmodule