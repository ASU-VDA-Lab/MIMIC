module fake_jpeg_20300_n_345 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_345);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_345;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_15),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_16),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

BUFx8_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

INVx8_ASAP7_75t_SL g32 ( 
.A(n_3),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_16),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_26),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_41),
.B(n_47),
.Y(n_66)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_23),
.Y(n_46)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_17),
.B(n_8),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_23),
.Y(n_49)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_37),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_51),
.B(n_18),
.Y(n_86)
);

BUFx4f_ASAP7_75t_SL g56 ( 
.A(n_38),
.Y(n_56)
);

BUFx2_ASAP7_75t_L g100 ( 
.A(n_56),
.Y(n_100)
);

BUFx12_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVx4_ASAP7_75t_SL g93 ( 
.A(n_59),
.Y(n_93)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_62),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_41),
.B(n_22),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_63),
.B(n_38),
.Y(n_96)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_67),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_51),
.A2(n_43),
.B1(n_54),
.B2(n_57),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g131 ( 
.A1(n_68),
.A2(n_80),
.B1(n_39),
.B2(n_35),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_66),
.B(n_47),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_69),
.B(n_85),
.Y(n_121)
);

AOI21xp33_ASAP7_75t_L g70 ( 
.A1(n_63),
.A2(n_37),
.B(n_32),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_70),
.A2(n_35),
.B(n_24),
.Y(n_113)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_71),
.Y(n_109)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_60),
.Y(n_72)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_72),
.Y(n_115)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_52),
.Y(n_74)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_74),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_57),
.A2(n_43),
.B1(n_18),
.B2(n_21),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_75),
.A2(n_89),
.B1(n_36),
.B2(n_24),
.Y(n_116)
);

OAI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_58),
.A2(n_43),
.B1(n_48),
.B2(n_45),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_76),
.A2(n_44),
.B1(n_42),
.B2(n_55),
.Y(n_102)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_60),
.Y(n_78)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_78),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_53),
.B(n_44),
.C(n_40),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_79),
.B(n_46),
.C(n_39),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_58),
.A2(n_48),
.B1(n_45),
.B2(n_42),
.Y(n_80)
);

HB1xp67_ASAP7_75t_L g81 ( 
.A(n_59),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_81),
.Y(n_129)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_53),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_82),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_64),
.B(n_38),
.Y(n_83)
);

FAx1_ASAP7_75t_SL g107 ( 
.A(n_83),
.B(n_59),
.CI(n_29),
.CON(n_107),
.SN(n_107)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_65),
.Y(n_84)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_84),
.Y(n_122)
);

OR2x2_ASAP7_75t_L g85 ( 
.A(n_50),
.B(n_21),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_86),
.B(n_94),
.Y(n_106)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_61),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_87),
.B(n_90),
.Y(n_110)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_50),
.Y(n_88)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_88),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_65),
.A2(n_17),
.B1(n_34),
.B2(n_36),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_67),
.B(n_34),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_55),
.Y(n_91)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_91),
.Y(n_133)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_61),
.Y(n_92)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_92),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_64),
.B(n_26),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_55),
.Y(n_95)
);

INVxp67_ASAP7_75t_SL g119 ( 
.A(n_95),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_96),
.B(n_49),
.Y(n_108)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_52),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_97),
.B(n_98),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_56),
.B(n_27),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_56),
.B(n_28),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_99),
.Y(n_132)
);

BUFx12f_ASAP7_75t_L g101 ( 
.A(n_52),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_101),
.A2(n_62),
.B1(n_59),
.B2(n_52),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_102),
.B(n_77),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_96),
.B(n_32),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_104),
.B(n_113),
.Y(n_155)
);

INVx13_ASAP7_75t_L g149 ( 
.A(n_105),
.Y(n_149)
);

NAND2xp67_ASAP7_75t_L g138 ( 
.A(n_107),
.B(n_83),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_108),
.B(n_114),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_71),
.B(n_70),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_116),
.B(n_131),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_79),
.A2(n_49),
.B1(n_46),
.B2(n_39),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_118),
.A2(n_73),
.B1(n_74),
.B2(n_77),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_88),
.A2(n_36),
.B1(n_27),
.B2(n_28),
.Y(n_123)
);

AOI21xp33_ASAP7_75t_L g148 ( 
.A1(n_123),
.A2(n_128),
.B(n_29),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_125),
.B(n_126),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_84),
.B(n_49),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_83),
.A2(n_0),
.B(n_1),
.Y(n_127)
);

NOR3xp33_ASAP7_75t_L g160 ( 
.A(n_127),
.B(n_25),
.C(n_20),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_93),
.A2(n_35),
.B1(n_20),
.B2(n_25),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_85),
.B(n_46),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_130),
.B(n_95),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_130),
.B(n_78),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_136),
.B(n_137),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_121),
.B(n_87),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_138),
.A2(n_148),
.B(n_152),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_108),
.A2(n_82),
.B1(n_92),
.B2(n_72),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_139),
.A2(n_142),
.B1(n_143),
.B2(n_145),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_121),
.B(n_132),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_140),
.B(n_144),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_114),
.A2(n_113),
.B1(n_126),
.B2(n_125),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_109),
.A2(n_73),
.B1(n_93),
.B2(n_91),
.Y(n_143)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_103),
.Y(n_146)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_146),
.Y(n_170)
);

AND2x6_ASAP7_75t_L g147 ( 
.A(n_107),
.B(n_100),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_147),
.B(n_159),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_106),
.B(n_15),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_150),
.B(n_156),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_132),
.B(n_100),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_151),
.B(n_154),
.Y(n_182)
);

OAI21xp33_ASAP7_75t_L g152 ( 
.A1(n_106),
.A2(n_97),
.B(n_14),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_122),
.Y(n_153)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_153),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_104),
.B(n_109),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_110),
.B(n_13),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_157),
.A2(n_118),
.B1(n_133),
.B2(n_124),
.Y(n_166)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_122),
.Y(n_158)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_158),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_127),
.B(n_22),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_160),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_111),
.B(n_22),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_161),
.B(n_101),
.Y(n_192)
);

OAI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_147),
.A2(n_116),
.B1(n_102),
.B2(n_120),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_164),
.A2(n_169),
.B1(n_173),
.B2(n_177),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_147),
.A2(n_129),
.B(n_115),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_165),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_166),
.B(n_150),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_155),
.B(n_107),
.C(n_129),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_167),
.B(n_161),
.C(n_137),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_135),
.A2(n_133),
.B1(n_115),
.B2(n_120),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_153),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_171),
.B(n_179),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_155),
.B(n_117),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_172),
.B(n_149),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_135),
.A2(n_145),
.B1(n_144),
.B2(n_141),
.Y(n_173)
);

INVx2_ASAP7_75t_SL g174 ( 
.A(n_146),
.Y(n_174)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_174),
.Y(n_198)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_158),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_175),
.B(n_191),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_142),
.A2(n_117),
.B1(n_124),
.B2(n_119),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_157),
.A2(n_103),
.B1(n_112),
.B2(n_12),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_178),
.A2(n_183),
.B1(n_188),
.B2(n_0),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_140),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_141),
.A2(n_112),
.B1(n_33),
.B2(n_30),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_139),
.Y(n_184)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_184),
.Y(n_208)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_136),
.Y(n_185)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_185),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_134),
.A2(n_112),
.B1(n_33),
.B2(n_30),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_134),
.A2(n_19),
.B(n_25),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_189),
.A2(n_193),
.B(n_0),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g191 ( 
.A(n_151),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_192),
.B(n_149),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_159),
.A2(n_19),
.B(n_20),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_194),
.B(n_201),
.Y(n_228)
);

O2A1O1Ixp33_ASAP7_75t_L g195 ( 
.A1(n_179),
.A2(n_138),
.B(n_154),
.C(n_143),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_195),
.B(n_203),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_196),
.A2(n_204),
.B1(n_215),
.B2(n_221),
.Y(n_230)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_174),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_197),
.B(n_218),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_172),
.B(n_101),
.C(n_156),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_180),
.B(n_31),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_167),
.A2(n_149),
.B1(n_33),
.B2(n_30),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_206),
.B(n_214),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_176),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_207),
.B(n_216),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_180),
.B(n_31),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_209),
.B(n_210),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_185),
.B(n_31),
.Y(n_210)
);

HB1xp67_ASAP7_75t_L g212 ( 
.A(n_165),
.Y(n_212)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_212),
.Y(n_242)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_176),
.Y(n_213)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_213),
.Y(n_233)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_181),
.Y(n_217)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_217),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_182),
.B(n_33),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_190),
.B(n_8),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_219),
.B(n_222),
.Y(n_241)
);

MAJx2_ASAP7_75t_L g220 ( 
.A(n_168),
.B(n_30),
.C(n_8),
.Y(n_220)
);

XNOR2x1_ASAP7_75t_L g227 ( 
.A(n_220),
.B(n_168),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_173),
.A2(n_7),
.B1(n_13),
.B2(n_11),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_174),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_182),
.B(n_16),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_223),
.B(n_224),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_183),
.B(n_11),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_187),
.B(n_10),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_225),
.B(n_194),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_227),
.A2(n_215),
.B1(n_220),
.B2(n_202),
.Y(n_263)
);

NOR2x1_ASAP7_75t_L g231 ( 
.A(n_200),
.B(n_171),
.Y(n_231)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_231),
.Y(n_256)
);

AOI32xp33_ASAP7_75t_L g236 ( 
.A1(n_202),
.A2(n_186),
.A3(n_189),
.B1(n_177),
.B2(n_184),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_236),
.B(n_237),
.Y(n_270)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_205),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_238),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_196),
.A2(n_163),
.B1(n_186),
.B2(n_166),
.Y(n_239)
);

CKINVDCx14_ASAP7_75t_R g262 ( 
.A(n_239),
.Y(n_262)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_211),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_240),
.Y(n_254)
);

BUFx2_ASAP7_75t_L g243 ( 
.A(n_197),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_243),
.Y(n_258)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_198),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_244),
.Y(n_269)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_198),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_245),
.B(n_251),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_208),
.A2(n_169),
.B1(n_163),
.B2(n_188),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_248),
.A2(n_199),
.B1(n_204),
.B2(n_178),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_210),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_249),
.Y(n_260)
);

AND2x2_ASAP7_75t_L g250 ( 
.A(n_214),
.B(n_181),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_L g264 ( 
.A1(n_250),
.A2(n_195),
.B(n_162),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_203),
.B(n_162),
.Y(n_251)
);

BUFx2_ASAP7_75t_L g252 ( 
.A(n_230),
.Y(n_252)
);

CKINVDCx14_ASAP7_75t_R g283 ( 
.A(n_252),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_228),
.B(n_201),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_255),
.B(n_263),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_257),
.A2(n_226),
.B1(n_231),
.B2(n_242),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_228),
.B(n_209),
.C(n_199),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_259),
.B(n_265),
.C(n_268),
.Y(n_278)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_264),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_237),
.B(n_206),
.C(n_225),
.Y(n_265)
);

CKINVDCx16_ASAP7_75t_R g266 ( 
.A(n_247),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_266),
.B(n_229),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_226),
.A2(n_175),
.B1(n_222),
.B2(n_221),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_267),
.B(n_248),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_250),
.B(n_193),
.C(n_170),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_250),
.B(n_170),
.C(n_10),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_271),
.B(n_272),
.C(n_246),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_234),
.B(n_9),
.C(n_7),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_261),
.Y(n_273)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_273),
.Y(n_302)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_274),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_275),
.A2(n_284),
.B1(n_269),
.B2(n_254),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g277 ( 
.A1(n_256),
.A2(n_264),
.B(n_262),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_277),
.Y(n_292)
);

XOR2x2_ASAP7_75t_L g279 ( 
.A(n_270),
.B(n_227),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_SL g298 ( 
.A1(n_279),
.A2(n_269),
.B(n_235),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_256),
.B(n_245),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_281),
.B(n_282),
.Y(n_300)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_261),
.Y(n_282)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_267),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_285),
.B(n_286),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_253),
.B(n_241),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_255),
.B(n_234),
.C(n_244),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_287),
.B(n_289),
.Y(n_306)
);

CKINVDCx16_ASAP7_75t_R g288 ( 
.A(n_257),
.Y(n_288)
);

BUFx2_ASAP7_75t_L g307 ( 
.A(n_288),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_259),
.B(n_238),
.C(n_251),
.Y(n_289)
);

NOR3xp33_ASAP7_75t_SL g290 ( 
.A(n_253),
.B(n_232),
.C(n_240),
.Y(n_290)
);

NOR3xp33_ASAP7_75t_L g294 ( 
.A(n_290),
.B(n_260),
.C(n_254),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_291),
.B(n_229),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_293),
.B(n_297),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_294),
.B(n_281),
.Y(n_308)
);

A2O1A1O1Ixp25_ASAP7_75t_L g295 ( 
.A1(n_279),
.A2(n_268),
.B(n_265),
.C(n_271),
.D(n_252),
.Y(n_295)
);

HB1xp67_ASAP7_75t_L g311 ( 
.A(n_295),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_280),
.B(n_272),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_296),
.B(n_298),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_278),
.B(n_235),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_301),
.B(n_303),
.C(n_287),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_278),
.B(n_233),
.Y(n_303)
);

AOI222xp33_ASAP7_75t_SL g304 ( 
.A1(n_276),
.A2(n_233),
.B1(n_258),
.B2(n_243),
.C1(n_7),
.C2(n_5),
.Y(n_304)
);

HB1xp67_ASAP7_75t_L g319 ( 
.A(n_304),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_308),
.Y(n_320)
);

BUFx6f_ASAP7_75t_L g309 ( 
.A(n_304),
.Y(n_309)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_309),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_294),
.B(n_275),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_310),
.B(n_314),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_299),
.B(n_289),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_292),
.A2(n_283),
.B1(n_284),
.B2(n_305),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_L g327 ( 
.A1(n_315),
.A2(n_282),
.B1(n_274),
.B2(n_295),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_316),
.B(n_296),
.C(n_312),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_306),
.B(n_280),
.C(n_285),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_317),
.B(n_318),
.Y(n_323)
);

INVx1_ASAP7_75t_SL g318 ( 
.A(n_302),
.Y(n_318)
);

AND2x2_ASAP7_75t_L g331 ( 
.A(n_321),
.B(n_290),
.Y(n_331)
);

AOI21xp5_ASAP7_75t_L g322 ( 
.A1(n_311),
.A2(n_292),
.B(n_277),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_322),
.B(n_325),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_311),
.A2(n_276),
.B(n_300),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_327),
.B(n_309),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_313),
.B(n_258),
.C(n_307),
.Y(n_328)
);

OR2x2_ASAP7_75t_L g333 ( 
.A(n_328),
.B(n_319),
.Y(n_333)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_330),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_SL g336 ( 
.A1(n_331),
.A2(n_333),
.B(n_334),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_320),
.A2(n_319),
.B1(n_307),
.B2(n_3),
.Y(n_332)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_332),
.Y(n_338)
);

A2O1A1Ixp33_ASAP7_75t_SL g334 ( 
.A1(n_324),
.A2(n_0),
.B(n_2),
.C(n_3),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_SL g335 ( 
.A1(n_323),
.A2(n_2),
.B(n_3),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_336),
.B(n_321),
.C(n_326),
.Y(n_339)
);

AOI322xp5_ASAP7_75t_L g340 ( 
.A1(n_339),
.A2(n_337),
.A3(n_335),
.B1(n_338),
.B2(n_329),
.C1(n_328),
.C2(n_334),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_340),
.B(n_2),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_341),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_342),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_343)
);

AOI21xp5_ASAP7_75t_L g344 ( 
.A1(n_343),
.A2(n_4),
.B(n_6),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g345 ( 
.A(n_344),
.B(n_4),
.Y(n_345)
);


endmodule