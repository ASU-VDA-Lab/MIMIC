module real_aes_16131_n_234 (n_17, n_28, n_226, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_230, n_165, n_51, n_195, n_176, n_27, n_163, n_222, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_86, n_93, n_182, n_154, n_127, n_199, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_38, n_155, n_118, n_143, n_139, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_107, n_184, n_53, n_36, n_234);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_230;
input n_165;
input n_51;
input n_195;
input n_176;
input n_27;
input n_163;
input n_222;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_38;
input n_155;
input n_118;
input n_143;
input n_139;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_107;
input n_184;
input n_53;
input n_36;
output n_234;
wire n_476;
wire n_599;
wire n_887;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_254;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_239;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_1423;
wire n_571;
wire n_549;
wire n_1034;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_260;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_870;
wire n_1248;
wire n_271;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_292;
wire n_1379;
wire n_400;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_553;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1382;
wire n_1225;
wire n_875;
wire n_951;
wire n_1199;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_281;
wire n_962;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_455;
wire n_682;
wire n_812;
wire n_817;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_363;
wire n_1317;
wire n_417;
wire n_323;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_947;
wire n_970;
wire n_1149;
wire n_368;
wire n_527;
wire n_1342;
wire n_552;
wire n_1346;
wire n_1383;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_805;
wire n_238;
wire n_619;
wire n_1095;
wire n_1284;
wire n_1250;
wire n_360;
wire n_859;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_246;
wire n_1247;
wire n_501;
wire n_488;
wire n_1380;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_404;
wire n_1073;
wire n_728;
wire n_1301;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_306;
wire n_1003;
wire n_346;
wire n_293;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_648;
wire n_939;
wire n_290;
wire n_928;
wire n_1384;
wire n_789;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_712;
wire n_266;
wire n_422;
wire n_861;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_258;
wire n_652;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_337;
wire n_247;
wire n_264;
wire n_237;
wire n_480;
wire n_684;
wire n_1178;
wire n_821;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_635;
wire n_792;
wire n_1392;
wire n_665;
wire n_991;
wire n_667;
wire n_580;
wire n_1004;
wire n_1370;
wire n_1417;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_328;
wire n_1260;
wire n_355;
wire n_1129;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_461;
wire n_1047;
wire n_1016;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_401;
wire n_538;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_704;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_948;
wire n_700;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_245;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1406;
wire n_550;
wire n_966;
wire n_333;
wire n_1368;
wire n_994;
wire n_384;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1401;
wire n_248;
wire n_1086;
wire n_1189;
wire n_1070;
wire n_535;
wire n_882;
wire n_1210;
wire n_746;
wire n_656;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_651;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_311;
wire n_278;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_277;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_1408;
wire n_428;
wire n_783;
wire n_1107;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1386;
wire n_406;
wire n_617;
wire n_733;
wire n_402;
wire n_1404;
wire n_602;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_255;
wire n_286;
wire n_1011;
wire n_416;
wire n_895;
wire n_799;
wire n_490;
wire n_261;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_645;
wire n_1145;
wire n_557;
wire n_777;
wire n_985;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_296;
wire n_1347;
wire n_1163;
wire n_1278;
wire n_734;
wire n_735;
wire n_334;
wire n_1179;
wire n_1171;
wire n_569;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_1026;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_643;
wire n_1403;
wire n_486;
wire n_291;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_268;
wire n_1194;
wire n_282;
wire n_389;
wire n_701;
wire n_809;
wire n_679;
wire n_520;
wire n_926;
wire n_942;
wire n_1374;
wire n_1120;
wire n_689;
wire n_946;
wire n_300;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_249;
wire n_1032;
wire n_1431;
wire n_721;
wire n_1133;
wire n_313;
wire n_739;
wire n_1322;
wire n_1162;
wire n_762;
wire n_325;
wire n_1298;
wire n_442;
wire n_740;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_253;
wire n_1172;
wire n_459;
wire n_998;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_279;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_473;
wire n_967;
wire n_1159;
wire n_474;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_307;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_257;
wire n_285;
wire n_1377;
wire n_800;
wire n_1175;
wire n_778;
wire n_1170;
wire n_522;
wire n_943;
wire n_977;
wire n_287;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1333;
wire n_577;
wire n_759;
wire n_1235;
wire n_299;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_766;
wire n_852;
wire n_1113;
wire n_1268;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_773;
wire n_353;
wire n_865;
wire n_594;
wire n_856;
wire n_1146;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_816;
wire n_625;
wire n_953;
wire n_289;
wire n_1373;
wire n_716;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_370;
wire n_352;
wire n_935;
wire n_467;
wire n_1213;
wire n_1053;
wire n_263;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_284;
wire n_316;
wire n_1168;
wire n_1309;
wire n_909;
wire n_996;
wire n_523;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1263;
wire n_1411;
wire n_1115;
wire n_310;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_1303;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_324;
wire n_664;
wire n_367;
wire n_267;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1414;
wire n_502;
wire n_434;
wire n_769;
wire n_250;
wire n_1212;
wire n_1054;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1134;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_251;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_945;
wire n_392;
wire n_288;
wire n_274;
wire n_303;
wire n_563;
wire n_891;
wire n_568;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1028;
wire n_366;
wire n_1083;
wire n_727;
wire n_397;
wire n_1056;
wire n_663;
wire n_588;
wire n_707;
wire n_915;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_273;
wire n_1038;
wire n_276;
wire n_1085;
wire n_295;
wire n_845;
wire n_1127;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_697;
wire n_978;
wire n_847;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_243;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1355;
wire n_309;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_262;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_252;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_1378;
wire n_524;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_525;
wire n_1226;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_929;
wire n_1143;
wire n_1190;
wire n_543;
wire n_305;
wire n_585;
wire n_465;
wire n_719;
wire n_1343;
wire n_1156;
wire n_988;
wire n_921;
wire n_1396;
wire n_640;
wire n_1176;
wire n_1151;
wire n_1254;
wire n_241;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1407;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1420;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1240;
wire n_987;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_319;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_242;
wire n_376;
wire n_308;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_460;
wire n_317;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_489;
wire n_1381;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_280;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_408;
wire n_372;
wire n_578;
wire n_892;
wire n_938;
wire n_327;
wire n_774;
wire n_466;
wire n_559;
wire n_1049;
wire n_1277;
wire n_984;
wire n_301;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_532;
wire n_1025;
wire n_298;
wire n_924;
wire n_1264;
wire n_297;
wire n_1245;
wire n_1152;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_304;
wire n_1307;
wire n_993;
wire n_236;
wire n_819;
wire n_737;
wire n_1290;
wire n_1318;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_425;
wire n_879;
wire n_331;
wire n_449;
wire n_1340;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_655;
wire n_654;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1334;
wire n_244;
wire n_1291;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1356;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1249;
wire n_1416;
wire n_387;
wire n_1239;
wire n_969;
wire n_256;
wire n_1009;
wire n_1202;
wire n_302;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_269;
wire n_430;
wire n_1252;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_385;
wire n_275;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1043;
wire n_435;
wire n_511;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1430;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1087;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1130;
wire n_794;
wire n_283;
wire n_314;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1253;
wire n_312;
wire n_1183;
wire n_335;
wire n_516;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_338;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_793;
wire n_1390;
wire n_272;
wire n_1412;
wire n_757;
wire n_803;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_340;
wire n_483;
wire n_394;
wire n_729;
wire n_1280;
wire n_1352;
wire n_1323;
wire n_703;
wire n_1097;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_342;
wire n_348;
wire n_603;
wire n_1288;
wire n_868;
wire n_240;
wire n_1024;
wire n_259;
wire n_1144;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_429;
AOI22xp5_ASAP7_75t_L g1224 ( .A1(n_0), .A2(n_178), .B1(n_1168), .B2(n_1172), .Y(n_1224) );
OAI22xp5_ASAP7_75t_L g641 ( .A1(n_1), .A2(n_71), .B1(n_642), .B2(n_644), .Y(n_641) );
OAI22xp33_ASAP7_75t_SL g681 ( .A1(n_1), .A2(n_229), .B1(n_682), .B2(n_684), .Y(n_681) );
CKINVDCx5p33_ASAP7_75t_R g459 ( .A(n_2), .Y(n_459) );
INVx1_ASAP7_75t_L g1084 ( .A(n_3), .Y(n_1084) );
AOI221xp5_ASAP7_75t_L g1122 ( .A1(n_4), .A2(n_181), .B1(n_532), .B2(n_623), .C(n_1123), .Y(n_1122) );
INVx1_ASAP7_75t_L g1150 ( .A(n_4), .Y(n_1150) );
AOI22xp33_ASAP7_75t_L g1192 ( .A1(n_5), .A2(n_45), .B1(n_1168), .B2(n_1172), .Y(n_1192) );
INVx1_ASAP7_75t_L g1124 ( .A(n_6), .Y(n_1124) );
AOI221xp5_ASAP7_75t_L g1152 ( .A1(n_6), .A2(n_131), .B1(n_419), .B2(n_678), .C(n_1153), .Y(n_1152) );
INVx1_ASAP7_75t_L g776 ( .A(n_7), .Y(n_776) );
AOI22xp33_ASAP7_75t_L g809 ( .A1(n_7), .A2(n_103), .B1(n_409), .B2(n_810), .Y(n_809) );
INVx1_ASAP7_75t_L g621 ( .A(n_8), .Y(n_621) );
OAI221xp5_ASAP7_75t_L g767 ( .A1(n_9), .A2(n_189), .B1(n_319), .B2(n_331), .C(n_595), .Y(n_767) );
OA222x2_ASAP7_75t_L g812 ( .A1(n_9), .A2(n_42), .B1(n_192), .B2(n_724), .C1(n_731), .C2(n_813), .Y(n_812) );
OAI22xp5_ASAP7_75t_L g943 ( .A1(n_10), .A2(n_17), .B1(n_944), .B2(n_947), .Y(n_943) );
OAI22xp33_ASAP7_75t_L g975 ( .A1(n_10), .A2(n_17), .B1(n_976), .B2(n_979), .Y(n_975) );
AOI221xp5_ASAP7_75t_L g529 ( .A1(n_11), .A2(n_167), .B1(n_530), .B2(n_532), .C(n_533), .Y(n_529) );
INVx1_ASAP7_75t_L g577 ( .A(n_11), .Y(n_577) );
INVx1_ASAP7_75t_L g249 ( .A(n_12), .Y(n_249) );
AND2x2_ASAP7_75t_L g275 ( .A(n_12), .B(n_276), .Y(n_275) );
AND2x2_ASAP7_75t_L g380 ( .A(n_12), .B(n_197), .Y(n_380) );
NOR2xp33_ASAP7_75t_L g417 ( .A(n_12), .B(n_259), .Y(n_417) );
INVx1_ASAP7_75t_L g914 ( .A(n_13), .Y(n_914) );
INVx1_ASAP7_75t_L g336 ( .A(n_14), .Y(n_336) );
AOI22xp5_ASAP7_75t_L g406 ( .A1(n_14), .A2(n_27), .B1(n_407), .B2(n_408), .Y(n_406) );
OAI22xp5_ASAP7_75t_L g698 ( .A1(n_15), .A2(n_109), .B1(n_282), .B2(n_293), .Y(n_698) );
INVxp67_ASAP7_75t_SL g743 ( .A(n_15), .Y(n_743) );
INVx2_ASAP7_75t_L g1171 ( .A(n_16), .Y(n_1171) );
AND2x2_ASAP7_75t_L g1173 ( .A(n_16), .B(n_97), .Y(n_1173) );
AND2x2_ASAP7_75t_L g1179 ( .A(n_16), .B(n_1177), .Y(n_1179) );
INVxp67_ASAP7_75t_SL g1004 ( .A(n_18), .Y(n_1004) );
AOI22xp33_ASAP7_75t_SL g1040 ( .A1(n_18), .A2(n_151), .B1(n_766), .B2(n_1041), .Y(n_1040) );
AOI22xp5_ASAP7_75t_L g1201 ( .A1(n_19), .A2(n_26), .B1(n_1175), .B2(n_1178), .Y(n_1201) );
XNOR2x2_ASAP7_75t_L g1117 ( .A(n_20), .B(n_1118), .Y(n_1117) );
INVx1_ASAP7_75t_L g709 ( .A(n_21), .Y(n_709) );
AOI22xp5_ASAP7_75t_L g1223 ( .A1(n_22), .A2(n_111), .B1(n_1175), .B2(n_1178), .Y(n_1223) );
INVx1_ASAP7_75t_L g1391 ( .A(n_23), .Y(n_1391) );
CKINVDCx5p33_ASAP7_75t_R g860 ( .A(n_24), .Y(n_860) );
AOI222xp33_ASAP7_75t_L g716 ( .A1(n_25), .A2(n_155), .B1(n_186), .B2(n_295), .C1(n_335), .C2(n_342), .Y(n_716) );
INVx1_ASAP7_75t_L g749 ( .A(n_25), .Y(n_749) );
XOR2x2_ASAP7_75t_L g987 ( .A(n_26), .B(n_988), .Y(n_987) );
INVx1_ASAP7_75t_L g359 ( .A(n_27), .Y(n_359) );
OAI22xp5_ASAP7_75t_SL g578 ( .A1(n_28), .A2(n_579), .B1(n_580), .B2(n_687), .Y(n_578) );
INVx1_ASAP7_75t_L g687 ( .A(n_28), .Y(n_687) );
AOI22xp5_ASAP7_75t_L g689 ( .A1(n_28), .A2(n_579), .B1(n_580), .B2(n_687), .Y(n_689) );
INVx1_ASAP7_75t_L g350 ( .A(n_29), .Y(n_350) );
AOI22xp33_ASAP7_75t_L g418 ( .A1(n_29), .A2(n_153), .B1(n_407), .B2(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g1125 ( .A(n_30), .Y(n_1125) );
AOI221xp5_ASAP7_75t_L g1145 ( .A1(n_30), .A2(n_69), .B1(n_1146), .B2(n_1147), .C(n_1149), .Y(n_1145) );
OAI22xp33_ASAP7_75t_L g1061 ( .A1(n_31), .A2(n_226), .B1(n_1062), .B2(n_1063), .Y(n_1061) );
OAI22xp5_ASAP7_75t_L g1107 ( .A1(n_31), .A2(n_226), .B1(n_1108), .B2(n_1110), .Y(n_1107) );
AOI22xp5_ASAP7_75t_L g1198 ( .A1(n_32), .A2(n_86), .B1(n_1168), .B2(n_1189), .Y(n_1198) );
AOI22xp33_ASAP7_75t_L g1261 ( .A1(n_33), .A2(n_96), .B1(n_1168), .B2(n_1262), .Y(n_1261) );
AOI211xp5_ASAP7_75t_L g517 ( .A1(n_34), .A2(n_518), .B(n_519), .C(n_521), .Y(n_517) );
INVx1_ASAP7_75t_L g568 ( .A(n_34), .Y(n_568) );
INVx1_ASAP7_75t_L g435 ( .A(n_35), .Y(n_435) );
OAI221xp5_ASAP7_75t_L g1135 ( .A1(n_36), .A2(n_59), .B1(n_324), .B2(n_476), .C(n_477), .Y(n_1135) );
INVxp67_ASAP7_75t_SL g1141 ( .A(n_36), .Y(n_1141) );
OAI22xp33_ASAP7_75t_L g475 ( .A1(n_37), .A2(n_146), .B1(n_476), .B2(n_477), .Y(n_475) );
OAI22xp5_ASAP7_75t_L g501 ( .A1(n_37), .A2(n_74), .B1(n_502), .B2(n_504), .Y(n_501) );
INVxp67_ASAP7_75t_SL g1000 ( .A(n_38), .Y(n_1000) );
AOI22xp33_ASAP7_75t_SL g1032 ( .A1(n_38), .A2(n_41), .B1(n_840), .B2(n_1033), .Y(n_1032) );
INVx1_ASAP7_75t_L g1087 ( .A(n_39), .Y(n_1087) );
INVx1_ASAP7_75t_L g290 ( .A(n_40), .Y(n_290) );
INVx1_ASAP7_75t_L g299 ( .A(n_40), .Y(n_299) );
AOI221xp5_ASAP7_75t_L g1007 ( .A1(n_41), .A2(n_151), .B1(n_742), .B2(n_796), .C(n_1008), .Y(n_1007) );
INVx1_ASAP7_75t_L g765 ( .A(n_42), .Y(n_765) );
AOI22xp5_ASAP7_75t_L g1188 ( .A1(n_43), .A2(n_115), .B1(n_1168), .B2(n_1189), .Y(n_1188) );
OAI221xp5_ASAP7_75t_L g514 ( .A1(n_44), .A2(n_212), .B1(n_324), .B2(n_476), .C(n_477), .Y(n_514) );
OAI22xp5_ASAP7_75t_L g548 ( .A1(n_44), .A2(n_113), .B1(n_397), .B2(n_401), .Y(n_548) );
INVx1_ASAP7_75t_L g1382 ( .A(n_46), .Y(n_1382) );
OAI221xp5_ASAP7_75t_L g588 ( .A1(n_47), .A2(n_150), .B1(n_589), .B2(n_592), .C(n_596), .Y(n_588) );
OAI211xp5_ASAP7_75t_L g647 ( .A1(n_47), .A2(n_648), .B(n_652), .C(n_662), .Y(n_647) );
OAI221xp5_ASAP7_75t_L g281 ( .A1(n_48), .A2(n_98), .B1(n_282), .B2(n_293), .C(n_300), .Y(n_281) );
INVxp67_ASAP7_75t_SL g382 ( .A(n_48), .Y(n_382) );
AOI221xp5_ASAP7_75t_L g700 ( .A1(n_49), .A2(n_138), .B1(n_701), .B2(n_703), .C(n_705), .Y(n_700) );
AOI221xp5_ASAP7_75t_L g744 ( .A1(n_49), .A2(n_191), .B1(n_745), .B2(n_747), .C(n_748), .Y(n_744) );
AOI22xp33_ASAP7_75t_L g1263 ( .A1(n_50), .A2(n_196), .B1(n_1175), .B2(n_1178), .Y(n_1263) );
OAI221xp5_ASAP7_75t_L g697 ( .A1(n_51), .A2(n_211), .B1(n_324), .B2(n_476), .C(n_477), .Y(n_697) );
OAI21xp33_ASAP7_75t_SL g730 ( .A1(n_51), .A2(n_375), .B(n_731), .Y(n_730) );
INVx1_ASAP7_75t_L g936 ( .A(n_52), .Y(n_936) );
INVx1_ASAP7_75t_L g242 ( .A(n_53), .Y(n_242) );
OAI22xp5_ASAP7_75t_L g1134 ( .A1(n_54), .A2(n_185), .B1(n_282), .B2(n_293), .Y(n_1134) );
INVx1_ASAP7_75t_L g1144 ( .A(n_54), .Y(n_1144) );
INVx2_ASAP7_75t_L g286 ( .A(n_55), .Y(n_286) );
OAI22xp5_ASAP7_75t_L g1121 ( .A1(n_56), .A2(n_162), .B1(n_527), .B2(n_528), .Y(n_1121) );
INVx1_ASAP7_75t_L g1142 ( .A(n_56), .Y(n_1142) );
INVx1_ASAP7_75t_L g1080 ( .A(n_57), .Y(n_1080) );
INVx1_ASAP7_75t_L g455 ( .A(n_58), .Y(n_455) );
AOI22xp33_ASAP7_75t_L g493 ( .A1(n_58), .A2(n_193), .B1(n_391), .B2(n_412), .Y(n_493) );
INVx1_ASAP7_75t_L g1159 ( .A(n_59), .Y(n_1159) );
CKINVDCx5p33_ASAP7_75t_R g471 ( .A(n_60), .Y(n_471) );
OAI22xp33_ASAP7_75t_L g710 ( .A1(n_61), .A2(n_66), .B1(n_527), .B2(n_528), .Y(n_710) );
INVxp67_ASAP7_75t_SL g722 ( .A(n_61), .Y(n_722) );
INVx1_ASAP7_75t_L g904 ( .A(n_62), .Y(n_904) );
INVx1_ASAP7_75t_L g903 ( .A(n_63), .Y(n_903) );
INVx1_ASAP7_75t_L g910 ( .A(n_64), .Y(n_910) );
AOI21xp33_ASAP7_75t_L g1386 ( .A1(n_65), .A2(n_458), .B(n_852), .Y(n_1386) );
INVxp67_ASAP7_75t_L g1405 ( .A(n_65), .Y(n_1405) );
INVx1_ASAP7_75t_L g728 ( .A(n_66), .Y(n_728) );
OAI211xp5_ASAP7_75t_L g931 ( .A1(n_67), .A2(n_498), .B(n_932), .C(n_935), .Y(n_931) );
INVx1_ASAP7_75t_L g974 ( .A(n_67), .Y(n_974) );
INVx1_ASAP7_75t_L g696 ( .A(n_68), .Y(n_696) );
OAI21xp33_ASAP7_75t_L g723 ( .A1(n_68), .A2(n_724), .B(n_725), .Y(n_723) );
AOI221xp5_ASAP7_75t_L g1126 ( .A1(n_69), .A2(n_182), .B1(n_532), .B2(n_1127), .C(n_1129), .Y(n_1126) );
CKINVDCx5p33_ASAP7_75t_R g771 ( .A(n_70), .Y(n_771) );
INVx1_ASAP7_75t_L g778 ( .A(n_72), .Y(n_778) );
AOI221x1_ASAP7_75t_SL g795 ( .A1(n_72), .A2(n_88), .B1(n_391), .B2(n_796), .C(n_800), .Y(n_795) );
INVx1_ASAP7_75t_L g1081 ( .A(n_73), .Y(n_1081) );
OAI221xp5_ASAP7_75t_L g465 ( .A1(n_74), .A2(n_145), .B1(n_466), .B2(n_468), .C(n_470), .Y(n_465) );
INVx1_ASAP7_75t_L g906 ( .A(n_75), .Y(n_906) );
INVx1_ASAP7_75t_L g354 ( .A(n_76), .Y(n_354) );
AOI22xp33_ASAP7_75t_L g411 ( .A1(n_76), .A2(n_199), .B1(n_391), .B2(n_412), .Y(n_411) );
XOR2x2_ASAP7_75t_L g509 ( .A(n_77), .B(n_510), .Y(n_509) );
AOI22xp5_ASAP7_75t_L g1174 ( .A1(n_78), .A2(n_112), .B1(n_1175), .B2(n_1178), .Y(n_1174) );
AOI22xp33_ASAP7_75t_L g1209 ( .A1(n_79), .A2(n_100), .B1(n_1168), .B2(n_1172), .Y(n_1209) );
INVx1_ASAP7_75t_L g1075 ( .A(n_80), .Y(n_1075) );
CKINVDCx5p33_ASAP7_75t_R g323 ( .A(n_81), .Y(n_323) );
INVx1_ASAP7_75t_L g761 ( .A(n_82), .Y(n_761) );
OAI22xp5_ASAP7_75t_L g811 ( .A1(n_82), .A2(n_189), .B1(n_502), .B2(n_504), .Y(n_811) );
INVx1_ASAP7_75t_L g1014 ( .A(n_83), .Y(n_1014) );
OAI22xp5_ASAP7_75t_L g1392 ( .A1(n_84), .A2(n_159), .B1(n_527), .B2(n_528), .Y(n_1392) );
INVxp67_ASAP7_75t_SL g1394 ( .A(n_84), .Y(n_1394) );
OAI22xp5_ASAP7_75t_L g526 ( .A1(n_85), .A2(n_113), .B1(n_527), .B2(n_528), .Y(n_526) );
OAI211xp5_ASAP7_75t_L g541 ( .A1(n_85), .A2(n_268), .B(n_542), .C(n_545), .Y(n_541) );
INVx1_ASAP7_75t_L g525 ( .A(n_87), .Y(n_525) );
INVx1_ASAP7_75t_L g790 ( .A(n_88), .Y(n_790) );
HB1xp67_ASAP7_75t_L g244 ( .A(n_89), .Y(n_244) );
AND2x2_ASAP7_75t_L g1169 ( .A(n_89), .B(n_242), .Y(n_1169) );
INVx1_ASAP7_75t_L g912 ( .A(n_90), .Y(n_912) );
INVx1_ASAP7_75t_L g536 ( .A(n_91), .Y(n_536) );
CKINVDCx5p33_ASAP7_75t_R g866 ( .A(n_92), .Y(n_866) );
OA22x2_ASAP7_75t_L g1045 ( .A1(n_93), .A2(n_1046), .B1(n_1114), .B2(n_1115), .Y(n_1045) );
INVxp67_ASAP7_75t_L g1115 ( .A(n_93), .Y(n_1115) );
AOI22xp33_ASAP7_75t_L g853 ( .A1(n_94), .A2(n_140), .B1(n_854), .B2(n_855), .Y(n_853) );
AOI22xp5_ASAP7_75t_L g885 ( .A1(n_94), .A2(n_95), .B1(n_886), .B2(n_888), .Y(n_885) );
INVx1_ASAP7_75t_L g868 ( .A(n_95), .Y(n_868) );
AND2x2_ASAP7_75t_L g1170 ( .A(n_97), .B(n_1171), .Y(n_1170) );
INVx1_ASAP7_75t_L g1177 ( .A(n_97), .Y(n_1177) );
INVx1_ASAP7_75t_L g434 ( .A(n_98), .Y(n_434) );
AOI22xp5_ASAP7_75t_L g824 ( .A1(n_99), .A2(n_825), .B1(n_826), .B2(n_894), .Y(n_824) );
INVx1_ASAP7_75t_L g894 ( .A(n_99), .Y(n_894) );
AOI22xp5_ASAP7_75t_L g1187 ( .A1(n_99), .A2(n_148), .B1(n_1175), .B2(n_1178), .Y(n_1187) );
CKINVDCx5p33_ASAP7_75t_R g1020 ( .A(n_101), .Y(n_1020) );
INVx1_ASAP7_75t_L g535 ( .A(n_102), .Y(n_535) );
INVx1_ASAP7_75t_L g782 ( .A(n_103), .Y(n_782) );
AOI22xp33_ASAP7_75t_L g1009 ( .A1(n_104), .A2(n_227), .B1(n_810), .B2(n_1010), .Y(n_1009) );
AOI22xp33_ASAP7_75t_L g1034 ( .A1(n_104), .A2(n_135), .B1(n_1035), .B2(n_1037), .Y(n_1034) );
INVx1_ASAP7_75t_L g1070 ( .A(n_105), .Y(n_1070) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_106), .B(n_286), .Y(n_285) );
INVx2_ASAP7_75t_L g315 ( .A(n_106), .Y(n_315) );
INVx1_ASAP7_75t_L g357 ( .A(n_106), .Y(n_357) );
CKINVDCx5p33_ASAP7_75t_R g448 ( .A(n_107), .Y(n_448) );
OAI22xp33_ASAP7_75t_L g1050 ( .A1(n_108), .A2(n_233), .B1(n_1051), .B2(n_1053), .Y(n_1050) );
OAI22xp33_ASAP7_75t_L g1112 ( .A1(n_108), .A2(n_233), .B1(n_251), .B2(n_1113), .Y(n_1112) );
INVxp67_ASAP7_75t_SL g719 ( .A(n_109), .Y(n_719) );
INVx1_ASAP7_75t_L g1384 ( .A(n_110), .Y(n_1384) );
XOR2xp5_ASAP7_75t_L g752 ( .A(n_111), .B(n_753), .Y(n_752) );
AOI22xp33_ASAP7_75t_L g1210 ( .A1(n_114), .A2(n_206), .B1(n_1175), .B2(n_1178), .Y(n_1210) );
AOI22xp5_ASAP7_75t_L g1167 ( .A1(n_116), .A2(n_119), .B1(n_1168), .B2(n_1172), .Y(n_1167) );
INVx1_ASAP7_75t_L g360 ( .A(n_117), .Y(n_360) );
AOI22xp33_ASAP7_75t_L g425 ( .A1(n_117), .A2(n_161), .B1(n_426), .B2(n_428), .Y(n_425) );
CKINVDCx5p33_ASAP7_75t_R g780 ( .A(n_118), .Y(n_780) );
OAI22xp33_ASAP7_75t_L g950 ( .A1(n_120), .A2(n_157), .B1(n_951), .B2(n_952), .Y(n_950) );
OAI22xp5_ASAP7_75t_L g958 ( .A1(n_120), .A2(n_157), .B1(n_959), .B2(n_960), .Y(n_958) );
OAI22xp33_ASAP7_75t_L g762 ( .A1(n_121), .A2(n_129), .B1(n_353), .B2(n_763), .Y(n_762) );
INVx1_ASAP7_75t_L g817 ( .A(n_121), .Y(n_817) );
INVx1_ASAP7_75t_L g1133 ( .A(n_122), .Y(n_1133) );
INVx1_ASAP7_75t_L g907 ( .A(n_123), .Y(n_907) );
AOI22xp33_ASAP7_75t_L g1191 ( .A1(n_124), .A2(n_126), .B1(n_1175), .B2(n_1178), .Y(n_1191) );
INVx1_ASAP7_75t_L g1078 ( .A(n_125), .Y(n_1078) );
XOR2x2_ASAP7_75t_L g1369 ( .A(n_126), .B(n_1370), .Y(n_1369) );
AOI22xp5_ASAP7_75t_L g1419 ( .A1(n_126), .A2(n_1420), .B1(n_1425), .B2(n_1428), .Y(n_1419) );
OAI22xp5_ASAP7_75t_L g451 ( .A1(n_127), .A2(n_293), .B1(n_452), .B2(n_456), .Y(n_451) );
INVx1_ASAP7_75t_L g484 ( .A(n_127), .Y(n_484) );
OAI22xp5_ASAP7_75t_L g515 ( .A1(n_128), .A2(n_130), .B1(n_282), .B2(n_293), .Y(n_515) );
INVxp67_ASAP7_75t_SL g546 ( .A(n_128), .Y(n_546) );
INVx1_ASAP7_75t_L g816 ( .A(n_129), .Y(n_816) );
INVxp67_ASAP7_75t_SL g543 ( .A(n_130), .Y(n_543) );
INVx1_ASAP7_75t_L g1130 ( .A(n_131), .Y(n_1130) );
INVx1_ASAP7_75t_L g995 ( .A(n_132), .Y(n_995) );
AOI22xp33_ASAP7_75t_SL g1038 ( .A1(n_132), .A2(n_227), .B1(n_1037), .B2(n_1039), .Y(n_1038) );
BUFx3_ASAP7_75t_L g292 ( .A(n_133), .Y(n_292) );
INVx1_ASAP7_75t_L g614 ( .A(n_134), .Y(n_614) );
INVx1_ASAP7_75t_L g996 ( .A(n_135), .Y(n_996) );
AOI22xp5_ASAP7_75t_L g1199 ( .A1(n_136), .A2(n_139), .B1(n_1175), .B2(n_1178), .Y(n_1199) );
INVx1_ASAP7_75t_L g1373 ( .A(n_137), .Y(n_1373) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_138), .B(n_734), .Y(n_733) );
AOI22xp33_ASAP7_75t_SL g878 ( .A1(n_140), .A2(n_202), .B1(n_879), .B2(n_880), .Y(n_878) );
INVx1_ASAP7_75t_L g520 ( .A(n_141), .Y(n_520) );
INVx1_ASAP7_75t_L g707 ( .A(n_142), .Y(n_707) );
AOI22xp5_ASAP7_75t_L g1202 ( .A1(n_143), .A2(n_198), .B1(n_1168), .B2(n_1172), .Y(n_1202) );
BUFx6f_ASAP7_75t_L g256 ( .A(n_144), .Y(n_256) );
OAI211xp5_ASAP7_75t_L g481 ( .A1(n_145), .A2(n_482), .B(n_483), .C(n_486), .Y(n_481) );
INVx1_ASAP7_75t_L g485 ( .A(n_146), .Y(n_485) );
OAI21xp5_ASAP7_75t_SL g1015 ( .A1(n_147), .A2(n_642), .B(n_1016), .Y(n_1015) );
CKINVDCx5p33_ASAP7_75t_R g447 ( .A(n_149), .Y(n_447) );
OAI221xp5_ASAP7_75t_SL g664 ( .A1(n_150), .A2(n_173), .B1(n_665), .B2(n_668), .C(n_672), .Y(n_664) );
AOI21xp5_ASAP7_75t_L g1378 ( .A1(n_152), .A2(n_840), .B(n_1379), .Y(n_1378) );
INVxp67_ASAP7_75t_SL g1402 ( .A(n_152), .Y(n_1402) );
INVx1_ASAP7_75t_L g333 ( .A(n_153), .Y(n_333) );
AOI22xp33_ASAP7_75t_L g622 ( .A1(n_154), .A2(n_216), .B1(n_623), .B2(n_625), .Y(n_622) );
INVxp67_ASAP7_75t_SL g676 ( .A(n_154), .Y(n_676) );
INVx1_ASAP7_75t_L g738 ( .A(n_155), .Y(n_738) );
INVx1_ASAP7_75t_L g845 ( .A(n_156), .Y(n_845) );
OAI221xp5_ASAP7_75t_L g881 ( .A1(n_156), .A2(n_731), .B1(n_804), .B2(n_882), .C(n_889), .Y(n_881) );
INVx1_ASAP7_75t_L g461 ( .A(n_158), .Y(n_461) );
AOI22xp33_ASAP7_75t_L g499 ( .A1(n_158), .A2(n_165), .B1(n_412), .B2(n_500), .Y(n_499) );
OAI221xp5_ASAP7_75t_L g1411 ( .A1(n_159), .A2(n_183), .B1(n_375), .B2(n_502), .C(n_504), .Y(n_1411) );
OAI211xp5_ASAP7_75t_SL g1054 ( .A1(n_160), .A2(n_964), .B(n_1055), .C(n_1057), .Y(n_1054) );
INVx1_ASAP7_75t_L g1104 ( .A(n_160), .Y(n_1104) );
INVx1_ASAP7_75t_L g344 ( .A(n_161), .Y(n_344) );
INVxp67_ASAP7_75t_SL g1157 ( .A(n_162), .Y(n_1157) );
INVx1_ASAP7_75t_L g1059 ( .A(n_163), .Y(n_1059) );
INVx1_ASAP7_75t_L g1390 ( .A(n_164), .Y(n_1390) );
AOI221xp5_ASAP7_75t_L g443 ( .A1(n_165), .A2(n_193), .B1(n_444), .B2(n_445), .C(n_446), .Y(n_443) );
INVxp67_ASAP7_75t_SL g601 ( .A(n_166), .Y(n_601) );
AOI221xp5_ASAP7_75t_L g677 ( .A1(n_166), .A2(n_204), .B1(n_659), .B2(n_678), .C(n_679), .Y(n_677) );
INVx1_ASAP7_75t_L g556 ( .A(n_167), .Y(n_556) );
BUFx6f_ASAP7_75t_L g255 ( .A(n_168), .Y(n_255) );
CKINVDCx5p33_ASAP7_75t_R g832 ( .A(n_169), .Y(n_832) );
OAI222xp33_ASAP7_75t_L g990 ( .A1(n_170), .A2(n_225), .B1(n_668), .B2(n_991), .C1(n_992), .C2(n_999), .Y(n_990) );
INVx1_ASAP7_75t_L g1023 ( .A(n_170), .Y(n_1023) );
INVx1_ASAP7_75t_L g1381 ( .A(n_171), .Y(n_1381) );
INVx1_ASAP7_75t_L g307 ( .A(n_172), .Y(n_307) );
OAI22xp5_ASAP7_75t_L g396 ( .A1(n_172), .A2(n_174), .B1(n_397), .B2(n_401), .Y(n_396) );
INVxp67_ASAP7_75t_SL g582 ( .A(n_173), .Y(n_582) );
INVx1_ASAP7_75t_L g320 ( .A(n_174), .Y(n_320) );
CKINVDCx5p33_ASAP7_75t_R g774 ( .A(n_175), .Y(n_774) );
INVx1_ASAP7_75t_L g523 ( .A(n_176), .Y(n_523) );
CKINVDCx5p33_ASAP7_75t_R g453 ( .A(n_177), .Y(n_453) );
INVx1_ASAP7_75t_L g1060 ( .A(n_179), .Y(n_1060) );
OAI211xp5_ASAP7_75t_SL g1100 ( .A1(n_179), .A2(n_932), .B(n_1101), .C(n_1102), .Y(n_1100) );
AOI22xp5_ASAP7_75t_L g1421 ( .A1(n_180), .A2(n_1422), .B1(n_1423), .B2(n_1424), .Y(n_1421) );
CKINVDCx5p33_ASAP7_75t_R g1422 ( .A(n_180), .Y(n_1422) );
INVx1_ASAP7_75t_L g1154 ( .A(n_181), .Y(n_1154) );
INVx1_ASAP7_75t_L g1155 ( .A(n_182), .Y(n_1155) );
OAI221xp5_ASAP7_75t_L g1374 ( .A1(n_183), .A2(n_201), .B1(n_324), .B2(n_476), .C(n_477), .Y(n_1374) );
INVx1_ASAP7_75t_L g1012 ( .A(n_184), .Y(n_1012) );
INVxp67_ASAP7_75t_SL g1137 ( .A(n_185), .Y(n_1137) );
AOI21xp33_ASAP7_75t_L g741 ( .A1(n_186), .A2(n_550), .B(n_742), .Y(n_741) );
OAI211xp5_ASAP7_75t_L g310 ( .A1(n_187), .A2(n_311), .B(n_316), .C(n_324), .Y(n_310) );
INVxp33_ASAP7_75t_SL g395 ( .A(n_187), .Y(n_395) );
INVx1_ASAP7_75t_L g513 ( .A(n_188), .Y(n_513) );
INVx1_ASAP7_75t_L g616 ( .A(n_190), .Y(n_616) );
AOI221xp5_ASAP7_75t_L g658 ( .A1(n_190), .A2(n_216), .B1(n_407), .B2(n_659), .C(n_661), .Y(n_658) );
AOI21xp33_ASAP7_75t_L g711 ( .A1(n_191), .A2(n_712), .B(n_715), .Y(n_711) );
INVx1_ASAP7_75t_L g758 ( .A(n_192), .Y(n_758) );
INVx1_ASAP7_75t_L g828 ( .A(n_194), .Y(n_828) );
INVxp67_ASAP7_75t_SL g833 ( .A(n_195), .Y(n_833) );
OAI221xp5_ASAP7_75t_L g856 ( .A1(n_195), .A2(n_282), .B1(n_324), .B2(n_857), .C(n_864), .Y(n_856) );
BUFx3_ASAP7_75t_L g259 ( .A(n_197), .Y(n_259) );
INVx1_ASAP7_75t_L g276 ( .A(n_197), .Y(n_276) );
INVx1_ASAP7_75t_L g340 ( .A(n_199), .Y(n_340) );
AOI21xp5_ASAP7_75t_L g849 ( .A1(n_200), .A2(n_850), .B(n_852), .Y(n_849) );
INVx1_ASAP7_75t_L g877 ( .A(n_200), .Y(n_877) );
INVxp67_ASAP7_75t_SL g1413 ( .A(n_201), .Y(n_1413) );
INVx1_ASAP7_75t_L g863 ( .A(n_202), .Y(n_863) );
CKINVDCx5p33_ASAP7_75t_R g841 ( .A(n_203), .Y(n_841) );
INVx1_ASAP7_75t_L g618 ( .A(n_204), .Y(n_618) );
OAI211xp5_ASAP7_75t_L g1005 ( .A1(n_205), .A2(n_684), .B(n_1006), .C(n_1011), .Y(n_1005) );
INVx1_ASAP7_75t_L g1027 ( .A(n_205), .Y(n_1027) );
INVx1_ASAP7_75t_L g273 ( .A(n_207), .Y(n_273) );
INVx2_ASAP7_75t_L g365 ( .A(n_207), .Y(n_365) );
INVx1_ASAP7_75t_L g373 ( .A(n_207), .Y(n_373) );
XOR2x2_ASAP7_75t_L g897 ( .A(n_208), .B(n_898), .Y(n_897) );
INVx1_ASAP7_75t_L g1131 ( .A(n_209), .Y(n_1131) );
AOI22xp33_ASAP7_75t_L g1387 ( .A1(n_210), .A2(n_220), .B1(n_295), .B2(n_445), .Y(n_1387) );
INVxp67_ASAP7_75t_SL g1409 ( .A(n_210), .Y(n_1409) );
INVx1_ASAP7_75t_L g726 ( .A(n_211), .Y(n_726) );
INVxp67_ASAP7_75t_SL g544 ( .A(n_212), .Y(n_544) );
INVx1_ASAP7_75t_L g438 ( .A(n_213), .Y(n_438) );
XOR2x2_ASAP7_75t_L g692 ( .A(n_214), .B(n_693), .Y(n_692) );
INVx1_ASAP7_75t_L g464 ( .A(n_215), .Y(n_464) );
INVx1_ASAP7_75t_L g640 ( .A(n_217), .Y(n_640) );
CKINVDCx5p33_ASAP7_75t_R g847 ( .A(n_218), .Y(n_847) );
INVx1_ASAP7_75t_L g1377 ( .A(n_219), .Y(n_1377) );
INVxp67_ASAP7_75t_SL g1400 ( .A(n_220), .Y(n_1400) );
NOR2xp33_ASAP7_75t_L g890 ( .A(n_221), .B(n_891), .Y(n_890) );
CKINVDCx5p33_ASAP7_75t_R g787 ( .A(n_222), .Y(n_787) );
OAI21xp33_ASAP7_75t_SL g267 ( .A1(n_223), .A2(n_268), .B(n_280), .Y(n_267) );
INVx1_ASAP7_75t_L g301 ( .A(n_223), .Y(n_301) );
INVx1_ASAP7_75t_L g915 ( .A(n_224), .Y(n_915) );
INVx1_ASAP7_75t_L g1025 ( .A(n_225), .Y(n_1025) );
INVx1_ASAP7_75t_L g604 ( .A(n_228), .Y(n_604) );
OAI322xp33_ASAP7_75t_SL g599 ( .A1(n_229), .A2(n_600), .A3(n_607), .B1(n_611), .B2(n_617), .C1(n_626), .C2(n_631), .Y(n_599) );
INVx1_ASAP7_75t_L g939 ( .A(n_230), .Y(n_939) );
OAI211xp5_ASAP7_75t_L g963 ( .A1(n_230), .A2(n_615), .B(n_964), .C(n_966), .Y(n_963) );
INVx1_ASAP7_75t_L g1077 ( .A(n_231), .Y(n_1077) );
INVx1_ASAP7_75t_L g844 ( .A(n_232), .Y(n_844) );
AOI21xp5_ASAP7_75t_L g234 ( .A1(n_235), .A2(n_260), .B(n_1161), .Y(n_234) );
INVx2_ASAP7_75t_SL g235 ( .A(n_236), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
INVx3_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
OR2x2_ASAP7_75t_L g238 ( .A(n_239), .B(n_245), .Y(n_238) );
NOR2xp33_ASAP7_75t_L g1418 ( .A(n_239), .B(n_248), .Y(n_1418) );
INVx1_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
NOR2xp33_ASAP7_75t_L g240 ( .A(n_241), .B(n_243), .Y(n_240) );
NOR2xp33_ASAP7_75t_L g1427 ( .A(n_241), .B(n_244), .Y(n_1427) );
INVx1_ASAP7_75t_L g1431 ( .A(n_241), .Y(n_1431) );
HB1xp67_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
INVx1_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
NOR2xp33_ASAP7_75t_L g1433 ( .A(n_244), .B(n_1431), .Y(n_1433) );
INVx1_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_247), .B(n_250), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
AND2x4_ASAP7_75t_L g955 ( .A(n_248), .B(n_956), .Y(n_955) );
INVx1_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
AND2x4_ASAP7_75t_L g421 ( .A(n_249), .B(n_259), .Y(n_421) );
AND2x4_ASAP7_75t_L g680 ( .A(n_249), .B(n_258), .Y(n_680) );
INVx1_ASAP7_75t_L g951 ( .A(n_250), .Y(n_951) );
AND2x4_ASAP7_75t_SL g1417 ( .A(n_250), .B(n_1418), .Y(n_1417) );
INVx3_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
OR2x6_ASAP7_75t_L g251 ( .A(n_252), .B(n_257), .Y(n_251) );
BUFx4f_ASAP7_75t_L g737 ( .A(n_252), .Y(n_737) );
OR2x6_ASAP7_75t_L g945 ( .A(n_252), .B(n_946), .Y(n_945) );
INVx1_ASAP7_75t_L g1074 ( .A(n_252), .Y(n_1074) );
INVx2_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
BUFx4f_ASAP7_75t_L g560 ( .A(n_253), .Y(n_560) );
INVx3_ASAP7_75t_L g575 ( .A(n_253), .Y(n_575) );
INVx3_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
OR2x2_ASAP7_75t_L g254 ( .A(n_255), .B(n_256), .Y(n_254) );
INVx2_ASAP7_75t_L g278 ( .A(n_255), .Y(n_278) );
NAND2x1_ASAP7_75t_L g371 ( .A(n_255), .B(n_256), .Y(n_371) );
AND2x2_ASAP7_75t_L g386 ( .A(n_255), .B(n_387), .Y(n_386) );
INVx2_ASAP7_75t_L g394 ( .A(n_255), .Y(n_394) );
INVx1_ASAP7_75t_L g404 ( .A(n_255), .Y(n_404) );
AND2x2_ASAP7_75t_L g410 ( .A(n_255), .B(n_256), .Y(n_410) );
INVx1_ASAP7_75t_L g279 ( .A(n_256), .Y(n_279) );
INVx2_ASAP7_75t_L g387 ( .A(n_256), .Y(n_387) );
AND2x2_ASAP7_75t_L g393 ( .A(n_256), .B(n_394), .Y(n_393) );
BUFx2_ASAP7_75t_L g400 ( .A(n_256), .Y(n_400) );
OR2x2_ASAP7_75t_L g491 ( .A(n_256), .B(n_278), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_256), .B(n_394), .Y(n_564) );
INVxp67_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
INVx1_ASAP7_75t_L g934 ( .A(n_258), .Y(n_934) );
INVx2_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
BUFx2_ASAP7_75t_L g938 ( .A(n_259), .Y(n_938) );
AND2x4_ASAP7_75t_L g942 ( .A(n_259), .B(n_403), .Y(n_942) );
OAI22xp33_ASAP7_75t_L g260 ( .A1(n_261), .A2(n_262), .B1(n_821), .B2(n_822), .Y(n_260) );
INVxp67_ASAP7_75t_SL g261 ( .A(n_262), .Y(n_261) );
AOI22xp33_ASAP7_75t_L g262 ( .A1(n_263), .A2(n_506), .B1(n_507), .B2(n_820), .Y(n_262) );
INVx1_ASAP7_75t_L g820 ( .A(n_263), .Y(n_820) );
OAI22xp5_ASAP7_75t_L g263 ( .A1(n_264), .A2(n_265), .B1(n_436), .B2(n_505), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
XOR2x2_ASAP7_75t_L g265 ( .A(n_266), .B(n_435), .Y(n_265) );
NOR2xp33_ASAP7_75t_L g266 ( .A(n_267), .B(n_366), .Y(n_266) );
INVx1_ASAP7_75t_L g1395 ( .A(n_268), .Y(n_1395) );
INVx3_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_269), .B(n_471), .Y(n_480) );
AOI211xp5_ASAP7_75t_L g721 ( .A1(n_269), .A2(n_722), .B(n_723), .C(n_730), .Y(n_721) );
AOI22xp33_ASAP7_75t_SL g815 ( .A1(n_269), .A2(n_383), .B1(n_816), .B2(n_817), .Y(n_815) );
AOI222xp33_ASAP7_75t_L g827 ( .A1(n_269), .A2(n_383), .B1(n_828), .B2(n_829), .C1(n_832), .C2(n_833), .Y(n_827) );
NAND2xp5_ASAP7_75t_L g1156 ( .A(n_269), .B(n_1157), .Y(n_1156) );
AND2x4_ASAP7_75t_L g269 ( .A(n_270), .B(n_274), .Y(n_269) );
AND2x4_ASAP7_75t_L g383 ( .A(n_270), .B(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
OR2x2_ASAP7_75t_L g401 ( .A(n_271), .B(n_402), .Y(n_401) );
OR2x2_ASAP7_75t_L g504 ( .A(n_271), .B(n_402), .Y(n_504) );
INVxp67_ASAP7_75t_L g645 ( .A(n_271), .Y(n_645) );
INVx1_ASAP7_75t_L g956 ( .A(n_271), .Y(n_956) );
BUFx2_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
INVx2_ASAP7_75t_L g424 ( .A(n_272), .Y(n_424) );
INVx1_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
BUFx6f_ASAP7_75t_L g683 ( .A(n_274), .Y(n_683) );
AND2x2_ASAP7_75t_L g274 ( .A(n_275), .B(n_277), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_275), .B(n_373), .Y(n_372) );
AND2x2_ASAP7_75t_L g384 ( .A(n_275), .B(n_385), .Y(n_384) );
AND2x4_ASAP7_75t_SL g651 ( .A(n_275), .B(n_409), .Y(n_651) );
AND2x4_ASAP7_75t_L g667 ( .A(n_275), .B(n_385), .Y(n_667) );
AND2x4_ASAP7_75t_L g685 ( .A(n_275), .B(n_500), .Y(n_685) );
HB1xp67_ASAP7_75t_L g946 ( .A(n_276), .Y(n_946) );
BUFx6f_ASAP7_75t_L g412 ( .A(n_277), .Y(n_412) );
INVx3_ASAP7_75t_L g427 ( .A(n_277), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_277), .B(n_380), .Y(n_433) );
AND2x2_ASAP7_75t_L g277 ( .A(n_278), .B(n_279), .Y(n_277) );
OAI31xp33_ASAP7_75t_SL g280 ( .A1(n_281), .A2(n_310), .A3(n_329), .B(n_364), .Y(n_280) );
CKINVDCx5p33_ASAP7_75t_R g1389 ( .A(n_282), .Y(n_1389) );
OR2x6_ASAP7_75t_SL g282 ( .A(n_283), .B(n_287), .Y(n_282) );
INVx2_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
AND2x4_ASAP7_75t_L g294 ( .A(n_284), .B(n_295), .Y(n_294) );
HB1xp67_ASAP7_75t_L g474 ( .A(n_284), .Y(n_474) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
INVx1_ASAP7_75t_L g306 ( .A(n_285), .Y(n_306) );
OR2x2_ASAP7_75t_L g587 ( .A(n_285), .B(n_424), .Y(n_587) );
INVx3_ASAP7_75t_L g313 ( .A(n_286), .Y(n_313) );
BUFx3_ASAP7_75t_L g338 ( .A(n_286), .Y(n_338) );
NAND2xp33_ASAP7_75t_SL g610 ( .A(n_286), .B(n_315), .Y(n_610) );
INVx3_ASAP7_75t_L g467 ( .A(n_287), .Y(n_467) );
INVx1_ASAP7_75t_L g603 ( .A(n_287), .Y(n_603) );
BUFx2_ASAP7_75t_L g909 ( .A(n_287), .Y(n_909) );
INVx2_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
BUFx8_ASAP7_75t_L g335 ( .A(n_288), .Y(n_335) );
BUFx6f_ASAP7_75t_L g450 ( .A(n_288), .Y(n_450) );
BUFx6f_ASAP7_75t_L g458 ( .A(n_288), .Y(n_458) );
AND2x4_ASAP7_75t_L g288 ( .A(n_289), .B(n_291), .Y(n_288) );
INVxp67_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
INVx1_ASAP7_75t_L g305 ( .A(n_290), .Y(n_305) );
AND2x4_ASAP7_75t_L g303 ( .A(n_291), .B(n_304), .Y(n_303) );
INVx2_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
BUFx6f_ASAP7_75t_L g296 ( .A(n_292), .Y(n_296) );
AND2x4_ASAP7_75t_L g309 ( .A(n_292), .B(n_298), .Y(n_309) );
OR2x2_ASAP7_75t_L g343 ( .A(n_292), .B(n_305), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_292), .B(n_299), .Y(n_348) );
INVx3_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g893 ( .A(n_294), .B(n_540), .Y(n_893) );
AOI221xp5_ASAP7_75t_L g1388 ( .A1(n_294), .A2(n_1389), .B1(n_1390), .B2(n_1391), .C(n_1392), .Y(n_1388) );
BUFx12f_ASAP7_75t_L g444 ( .A(n_295), .Y(n_444) );
BUFx3_ASAP7_75t_L g532 ( .A(n_295), .Y(n_532) );
INVx5_ASAP7_75t_L g706 ( .A(n_295), .Y(n_706) );
BUFx3_ASAP7_75t_L g1037 ( .A(n_295), .Y(n_1037) );
AND2x4_ASAP7_75t_L g295 ( .A(n_296), .B(n_297), .Y(n_295) );
INVx2_ASAP7_75t_L g319 ( .A(n_296), .Y(n_319) );
NAND2x1p5_ASAP7_75t_L g326 ( .A(n_296), .B(n_327), .Y(n_326) );
BUFx2_ASAP7_75t_L g970 ( .A(n_296), .Y(n_970) );
INVx1_ASAP7_75t_L g322 ( .A(n_297), .Y(n_322) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
INVx2_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
INVx1_ASAP7_75t_L g327 ( .A(n_299), .Y(n_327) );
AOI22xp5_ASAP7_75t_L g300 ( .A1(n_301), .A2(n_302), .B1(n_307), .B2(n_308), .Y(n_300) );
INVx2_ASAP7_75t_L g527 ( .A(n_302), .Y(n_527) );
AND2x2_ASAP7_75t_L g302 ( .A(n_303), .B(n_306), .Y(n_302) );
NAND2x1p5_ASAP7_75t_L g311 ( .A(n_303), .B(n_312), .Y(n_311) );
BUFx3_ASAP7_75t_L g445 ( .A(n_303), .Y(n_445) );
BUFx3_ASAP7_75t_L g472 ( .A(n_303), .Y(n_472) );
INVx8_ASAP7_75t_L g624 ( .A(n_303), .Y(n_624) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
AND2x2_ASAP7_75t_L g308 ( .A(n_306), .B(n_309), .Y(n_308) );
INVx1_ASAP7_75t_L g528 ( .A(n_308), .Y(n_528) );
BUFx3_ASAP7_75t_L g518 ( .A(n_309), .Y(n_518) );
BUFx2_ASAP7_75t_L g598 ( .A(n_309), .Y(n_598) );
BUFx2_ASAP7_75t_L g625 ( .A(n_309), .Y(n_625) );
INVx2_ASAP7_75t_L g760 ( .A(n_309), .Y(n_760) );
BUFx2_ASAP7_75t_L g842 ( .A(n_309), .Y(n_842) );
AND2x4_ASAP7_75t_L g965 ( .A(n_309), .B(n_313), .Y(n_965) );
BUFx2_ASAP7_75t_L g1041 ( .A(n_309), .Y(n_1041) );
INVx2_ASAP7_75t_L g463 ( .A(n_311), .Y(n_463) );
OR2x6_ASAP7_75t_L g644 ( .A(n_311), .B(n_645), .Y(n_644) );
OR2x2_ASAP7_75t_L g830 ( .A(n_311), .B(n_645), .Y(n_830) );
AND2x6_ASAP7_75t_L g317 ( .A(n_312), .B(n_318), .Y(n_317) );
AND2x2_ASAP7_75t_L g321 ( .A(n_312), .B(n_322), .Y(n_321) );
INVx1_ASAP7_75t_L g328 ( .A(n_312), .Y(n_328) );
AND2x4_ASAP7_75t_L g591 ( .A(n_312), .B(n_431), .Y(n_591) );
AND2x4_ASAP7_75t_L g312 ( .A(n_313), .B(n_314), .Y(n_312) );
NAND2x1p5_ASAP7_75t_L g356 ( .A(n_313), .B(n_357), .Y(n_356) );
NAND3x1_ASAP7_75t_L g629 ( .A(n_313), .B(n_357), .C(n_630), .Y(n_629) );
OR2x4_ASAP7_75t_L g959 ( .A(n_313), .B(n_343), .Y(n_959) );
INVx1_ASAP7_75t_L g962 ( .A(n_313), .Y(n_962) );
OR2x6_ASAP7_75t_L g980 ( .A(n_313), .B(n_606), .Y(n_980) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
AND2x2_ASAP7_75t_L g337 ( .A(n_315), .B(n_338), .Y(n_337) );
HB1xp67_ASAP7_75t_L g984 ( .A(n_315), .Y(n_984) );
AND3x4_ASAP7_75t_L g1031 ( .A(n_315), .B(n_338), .C(n_364), .Y(n_1031) );
AOI22xp33_ASAP7_75t_L g316 ( .A1(n_317), .A2(n_320), .B1(n_321), .B2(n_323), .Y(n_316) );
INVx4_ASAP7_75t_L g476 ( .A(n_317), .Y(n_476) );
AOI22xp33_ASAP7_75t_L g843 ( .A1(n_317), .A2(n_321), .B1(n_844), .B2(n_845), .Y(n_843) );
AND2x2_ASAP7_75t_L g590 ( .A(n_318), .B(n_591), .Y(n_590) );
AND2x2_ASAP7_75t_L g1024 ( .A(n_318), .B(n_591), .Y(n_1024) );
INVx3_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
INVx2_ASAP7_75t_L g477 ( .A(n_321), .Y(n_477) );
INVx1_ASAP7_75t_L g595 ( .A(n_322), .Y(n_595) );
AOI21xp5_ASAP7_75t_L g367 ( .A1(n_323), .A2(n_368), .B(n_374), .Y(n_367) );
CKINVDCx5p33_ASAP7_75t_R g442 ( .A(n_324), .Y(n_442) );
OR2x6_ASAP7_75t_L g324 ( .A(n_325), .B(n_328), .Y(n_324) );
OAI221xp5_ASAP7_75t_L g452 ( .A1(n_325), .A2(n_355), .B1(n_453), .B2(n_454), .C(n_455), .Y(n_452) );
INVx1_ASAP7_75t_L g714 ( .A(n_325), .Y(n_714) );
INVx1_ASAP7_75t_L g1056 ( .A(n_325), .Y(n_1056) );
BUFx2_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
BUFx6f_ASAP7_75t_L g332 ( .A(n_326), .Y(n_332) );
BUFx3_ASAP7_75t_L g534 ( .A(n_326), .Y(n_534) );
BUFx2_ASAP7_75t_L g973 ( .A(n_327), .Y(n_973) );
INVx1_ASAP7_75t_L g768 ( .A(n_328), .Y(n_768) );
OAI22xp5_ASAP7_75t_L g329 ( .A1(n_330), .A2(n_339), .B1(n_349), .B2(n_358), .Y(n_329) );
OAI221xp5_ASAP7_75t_L g330 ( .A1(n_331), .A2(n_333), .B1(n_334), .B2(n_336), .C(n_337), .Y(n_330) );
OAI22xp33_ASAP7_75t_L g902 ( .A1(n_331), .A2(n_861), .B1(n_903), .B2(n_904), .Y(n_902) );
HB1xp67_ASAP7_75t_L g1090 ( .A(n_331), .Y(n_1090) );
BUFx6f_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
INVx4_ASAP7_75t_L g352 ( .A(n_332), .Y(n_352) );
OAI221xp5_ASAP7_75t_L g446 ( .A1(n_332), .A2(n_337), .B1(n_447), .B2(n_448), .C(n_449), .Y(n_446) );
INVx3_ASAP7_75t_L g469 ( .A(n_332), .Y(n_469) );
OR2x2_ASAP7_75t_L g643 ( .A(n_332), .B(n_587), .Y(n_643) );
OAI22xp5_ASAP7_75t_L g358 ( .A1(n_334), .A2(n_359), .B1(n_360), .B2(n_361), .Y(n_358) );
OAI21xp33_ASAP7_75t_L g519 ( .A1(n_334), .A2(n_337), .B(n_520), .Y(n_519) );
INVx3_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
AND2x4_ASAP7_75t_L g585 ( .A(n_335), .B(n_586), .Y(n_585) );
INVx3_ASAP7_75t_L g851 ( .A(n_335), .Y(n_851) );
INVx2_ASAP7_75t_SL g865 ( .A(n_335), .Y(n_865) );
HB1xp67_ASAP7_75t_L g1039 ( .A(n_335), .Y(n_1039) );
INVx2_ASAP7_75t_SL g1128 ( .A(n_335), .Y(n_1128) );
OAI221xp5_ASAP7_75t_L g705 ( .A1(n_337), .A2(n_706), .B1(n_707), .B2(n_708), .C(n_709), .Y(n_705) );
OAI221xp5_ASAP7_75t_L g786 ( .A1(n_337), .A2(n_351), .B1(n_787), .B2(n_788), .C(n_790), .Y(n_786) );
OAI221xp5_ASAP7_75t_L g1123 ( .A1(n_337), .A2(n_534), .B1(n_763), .B2(n_1124), .C(n_1125), .Y(n_1123) );
INVx3_ASAP7_75t_L g969 ( .A(n_338), .Y(n_969) );
OAI22xp5_ASAP7_75t_L g339 ( .A1(n_340), .A2(n_341), .B1(n_344), .B2(n_345), .Y(n_339) );
BUFx4f_ASAP7_75t_SL g781 ( .A(n_341), .Y(n_781) );
INVx3_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
INVx2_ASAP7_75t_SL g632 ( .A(n_342), .Y(n_632) );
INVx2_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
BUFx3_ASAP7_75t_L g353 ( .A(n_343), .Y(n_353) );
BUFx4f_ASAP7_75t_L g454 ( .A(n_343), .Y(n_454) );
BUFx3_ASAP7_75t_L g522 ( .A(n_343), .Y(n_522) );
OR2x4_ASAP7_75t_L g978 ( .A(n_343), .B(n_962), .Y(n_978) );
INVx3_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
INVx3_ASAP7_75t_L g460 ( .A(n_346), .Y(n_460) );
INVx1_ASAP7_75t_L g524 ( .A(n_346), .Y(n_524) );
CKINVDCx8_ASAP7_75t_R g867 ( .A(n_346), .Y(n_867) );
INVx3_ASAP7_75t_L g1092 ( .A(n_346), .Y(n_1092) );
BUFx6f_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
INVx1_ASAP7_75t_L g363 ( .A(n_347), .Y(n_363) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
BUFx2_ASAP7_75t_L g606 ( .A(n_348), .Y(n_606) );
OAI221xp5_ASAP7_75t_L g349 ( .A1(n_350), .A2(n_351), .B1(n_353), .B2(n_354), .C(n_355), .Y(n_349) );
OAI21xp33_ASAP7_75t_L g1376 ( .A1(n_351), .A2(n_1377), .B(n_1378), .Y(n_1376) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx2_ASAP7_75t_L g704 ( .A(n_352), .Y(n_704) );
INVx1_ASAP7_75t_L g777 ( .A(n_352), .Y(n_777) );
OAI221xp5_ASAP7_75t_L g533 ( .A1(n_353), .A2(n_355), .B1(n_534), .B2(n_535), .C(n_536), .Y(n_533) );
INVx1_ASAP7_75t_L g613 ( .A(n_353), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_355), .B(n_716), .Y(n_715) );
OAI221xp5_ASAP7_75t_L g775 ( .A1(n_355), .A2(n_522), .B1(n_776), .B2(n_777), .C(n_778), .Y(n_775) );
OAI221xp5_ASAP7_75t_L g857 ( .A1(n_355), .A2(n_858), .B1(n_860), .B2(n_861), .C(n_863), .Y(n_857) );
OAI221xp5_ASAP7_75t_L g1129 ( .A1(n_355), .A2(n_454), .B1(n_534), .B2(n_1130), .C(n_1131), .Y(n_1129) );
INVx3_ASAP7_75t_L g1379 ( .A(n_355), .Y(n_1379) );
INVx3_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
OAI22xp5_ASAP7_75t_L g1380 ( .A1(n_361), .A2(n_1128), .B1(n_1381), .B2(n_1382), .Y(n_1380) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
OR2x2_ASAP7_75t_L g638 ( .A(n_363), .B(n_587), .Y(n_638) );
BUFx3_ASAP7_75t_L g911 ( .A(n_363), .Y(n_911) );
INVx1_ASAP7_75t_L g479 ( .A(n_364), .Y(n_479) );
INVx2_ASAP7_75t_SL g717 ( .A(n_364), .Y(n_717) );
INVx2_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_365), .B(n_380), .Y(n_379) );
BUFx2_ASAP7_75t_L g416 ( .A(n_365), .Y(n_416) );
NAND4xp25_ASAP7_75t_SL g366 ( .A(n_367), .B(n_381), .C(n_388), .D(n_405), .Y(n_366) );
AOI332xp33_ASAP7_75t_L g483 ( .A1(n_368), .A2(n_390), .A3(n_391), .B1(n_430), .B2(n_432), .B3(n_464), .C1(n_484), .C2(n_485), .Y(n_483) );
AOI222xp33_ASAP7_75t_L g542 ( .A1(n_368), .A2(n_389), .B1(n_429), .B2(n_513), .C1(n_543), .C2(n_544), .Y(n_542) );
AOI21xp5_ASAP7_75t_L g1158 ( .A1(n_368), .A2(n_374), .B(n_1159), .Y(n_1158) );
AOI222xp33_ASAP7_75t_L g1412 ( .A1(n_368), .A2(n_389), .B1(n_429), .B2(n_1373), .C1(n_1391), .C2(n_1413), .Y(n_1412) );
INVx2_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
OR2x2_ASAP7_75t_L g369 ( .A(n_370), .B(n_372), .Y(n_369) );
OR2x2_ASAP7_75t_L g731 ( .A(n_370), .B(n_372), .Y(n_731) );
BUFx3_ASAP7_75t_L g802 ( .A(n_370), .Y(n_802) );
INVx2_ASAP7_75t_SL g994 ( .A(n_370), .Y(n_994) );
BUFx3_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
BUFx6f_ASAP7_75t_L g376 ( .A(n_371), .Y(n_376) );
INVx1_ASAP7_75t_L g390 ( .A(n_372), .Y(n_390) );
INVx1_ASAP7_75t_L g431 ( .A(n_373), .Y(n_431) );
INVx1_ASAP7_75t_L g630 ( .A(n_373), .Y(n_630) );
NOR3xp33_ASAP7_75t_L g486 ( .A(n_374), .B(n_487), .C(n_501), .Y(n_486) );
OR3x1_ASAP7_75t_L g547 ( .A(n_374), .B(n_548), .C(n_549), .Y(n_547) );
CKINVDCx5p33_ASAP7_75t_R g374 ( .A(n_375), .Y(n_374) );
OAI21xp5_ASAP7_75t_L g803 ( .A1(n_375), .A2(n_804), .B(n_805), .Y(n_803) );
OAI21xp5_ASAP7_75t_SL g872 ( .A1(n_375), .A2(n_873), .B(n_875), .Y(n_872) );
OR2x6_ASAP7_75t_L g375 ( .A(n_376), .B(n_377), .Y(n_375) );
BUFx4f_ASAP7_75t_L g492 ( .A(n_376), .Y(n_492) );
BUFx6f_ASAP7_75t_L g498 ( .A(n_376), .Y(n_498) );
BUFx4f_ASAP7_75t_L g555 ( .A(n_376), .Y(n_555) );
INVx4_ASAP7_75t_L g570 ( .A(n_376), .Y(n_570) );
BUFx4f_ASAP7_75t_L g884 ( .A(n_376), .Y(n_884) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
NAND2x2_ASAP7_75t_L g397 ( .A(n_378), .B(n_398), .Y(n_397) );
INVx2_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_380), .B(n_403), .Y(n_402) );
AND2x6_ASAP7_75t_L g663 ( .A(n_380), .B(n_409), .Y(n_663) );
INVx1_ASAP7_75t_L g671 ( .A(n_380), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_382), .B(n_383), .Y(n_381) );
INVx1_ASAP7_75t_L g482 ( .A(n_383), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_383), .B(n_546), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_383), .B(n_719), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g1414 ( .A(n_383), .B(n_1390), .Y(n_1414) );
BUFx6f_ASAP7_75t_L g407 ( .A(n_385), .Y(n_407) );
BUFx6f_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
BUFx3_ASAP7_75t_L g678 ( .A(n_386), .Y(n_678) );
INVx2_ASAP7_75t_L g799 ( .A(n_386), .Y(n_799) );
AND2x4_ASAP7_75t_L g953 ( .A(n_386), .B(n_946), .Y(n_953) );
AOI21xp33_ASAP7_75t_L g388 ( .A1(n_389), .A2(n_395), .B(n_396), .Y(n_388) );
INVx1_ASAP7_75t_L g724 ( .A(n_389), .Y(n_724) );
INVx1_ASAP7_75t_L g831 ( .A(n_389), .Y(n_831) );
AOI222xp33_ASAP7_75t_L g1140 ( .A1(n_389), .A2(n_727), .B1(n_729), .B2(n_1133), .C1(n_1141), .C2(n_1142), .Y(n_1140) );
AND2x4_ASAP7_75t_L g389 ( .A(n_390), .B(n_391), .Y(n_389) );
INVx3_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
INVx2_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
BUFx3_ASAP7_75t_L g428 ( .A(n_393), .Y(n_428) );
BUFx6f_ASAP7_75t_L g500 ( .A(n_393), .Y(n_500) );
BUFx3_ASAP7_75t_L g888 ( .A(n_393), .Y(n_888) );
INVx2_ASAP7_75t_SL g503 ( .A(n_397), .Y(n_503) );
INVx1_ASAP7_75t_L g727 ( .A(n_397), .Y(n_727) );
INVx2_ASAP7_75t_SL g398 ( .A(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g670 ( .A(n_400), .Y(n_670) );
AND2x4_ASAP7_75t_L g937 ( .A(n_400), .B(n_938), .Y(n_937) );
AND2x4_ASAP7_75t_L g642 ( .A(n_401), .B(n_643), .Y(n_642) );
INVx2_ASAP7_75t_SL g729 ( .A(n_401), .Y(n_729) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
AOI332xp33_ASAP7_75t_L g405 ( .A1(n_406), .A2(n_411), .A3(n_413), .B1(n_418), .B2(n_420), .B3(n_425), .C1(n_429), .C2(n_434), .Y(n_405) );
BUFx3_ASAP7_75t_L g734 ( .A(n_407), .Y(n_734) );
BUFx3_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
BUFx3_ASAP7_75t_L g419 ( .A(n_409), .Y(n_419) );
INVx1_ASAP7_75t_L g660 ( .A(n_409), .Y(n_660) );
BUFx3_ASAP7_75t_L g742 ( .A(n_409), .Y(n_742) );
BUFx6f_ASAP7_75t_L g746 ( .A(n_409), .Y(n_746) );
AND2x2_ASAP7_75t_L g933 ( .A(n_409), .B(n_934), .Y(n_933) );
BUFx6f_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx3_ASAP7_75t_L g887 ( .A(n_412), .Y(n_887) );
HB1xp67_ASAP7_75t_L g874 ( .A(n_413), .Y(n_874) );
INVx2_ASAP7_75t_SL g413 ( .A(n_414), .Y(n_413) );
INVx4_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx2_ASAP7_75t_L g488 ( .A(n_415), .Y(n_488) );
INVx2_ASAP7_75t_L g550 ( .A(n_415), .Y(n_550) );
HB1xp67_ASAP7_75t_L g794 ( .A(n_415), .Y(n_794) );
INVx2_ASAP7_75t_L g1068 ( .A(n_415), .Y(n_1068) );
AOI222xp33_ASAP7_75t_L g1143 ( .A1(n_415), .A2(n_420), .B1(n_429), .B2(n_1144), .C1(n_1145), .C2(n_1152), .Y(n_1143) );
AND2x4_ASAP7_75t_L g415 ( .A(n_416), .B(n_417), .Y(n_415) );
INVx1_ASAP7_75t_L g540 ( .A(n_416), .Y(n_540) );
AOI322xp5_ASAP7_75t_L g732 ( .A1(n_420), .A2(n_429), .A3(n_733), .B1(n_735), .B2(n_741), .C1(n_743), .C2(n_744), .Y(n_732) );
CKINVDCx5p33_ASAP7_75t_R g804 ( .A(n_420), .Y(n_804) );
AND2x4_ASAP7_75t_L g420 ( .A(n_421), .B(n_422), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_421), .B(n_422), .Y(n_494) );
AND2x2_ASAP7_75t_SL g572 ( .A(n_421), .B(n_424), .Y(n_572) );
INVx4_ASAP7_75t_L g661 ( .A(n_421), .Y(n_661) );
INVx4_ASAP7_75t_L g1008 ( .A(n_421), .Y(n_1008) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
OR2x2_ASAP7_75t_L g609 ( .A(n_424), .B(n_610), .Y(n_609) );
HB1xp67_ASAP7_75t_L g986 ( .A(n_424), .Y(n_986) );
INVx2_ASAP7_75t_SL g426 ( .A(n_427), .Y(n_426) );
INVx2_ASAP7_75t_L g810 ( .A(n_427), .Y(n_810) );
INVx2_ASAP7_75t_L g879 ( .A(n_427), .Y(n_879) );
HB1xp67_ASAP7_75t_L g1010 ( .A(n_428), .Y(n_1010) );
AND2x4_ASAP7_75t_L g429 ( .A(n_430), .B(n_432), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
OR2x2_ASAP7_75t_L g639 ( .A(n_431), .B(n_433), .Y(n_639) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g505 ( .A(n_436), .Y(n_505) );
HB1xp67_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
XNOR2x1_ASAP7_75t_L g437 ( .A(n_438), .B(n_439), .Y(n_437) );
OR2x2_ASAP7_75t_L g439 ( .A(n_440), .B(n_481), .Y(n_439) );
A2O1A1Ixp33_ASAP7_75t_L g440 ( .A1(n_441), .A2(n_462), .B(n_478), .C(n_480), .Y(n_440) );
NOR3xp33_ASAP7_75t_L g441 ( .A(n_442), .B(n_443), .C(n_451), .Y(n_441) );
BUFx2_ASAP7_75t_L g854 ( .A(n_445), .Y(n_854) );
OAI221xp5_ASAP7_75t_L g495 ( .A1(n_447), .A2(n_453), .B1(n_496), .B2(n_498), .C(n_499), .Y(n_495) );
OAI221xp5_ASAP7_75t_L g489 ( .A1(n_448), .A2(n_459), .B1(n_490), .B2(n_492), .C(n_493), .Y(n_489) );
INVx2_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx2_ASAP7_75t_L g531 ( .A(n_450), .Y(n_531) );
INVx1_ASAP7_75t_L g702 ( .A(n_450), .Y(n_702) );
BUFx6f_ASAP7_75t_L g789 ( .A(n_450), .Y(n_789) );
AND2x4_ASAP7_75t_L g961 ( .A(n_450), .B(n_962), .Y(n_961) );
INVx1_ASAP7_75t_L g862 ( .A(n_454), .Y(n_862) );
OAI22xp5_ASAP7_75t_L g456 ( .A1(n_457), .A2(n_459), .B1(n_460), .B2(n_461), .Y(n_456) );
INVx2_ASAP7_75t_L g620 ( .A(n_457), .Y(n_620) );
INVx3_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx2_ASAP7_75t_SL g763 ( .A(n_458), .Y(n_763) );
HB1xp67_ASAP7_75t_L g773 ( .A(n_458), .Y(n_773) );
INVx5_ASAP7_75t_L g1036 ( .A(n_458), .Y(n_1036) );
OAI22xp5_ASAP7_75t_L g905 ( .A1(n_460), .A2(n_531), .B1(n_906), .B2(n_907), .Y(n_905) );
AOI221xp5_ASAP7_75t_L g462 ( .A1(n_463), .A2(n_464), .B1(n_465), .B2(n_473), .C(n_475), .Y(n_462) );
AOI211xp5_ASAP7_75t_L g512 ( .A1(n_463), .A2(n_513), .B(n_514), .C(n_515), .Y(n_512) );
AOI211xp5_ASAP7_75t_SL g695 ( .A1(n_463), .A2(n_696), .B(n_697), .C(n_698), .Y(n_695) );
AOI211xp5_ASAP7_75t_SL g1132 ( .A1(n_463), .A2(n_1133), .B(n_1134), .C(n_1135), .Y(n_1132) );
AOI211xp5_ASAP7_75t_L g1372 ( .A1(n_463), .A2(n_1373), .B(n_1374), .C(n_1375), .Y(n_1372) );
INVx2_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVx2_ASAP7_75t_L g1094 ( .A(n_467), .Y(n_1094) );
HB1xp67_ASAP7_75t_L g848 ( .A(n_468), .Y(n_848) );
INVx2_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVx2_ASAP7_75t_L g1098 ( .A(n_469), .Y(n_1098) );
INVx3_ASAP7_75t_L g1385 ( .A(n_469), .Y(n_1385) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_471), .B(n_472), .Y(n_470) );
INVx2_ASAP7_75t_SL g708 ( .A(n_472), .Y(n_708) );
INVx1_ASAP7_75t_L g756 ( .A(n_473), .Y(n_756) );
BUFx2_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
INVx1_ASAP7_75t_L g838 ( .A(n_474), .Y(n_838) );
HB1xp67_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
BUFx2_ASAP7_75t_L g870 ( .A(n_479), .Y(n_870) );
INVx1_ASAP7_75t_L g1138 ( .A(n_482), .Y(n_1138) );
OAI22xp5_ASAP7_75t_SL g487 ( .A1(n_488), .A2(n_489), .B1(n_494), .B2(n_495), .Y(n_487) );
OAI33xp33_ASAP7_75t_L g1398 ( .A1(n_488), .A2(n_1399), .A3(n_1404), .B1(n_1406), .B2(n_1408), .B3(n_1410), .Y(n_1398) );
INVx2_ASAP7_75t_L g926 ( .A(n_490), .Y(n_926) );
BUFx3_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
INVx2_ASAP7_75t_L g497 ( .A(n_491), .Y(n_497) );
BUFx2_ASAP7_75t_L g554 ( .A(n_491), .Y(n_554) );
INVx1_ASAP7_75t_L g807 ( .A(n_491), .Y(n_807) );
BUFx2_ASAP7_75t_L g1407 ( .A(n_491), .Y(n_1407) );
OAI221xp5_ASAP7_75t_L g875 ( .A1(n_492), .A2(n_866), .B1(n_876), .B2(n_877), .C(n_878), .Y(n_875) );
INVx1_ASAP7_75t_L g928 ( .A(n_494), .Y(n_928) );
OAI221xp5_ASAP7_75t_L g992 ( .A1(n_496), .A2(n_993), .B1(n_995), .B2(n_996), .C(n_997), .Y(n_992) );
INVx2_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
BUFx2_ASAP7_75t_L g567 ( .A(n_497), .Y(n_567) );
INVx2_ASAP7_75t_L g876 ( .A(n_497), .Y(n_876) );
OAI22xp5_ASAP7_75t_L g1076 ( .A1(n_498), .A2(n_883), .B1(n_1077), .B2(n_1078), .Y(n_1076) );
OAI22xp5_ASAP7_75t_L g1406 ( .A1(n_498), .A2(n_1377), .B1(n_1384), .B2(n_1407), .Y(n_1406) );
BUFx2_ASAP7_75t_L g880 ( .A(n_500), .Y(n_880) );
INVx2_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
INVx1_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
OAI22xp33_ASAP7_75t_L g507 ( .A1(n_508), .A2(n_690), .B1(n_691), .B2(n_819), .Y(n_507) );
INVx1_ASAP7_75t_L g819 ( .A(n_508), .Y(n_819) );
OAI22xp5_ASAP7_75t_L g508 ( .A1(n_509), .A2(n_578), .B1(n_688), .B2(n_689), .Y(n_508) );
INVx2_ASAP7_75t_L g688 ( .A(n_509), .Y(n_688) );
AOI211x1_ASAP7_75t_L g510 ( .A1(n_511), .A2(n_537), .B(n_541), .C(n_547), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_512), .B(n_516), .Y(n_511) );
NOR3xp33_ASAP7_75t_L g516 ( .A(n_517), .B(n_526), .C(n_529), .Y(n_516) );
OAI22xp5_ASAP7_75t_L g551 ( .A1(n_520), .A2(n_552), .B1(n_555), .B2(n_556), .Y(n_551) );
OAI22xp5_ASAP7_75t_L g521 ( .A1(n_522), .A2(n_523), .B1(n_524), .B2(n_525), .Y(n_521) );
OAI22xp5_ASAP7_75t_L g557 ( .A1(n_523), .A2(n_536), .B1(n_558), .B2(n_561), .Y(n_557) );
OAI22xp5_ASAP7_75t_L g573 ( .A1(n_525), .A2(n_574), .B1(n_576), .B2(n_577), .Y(n_573) );
INVx1_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
AOI221xp5_ASAP7_75t_SL g757 ( .A1(n_532), .A2(n_758), .B1(n_759), .B2(n_761), .C(n_762), .Y(n_757) );
BUFx6f_ASAP7_75t_L g615 ( .A(n_534), .Y(n_615) );
INVx2_ASAP7_75t_L g859 ( .A(n_534), .Y(n_859) );
OAI22xp5_ASAP7_75t_L g565 ( .A1(n_535), .A2(n_566), .B1(n_568), .B2(n_569), .Y(n_565) );
INVx1_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
A2O1A1Ixp33_ASAP7_75t_L g1119 ( .A1(n_538), .A2(n_1120), .B(n_1132), .C(n_1136), .Y(n_1119) );
INVx2_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
INVx1_ASAP7_75t_L g686 ( .A(n_539), .Y(n_686) );
BUFx2_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
INVx1_ASAP7_75t_L g792 ( .A(n_540), .Y(n_792) );
OAI33xp33_ASAP7_75t_L g549 ( .A1(n_550), .A2(n_551), .A3(n_557), .B1(n_565), .B2(n_571), .B3(n_573), .Y(n_549) );
OAI33xp33_ASAP7_75t_L g916 ( .A1(n_550), .A2(n_917), .A3(n_921), .B1(n_924), .B2(n_927), .B3(n_929), .Y(n_916) );
INVx2_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
INVx2_ASAP7_75t_L g883 ( .A(n_553), .Y(n_883) );
INVx4_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
INVx3_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
INVx2_ASAP7_75t_SL g1083 ( .A(n_559), .Y(n_1083) );
BUFx6f_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
INVx3_ASAP7_75t_L g675 ( .A(n_560), .Y(n_675) );
INVx4_ASAP7_75t_L g1151 ( .A(n_560), .Y(n_1151) );
OAI22xp5_ASAP7_75t_L g748 ( .A1(n_561), .A2(n_574), .B1(n_707), .B2(n_749), .Y(n_748) );
INVx2_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
INVx2_ASAP7_75t_SL g576 ( .A(n_562), .Y(n_576) );
INVx4_ASAP7_75t_L g657 ( .A(n_562), .Y(n_657) );
BUFx6f_ASAP7_75t_L g740 ( .A(n_562), .Y(n_740) );
INVx2_ASAP7_75t_L g1003 ( .A(n_562), .Y(n_1003) );
INVx1_ASAP7_75t_L g1086 ( .A(n_562), .Y(n_1086) );
INVx8_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
OR2x2_ASAP7_75t_L g949 ( .A(n_563), .B(n_938), .Y(n_949) );
BUFx2_ASAP7_75t_L g1403 ( .A(n_563), .Y(n_1403) );
BUFx6f_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
INVx4_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
INVx1_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
INVx2_ASAP7_75t_L g923 ( .A(n_570), .Y(n_923) );
INVx2_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
INVx2_ASAP7_75t_L g1410 ( .A(n_572), .Y(n_1410) );
BUFx3_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
INVx2_ASAP7_75t_SL g654 ( .A(n_575), .Y(n_654) );
BUFx3_ASAP7_75t_L g801 ( .A(n_575), .Y(n_801) );
BUFx6f_ASAP7_75t_L g1401 ( .A(n_575), .Y(n_1401) );
OAI22xp5_ASAP7_75t_L g1153 ( .A1(n_576), .A2(n_1073), .B1(n_1154), .B2(n_1155), .Y(n_1153) );
INVx2_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
AND3x2_ASAP7_75t_L g580 ( .A(n_581), .B(n_635), .C(n_646), .Y(n_580) );
AOI211xp5_ASAP7_75t_SL g581 ( .A1(n_582), .A2(n_583), .B(n_588), .C(n_599), .Y(n_581) );
INVxp67_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
INVx2_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
AOI22xp33_ASAP7_75t_L g1016 ( .A1(n_585), .A2(n_1012), .B1(n_1014), .B2(n_1017), .Y(n_1016) );
AND2x4_ASAP7_75t_L g1017 ( .A(n_586), .B(n_1018), .Y(n_1017) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
INVx1_ASAP7_75t_L g634 ( .A(n_587), .Y(n_634) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
AND2x4_ASAP7_75t_L g593 ( .A(n_591), .B(n_594), .Y(n_593) );
AND2x4_ASAP7_75t_L g597 ( .A(n_591), .B(n_598), .Y(n_597) );
INVx1_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
AOI22xp5_ASAP7_75t_L g1022 ( .A1(n_593), .A2(n_1023), .B1(n_1024), .B2(n_1025), .Y(n_1022) );
INVx2_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
AND4x1_ASAP7_75t_SL g1021 ( .A(n_596), .B(n_1022), .C(n_1026), .D(n_1029), .Y(n_1021) );
INVx3_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
BUFx2_ASAP7_75t_L g1033 ( .A(n_598), .Y(n_1033) );
OAI22xp5_ASAP7_75t_L g600 ( .A1(n_601), .A2(n_602), .B1(n_604), .B2(n_605), .Y(n_600) );
INVx1_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
OAI221xp5_ASAP7_75t_L g652 ( .A1(n_604), .A2(n_621), .B1(n_653), .B2(n_655), .C(n_658), .Y(n_652) );
OAI221xp5_ASAP7_75t_L g617 ( .A1(n_605), .A2(n_618), .B1(n_619), .B2(n_621), .C(n_622), .Y(n_617) );
OAI22xp5_ASAP7_75t_L g770 ( .A1(n_605), .A2(n_771), .B1(n_772), .B2(n_774), .Y(n_770) );
OAI22xp5_ASAP7_75t_L g1093 ( .A1(n_605), .A2(n_1078), .B1(n_1087), .B2(n_1094), .Y(n_1093) );
BUFx3_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
INVx1_ASAP7_75t_L g785 ( .A(n_606), .Y(n_785) );
OAI33xp33_ASAP7_75t_L g1088 ( .A1(n_607), .A2(n_1089), .A3(n_1091), .B1(n_1093), .B2(n_1095), .B3(n_1097), .Y(n_1088) );
BUFx3_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
BUFx4f_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
BUFx2_ASAP7_75t_L g901 ( .A(n_609), .Y(n_901) );
BUFx2_ASAP7_75t_L g852 ( .A(n_610), .Y(n_852) );
OAI22xp5_ASAP7_75t_L g611 ( .A1(n_612), .A2(n_614), .B1(n_615), .B2(n_616), .Y(n_611) );
OAI22xp33_ASAP7_75t_L g1089 ( .A1(n_612), .A2(n_1070), .B1(n_1080), .B2(n_1090), .Y(n_1089) );
INVx2_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
OAI221xp5_ASAP7_75t_L g672 ( .A1(n_614), .A2(n_655), .B1(n_673), .B2(n_676), .C(n_677), .Y(n_672) );
OAI22xp33_ASAP7_75t_L g913 ( .A1(n_615), .A2(n_861), .B1(n_914), .B2(n_915), .Y(n_913) );
INVx2_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
INVx2_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
INVx3_ASAP7_75t_L g766 ( .A(n_624), .Y(n_766) );
INVx8_ASAP7_75t_L g840 ( .A(n_624), .Y(n_840) );
INVx2_ASAP7_75t_L g1018 ( .A(n_624), .Y(n_1018) );
OAI33xp33_ASAP7_75t_L g900 ( .A1(n_626), .A2(n_901), .A3(n_902), .B1(n_905), .B2(n_908), .B3(n_913), .Y(n_900) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
AOI33xp33_ASAP7_75t_L g1029 ( .A1(n_627), .A2(n_1030), .A3(n_1032), .B1(n_1034), .B2(n_1038), .B3(n_1040), .Y(n_1029) );
BUFx2_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
INVx3_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
INVx3_ASAP7_75t_L g1096 ( .A(n_629), .Y(n_1096) );
OR2x2_ASAP7_75t_L g631 ( .A(n_632), .B(n_633), .Y(n_631) );
OAI22xp5_ASAP7_75t_L g1097 ( .A1(n_632), .A2(n_1075), .B1(n_1081), .B2(n_1098), .Y(n_1097) );
INVxp67_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
AOI21xp5_ASAP7_75t_L g635 ( .A1(n_636), .A2(n_640), .B(n_641), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g1019 ( .A(n_636), .B(n_1020), .Y(n_1019) );
INVx8_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
AND2x4_ASAP7_75t_L g637 ( .A(n_638), .B(n_639), .Y(n_637) );
INVx1_ASAP7_75t_L g814 ( .A(n_639), .Y(n_814) );
NAND2xp5_ASAP7_75t_L g892 ( .A(n_639), .B(n_893), .Y(n_892) );
INVx5_ASAP7_75t_L g1028 ( .A(n_644), .Y(n_1028) );
OAI31xp33_ASAP7_75t_L g646 ( .A1(n_647), .A2(n_664), .A3(n_681), .B(n_686), .Y(n_646) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
INVx2_ASAP7_75t_L g991 ( .A(n_649), .Y(n_991) );
INVx4_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
INVx2_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
OAI22xp5_ASAP7_75t_L g999 ( .A1(n_653), .A2(n_1000), .B1(n_1001), .B2(n_1004), .Y(n_999) );
OAI22xp5_ASAP7_75t_L g1408 ( .A1(n_653), .A2(n_1382), .B1(n_1403), .B2(n_1409), .Y(n_1408) );
INVx2_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
OAI22xp5_ASAP7_75t_L g929 ( .A1(n_655), .A2(n_907), .B1(n_912), .B2(n_918), .Y(n_929) );
INVx2_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
INVx2_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
HB1xp67_ASAP7_75t_L g920 ( .A(n_657), .Y(n_920) );
OAI22xp5_ASAP7_75t_L g1149 ( .A1(n_657), .A2(n_1131), .B1(n_1150), .B2(n_1151), .Y(n_1149) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
INVx1_ASAP7_75t_L g1146 ( .A(n_660), .Y(n_1146) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
AOI21xp5_ASAP7_75t_L g1006 ( .A1(n_663), .A2(n_1007), .B(n_1009), .Y(n_1006) );
INVxp67_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
HB1xp67_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
BUFx6f_ASAP7_75t_L g1013 ( .A(n_667), .Y(n_1013) );
INVx2_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
NOR2x1_ASAP7_75t_L g669 ( .A(n_670), .B(n_671), .Y(n_669) );
INVx2_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
INVx2_ASAP7_75t_SL g674 ( .A(n_675), .Y(n_674) );
BUFx2_ASAP7_75t_L g747 ( .A(n_678), .Y(n_747) );
INVx1_ASAP7_75t_L g1148 ( .A(n_678), .Y(n_1148) );
INVx3_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
INVx2_ASAP7_75t_L g998 ( .A(n_680), .Y(n_998) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
AOI22xp33_ASAP7_75t_L g1011 ( .A1(n_683), .A2(n_1012), .B1(n_1013), .B2(n_1014), .Y(n_1011) );
INVx3_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
AOI22xp5_ASAP7_75t_L g691 ( .A1(n_692), .A2(n_750), .B1(n_751), .B2(n_818), .Y(n_691) );
INVx2_ASAP7_75t_L g818 ( .A(n_692), .Y(n_818) );
NOR2x1_ASAP7_75t_L g693 ( .A(n_694), .B(n_720), .Y(n_693) );
A2O1A1Ixp33_ASAP7_75t_L g694 ( .A1(n_695), .A2(n_699), .B(n_717), .C(n_718), .Y(n_694) );
NOR3xp33_ASAP7_75t_SL g699 ( .A(n_700), .B(n_710), .C(n_711), .Y(n_699) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
INVx1_ASAP7_75t_L g855 ( .A(n_706), .Y(n_855) );
OAI22xp5_ASAP7_75t_L g736 ( .A1(n_709), .A2(n_737), .B1(n_738), .B2(n_739), .Y(n_736) );
INVx1_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
O2A1O1Ixp5_ASAP7_75t_L g989 ( .A1(n_717), .A2(n_990), .B(n_1005), .C(n_1015), .Y(n_989) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_721), .B(n_732), .Y(n_720) );
AOI22xp5_ASAP7_75t_L g725 ( .A1(n_726), .A2(n_727), .B1(n_728), .B2(n_729), .Y(n_725) );
AOI22xp5_ASAP7_75t_L g889 ( .A1(n_727), .A2(n_729), .B1(n_841), .B2(n_844), .Y(n_889) );
INVx1_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
OAI22xp33_ASAP7_75t_L g1069 ( .A1(n_739), .A2(n_1070), .B1(n_1071), .B2(n_1075), .Y(n_1069) );
INVx5_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
INVx6_ASAP7_75t_L g808 ( .A(n_740), .Y(n_808) );
BUFx2_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
INVx2_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
INVx1_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
NAND4xp75_ASAP7_75t_L g753 ( .A(n_754), .B(n_793), .C(n_812), .D(n_815), .Y(n_753) );
OAI21x1_ASAP7_75t_L g754 ( .A1(n_755), .A2(n_769), .B(n_791), .Y(n_754) );
OAI21xp5_ASAP7_75t_L g755 ( .A1(n_756), .A2(n_757), .B(n_764), .Y(n_755) );
INVx1_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
OAI22xp5_ASAP7_75t_L g1091 ( .A1(n_763), .A2(n_1077), .B1(n_1084), .B2(n_1092), .Y(n_1091) );
A2O1A1Ixp33_ASAP7_75t_L g764 ( .A1(n_765), .A2(n_766), .B(n_767), .C(n_768), .Y(n_764) );
OAI22xp5_ASAP7_75t_L g769 ( .A1(n_770), .A2(n_775), .B1(n_779), .B2(n_786), .Y(n_769) );
OAI22xp5_ASAP7_75t_L g800 ( .A1(n_771), .A2(n_780), .B1(n_801), .B2(n_802), .Y(n_800) );
INVx1_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
OAI221xp5_ASAP7_75t_L g805 ( .A1(n_774), .A2(n_787), .B1(n_806), .B2(n_808), .C(n_809), .Y(n_805) );
OAI22xp5_ASAP7_75t_L g779 ( .A1(n_780), .A2(n_781), .B1(n_782), .B2(n_783), .Y(n_779) );
INVx3_ASAP7_75t_L g783 ( .A(n_784), .Y(n_783) );
BUFx2_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
INVx2_ASAP7_75t_L g788 ( .A(n_789), .Y(n_788) );
INVx1_ASAP7_75t_L g791 ( .A(n_792), .Y(n_791) );
AOI211x1_ASAP7_75t_L g793 ( .A1(n_794), .A2(n_795), .B(n_803), .C(n_811), .Y(n_793) );
INVx2_ASAP7_75t_L g796 ( .A(n_797), .Y(n_796) );
INVx2_ASAP7_75t_L g797 ( .A(n_798), .Y(n_797) );
INVx2_ASAP7_75t_L g798 ( .A(n_799), .Y(n_798) );
INVx1_ASAP7_75t_L g919 ( .A(n_801), .Y(n_919) );
BUFx2_ASAP7_75t_L g1101 ( .A(n_802), .Y(n_1101) );
OAI22xp5_ASAP7_75t_L g1404 ( .A1(n_802), .A2(n_806), .B1(n_1381), .B2(n_1405), .Y(n_1404) );
INVx2_ASAP7_75t_L g806 ( .A(n_807), .Y(n_806) );
INVx1_ASAP7_75t_L g813 ( .A(n_814), .Y(n_813) );
INVx1_ASAP7_75t_L g821 ( .A(n_822), .Y(n_821) );
XNOR2xp5_ASAP7_75t_L g822 ( .A(n_823), .B(n_895), .Y(n_822) );
HB1xp67_ASAP7_75t_L g823 ( .A(n_824), .Y(n_823) );
INVx1_ASAP7_75t_L g825 ( .A(n_826), .Y(n_825) );
NAND3xp33_ASAP7_75t_L g826 ( .A(n_827), .B(n_834), .C(n_871), .Y(n_826) );
NAND2xp5_ASAP7_75t_L g829 ( .A(n_830), .B(n_831), .Y(n_829) );
AOI22xp33_ASAP7_75t_L g839 ( .A1(n_832), .A2(n_840), .B1(n_841), .B2(n_842), .Y(n_839) );
OAI21xp33_ASAP7_75t_L g834 ( .A1(n_835), .A2(n_856), .B(n_869), .Y(n_834) );
OAI211xp5_ASAP7_75t_L g835 ( .A1(n_836), .A2(n_839), .B(n_843), .C(n_846), .Y(n_835) );
INVxp67_ASAP7_75t_L g836 ( .A(n_837), .Y(n_836) );
INVx1_ASAP7_75t_L g837 ( .A(n_838), .Y(n_837) );
OAI211xp5_ASAP7_75t_L g846 ( .A1(n_847), .A2(n_848), .B(n_849), .C(n_853), .Y(n_846) );
OAI221xp5_ASAP7_75t_L g882 ( .A1(n_847), .A2(n_860), .B1(n_883), .B2(n_884), .C(n_885), .Y(n_882) );
INVx1_ASAP7_75t_L g850 ( .A(n_851), .Y(n_850) );
INVx1_ASAP7_75t_L g858 ( .A(n_859), .Y(n_858) );
INVx2_ASAP7_75t_L g861 ( .A(n_862), .Y(n_861) );
OAI22xp5_ASAP7_75t_L g864 ( .A1(n_865), .A2(n_866), .B1(n_867), .B2(n_868), .Y(n_864) );
INVx1_ASAP7_75t_L g869 ( .A(n_870), .Y(n_869) );
A2O1A1Ixp33_ASAP7_75t_SL g1371 ( .A1(n_870), .A2(n_1372), .B(n_1388), .C(n_1393), .Y(n_1371) );
NOR3xp33_ASAP7_75t_L g871 ( .A(n_872), .B(n_881), .C(n_890), .Y(n_871) );
INVxp67_ASAP7_75t_L g873 ( .A(n_874), .Y(n_873) );
OAI22xp5_ASAP7_75t_L g921 ( .A1(n_876), .A2(n_906), .B1(n_910), .B2(n_922), .Y(n_921) );
OAI22xp5_ASAP7_75t_L g1079 ( .A1(n_883), .A2(n_993), .B1(n_1080), .B2(n_1081), .Y(n_1079) );
OAI22xp5_ASAP7_75t_L g924 ( .A1(n_884), .A2(n_904), .B1(n_915), .B2(n_925), .Y(n_924) );
INVx2_ASAP7_75t_L g886 ( .A(n_887), .Y(n_886) );
INVx1_ASAP7_75t_L g891 ( .A(n_892), .Y(n_891) );
AO22x2_ASAP7_75t_L g895 ( .A1(n_896), .A2(n_1042), .B1(n_1043), .B2(n_1160), .Y(n_895) );
INVx1_ASAP7_75t_L g1160 ( .A(n_896), .Y(n_1160) );
XNOR2xp5_ASAP7_75t_L g896 ( .A(n_897), .B(n_987), .Y(n_896) );
NAND3xp33_ASAP7_75t_L g898 ( .A(n_899), .B(n_930), .C(n_957), .Y(n_898) );
NOR2xp33_ASAP7_75t_L g899 ( .A(n_900), .B(n_916), .Y(n_899) );
OAI22xp5_ASAP7_75t_SL g917 ( .A1(n_903), .A2(n_914), .B1(n_918), .B2(n_920), .Y(n_917) );
OAI22xp5_ASAP7_75t_L g908 ( .A1(n_909), .A2(n_910), .B1(n_911), .B2(n_912), .Y(n_908) );
INVx2_ASAP7_75t_L g918 ( .A(n_919), .Y(n_918) );
HB1xp67_ASAP7_75t_L g922 ( .A(n_923), .Y(n_922) );
INVx3_ASAP7_75t_L g925 ( .A(n_926), .Y(n_925) );
OAI33xp33_ASAP7_75t_L g1066 ( .A1(n_927), .A2(n_1067), .A3(n_1069), .B1(n_1076), .B2(n_1079), .B3(n_1082), .Y(n_1066) );
INVx2_ASAP7_75t_L g927 ( .A(n_928), .Y(n_927) );
OAI31xp33_ASAP7_75t_L g930 ( .A1(n_931), .A2(n_943), .A3(n_950), .B(n_954), .Y(n_930) );
INVx3_ASAP7_75t_L g932 ( .A(n_933), .Y(n_932) );
AOI22xp33_ASAP7_75t_L g935 ( .A1(n_936), .A2(n_937), .B1(n_939), .B2(n_940), .Y(n_935) );
AOI22xp33_ASAP7_75t_L g966 ( .A1(n_936), .A2(n_967), .B1(n_971), .B2(n_974), .Y(n_966) );
BUFx3_ASAP7_75t_L g1103 ( .A(n_937), .Y(n_1103) );
INVx2_ASAP7_75t_L g940 ( .A(n_941), .Y(n_940) );
INVx2_ASAP7_75t_L g941 ( .A(n_942), .Y(n_941) );
INVx2_ASAP7_75t_L g1106 ( .A(n_942), .Y(n_1106) );
HB1xp67_ASAP7_75t_L g944 ( .A(n_945), .Y(n_944) );
INVx1_ASAP7_75t_L g1109 ( .A(n_945), .Y(n_1109) );
INVx2_ASAP7_75t_L g947 ( .A(n_948), .Y(n_947) );
INVx2_ASAP7_75t_L g948 ( .A(n_949), .Y(n_948) );
BUFx2_ASAP7_75t_L g1111 ( .A(n_949), .Y(n_1111) );
INVx3_ASAP7_75t_SL g952 ( .A(n_953), .Y(n_952) );
CKINVDCx16_ASAP7_75t_R g1113 ( .A(n_953), .Y(n_1113) );
OAI31xp33_ASAP7_75t_L g1099 ( .A1(n_954), .A2(n_1100), .A3(n_1107), .B(n_1112), .Y(n_1099) );
BUFx3_ASAP7_75t_L g954 ( .A(n_955), .Y(n_954) );
OAI31xp33_ASAP7_75t_L g957 ( .A1(n_958), .A2(n_963), .A3(n_975), .B(n_981), .Y(n_957) );
INVx2_ASAP7_75t_SL g1052 ( .A(n_959), .Y(n_1052) );
INVx2_ASAP7_75t_L g960 ( .A(n_961), .Y(n_960) );
INVx1_ASAP7_75t_L g1053 ( .A(n_961), .Y(n_1053) );
CKINVDCx8_ASAP7_75t_R g964 ( .A(n_965), .Y(n_964) );
BUFx3_ASAP7_75t_L g967 ( .A(n_968), .Y(n_967) );
BUFx3_ASAP7_75t_L g1058 ( .A(n_968), .Y(n_1058) );
AND2x2_ASAP7_75t_L g968 ( .A(n_969), .B(n_970), .Y(n_968) );
AND2x4_ASAP7_75t_L g972 ( .A(n_969), .B(n_973), .Y(n_972) );
AOI22xp33_ASAP7_75t_L g1057 ( .A1(n_971), .A2(n_1058), .B1(n_1059), .B2(n_1060), .Y(n_1057) );
BUFx6f_ASAP7_75t_L g971 ( .A(n_972), .Y(n_971) );
INVx1_ASAP7_75t_L g976 ( .A(n_977), .Y(n_976) );
INVx2_ASAP7_75t_SL g977 ( .A(n_978), .Y(n_977) );
BUFx2_ASAP7_75t_L g1062 ( .A(n_978), .Y(n_1062) );
BUFx3_ASAP7_75t_L g979 ( .A(n_980), .Y(n_979) );
INVx2_ASAP7_75t_L g1064 ( .A(n_980), .Y(n_1064) );
BUFx2_ASAP7_75t_L g981 ( .A(n_982), .Y(n_981) );
AND2x2_ASAP7_75t_SL g982 ( .A(n_983), .B(n_985), .Y(n_982) );
AND2x4_ASAP7_75t_L g1048 ( .A(n_983), .B(n_985), .Y(n_1048) );
INVx1_ASAP7_75t_SL g983 ( .A(n_984), .Y(n_983) );
INVx1_ASAP7_75t_L g985 ( .A(n_986), .Y(n_985) );
NAND3x1_ASAP7_75t_L g988 ( .A(n_989), .B(n_1019), .C(n_1021), .Y(n_988) );
INVx5_ASAP7_75t_L g993 ( .A(n_994), .Y(n_993) );
INVx1_ASAP7_75t_L g997 ( .A(n_998), .Y(n_997) );
BUFx2_ASAP7_75t_L g1001 ( .A(n_1002), .Y(n_1001) );
BUFx6f_ASAP7_75t_L g1002 ( .A(n_1003), .Y(n_1002) );
NAND2xp5_ASAP7_75t_L g1026 ( .A(n_1027), .B(n_1028), .Y(n_1026) );
BUFx3_ASAP7_75t_L g1030 ( .A(n_1031), .Y(n_1030) );
INVx8_ASAP7_75t_L g1035 ( .A(n_1036), .Y(n_1035) );
INVx1_ASAP7_75t_L g1042 ( .A(n_1043), .Y(n_1042) );
AOI22xp5_ASAP7_75t_L g1043 ( .A1(n_1044), .A2(n_1045), .B1(n_1116), .B2(n_1117), .Y(n_1043) );
INVx2_ASAP7_75t_L g1044 ( .A(n_1045), .Y(n_1044) );
INVx1_ASAP7_75t_L g1114 ( .A(n_1046), .Y(n_1114) );
OAI211xp5_ASAP7_75t_L g1046 ( .A1(n_1047), .A2(n_1049), .B(n_1065), .C(n_1099), .Y(n_1046) );
CKINVDCx14_ASAP7_75t_R g1047 ( .A(n_1048), .Y(n_1047) );
NOR3xp33_ASAP7_75t_SL g1049 ( .A(n_1050), .B(n_1054), .C(n_1061), .Y(n_1049) );
INVx2_ASAP7_75t_L g1051 ( .A(n_1052), .Y(n_1051) );
INVx1_ASAP7_75t_L g1055 ( .A(n_1056), .Y(n_1055) );
AOI22xp33_ASAP7_75t_L g1102 ( .A1(n_1059), .A2(n_1103), .B1(n_1104), .B2(n_1105), .Y(n_1102) );
INVx1_ASAP7_75t_L g1063 ( .A(n_1064), .Y(n_1063) );
NOR2xp33_ASAP7_75t_L g1065 ( .A(n_1066), .B(n_1088), .Y(n_1065) );
BUFx6f_ASAP7_75t_L g1067 ( .A(n_1068), .Y(n_1067) );
INVx1_ASAP7_75t_L g1071 ( .A(n_1072), .Y(n_1071) );
INVx1_ASAP7_75t_L g1072 ( .A(n_1073), .Y(n_1072) );
INVx1_ASAP7_75t_L g1073 ( .A(n_1074), .Y(n_1073) );
OAI22xp5_ASAP7_75t_L g1082 ( .A1(n_1083), .A2(n_1084), .B1(n_1085), .B2(n_1087), .Y(n_1082) );
BUFx3_ASAP7_75t_L g1085 ( .A(n_1086), .Y(n_1085) );
INVx2_ASAP7_75t_L g1095 ( .A(n_1096), .Y(n_1095) );
INVx2_ASAP7_75t_L g1105 ( .A(n_1106), .Y(n_1105) );
INVx1_ASAP7_75t_L g1108 ( .A(n_1109), .Y(n_1108) );
HB1xp67_ASAP7_75t_L g1110 ( .A(n_1111), .Y(n_1110) );
INVx1_ASAP7_75t_L g1116 ( .A(n_1117), .Y(n_1116) );
OR2x2_ASAP7_75t_L g1118 ( .A(n_1119), .B(n_1139), .Y(n_1118) );
NOR3xp33_ASAP7_75t_L g1120 ( .A(n_1121), .B(n_1122), .C(n_1126), .Y(n_1120) );
INVx1_ASAP7_75t_L g1127 ( .A(n_1128), .Y(n_1127) );
NAND2xp5_ASAP7_75t_L g1136 ( .A(n_1137), .B(n_1138), .Y(n_1136) );
NAND4xp25_ASAP7_75t_L g1139 ( .A(n_1140), .B(n_1143), .C(n_1156), .D(n_1158), .Y(n_1139) );
INVx1_ASAP7_75t_L g1147 ( .A(n_1148), .Y(n_1147) );
OAI221xp5_ASAP7_75t_L g1161 ( .A1(n_1162), .A2(n_1365), .B1(n_1368), .B2(n_1415), .C(n_1419), .Y(n_1161) );
NOR2xp67_ASAP7_75t_SL g1162 ( .A(n_1163), .B(n_1303), .Y(n_1162) );
NAND2xp5_ASAP7_75t_L g1163 ( .A(n_1164), .B(n_1264), .Y(n_1163) );
A2O1A1Ixp33_ASAP7_75t_SL g1164 ( .A1(n_1165), .A2(n_1180), .B(n_1213), .C(n_1259), .Y(n_1164) );
AND2x2_ASAP7_75t_L g1229 ( .A(n_1165), .B(n_1230), .Y(n_1229) );
INVx1_ASAP7_75t_L g1274 ( .A(n_1165), .Y(n_1274) );
NAND2xp5_ASAP7_75t_L g1301 ( .A(n_1165), .B(n_1302), .Y(n_1301) );
AND2x2_ASAP7_75t_L g1326 ( .A(n_1165), .B(n_1251), .Y(n_1326) );
INVx1_ASAP7_75t_L g1357 ( .A(n_1165), .Y(n_1357) );
AND2x2_ASAP7_75t_L g1362 ( .A(n_1165), .B(n_1197), .Y(n_1362) );
INVx1_ASAP7_75t_L g1165 ( .A(n_1166), .Y(n_1165) );
INVx1_ASAP7_75t_L g1216 ( .A(n_1166), .Y(n_1216) );
INVx1_ASAP7_75t_L g1288 ( .A(n_1166), .Y(n_1288) );
AND2x2_ASAP7_75t_L g1294 ( .A(n_1166), .B(n_1211), .Y(n_1294) );
NAND2xp5_ASAP7_75t_L g1321 ( .A(n_1166), .B(n_1258), .Y(n_1321) );
AND2x2_ASAP7_75t_L g1353 ( .A(n_1166), .B(n_1197), .Y(n_1353) );
NAND2xp5_ASAP7_75t_L g1166 ( .A(n_1167), .B(n_1174), .Y(n_1166) );
AND2x6_ASAP7_75t_L g1168 ( .A(n_1169), .B(n_1170), .Y(n_1168) );
AND2x2_ASAP7_75t_L g1172 ( .A(n_1169), .B(n_1173), .Y(n_1172) );
AND2x4_ASAP7_75t_L g1175 ( .A(n_1169), .B(n_1176), .Y(n_1175) );
AND2x6_ASAP7_75t_L g1178 ( .A(n_1169), .B(n_1179), .Y(n_1178) );
AND2x2_ASAP7_75t_L g1189 ( .A(n_1169), .B(n_1173), .Y(n_1189) );
AND2x2_ASAP7_75t_L g1262 ( .A(n_1169), .B(n_1173), .Y(n_1262) );
AND2x2_ASAP7_75t_L g1176 ( .A(n_1171), .B(n_1177), .Y(n_1176) );
INVx2_ASAP7_75t_L g1367 ( .A(n_1178), .Y(n_1367) );
HB1xp67_ASAP7_75t_L g1430 ( .A(n_1179), .Y(n_1430) );
OAI22xp5_ASAP7_75t_L g1180 ( .A1(n_1181), .A2(n_1196), .B1(n_1203), .B2(n_1212), .Y(n_1180) );
INVx1_ASAP7_75t_L g1181 ( .A(n_1182), .Y(n_1181) );
NOR2xp33_ASAP7_75t_L g1182 ( .A(n_1183), .B(n_1193), .Y(n_1182) );
NAND2xp5_ASAP7_75t_L g1313 ( .A(n_1183), .B(n_1200), .Y(n_1313) );
INVx1_ASAP7_75t_L g1183 ( .A(n_1184), .Y(n_1183) );
OR2x2_ASAP7_75t_L g1225 ( .A(n_1184), .B(n_1222), .Y(n_1225) );
OR2x2_ASAP7_75t_L g1277 ( .A(n_1184), .B(n_1228), .Y(n_1277) );
OR2x2_ASAP7_75t_L g1184 ( .A(n_1185), .B(n_1190), .Y(n_1184) );
AND2x2_ASAP7_75t_L g1221 ( .A(n_1185), .B(n_1222), .Y(n_1221) );
AND2x2_ASAP7_75t_L g1244 ( .A(n_1185), .B(n_1245), .Y(n_1244) );
A2O1A1Ixp33_ASAP7_75t_L g1306 ( .A1(n_1185), .A2(n_1288), .B(n_1307), .C(n_1309), .Y(n_1306) );
INVx1_ASAP7_75t_L g1185 ( .A(n_1186), .Y(n_1185) );
OR2x2_ASAP7_75t_L g1194 ( .A(n_1186), .B(n_1195), .Y(n_1194) );
AND2x2_ASAP7_75t_L g1237 ( .A(n_1186), .B(n_1190), .Y(n_1237) );
OR2x2_ASAP7_75t_L g1332 ( .A(n_1186), .B(n_1222), .Y(n_1332) );
NOR2xp33_ASAP7_75t_L g1337 ( .A(n_1186), .B(n_1338), .Y(n_1337) );
AND2x2_ASAP7_75t_L g1186 ( .A(n_1187), .B(n_1188), .Y(n_1186) );
INVx1_ASAP7_75t_L g1195 ( .A(n_1190), .Y(n_1195) );
INVx1_ASAP7_75t_L g1212 ( .A(n_1190), .Y(n_1212) );
INVx1_ASAP7_75t_L g1245 ( .A(n_1190), .Y(n_1245) );
NAND2xp5_ASAP7_75t_L g1297 ( .A(n_1190), .B(n_1228), .Y(n_1297) );
NAND2x1_ASAP7_75t_L g1190 ( .A(n_1191), .B(n_1192), .Y(n_1190) );
AND2x2_ASAP7_75t_L g1329 ( .A(n_1193), .B(n_1228), .Y(n_1329) );
INVx1_ASAP7_75t_L g1193 ( .A(n_1194), .Y(n_1193) );
OR2x2_ASAP7_75t_L g1227 ( .A(n_1194), .B(n_1228), .Y(n_1227) );
NAND2xp5_ASAP7_75t_L g1196 ( .A(n_1197), .B(n_1200), .Y(n_1196) );
CKINVDCx5p33_ASAP7_75t_R g1211 ( .A(n_1197), .Y(n_1211) );
OR2x2_ASAP7_75t_L g1231 ( .A(n_1197), .B(n_1208), .Y(n_1231) );
NAND2xp5_ASAP7_75t_L g1247 ( .A(n_1197), .B(n_1248), .Y(n_1247) );
OAI22xp5_ASAP7_75t_L g1327 ( .A1(n_1197), .A2(n_1291), .B1(n_1310), .B2(n_1328), .Y(n_1327) );
AND2x4_ASAP7_75t_L g1197 ( .A(n_1198), .B(n_1199), .Y(n_1197) );
INVx3_ASAP7_75t_L g1205 ( .A(n_1200), .Y(n_1205) );
CKINVDCx5p33_ASAP7_75t_R g1220 ( .A(n_1200), .Y(n_1220) );
AND2x2_ASAP7_75t_L g1246 ( .A(n_1200), .B(n_1222), .Y(n_1246) );
NAND2xp5_ASAP7_75t_L g1270 ( .A(n_1200), .B(n_1244), .Y(n_1270) );
AND2x2_ASAP7_75t_L g1298 ( .A(n_1200), .B(n_1274), .Y(n_1298) );
AND2x4_ASAP7_75t_SL g1200 ( .A(n_1201), .B(n_1202), .Y(n_1200) );
INVx1_ASAP7_75t_L g1203 ( .A(n_1204), .Y(n_1203) );
NOR2xp33_ASAP7_75t_L g1204 ( .A(n_1205), .B(n_1206), .Y(n_1204) );
NAND2xp5_ASAP7_75t_L g1254 ( .A(n_1205), .B(n_1228), .Y(n_1254) );
AND2x2_ASAP7_75t_L g1258 ( .A(n_1205), .B(n_1207), .Y(n_1258) );
NOR2xp33_ASAP7_75t_L g1316 ( .A(n_1205), .B(n_1317), .Y(n_1316) );
NAND2xp5_ASAP7_75t_L g1324 ( .A(n_1205), .B(n_1237), .Y(n_1324) );
CKINVDCx14_ASAP7_75t_R g1343 ( .A(n_1205), .Y(n_1343) );
AND2x2_ASAP7_75t_L g1346 ( .A(n_1205), .B(n_1226), .Y(n_1346) );
AOI211xp5_ASAP7_75t_L g1272 ( .A1(n_1206), .A2(n_1273), .B(n_1275), .C(n_1278), .Y(n_1272) );
OR2x2_ASAP7_75t_L g1206 ( .A(n_1207), .B(n_1211), .Y(n_1206) );
AND2x2_ASAP7_75t_L g1267 ( .A(n_1207), .B(n_1268), .Y(n_1267) );
INVx2_ASAP7_75t_L g1317 ( .A(n_1207), .Y(n_1317) );
NOR2xp33_ASAP7_75t_L g1340 ( .A(n_1207), .B(n_1269), .Y(n_1340) );
NAND2xp5_ASAP7_75t_L g1341 ( .A(n_1207), .B(n_1342), .Y(n_1341) );
INVx2_ASAP7_75t_SL g1207 ( .A(n_1208), .Y(n_1207) );
NAND2xp5_ASAP7_75t_L g1241 ( .A(n_1208), .B(n_1211), .Y(n_1241) );
INVx1_ASAP7_75t_L g1248 ( .A(n_1208), .Y(n_1248) );
AND2x2_ASAP7_75t_L g1208 ( .A(n_1209), .B(n_1210), .Y(n_1208) );
AND2x2_ASAP7_75t_L g1215 ( .A(n_1211), .B(n_1216), .Y(n_1215) );
NAND3xp33_ASAP7_75t_L g1315 ( .A(n_1211), .B(n_1237), .C(n_1316), .Y(n_1315) );
AND2x2_ASAP7_75t_L g1320 ( .A(n_1212), .B(n_1228), .Y(n_1320) );
NAND4xp25_ASAP7_75t_SL g1213 ( .A(n_1214), .B(n_1232), .C(n_1249), .D(n_1255), .Y(n_1213) );
AOI22xp5_ASAP7_75t_L g1214 ( .A1(n_1215), .A2(n_1217), .B1(n_1226), .B2(n_1229), .Y(n_1214) );
INVx1_ASAP7_75t_L g1271 ( .A(n_1216), .Y(n_1271) );
OAI211xp5_ASAP7_75t_L g1335 ( .A1(n_1216), .A2(n_1336), .B(n_1339), .C(n_1341), .Y(n_1335) );
NAND2xp5_ASAP7_75t_L g1217 ( .A(n_1218), .B(n_1225), .Y(n_1217) );
INVx1_ASAP7_75t_L g1218 ( .A(n_1219), .Y(n_1218) );
OAI21xp5_ASAP7_75t_L g1283 ( .A1(n_1219), .A2(n_1230), .B(n_1284), .Y(n_1283) );
AND2x2_ASAP7_75t_L g1219 ( .A(n_1220), .B(n_1221), .Y(n_1219) );
NAND2xp5_ASAP7_75t_L g1239 ( .A(n_1220), .B(n_1240), .Y(n_1239) );
INVx1_ASAP7_75t_L g1276 ( .A(n_1220), .Y(n_1276) );
AND2x2_ASAP7_75t_L g1292 ( .A(n_1220), .B(n_1290), .Y(n_1292) );
OR2x2_ASAP7_75t_L g1308 ( .A(n_1220), .B(n_1247), .Y(n_1308) );
NOR2xp33_ASAP7_75t_L g1309 ( .A(n_1220), .B(n_1310), .Y(n_1309) );
INVx2_ASAP7_75t_L g1228 ( .A(n_1222), .Y(n_1228) );
OR2x2_ASAP7_75t_L g1269 ( .A(n_1222), .B(n_1270), .Y(n_1269) );
AND2x2_ASAP7_75t_L g1290 ( .A(n_1222), .B(n_1245), .Y(n_1290) );
AOI22xp33_ASAP7_75t_L g1330 ( .A1(n_1222), .A2(n_1331), .B1(n_1333), .B2(n_1334), .Y(n_1330) );
AND2x2_ASAP7_75t_L g1222 ( .A(n_1223), .B(n_1224), .Y(n_1222) );
INVx1_ASAP7_75t_L g1233 ( .A(n_1225), .Y(n_1233) );
INVx1_ASAP7_75t_L g1226 ( .A(n_1227), .Y(n_1226) );
NOR2xp33_ASAP7_75t_L g1256 ( .A(n_1227), .B(n_1257), .Y(n_1256) );
OR2x2_ASAP7_75t_L g1235 ( .A(n_1228), .B(n_1236), .Y(n_1235) );
NAND2xp5_ASAP7_75t_L g1300 ( .A(n_1228), .B(n_1244), .Y(n_1300) );
OR2x2_ASAP7_75t_L g1360 ( .A(n_1228), .B(n_1324), .Y(n_1360) );
NAND2xp5_ASAP7_75t_L g1286 ( .A(n_1230), .B(n_1287), .Y(n_1286) );
INVx2_ASAP7_75t_L g1230 ( .A(n_1231), .Y(n_1230) );
O2A1O1Ixp33_ASAP7_75t_L g1232 ( .A1(n_1233), .A2(n_1234), .B(n_1238), .C(n_1242), .Y(n_1232) );
AOI22xp5_ASAP7_75t_L g1336 ( .A1(n_1233), .A2(n_1241), .B1(n_1317), .B2(n_1337), .Y(n_1336) );
INVx1_ASAP7_75t_L g1234 ( .A(n_1235), .Y(n_1234) );
AOI21xp5_ASAP7_75t_L g1242 ( .A1(n_1235), .A2(n_1243), .B(n_1247), .Y(n_1242) );
OR2x2_ASAP7_75t_L g1253 ( .A(n_1236), .B(n_1254), .Y(n_1253) );
INVx1_ASAP7_75t_L g1236 ( .A(n_1237), .Y(n_1236) );
AND2x2_ASAP7_75t_L g1268 ( .A(n_1237), .B(n_1246), .Y(n_1268) );
OAI211xp5_ASAP7_75t_L g1295 ( .A1(n_1237), .A2(n_1240), .B(n_1296), .C(n_1298), .Y(n_1295) );
INVx1_ASAP7_75t_L g1238 ( .A(n_1239), .Y(n_1238) );
INVx1_ASAP7_75t_L g1310 ( .A(n_1240), .Y(n_1310) );
INVx1_ASAP7_75t_L g1240 ( .A(n_1241), .Y(n_1240) );
OR2x2_ASAP7_75t_L g1356 ( .A(n_1241), .B(n_1357), .Y(n_1356) );
NAND2xp5_ASAP7_75t_L g1243 ( .A(n_1244), .B(n_1246), .Y(n_1243) );
AND2x2_ASAP7_75t_L g1348 ( .A(n_1244), .B(n_1349), .Y(n_1348) );
INVx1_ASAP7_75t_L g1338 ( .A(n_1246), .Y(n_1338) );
INVx1_ASAP7_75t_L g1282 ( .A(n_1247), .Y(n_1282) );
INVx1_ASAP7_75t_L g1302 ( .A(n_1247), .Y(n_1302) );
INVx2_ASAP7_75t_L g1251 ( .A(n_1248), .Y(n_1251) );
NAND2xp5_ASAP7_75t_L g1249 ( .A(n_1250), .B(n_1252), .Y(n_1249) );
INVx1_ASAP7_75t_L g1250 ( .A(n_1251), .Y(n_1250) );
OR2x2_ASAP7_75t_L g1273 ( .A(n_1251), .B(n_1274), .Y(n_1273) );
AOI21xp5_ASAP7_75t_L g1347 ( .A1(n_1251), .A2(n_1348), .B(n_1350), .Y(n_1347) );
INVx1_ASAP7_75t_L g1252 ( .A(n_1253), .Y(n_1252) );
A2O1A1Ixp33_ASAP7_75t_L g1279 ( .A1(n_1253), .A2(n_1280), .B(n_1281), .C(n_1283), .Y(n_1279) );
INVx1_ASAP7_75t_L g1349 ( .A(n_1254), .Y(n_1349) );
INVx1_ASAP7_75t_L g1255 ( .A(n_1256), .Y(n_1255) );
INVx1_ASAP7_75t_L g1257 ( .A(n_1258), .Y(n_1257) );
CKINVDCx14_ASAP7_75t_R g1278 ( .A(n_1259), .Y(n_1278) );
A2O1A1Ixp33_ASAP7_75t_L g1344 ( .A1(n_1259), .A2(n_1345), .B(n_1347), .C(n_1352), .Y(n_1344) );
INVx3_ASAP7_75t_L g1259 ( .A(n_1260), .Y(n_1259) );
OAI221xp5_ASAP7_75t_L g1318 ( .A1(n_1260), .A2(n_1289), .B1(n_1293), .B2(n_1319), .C(n_1321), .Y(n_1318) );
AND2x2_ASAP7_75t_L g1260 ( .A(n_1261), .B(n_1263), .Y(n_1260) );
NOR5xp2_ASAP7_75t_L g1264 ( .A(n_1265), .B(n_1272), .C(n_1279), .D(n_1285), .E(n_1299), .Y(n_1264) );
AOI21xp33_ASAP7_75t_L g1265 ( .A1(n_1266), .A2(n_1269), .B(n_1271), .Y(n_1265) );
INVx1_ASAP7_75t_L g1266 ( .A(n_1267), .Y(n_1266) );
INVxp67_ASAP7_75t_L g1280 ( .A(n_1268), .Y(n_1280) );
OR2x2_ASAP7_75t_L g1275 ( .A(n_1276), .B(n_1277), .Y(n_1275) );
INVx2_ASAP7_75t_L g1284 ( .A(n_1277), .Y(n_1284) );
INVx1_ASAP7_75t_L g1281 ( .A(n_1282), .Y(n_1281) );
AOI211xp5_ASAP7_75t_L g1311 ( .A1(n_1282), .A2(n_1312), .B(n_1314), .C(n_1318), .Y(n_1311) );
NAND2xp5_ASAP7_75t_L g1351 ( .A(n_1284), .B(n_1343), .Y(n_1351) );
OAI221xp5_ASAP7_75t_SL g1285 ( .A1(n_1286), .A2(n_1289), .B1(n_1291), .B2(n_1293), .C(n_1295), .Y(n_1285) );
INVx1_ASAP7_75t_L g1334 ( .A(n_1286), .Y(n_1334) );
INVx1_ASAP7_75t_L g1287 ( .A(n_1288), .Y(n_1287) );
INVx1_ASAP7_75t_L g1289 ( .A(n_1290), .Y(n_1289) );
INVx1_ASAP7_75t_L g1291 ( .A(n_1292), .Y(n_1291) );
INVx1_ASAP7_75t_L g1293 ( .A(n_1294), .Y(n_1293) );
INVx1_ASAP7_75t_L g1296 ( .A(n_1297), .Y(n_1296) );
NOR2xp33_ASAP7_75t_L g1299 ( .A(n_1300), .B(n_1301), .Y(n_1299) );
INVx1_ASAP7_75t_L g1325 ( .A(n_1300), .Y(n_1325) );
INVx1_ASAP7_75t_L g1333 ( .A(n_1301), .Y(n_1333) );
NAND2xp5_ASAP7_75t_L g1303 ( .A(n_1304), .B(n_1354), .Y(n_1303) );
OAI21xp5_ASAP7_75t_L g1304 ( .A1(n_1305), .A2(n_1335), .B(n_1344), .Y(n_1304) );
NAND4xp25_ASAP7_75t_L g1305 ( .A(n_1306), .B(n_1311), .C(n_1322), .D(n_1330), .Y(n_1305) );
INVx1_ASAP7_75t_L g1307 ( .A(n_1308), .Y(n_1307) );
INVx1_ASAP7_75t_L g1312 ( .A(n_1313), .Y(n_1312) );
INVx1_ASAP7_75t_L g1314 ( .A(n_1315), .Y(n_1314) );
OAI21xp5_ASAP7_75t_SL g1355 ( .A1(n_1319), .A2(n_1356), .B(n_1358), .Y(n_1355) );
INVx1_ASAP7_75t_L g1319 ( .A(n_1320), .Y(n_1319) );
O2A1O1Ixp33_ASAP7_75t_L g1322 ( .A1(n_1323), .A2(n_1325), .B(n_1326), .C(n_1327), .Y(n_1322) );
AOI22xp5_ASAP7_75t_L g1354 ( .A1(n_1323), .A2(n_1343), .B1(n_1355), .B2(n_1363), .Y(n_1354) );
INVx1_ASAP7_75t_L g1323 ( .A(n_1324), .Y(n_1323) );
INVx2_ASAP7_75t_L g1328 ( .A(n_1329), .Y(n_1328) );
AND2x2_ASAP7_75t_L g1342 ( .A(n_1329), .B(n_1343), .Y(n_1342) );
OAI31xp33_ASAP7_75t_L g1358 ( .A1(n_1331), .A2(n_1359), .A3(n_1361), .B(n_1362), .Y(n_1358) );
INVx1_ASAP7_75t_L g1331 ( .A(n_1332), .Y(n_1331) );
A2O1A1Ixp33_ASAP7_75t_L g1363 ( .A1(n_1332), .A2(n_1356), .B(n_1360), .C(n_1364), .Y(n_1363) );
INVxp67_ASAP7_75t_SL g1339 ( .A(n_1340), .Y(n_1339) );
INVx1_ASAP7_75t_L g1345 ( .A(n_1346), .Y(n_1345) );
INVx1_ASAP7_75t_L g1350 ( .A(n_1351), .Y(n_1350) );
INVx1_ASAP7_75t_L g1352 ( .A(n_1353), .Y(n_1352) );
INVx1_ASAP7_75t_L g1361 ( .A(n_1356), .Y(n_1361) );
INVx1_ASAP7_75t_L g1359 ( .A(n_1360), .Y(n_1359) );
INVx1_ASAP7_75t_L g1364 ( .A(n_1362), .Y(n_1364) );
CKINVDCx20_ASAP7_75t_R g1365 ( .A(n_1366), .Y(n_1365) );
CKINVDCx20_ASAP7_75t_R g1366 ( .A(n_1367), .Y(n_1366) );
BUFx2_ASAP7_75t_SL g1368 ( .A(n_1369), .Y(n_1368) );
HB1xp67_ASAP7_75t_L g1424 ( .A(n_1370), .Y(n_1424) );
OR2x2_ASAP7_75t_L g1370 ( .A(n_1371), .B(n_1396), .Y(n_1370) );
OAI21xp33_ASAP7_75t_L g1375 ( .A1(n_1376), .A2(n_1380), .B(n_1383), .Y(n_1375) );
OAI211xp5_ASAP7_75t_L g1383 ( .A1(n_1384), .A2(n_1385), .B(n_1386), .C(n_1387), .Y(n_1383) );
NAND2xp5_ASAP7_75t_L g1393 ( .A(n_1394), .B(n_1395), .Y(n_1393) );
NAND3xp33_ASAP7_75t_L g1396 ( .A(n_1397), .B(n_1412), .C(n_1414), .Y(n_1396) );
NOR2xp33_ASAP7_75t_SL g1397 ( .A(n_1398), .B(n_1411), .Y(n_1397) );
OAI22xp5_ASAP7_75t_L g1399 ( .A1(n_1400), .A2(n_1401), .B1(n_1402), .B2(n_1403), .Y(n_1399) );
INVx2_ASAP7_75t_L g1415 ( .A(n_1416), .Y(n_1415) );
BUFx3_ASAP7_75t_L g1416 ( .A(n_1417), .Y(n_1416) );
INVxp33_ASAP7_75t_SL g1420 ( .A(n_1421), .Y(n_1420) );
INVx1_ASAP7_75t_L g1423 ( .A(n_1424), .Y(n_1423) );
BUFx2_ASAP7_75t_SL g1425 ( .A(n_1426), .Y(n_1425) );
BUFx3_ASAP7_75t_L g1426 ( .A(n_1427), .Y(n_1426) );
HB1xp67_ASAP7_75t_L g1428 ( .A(n_1429), .Y(n_1428) );
OAI21xp5_ASAP7_75t_L g1429 ( .A1(n_1430), .A2(n_1431), .B(n_1432), .Y(n_1429) );
INVx1_ASAP7_75t_L g1432 ( .A(n_1433), .Y(n_1432) );
endmodule