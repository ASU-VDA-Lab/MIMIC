module fake_jpeg_22898_n_348 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_348);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_348;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_12),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_16),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_12),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_15),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx2_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_6),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_10),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_27),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_37),
.B(n_46),
.Y(n_55)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g39 ( 
.A1(n_26),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_39),
.A2(n_26),
.B1(n_33),
.B2(n_20),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

CKINVDCx14_ASAP7_75t_R g65 ( 
.A(n_44),
.Y(n_65)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_19),
.Y(n_46)
);

BUFx16f_ASAP7_75t_L g47 ( 
.A(n_19),
.Y(n_47)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_26),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_48),
.A2(n_22),
.B1(n_23),
.B2(n_20),
.Y(n_72)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_49),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_23),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_50),
.Y(n_66)
);

A2O1A1Ixp33_ASAP7_75t_L g51 ( 
.A1(n_37),
.A2(n_24),
.B(n_23),
.C(n_34),
.Y(n_51)
);

A2O1A1Ixp33_ASAP7_75t_L g102 ( 
.A1(n_51),
.A2(n_53),
.B(n_69),
.C(n_34),
.Y(n_102)
);

A2O1A1Ixp33_ASAP7_75t_L g53 ( 
.A1(n_37),
.A2(n_24),
.B(n_23),
.C(n_34),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_54),
.A2(n_42),
.B1(n_49),
.B2(n_21),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_33),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_56),
.B(n_67),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_48),
.A2(n_26),
.B1(n_22),
.B2(n_24),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_57),
.A2(n_46),
.B1(n_45),
.B2(n_43),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_40),
.B(n_23),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_59),
.B(n_61),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_42),
.B(n_29),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_41),
.B(n_33),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_41),
.A2(n_22),
.B1(n_30),
.B2(n_25),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_38),
.B(n_20),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_70),
.B(n_22),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_72),
.A2(n_38),
.B1(n_23),
.B2(n_40),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_71),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_74),
.B(n_77),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_71),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_76),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_71),
.Y(n_78)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_78),
.Y(n_132)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_67),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_79),
.B(n_85),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_61),
.B(n_40),
.C(n_50),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_80),
.B(n_44),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_56),
.A2(n_48),
.B1(n_49),
.B2(n_42),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_81),
.A2(n_91),
.B1(n_99),
.B2(n_58),
.Y(n_111)
);

OAI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_82),
.A2(n_90),
.B1(n_102),
.B2(n_104),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_55),
.B(n_49),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_83),
.B(n_84),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_55),
.B(n_61),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_70),
.Y(n_85)
);

CKINVDCx5p33_ASAP7_75t_R g86 ( 
.A(n_71),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_86),
.B(n_87),
.Y(n_136)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_69),
.Y(n_87)
);

HB1xp67_ASAP7_75t_L g88 ( 
.A(n_58),
.Y(n_88)
);

INVx1_ASAP7_75t_SL g134 ( 
.A(n_88),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_69),
.B(n_17),
.Y(n_89)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_89),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_51),
.A2(n_46),
.B1(n_45),
.B2(n_43),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_52),
.Y(n_92)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_92),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_71),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_93),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_66),
.B(n_21),
.Y(n_94)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_94),
.Y(n_110)
);

AND2x4_ASAP7_75t_L g95 ( 
.A(n_59),
.B(n_40),
.Y(n_95)
);

NOR2x1_ASAP7_75t_R g117 ( 
.A(n_95),
.B(n_101),
.Y(n_117)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_52),
.Y(n_96)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_96),
.Y(n_109)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_52),
.Y(n_97)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_97),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_71),
.Y(n_98)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_98),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_64),
.B(n_40),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_100),
.B(n_62),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_59),
.B(n_50),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_66),
.B(n_17),
.Y(n_103)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_103),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_66),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_63),
.Y(n_105)
);

OAI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_105),
.A2(n_106),
.B1(n_60),
.B2(n_44),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_58),
.A2(n_17),
.B1(n_21),
.B2(n_25),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_111),
.A2(n_114),
.B1(n_128),
.B2(n_65),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_87),
.A2(n_54),
.B1(n_59),
.B2(n_52),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_102),
.A2(n_53),
.B1(n_51),
.B2(n_57),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_119),
.A2(n_121),
.B1(n_129),
.B2(n_135),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_120),
.B(n_100),
.C(n_101),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_89),
.A2(n_53),
.B1(n_72),
.B2(n_68),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_84),
.A2(n_64),
.B(n_31),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_124),
.A2(n_127),
.B(n_130),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_126),
.B(n_81),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_95),
.B(n_50),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_91),
.A2(n_62),
.B1(n_68),
.B2(n_60),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_95),
.A2(n_68),
.B1(n_60),
.B2(n_62),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_73),
.A2(n_64),
.B(n_35),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_131),
.A2(n_78),
.B1(n_18),
.B2(n_30),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_95),
.A2(n_75),
.B1(n_73),
.B2(n_80),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_135),
.B(n_95),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_137),
.B(n_120),
.Y(n_185)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_133),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_138),
.B(n_140),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_124),
.B(n_83),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_139),
.B(n_142),
.Y(n_175)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_133),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_141),
.B(n_117),
.C(n_127),
.Y(n_173)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_125),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_143),
.B(n_150),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_125),
.B(n_75),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_144),
.B(n_164),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_136),
.A2(n_101),
.B(n_75),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_146),
.A2(n_161),
.B(n_118),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_119),
.A2(n_99),
.B1(n_85),
.B2(n_79),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_147),
.A2(n_149),
.B1(n_153),
.B2(n_157),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_110),
.B(n_104),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_148),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_121),
.A2(n_77),
.B1(n_97),
.B2(n_96),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_136),
.Y(n_150)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_132),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_151),
.B(n_158),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_110),
.B(n_103),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_152),
.B(n_155),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_129),
.A2(n_92),
.B1(n_65),
.B2(n_44),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_122),
.B(n_94),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_156),
.A2(n_159),
.B1(n_165),
.B2(n_134),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_123),
.A2(n_63),
.B1(n_105),
.B2(n_25),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_126),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_114),
.A2(n_63),
.B1(n_105),
.B2(n_36),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_122),
.B(n_30),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_160),
.B(n_18),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_117),
.A2(n_78),
.B(n_86),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_L g183 ( 
.A1(n_162),
.A2(n_127),
.B1(n_134),
.B2(n_115),
.Y(n_183)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_112),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_163),
.B(n_167),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_120),
.B(n_47),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_108),
.A2(n_18),
.B1(n_31),
.B2(n_28),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_120),
.B(n_47),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_166),
.B(n_47),
.Y(n_200)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_112),
.Y(n_167)
);

XOR2x2_ASAP7_75t_SL g171 ( 
.A(n_154),
.B(n_117),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_171),
.B(n_165),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_148),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_172),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_173),
.B(n_196),
.C(n_150),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_174),
.B(n_190),
.Y(n_223)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_152),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_176),
.B(n_178),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_161),
.A2(n_108),
.B(n_130),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_177),
.A2(n_154),
.B(n_139),
.Y(n_211)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_155),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_180),
.B(n_192),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_164),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_181),
.B(n_184),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_183),
.A2(n_98),
.B1(n_76),
.B2(n_34),
.Y(n_231)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_153),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_185),
.B(n_186),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_137),
.B(n_127),
.Y(n_186)
);

OAI32xp33_ASAP7_75t_L g188 ( 
.A1(n_144),
.A2(n_156),
.A3(n_145),
.B1(n_143),
.B2(n_159),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_188),
.B(n_29),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_141),
.B(n_111),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_189),
.B(n_32),
.Y(n_224)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_149),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_147),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_191),
.B(n_194),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_138),
.B(n_132),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_142),
.A2(n_128),
.B1(n_134),
.B2(n_118),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_193),
.A2(n_199),
.B1(n_157),
.B2(n_163),
.Y(n_205)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_142),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_195),
.A2(n_200),
.B(n_146),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_145),
.B(n_47),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_160),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_197),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_166),
.A2(n_109),
.B1(n_107),
.B2(n_113),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_202),
.A2(n_231),
.B1(n_168),
.B2(n_178),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_204),
.B(n_208),
.C(n_212),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_205),
.A2(n_216),
.B1(n_219),
.B2(n_221),
.Y(n_251)
);

AOI21x1_ASAP7_75t_SL g207 ( 
.A1(n_171),
.A2(n_195),
.B(n_177),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_207),
.B(n_217),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_173),
.B(n_187),
.C(n_194),
.Y(n_208)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_182),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_210),
.B(n_220),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_211),
.B(n_188),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_187),
.B(n_158),
.C(n_167),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_SL g256 ( 
.A(n_213),
.B(n_205),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_191),
.A2(n_140),
.B1(n_109),
.B2(n_107),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_199),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_190),
.A2(n_151),
.B1(n_116),
.B2(n_115),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_218),
.A2(n_230),
.B1(n_193),
.B2(n_184),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_175),
.A2(n_116),
.B1(n_27),
.B2(n_36),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_169),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_175),
.A2(n_27),
.B1(n_28),
.B2(n_36),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_201),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_222),
.B(n_220),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_224),
.B(n_225),
.C(n_227),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_196),
.B(n_185),
.C(n_186),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_200),
.B(n_98),
.C(n_76),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_198),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_228),
.Y(n_232)
);

OR2x2_ASAP7_75t_L g233 ( 
.A(n_214),
.B(n_197),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_233),
.B(n_236),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_234),
.B(n_255),
.Y(n_264)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_218),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_237),
.B(n_247),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_214),
.B(n_215),
.Y(n_238)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_238),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_230),
.A2(n_174),
.B1(n_181),
.B2(n_170),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_239),
.A2(n_240),
.B1(n_245),
.B2(n_221),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_210),
.Y(n_242)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_242),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_217),
.A2(n_176),
.B1(n_179),
.B2(n_170),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_243),
.A2(n_249),
.B1(n_15),
.B2(n_14),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_209),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_244),
.B(n_222),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_229),
.A2(n_189),
.B1(n_35),
.B2(n_31),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_216),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_246),
.B(n_250),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_203),
.B(n_32),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_223),
.A2(n_231),
.B1(n_226),
.B2(n_228),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_212),
.Y(n_250)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_252),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_203),
.B(n_32),
.C(n_35),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_253),
.B(n_225),
.C(n_224),
.Y(n_262)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_227),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_SL g276 ( 
.A(n_256),
.B(n_1),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_219),
.B(n_0),
.Y(n_257)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_257),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_258),
.B(n_251),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_259),
.B(n_267),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_246),
.A2(n_208),
.B1(n_204),
.B2(n_207),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_260),
.A2(n_269),
.B1(n_271),
.B2(n_254),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_262),
.B(n_270),
.C(n_241),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_252),
.B(n_206),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_263),
.B(n_272),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_232),
.B(n_213),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_239),
.A2(n_202),
.B1(n_211),
.B2(n_28),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_241),
.B(n_32),
.C(n_2),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_234),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_232),
.B(n_16),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_256),
.B(n_16),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_275),
.B(n_276),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_277),
.B(n_278),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_248),
.B(n_15),
.Y(n_278)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_280),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_266),
.A2(n_236),
.B(n_255),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_282),
.B(n_264),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_268),
.A2(n_265),
.B(n_261),
.Y(n_283)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_283),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_284),
.B(n_294),
.C(n_270),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_286),
.B(n_295),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_262),
.B(n_235),
.C(n_250),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_288),
.B(n_292),
.C(n_284),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_271),
.B(n_251),
.Y(n_290)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_290),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_266),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_291),
.B(n_297),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_261),
.B(n_235),
.C(n_247),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_279),
.B(n_237),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_293),
.B(n_296),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_268),
.A2(n_248),
.B(n_233),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_258),
.B(n_245),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_260),
.B(n_253),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_274),
.B(n_242),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_298),
.A2(n_299),
.B(n_303),
.Y(n_323)
);

A2O1A1Ixp33_ASAP7_75t_L g303 ( 
.A1(n_294),
.A2(n_269),
.B(n_257),
.C(n_276),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_304),
.B(n_307),
.C(n_312),
.Y(n_317)
);

HB1xp67_ASAP7_75t_L g305 ( 
.A(n_282),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_305),
.B(n_287),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_293),
.B(n_279),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_306),
.B(n_309),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_288),
.B(n_273),
.C(n_274),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_SL g309 ( 
.A(n_280),
.B(n_275),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_292),
.B(n_13),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_L g329 ( 
.A1(n_313),
.A2(n_315),
.B(n_316),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_311),
.B(n_285),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_314),
.B(n_321),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_L g315 ( 
.A1(n_300),
.A2(n_289),
.B(n_296),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_301),
.A2(n_281),
.B(n_14),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_303),
.A2(n_281),
.B1(n_2),
.B2(n_3),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_318),
.B(n_320),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_L g319 ( 
.A1(n_310),
.A2(n_1),
.B(n_3),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_SL g327 ( 
.A1(n_319),
.A2(n_4),
.B(n_5),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_308),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_312),
.B(n_14),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_302),
.B(n_13),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_322),
.B(n_309),
.C(n_304),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_325),
.B(n_317),
.C(n_324),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_327),
.Y(n_336)
);

NAND2xp33_ASAP7_75t_L g330 ( 
.A(n_318),
.B(n_302),
.Y(n_330)
);

A2O1A1Ixp33_ASAP7_75t_SL g337 ( 
.A1(n_330),
.A2(n_324),
.B(n_320),
.C(n_8),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_319),
.B(n_306),
.Y(n_331)
);

AOI21xp5_ASAP7_75t_L g340 ( 
.A1(n_331),
.A2(n_6),
.B(n_8),
.Y(n_340)
);

AOI31xp33_ASAP7_75t_L g332 ( 
.A1(n_322),
.A2(n_13),
.A3(n_11),
.B(n_7),
.Y(n_332)
);

AOI21xp33_ASAP7_75t_L g339 ( 
.A1(n_332),
.A2(n_5),
.B(n_6),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_SL g333 ( 
.A(n_323),
.B(n_11),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_333),
.B(n_328),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_SL g334 ( 
.A1(n_329),
.A2(n_317),
.B(n_315),
.Y(n_334)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_334),
.Y(n_341)
);

OAI21xp5_ASAP7_75t_L g343 ( 
.A1(n_335),
.A2(n_338),
.B(n_339),
.Y(n_343)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_337),
.Y(n_342)
);

AOI21xp5_ASAP7_75t_L g344 ( 
.A1(n_341),
.A2(n_343),
.B(n_331),
.Y(n_344)
);

OAI321xp33_ASAP7_75t_L g345 ( 
.A1(n_344),
.A2(n_340),
.A3(n_337),
.B1(n_342),
.B2(n_336),
.C(n_326),
.Y(n_345)
);

OAI21x1_ASAP7_75t_SL g346 ( 
.A1(n_345),
.A2(n_9),
.B(n_10),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_L g347 ( 
.A1(n_346),
.A2(n_9),
.B(n_10),
.Y(n_347)
);

OAI21xp5_ASAP7_75t_SL g348 ( 
.A1(n_347),
.A2(n_9),
.B(n_10),
.Y(n_348)
);


endmodule