module fake_netlist_6_3909_n_451 (n_41, n_52, n_16, n_45, n_1, n_46, n_34, n_42, n_9, n_8, n_70, n_18, n_10, n_21, n_24, n_71, n_37, n_6, n_15, n_33, n_54, n_67, n_27, n_3, n_14, n_38, n_72, n_0, n_61, n_39, n_63, n_60, n_59, n_32, n_4, n_66, n_36, n_22, n_26, n_68, n_55, n_13, n_35, n_11, n_28, n_17, n_23, n_58, n_12, n_69, n_20, n_50, n_49, n_7, n_30, n_64, n_2, n_43, n_5, n_19, n_47, n_48, n_29, n_62, n_31, n_65, n_25, n_40, n_57, n_53, n_51, n_44, n_56, n_451);

input n_41;
input n_52;
input n_16;
input n_45;
input n_1;
input n_46;
input n_34;
input n_42;
input n_9;
input n_8;
input n_70;
input n_18;
input n_10;
input n_21;
input n_24;
input n_71;
input n_37;
input n_6;
input n_15;
input n_33;
input n_54;
input n_67;
input n_27;
input n_3;
input n_14;
input n_38;
input n_72;
input n_0;
input n_61;
input n_39;
input n_63;
input n_60;
input n_59;
input n_32;
input n_4;
input n_66;
input n_36;
input n_22;
input n_26;
input n_68;
input n_55;
input n_13;
input n_35;
input n_11;
input n_28;
input n_17;
input n_23;
input n_58;
input n_12;
input n_69;
input n_20;
input n_50;
input n_49;
input n_7;
input n_30;
input n_64;
input n_2;
input n_43;
input n_5;
input n_19;
input n_47;
input n_48;
input n_29;
input n_62;
input n_31;
input n_65;
input n_25;
input n_40;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_451;

wire n_435;
wire n_91;
wire n_326;
wire n_256;
wire n_440;
wire n_209;
wire n_367;
wire n_223;
wire n_278;
wire n_362;
wire n_341;
wire n_148;
wire n_226;
wire n_161;
wire n_208;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_144;
wire n_365;
wire n_125;
wire n_168;
wire n_384;
wire n_297;
wire n_342;
wire n_77;
wire n_106;
wire n_358;
wire n_160;
wire n_449;
wire n_131;
wire n_188;
wire n_310;
wire n_186;
wire n_245;
wire n_368;
wire n_396;
wire n_350;
wire n_78;
wire n_84;
wire n_392;
wire n_442;
wire n_142;
wire n_143;
wire n_382;
wire n_180;
wire n_349;
wire n_233;
wire n_255;
wire n_284;
wire n_400;
wire n_140;
wire n_337;
wire n_214;
wire n_443;
wire n_246;
wire n_289;
wire n_421;
wire n_424;
wire n_181;
wire n_182;
wire n_238;
wire n_202;
wire n_320;
wire n_108;
wire n_327;
wire n_369;
wire n_280;
wire n_287;
wire n_353;
wire n_389;
wire n_415;
wire n_230;
wire n_141;
wire n_383;
wire n_200;
wire n_447;
wire n_176;
wire n_114;
wire n_86;
wire n_198;
wire n_104;
wire n_222;
wire n_179;
wire n_248;
wire n_300;
wire n_74;
wire n_229;
wire n_305;
wire n_173;
wire n_250;
wire n_372;
wire n_111;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_183;
wire n_79;
wire n_375;
wire n_338;
wire n_360;
wire n_119;
wire n_235;
wire n_147;
wire n_191;
wire n_340;
wire n_387;
wire n_344;
wire n_73;
wire n_428;
wire n_432;
wire n_101;
wire n_167;
wire n_174;
wire n_127;
wire n_153;
wire n_156;
wire n_145;
wire n_133;
wire n_96;
wire n_371;
wire n_189;
wire n_405;
wire n_213;
wire n_294;
wire n_302;
wire n_380;
wire n_129;
wire n_197;
wire n_137;
wire n_343;
wire n_448;
wire n_397;
wire n_155;
wire n_109;
wire n_445;
wire n_425;
wire n_122;
wire n_218;
wire n_234;
wire n_381;
wire n_82;
wire n_236;
wire n_112;
wire n_172;
wire n_270;
wire n_239;
wire n_126;
wire n_414;
wire n_97;
wire n_290;
wire n_220;
wire n_118;
wire n_224;
wire n_93;
wire n_80;
wire n_196;
wire n_402;
wire n_352;
wire n_107;
wire n_417;
wire n_446;
wire n_89;
wire n_374;
wire n_366;
wire n_407;
wire n_450;
wire n_103;
wire n_272;
wire n_185;
wire n_348;
wire n_376;
wire n_390;
wire n_293;
wire n_334;
wire n_370;
wire n_232;
wire n_163;
wire n_330;
wire n_298;
wire n_281;
wire n_258;
wire n_154;
wire n_98;
wire n_260;
wire n_265;
wire n_313;
wire n_279;
wire n_252;
wire n_228;
wire n_356;
wire n_166;
wire n_184;
wire n_216;
wire n_83;
wire n_363;
wire n_395;
wire n_323;
wire n_393;
wire n_411;
wire n_152;
wire n_92;
wire n_321;
wire n_331;
wire n_105;
wire n_227;
wire n_132;
wire n_406;
wire n_102;
wire n_204;
wire n_261;
wire n_420;
wire n_312;
wire n_394;
wire n_130;
wire n_164;
wire n_292;
wire n_100;
wire n_121;
wire n_307;
wire n_433;
wire n_291;
wire n_219;
wire n_357;
wire n_150;
wire n_264;
wire n_263;
wire n_325;
wire n_329;
wire n_408;
wire n_237;
wire n_244;
wire n_399;
wire n_76;
wire n_243;
wire n_124;
wire n_94;
wire n_282;
wire n_436;
wire n_116;
wire n_211;
wire n_117;
wire n_175;
wire n_322;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_240;
wire n_139;
wire n_319;
wire n_134;
wire n_273;
wire n_95;
wire n_311;
wire n_403;
wire n_253;
wire n_123;
wire n_136;
wire n_249;
wire n_201;
wire n_386;
wire n_159;
wire n_157;
wire n_162;
wire n_115;
wire n_128;
wire n_241;
wire n_275;
wire n_276;
wire n_441;
wire n_221;
wire n_444;
wire n_423;
wire n_146;
wire n_318;
wire n_303;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_346;
wire n_88;
wire n_416;
wire n_277;
wire n_418;
wire n_113;
wire n_199;
wire n_138;
wire n_266;
wire n_296;
wire n_268;
wire n_271;
wire n_404;
wire n_439;
wire n_158;
wire n_217;
wire n_210;
wire n_299;
wire n_206;
wire n_333;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_355;
wire n_426;
wire n_317;
wire n_149;
wire n_431;
wire n_90;
wire n_347;
wire n_328;
wire n_429;
wire n_373;
wire n_87;
wire n_195;
wire n_285;
wire n_257;
wire n_99;
wire n_85;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_242;
wire n_75;
wire n_401;
wire n_324;
wire n_335;
wire n_430;
wire n_205;
wire n_120;
wire n_251;
wire n_301;
wire n_274;
wire n_110;
wire n_151;
wire n_412;
wire n_81;
wire n_267;
wire n_438;
wire n_339;
wire n_315;
wire n_434;
wire n_288;
wire n_427;
wire n_422;
wire n_135;
wire n_165;
wire n_351;
wire n_437;
wire n_259;
wire n_177;
wire n_391;
wire n_364;
wire n_295;
wire n_385;
wire n_388;
wire n_190;
wire n_262;
wire n_187;
wire n_361;
wire n_379;
wire n_170;
wire n_332;
wire n_336;
wire n_398;
wire n_410;
wire n_194;
wire n_171;
wire n_192;
wire n_169;
wire n_283;

INVx1_ASAP7_75t_L g73 ( 
.A(n_3),
.Y(n_73)
);

INVxp33_ASAP7_75t_SL g74 ( 
.A(n_25),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_48),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_70),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_33),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_19),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_68),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_13),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_56),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_50),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_46),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_8),
.Y(n_84)
);

INVxp67_ASAP7_75t_SL g85 ( 
.A(n_45),
.Y(n_85)
);

OR2x2_ASAP7_75t_L g86 ( 
.A(n_40),
.B(n_67),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_54),
.Y(n_87)
);

INVxp67_ASAP7_75t_SL g88 ( 
.A(n_36),
.Y(n_88)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_72),
.Y(n_89)
);

INVxp67_ASAP7_75t_SL g90 ( 
.A(n_10),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_24),
.Y(n_91)
);

BUFx2_ASAP7_75t_L g92 ( 
.A(n_23),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_9),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_21),
.Y(n_94)
);

CKINVDCx14_ASAP7_75t_R g95 ( 
.A(n_44),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_5),
.Y(n_96)
);

CKINVDCx5p33_ASAP7_75t_R g97 ( 
.A(n_47),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_37),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_34),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_5),
.B(n_69),
.Y(n_100)
);

INVxp67_ASAP7_75t_SL g101 ( 
.A(n_51),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_15),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_11),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_63),
.Y(n_104)
);

INVxp33_ASAP7_75t_SL g105 ( 
.A(n_7),
.Y(n_105)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_35),
.Y(n_106)
);

CKINVDCx5p33_ASAP7_75t_R g107 ( 
.A(n_16),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_66),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_7),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_32),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_38),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_57),
.Y(n_112)
);

INVxp33_ASAP7_75t_SL g113 ( 
.A(n_52),
.Y(n_113)
);

INVxp33_ASAP7_75t_L g114 ( 
.A(n_18),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_28),
.Y(n_115)
);

INVxp67_ASAP7_75t_SL g116 ( 
.A(n_61),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_58),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_1),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_43),
.Y(n_119)
);

INVxp33_ASAP7_75t_SL g120 ( 
.A(n_60),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_55),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_65),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_27),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_0),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_20),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_64),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_62),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_22),
.Y(n_128)
);

CKINVDCx5p33_ASAP7_75t_R g129 ( 
.A(n_30),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_12),
.Y(n_130)
);

INVxp33_ASAP7_75t_SL g131 ( 
.A(n_29),
.Y(n_131)
);

INVxp33_ASAP7_75t_L g132 ( 
.A(n_0),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_17),
.Y(n_133)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_71),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_31),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_26),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_2),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_1),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_53),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_73),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_118),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_124),
.Y(n_142)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_139),
.Y(n_143)
);

OA21x2_ASAP7_75t_L g144 ( 
.A1(n_137),
.A2(n_2),
.B(n_3),
.Y(n_144)
);

AND2x4_ASAP7_75t_L g145 ( 
.A(n_92),
.B(n_41),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_75),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_76),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_98),
.B(n_4),
.Y(n_148)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_139),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_77),
.Y(n_150)
);

HB1xp67_ASAP7_75t_L g151 ( 
.A(n_96),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_78),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_95),
.A2(n_4),
.B1(n_6),
.B2(n_14),
.Y(n_153)
);

INVx1_ASAP7_75t_SL g154 ( 
.A(n_138),
.Y(n_154)
);

AND2x4_ASAP7_75t_L g155 ( 
.A(n_106),
.B(n_39),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_80),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_81),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_89),
.B(n_6),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_82),
.Y(n_159)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_139),
.Y(n_160)
);

AND2x6_ASAP7_75t_L g161 ( 
.A(n_134),
.B(n_108),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_83),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_84),
.Y(n_163)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_87),
.Y(n_164)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_91),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_93),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_99),
.Y(n_167)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_102),
.Y(n_168)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_103),
.Y(n_169)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_110),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_112),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_94),
.B(n_42),
.Y(n_172)
);

HB1xp67_ASAP7_75t_L g173 ( 
.A(n_96),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_115),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_104),
.B(n_49),
.Y(n_175)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_117),
.Y(n_176)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_122),
.Y(n_177)
);

HB1xp67_ASAP7_75t_L g178 ( 
.A(n_109),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_123),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_132),
.B(n_59),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_114),
.B(n_109),
.Y(n_181)
);

BUFx3_ASAP7_75t_L g182 ( 
.A(n_126),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_127),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_105),
.B(n_100),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_128),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_130),
.Y(n_186)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_133),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_135),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_94),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_85),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_85),
.Y(n_191)
);

OA21x2_ASAP7_75t_L g192 ( 
.A1(n_88),
.A2(n_90),
.B(n_101),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_88),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_90),
.B(n_101),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_97),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_107),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_129),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_86),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_116),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_79),
.B(n_111),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_74),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_113),
.Y(n_202)
);

AND2x4_ASAP7_75t_L g203 ( 
.A(n_119),
.B(n_121),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_195),
.B(n_120),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_198),
.B(n_131),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_195),
.B(n_125),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_143),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_164),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_198),
.B(n_136),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_190),
.B(n_194),
.Y(n_210)
);

BUFx3_ASAP7_75t_L g211 ( 
.A(n_182),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_196),
.B(n_197),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_181),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_143),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_201),
.B(n_202),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_164),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_191),
.B(n_193),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_199),
.B(n_155),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_168),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_199),
.B(n_189),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_155),
.B(n_145),
.Y(n_221)
);

OR2x2_ASAP7_75t_L g222 ( 
.A(n_151),
.B(n_178),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_149),
.Y(n_223)
);

INVx2_ASAP7_75t_SL g224 ( 
.A(n_151),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_168),
.Y(n_225)
);

OAI221xp5_ASAP7_75t_L g226 ( 
.A1(n_173),
.A2(n_178),
.B1(n_158),
.B2(n_142),
.C(n_140),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_169),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_180),
.B(n_175),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_145),
.B(n_175),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_145),
.B(n_158),
.Y(n_230)
);

NAND3xp33_ASAP7_75t_SL g231 ( 
.A(n_153),
.B(n_184),
.C(n_154),
.Y(n_231)
);

OR2x2_ASAP7_75t_L g232 ( 
.A(n_173),
.B(n_182),
.Y(n_232)
);

OR2x2_ASAP7_75t_SL g233 ( 
.A(n_144),
.B(n_148),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_155),
.B(n_160),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_149),
.B(n_160),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_149),
.B(n_160),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_L g237 ( 
.A1(n_192),
.A2(n_144),
.B1(n_141),
.B2(n_184),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_167),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_172),
.B(n_166),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_146),
.B(n_171),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_176),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_147),
.B(n_163),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_150),
.B(n_174),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_200),
.Y(n_244)
);

INVx8_ASAP7_75t_L g245 ( 
.A(n_203),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_179),
.Y(n_246)
);

NAND2xp33_ASAP7_75t_L g247 ( 
.A(n_161),
.B(n_167),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_203),
.B(n_167),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_152),
.B(n_188),
.Y(n_249)
);

OR2x2_ASAP7_75t_L g250 ( 
.A(n_156),
.B(n_185),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_L g251 ( 
.A1(n_192),
.A2(n_144),
.B1(n_157),
.B2(n_159),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_203),
.B(n_186),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_162),
.B(n_183),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_228),
.B(n_187),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_250),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_235),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_221),
.B(n_192),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_228),
.B(n_165),
.Y(n_258)
);

AND2x4_ASAP7_75t_L g259 ( 
.A(n_211),
.B(n_177),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_207),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_251),
.B(n_165),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_214),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_236),
.Y(n_263)
);

AND2x4_ASAP7_75t_L g264 ( 
.A(n_248),
.B(n_170),
.Y(n_264)
);

INVx3_ASAP7_75t_L g265 ( 
.A(n_223),
.Y(n_265)
);

BUFx12f_ASAP7_75t_L g266 ( 
.A(n_244),
.Y(n_266)
);

AND2x4_ASAP7_75t_L g267 ( 
.A(n_220),
.B(n_165),
.Y(n_267)
);

BUFx12f_ASAP7_75t_L g268 ( 
.A(n_232),
.Y(n_268)
);

OAI21xp33_ASAP7_75t_L g269 ( 
.A1(n_229),
.A2(n_161),
.B(n_230),
.Y(n_269)
);

BUFx8_ASAP7_75t_L g270 ( 
.A(n_224),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_208),
.Y(n_271)
);

BUFx3_ASAP7_75t_L g272 ( 
.A(n_242),
.Y(n_272)
);

INVx3_ASAP7_75t_L g273 ( 
.A(n_216),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_213),
.B(n_161),
.Y(n_274)
);

BUFx2_ASAP7_75t_L g275 ( 
.A(n_222),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_206),
.B(n_161),
.Y(n_276)
);

OR2x6_ASAP7_75t_L g277 ( 
.A(n_245),
.B(n_209),
.Y(n_277)
);

BUFx4f_ASAP7_75t_L g278 ( 
.A(n_245),
.Y(n_278)
);

INVx5_ASAP7_75t_L g279 ( 
.A(n_245),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_R g280 ( 
.A(n_231),
.B(n_215),
.Y(n_280)
);

BUFx3_ASAP7_75t_L g281 ( 
.A(n_243),
.Y(n_281)
);

AND2x2_ASAP7_75t_L g282 ( 
.A(n_210),
.B(n_239),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_226),
.A2(n_237),
.B1(n_205),
.B2(n_218),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_219),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_225),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_251),
.B(n_239),
.Y(n_286)
);

INVx3_ASAP7_75t_L g287 ( 
.A(n_227),
.Y(n_287)
);

HB1xp67_ASAP7_75t_L g288 ( 
.A(n_234),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_231),
.A2(n_237),
.B1(n_252),
.B2(n_217),
.Y(n_289)
);

AND2x4_ASAP7_75t_L g290 ( 
.A(n_217),
.B(n_212),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_241),
.B(n_246),
.Y(n_291)
);

AO21x1_ASAP7_75t_L g292 ( 
.A1(n_204),
.A2(n_233),
.B(n_247),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_249),
.Y(n_293)
);

AND2x2_ASAP7_75t_L g294 ( 
.A(n_240),
.B(n_253),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_240),
.Y(n_295)
);

AND2x4_ASAP7_75t_L g296 ( 
.A(n_211),
.B(n_248),
.Y(n_296)
);

BUFx6f_ASAP7_75t_L g297 ( 
.A(n_211),
.Y(n_297)
);

INVx3_ASAP7_75t_L g298 ( 
.A(n_238),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_284),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_273),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_286),
.B(n_282),
.Y(n_301)
);

AND2x2_ASAP7_75t_L g302 ( 
.A(n_294),
.B(n_290),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_289),
.A2(n_286),
.B1(n_283),
.B2(n_269),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_258),
.B(n_288),
.Y(n_304)
);

BUFx4f_ASAP7_75t_SL g305 ( 
.A(n_266),
.Y(n_305)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_273),
.Y(n_306)
);

HB1xp67_ASAP7_75t_L g307 ( 
.A(n_275),
.Y(n_307)
);

AND2x4_ASAP7_75t_L g308 ( 
.A(n_259),
.B(n_267),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_287),
.Y(n_309)
);

OR2x2_ASAP7_75t_L g310 ( 
.A(n_255),
.B(n_290),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_272),
.B(n_281),
.Y(n_311)
);

AND2x2_ASAP7_75t_L g312 ( 
.A(n_288),
.B(n_293),
.Y(n_312)
);

BUFx4f_ASAP7_75t_SL g313 ( 
.A(n_268),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_L g314 ( 
.A1(n_289),
.A2(n_283),
.B1(n_258),
.B2(n_295),
.Y(n_314)
);

INVx5_ASAP7_75t_L g315 ( 
.A(n_277),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_291),
.Y(n_316)
);

NAND2xp33_ASAP7_75t_L g317 ( 
.A(n_280),
.B(n_256),
.Y(n_317)
);

AND2x4_ASAP7_75t_L g318 ( 
.A(n_259),
.B(n_296),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_263),
.B(n_264),
.Y(n_319)
);

BUFx2_ASAP7_75t_L g320 ( 
.A(n_270),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_264),
.A2(n_254),
.B1(n_274),
.B2(n_296),
.Y(n_321)
);

OR2x2_ASAP7_75t_L g322 ( 
.A(n_297),
.B(n_291),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_271),
.Y(n_323)
);

AND2x2_ASAP7_75t_L g324 ( 
.A(n_297),
.B(n_277),
.Y(n_324)
);

AO22x2_ASAP7_75t_L g325 ( 
.A1(n_276),
.A2(n_277),
.B1(n_292),
.B2(n_285),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_260),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_262),
.Y(n_327)
);

HB1xp67_ASAP7_75t_L g328 ( 
.A(n_297),
.Y(n_328)
);

BUFx6f_ASAP7_75t_L g329 ( 
.A(n_298),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_265),
.Y(n_330)
);

AOI21xp5_ASAP7_75t_L g331 ( 
.A1(n_278),
.A2(n_279),
.B(n_270),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_279),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_279),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_278),
.B(n_228),
.Y(n_334)
);

BUFx10_ASAP7_75t_L g335 ( 
.A(n_259),
.Y(n_335)
);

HB1xp67_ASAP7_75t_L g336 ( 
.A(n_275),
.Y(n_336)
);

AND2x4_ASAP7_75t_L g337 ( 
.A(n_259),
.B(n_267),
.Y(n_337)
);

BUFx2_ASAP7_75t_L g338 ( 
.A(n_268),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_272),
.B(n_281),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_289),
.A2(n_228),
.B1(n_229),
.B2(n_283),
.Y(n_340)
);

OR2x6_ASAP7_75t_L g341 ( 
.A(n_268),
.B(n_245),
.Y(n_341)
);

AOI222xp33_ASAP7_75t_L g342 ( 
.A1(n_282),
.A2(n_184),
.B1(n_231),
.B2(n_226),
.C1(n_190),
.C2(n_158),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_266),
.Y(n_343)
);

AOI21xp5_ASAP7_75t_L g344 ( 
.A1(n_257),
.A2(n_261),
.B(n_221),
.Y(n_344)
);

AOI21xp5_ASAP7_75t_L g345 ( 
.A1(n_257),
.A2(n_261),
.B(n_221),
.Y(n_345)
);

AND2x4_ASAP7_75t_L g346 ( 
.A(n_259),
.B(n_267),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_L g347 ( 
.A1(n_257),
.A2(n_286),
.B(n_261),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_323),
.Y(n_348)
);

OA21x2_ASAP7_75t_L g349 ( 
.A1(n_347),
.A2(n_344),
.B(n_345),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_300),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_323),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_302),
.B(n_301),
.Y(n_352)
);

AO21x2_ASAP7_75t_L g353 ( 
.A1(n_340),
.A2(n_314),
.B(n_303),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_306),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_326),
.Y(n_355)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_309),
.Y(n_356)
);

INVx2_ASAP7_75t_SL g357 ( 
.A(n_322),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_327),
.Y(n_358)
);

AOI221xp5_ASAP7_75t_L g359 ( 
.A1(n_312),
.A2(n_311),
.B1(n_339),
.B2(n_304),
.C(n_310),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_299),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_305),
.Y(n_361)
);

INVx2_ASAP7_75t_SL g362 ( 
.A(n_307),
.Y(n_362)
);

OR2x2_ASAP7_75t_L g363 ( 
.A(n_336),
.B(n_319),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_343),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_316),
.B(n_334),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_330),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_308),
.Y(n_367)
);

AND2x2_ASAP7_75t_L g368 ( 
.A(n_342),
.B(n_318),
.Y(n_368)
);

AND2x4_ASAP7_75t_L g369 ( 
.A(n_308),
.B(n_346),
.Y(n_369)
);

OA21x2_ASAP7_75t_L g370 ( 
.A1(n_321),
.A2(n_332),
.B(n_333),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_337),
.Y(n_371)
);

AND2x2_ASAP7_75t_L g372 ( 
.A(n_318),
.B(n_346),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_337),
.Y(n_373)
);

CKINVDCx6p67_ASAP7_75t_R g374 ( 
.A(n_315),
.Y(n_374)
);

OAI21x1_ASAP7_75t_L g375 ( 
.A1(n_332),
.A2(n_324),
.B(n_331),
.Y(n_375)
);

NAND2x1p5_ASAP7_75t_L g376 ( 
.A(n_315),
.B(n_329),
.Y(n_376)
);

OR2x2_ASAP7_75t_L g377 ( 
.A(n_328),
.B(n_338),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_335),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_348),
.Y(n_379)
);

AND2x2_ASAP7_75t_L g380 ( 
.A(n_368),
.B(n_352),
.Y(n_380)
);

AND2x2_ASAP7_75t_L g381 ( 
.A(n_352),
.B(n_335),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_365),
.B(n_317),
.Y(n_382)
);

INVxp67_ASAP7_75t_L g383 ( 
.A(n_363),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_351),
.Y(n_384)
);

INVx2_ASAP7_75t_SL g385 ( 
.A(n_362),
.Y(n_385)
);

AND2x4_ASAP7_75t_L g386 ( 
.A(n_369),
.B(n_315),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_355),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_358),
.Y(n_388)
);

NOR2x1_ASAP7_75t_L g389 ( 
.A(n_365),
.B(n_341),
.Y(n_389)
);

INVx2_ASAP7_75t_SL g390 ( 
.A(n_377),
.Y(n_390)
);

OR2x2_ASAP7_75t_L g391 ( 
.A(n_357),
.B(n_341),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_350),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_350),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_354),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_354),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_357),
.B(n_313),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_356),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_379),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_384),
.Y(n_399)
);

AND2x2_ASAP7_75t_L g400 ( 
.A(n_380),
.B(n_353),
.Y(n_400)
);

AND2x2_ASAP7_75t_L g401 ( 
.A(n_381),
.B(n_353),
.Y(n_401)
);

OAI221xp5_ASAP7_75t_L g402 ( 
.A1(n_383),
.A2(n_359),
.B1(n_373),
.B2(n_371),
.C(n_367),
.Y(n_402)
);

HB1xp67_ASAP7_75t_L g403 ( 
.A(n_390),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_392),
.Y(n_404)
);

BUFx2_ASAP7_75t_L g405 ( 
.A(n_385),
.Y(n_405)
);

AND2x4_ASAP7_75t_L g406 ( 
.A(n_386),
.B(n_369),
.Y(n_406)
);

AOI22xp33_ASAP7_75t_L g407 ( 
.A1(n_382),
.A2(n_325),
.B1(n_349),
.B2(n_370),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_396),
.A2(n_372),
.B1(n_369),
.B2(n_361),
.Y(n_408)
);

INVx1_ASAP7_75t_SL g409 ( 
.A(n_385),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_393),
.Y(n_410)
);

INVxp67_ASAP7_75t_L g411 ( 
.A(n_383),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_394),
.Y(n_412)
);

INVx1_ASAP7_75t_SL g413 ( 
.A(n_391),
.Y(n_413)
);

AND2x2_ASAP7_75t_L g414 ( 
.A(n_395),
.B(n_397),
.Y(n_414)
);

OAI32xp33_ASAP7_75t_L g415 ( 
.A1(n_402),
.A2(n_388),
.A3(n_387),
.B1(n_396),
.B2(n_376),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_398),
.Y(n_416)
);

AND2x4_ASAP7_75t_L g417 ( 
.A(n_406),
.B(n_386),
.Y(n_417)
);

AOI22xp33_ASAP7_75t_L g418 ( 
.A1(n_400),
.A2(n_389),
.B1(n_349),
.B2(n_360),
.Y(n_418)
);

AND2x2_ASAP7_75t_L g419 ( 
.A(n_401),
.B(n_386),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_414),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_399),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_400),
.B(n_366),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_414),
.Y(n_423)
);

INVx2_ASAP7_75t_SL g424 ( 
.A(n_403),
.Y(n_424)
);

NAND3xp33_ASAP7_75t_L g425 ( 
.A(n_418),
.B(n_408),
.C(n_411),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_416),
.Y(n_426)
);

INVx3_ASAP7_75t_L g427 ( 
.A(n_417),
.Y(n_427)
);

AND2x2_ASAP7_75t_L g428 ( 
.A(n_419),
.B(n_401),
.Y(n_428)
);

NOR2x1_ASAP7_75t_L g429 ( 
.A(n_422),
.B(n_405),
.Y(n_429)
);

AND2x2_ASAP7_75t_L g430 ( 
.A(n_420),
.B(n_413),
.Y(n_430)
);

AND2x2_ASAP7_75t_L g431 ( 
.A(n_428),
.B(n_423),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_426),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_430),
.B(n_420),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_429),
.Y(n_434)
);

AND2x2_ASAP7_75t_L g435 ( 
.A(n_427),
.B(n_423),
.Y(n_435)
);

OR2x2_ASAP7_75t_L g436 ( 
.A(n_427),
.B(n_421),
.Y(n_436)
);

OAI211xp5_ASAP7_75t_L g437 ( 
.A1(n_434),
.A2(n_415),
.B(n_425),
.C(n_418),
.Y(n_437)
);

NOR3xp33_ASAP7_75t_L g438 ( 
.A(n_434),
.B(n_425),
.C(n_375),
.Y(n_438)
);

AOI21xp5_ASAP7_75t_L g439 ( 
.A1(n_436),
.A2(n_349),
.B(n_407),
.Y(n_439)
);

NOR3xp33_ASAP7_75t_L g440 ( 
.A(n_433),
.B(n_375),
.C(n_424),
.Y(n_440)
);

AND3x1_ASAP7_75t_L g441 ( 
.A(n_431),
.B(n_364),
.C(n_378),
.Y(n_441)
);

OAI211xp5_ASAP7_75t_L g442 ( 
.A1(n_432),
.A2(n_409),
.B(n_320),
.C(n_407),
.Y(n_442)
);

A2O1A1Ixp33_ASAP7_75t_L g443 ( 
.A1(n_437),
.A2(n_435),
.B(n_417),
.C(n_364),
.Y(n_443)
);

OAI32xp33_ASAP7_75t_L g444 ( 
.A1(n_438),
.A2(n_404),
.A3(n_410),
.B1(n_412),
.B2(n_376),
.Y(n_444)
);

AND2x4_ASAP7_75t_L g445 ( 
.A(n_443),
.B(n_440),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_445),
.Y(n_446)
);

NAND5xp2_ASAP7_75t_L g447 ( 
.A(n_446),
.B(n_442),
.C(n_439),
.D(n_445),
.E(n_441),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_447),
.B(n_361),
.Y(n_448)
);

AOI21xp5_ASAP7_75t_L g449 ( 
.A1(n_448),
.A2(n_444),
.B(n_417),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_449),
.Y(n_450)
);

AOI21xp33_ASAP7_75t_SL g451 ( 
.A1(n_450),
.A2(n_374),
.B(n_406),
.Y(n_451)
);


endmodule