module fake_jpeg_9007_n_331 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_331);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_331;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_13),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_6),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_7),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_40),
.Y(n_51)
);

CKINVDCx16_ASAP7_75t_R g40 ( 
.A(n_23),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_31),
.B(n_0),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_41),
.B(n_28),
.Y(n_54)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_42),
.B(n_31),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_16),
.B(n_15),
.Y(n_43)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_24),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_46),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_45),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_48),
.B(n_53),
.Y(n_83)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_52),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_43),
.B(n_16),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_54),
.B(n_32),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_44),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_55),
.B(n_61),
.Y(n_103)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

HB1xp67_ASAP7_75t_L g93 ( 
.A(n_56),
.Y(n_93)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_57),
.Y(n_94)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_41),
.B(n_16),
.Y(n_62)
);

CKINVDCx14_ASAP7_75t_R g80 ( 
.A(n_62),
.Y(n_80)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_63),
.B(n_67),
.Y(n_77)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

INVx1_ASAP7_75t_SL g84 ( 
.A(n_65),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

INVx1_ASAP7_75t_SL g92 ( 
.A(n_66),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_44),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_44),
.A2(n_31),
.B1(n_18),
.B2(n_22),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_68),
.A2(n_32),
.B1(n_28),
.B2(n_29),
.Y(n_86)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_36),
.Y(n_69)
);

BUFx2_ASAP7_75t_L g74 ( 
.A(n_69),
.Y(n_74)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_70),
.B(n_46),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_66),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_71),
.B(n_88),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_49),
.A2(n_18),
.B1(n_22),
.B2(n_20),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_72),
.A2(n_73),
.B1(n_76),
.B2(n_82),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_49),
.A2(n_18),
.B1(n_22),
.B2(n_42),
.Y(n_73)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_50),
.Y(n_75)
);

INVx11_ASAP7_75t_L g127 ( 
.A(n_75),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_50),
.A2(n_42),
.B1(n_37),
.B2(n_19),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_78),
.B(n_10),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_61),
.A2(n_37),
.B1(n_39),
.B2(n_38),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_81),
.A2(n_86),
.B1(n_91),
.B2(n_96),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_64),
.A2(n_19),
.B1(n_21),
.B2(n_29),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_64),
.A2(n_19),
.B1(n_21),
.B2(n_29),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_85),
.Y(n_114)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_87),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_66),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_68),
.B(n_21),
.Y(n_89)
);

CKINVDCx14_ASAP7_75t_R g126 ( 
.A(n_89),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_51),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_90),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_67),
.A2(n_39),
.B1(n_38),
.B2(n_46),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_66),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_95),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_59),
.A2(n_39),
.B1(n_38),
.B2(n_28),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_59),
.A2(n_32),
.B1(n_35),
.B2(n_26),
.Y(n_97)
);

O2A1O1Ixp33_ASAP7_75t_L g117 ( 
.A1(n_97),
.A2(n_104),
.B(n_109),
.C(n_96),
.Y(n_117)
);

OAI22xp33_ASAP7_75t_L g98 ( 
.A1(n_58),
.A2(n_27),
.B1(n_34),
.B2(n_35),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_98),
.A2(n_102),
.B1(n_106),
.B2(n_108),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_48),
.A2(n_27),
.B1(n_34),
.B2(n_35),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_99),
.B(n_100),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_63),
.B(n_0),
.Y(n_100)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_60),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_101),
.B(n_107),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_58),
.A2(n_25),
.B1(n_33),
.B2(n_17),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_47),
.A2(n_17),
.B1(n_33),
.B2(n_25),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_56),
.B(n_35),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_105),
.B(n_1),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_47),
.A2(n_33),
.B1(n_17),
.B2(n_26),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_60),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_57),
.A2(n_34),
.B1(n_26),
.B2(n_30),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_69),
.A2(n_34),
.B1(n_26),
.B2(n_30),
.Y(n_109)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_65),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_110),
.B(n_1),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_80),
.B(n_10),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_115),
.B(n_118),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_117),
.A2(n_109),
.B1(n_86),
.B2(n_75),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_80),
.B(n_10),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_77),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_119),
.B(n_137),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_120),
.B(n_12),
.Y(n_162)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_87),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_121),
.B(n_123),
.Y(n_145)
);

AO22x1_ASAP7_75t_L g122 ( 
.A1(n_89),
.A2(n_70),
.B1(n_30),
.B2(n_23),
.Y(n_122)
);

AO22x1_ASAP7_75t_L g172 ( 
.A1(n_122),
.A2(n_129),
.B1(n_94),
.B2(n_74),
.Y(n_172)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_77),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_128),
.B(n_130),
.Y(n_165)
);

AO21x2_ASAP7_75t_L g129 ( 
.A1(n_81),
.A2(n_23),
.B(n_2),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_105),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_78),
.B(n_1),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_131),
.B(n_134),
.Y(n_143)
);

OR2x2_ASAP7_75t_L g134 ( 
.A(n_83),
.B(n_1),
.Y(n_134)
);

A2O1A1Ixp33_ASAP7_75t_L g135 ( 
.A1(n_78),
.A2(n_83),
.B(n_89),
.C(n_100),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_135),
.B(n_131),
.Y(n_149)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_103),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_103),
.B(n_15),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_138),
.B(n_139),
.Y(n_154)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_91),
.Y(n_139)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_140),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_139),
.A2(n_99),
.B1(n_102),
.B2(n_79),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_141),
.A2(n_172),
.B1(n_122),
.B2(n_138),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_126),
.A2(n_100),
.B(n_79),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_144),
.A2(n_149),
.B(n_156),
.Y(n_184)
);

INVx13_ASAP7_75t_L g146 ( 
.A(n_136),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_146),
.B(n_148),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_147),
.A2(n_113),
.B1(n_133),
.B2(n_122),
.Y(n_203)
);

HB1xp67_ASAP7_75t_L g148 ( 
.A(n_129),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_111),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_150),
.B(n_151),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_112),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_117),
.A2(n_84),
.B1(n_110),
.B2(n_94),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_152),
.A2(n_157),
.B1(n_173),
.B2(n_132),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_111),
.B(n_127),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_155),
.B(n_163),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_114),
.A2(n_71),
.B(n_88),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_117),
.A2(n_84),
.B1(n_94),
.B2(n_104),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_126),
.A2(n_92),
.B(n_97),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_SL g179 ( 
.A(n_158),
.B(n_162),
.C(n_129),
.Y(n_179)
);

INVx4_ASAP7_75t_SL g159 ( 
.A(n_129),
.Y(n_159)
);

INVx1_ASAP7_75t_SL g192 ( 
.A(n_159),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_119),
.B(n_92),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_160),
.B(n_161),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_128),
.B(n_107),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_127),
.B(n_112),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_SL g166 ( 
.A(n_124),
.B(n_95),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_166),
.B(n_124),
.C(n_130),
.Y(n_186)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_123),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_167),
.B(n_168),
.Y(n_202)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_140),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_127),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_169),
.Y(n_193)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_129),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_170),
.B(n_93),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_116),
.B(n_101),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_171),
.B(n_116),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_129),
.A2(n_93),
.B1(n_74),
.B2(n_95),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_174),
.A2(n_187),
.B1(n_203),
.B2(n_205),
.Y(n_211)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_161),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_175),
.B(n_180),
.Y(n_223)
);

AOI22x1_ASAP7_75t_SL g176 ( 
.A1(n_166),
.A2(n_132),
.B1(n_129),
.B2(n_135),
.Y(n_176)
);

OAI21xp33_ASAP7_75t_SL g224 ( 
.A1(n_176),
.A2(n_179),
.B(n_189),
.Y(n_224)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_171),
.Y(n_180)
);

AND2x6_ASAP7_75t_L g181 ( 
.A(n_156),
.B(n_135),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_181),
.Y(n_218)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_160),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_182),
.B(n_188),
.Y(n_213)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_185),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_186),
.B(n_167),
.C(n_150),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_159),
.A2(n_113),
.B1(n_133),
.B2(n_121),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_165),
.Y(n_188)
);

NOR4xp25_ASAP7_75t_SL g189 ( 
.A(n_144),
.B(n_122),
.C(n_120),
.D(n_125),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_165),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_190),
.B(n_195),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_153),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_191),
.B(n_198),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_145),
.B(n_137),
.Y(n_194)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_194),
.Y(n_226)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_173),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_152),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_196),
.B(n_200),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_145),
.B(n_134),
.Y(n_197)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_197),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_169),
.Y(n_198)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_157),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_201),
.A2(n_164),
.B1(n_134),
.B2(n_162),
.Y(n_230)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_154),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_204),
.A2(n_168),
.B1(n_142),
.B2(n_151),
.Y(n_214)
);

AND2x6_ASAP7_75t_L g206 ( 
.A(n_158),
.B(n_133),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_206),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_186),
.B(n_149),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_208),
.B(n_210),
.C(n_216),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_195),
.A2(n_159),
.B1(n_170),
.B2(n_147),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_209),
.A2(n_192),
.B1(n_200),
.B2(n_188),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_178),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_212),
.B(n_219),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_214),
.B(n_227),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_184),
.B(n_141),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_179),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_184),
.B(n_143),
.C(n_142),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_220),
.B(n_222),
.C(n_194),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_176),
.A2(n_177),
.B(n_181),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_221),
.A2(n_234),
.B(n_169),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_183),
.B(n_143),
.C(n_172),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_199),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_225),
.B(n_228),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_187),
.A2(n_172),
.B1(n_115),
.B2(n_118),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_227),
.A2(n_233),
.B1(n_190),
.B2(n_197),
.Y(n_243)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_193),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_230),
.B(n_193),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_174),
.A2(n_146),
.B1(n_162),
.B2(n_74),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_182),
.A2(n_196),
.B(n_183),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_229),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_235),
.B(n_245),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_L g276 ( 
.A1(n_236),
.A2(n_238),
.B(n_241),
.Y(n_276)
);

AND2x4_ASAP7_75t_L g238 ( 
.A(n_219),
.B(n_192),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_SL g239 ( 
.A(n_208),
.B(n_185),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_239),
.B(n_213),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_216),
.B(n_201),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_240),
.B(n_249),
.C(n_251),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_217),
.A2(n_175),
.B(n_180),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_242),
.A2(n_255),
.B1(n_256),
.B2(n_257),
.Y(n_274)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_243),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_214),
.B(n_204),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_223),
.Y(n_246)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_246),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_232),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_247),
.B(n_252),
.Y(n_260)
);

AND2x6_ASAP7_75t_L g248 ( 
.A(n_218),
.B(n_206),
.Y(n_248)
);

INVxp33_ASAP7_75t_SL g271 ( 
.A(n_248),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_220),
.B(n_202),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_217),
.Y(n_250)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_250),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_210),
.B(n_226),
.Y(n_254)
);

CKINVDCx16_ASAP7_75t_R g259 ( 
.A(n_254),
.Y(n_259)
);

AO21x2_ASAP7_75t_L g256 ( 
.A1(n_209),
.A2(n_2),
.B(n_3),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_224),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_238),
.Y(n_258)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_258),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_247),
.B(n_226),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_261),
.B(n_265),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_238),
.A2(n_218),
.B1(n_207),
.B2(n_256),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_264),
.A2(n_256),
.B1(n_231),
.B2(n_211),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_237),
.B(n_213),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_244),
.B(n_222),
.C(n_234),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_266),
.B(n_267),
.C(n_270),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_244),
.B(n_215),
.C(n_221),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_269),
.B(n_239),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_251),
.B(n_215),
.C(n_231),
.Y(n_270)
);

HB1xp67_ASAP7_75t_L g273 ( 
.A(n_238),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_273),
.B(n_228),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_271),
.A2(n_255),
.B(n_276),
.Y(n_280)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_280),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_266),
.B(n_240),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_281),
.B(n_287),
.C(n_289),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_272),
.A2(n_256),
.B1(n_211),
.B2(n_248),
.Y(n_282)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_282),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_265),
.B(n_253),
.Y(n_283)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_283),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_284),
.B(n_290),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_SL g285 ( 
.A(n_276),
.B(n_249),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_SL g293 ( 
.A(n_285),
.B(n_288),
.Y(n_293)
);

CKINVDCx14_ASAP7_75t_R g286 ( 
.A(n_263),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_286),
.B(n_291),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_262),
.B(n_241),
.C(n_242),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_262),
.B(n_232),
.C(n_233),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_267),
.B(n_257),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_L g292 ( 
.A1(n_264),
.A2(n_15),
.B(n_14),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_292),
.A2(n_274),
.B(n_260),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_277),
.A2(n_274),
.B1(n_275),
.B2(n_259),
.Y(n_298)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_298),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_279),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_299),
.B(n_301),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_288),
.B(n_268),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_287),
.B(n_270),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g313 ( 
.A(n_303),
.B(n_305),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_285),
.A2(n_275),
.B1(n_268),
.B2(n_258),
.Y(n_304)
);

AND2x2_ASAP7_75t_L g306 ( 
.A(n_304),
.B(n_290),
.Y(n_306)
);

AOI322xp5_ASAP7_75t_L g318 ( 
.A1(n_306),
.A2(n_308),
.A3(n_293),
.B1(n_300),
.B2(n_294),
.C1(n_14),
.C2(n_11),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_297),
.B(n_278),
.C(n_289),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_SL g321 ( 
.A(n_307),
.B(n_309),
.Y(n_321)
);

AOI22xp33_ASAP7_75t_SL g308 ( 
.A1(n_295),
.A2(n_261),
.B1(n_260),
.B2(n_292),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_297),
.B(n_278),
.C(n_281),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_296),
.A2(n_269),
.B(n_284),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_310),
.A2(n_314),
.B(n_298),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_302),
.A2(n_14),
.B(n_13),
.Y(n_314)
);

HB1xp67_ASAP7_75t_L g315 ( 
.A(n_308),
.Y(n_315)
);

NAND3xp33_ASAP7_75t_SL g323 ( 
.A(n_315),
.B(n_317),
.C(n_318),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_316),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_324)
);

NOR3xp33_ASAP7_75t_SL g317 ( 
.A(n_306),
.B(n_304),
.C(n_313),
.Y(n_317)
);

AOI322xp5_ASAP7_75t_L g319 ( 
.A1(n_311),
.A2(n_293),
.A3(n_294),
.B1(n_11),
.B2(n_7),
.C1(n_3),
.C2(n_9),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_L g322 ( 
.A1(n_319),
.A2(n_320),
.B(n_6),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_SL g320 ( 
.A1(n_312),
.A2(n_3),
.B(n_5),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_322),
.B(n_324),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_SL g325 ( 
.A(n_321),
.B(n_8),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_325),
.B(n_9),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_SL g328 ( 
.A1(n_327),
.A2(n_326),
.B(n_323),
.Y(n_328)
);

OR2x2_ASAP7_75t_L g329 ( 
.A(n_328),
.B(n_9),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_329),
.B(n_9),
.Y(n_330)
);

BUFx24_ASAP7_75t_SL g331 ( 
.A(n_330),
.Y(n_331)
);


endmodule