module fake_jpeg_16725_n_31 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_31);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_31;

wire n_13;
wire n_21;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_20;
wire n_18;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_11;
wire n_17;
wire n_25;
wire n_29;
wire n_12;
wire n_15;

INVx2_ASAP7_75t_L g10 ( 
.A(n_4),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_2),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_L g12 ( 
.A(n_0),
.B(n_2),
.Y(n_12)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_SL g14 ( 
.A(n_4),
.B(n_3),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_7),
.B(n_3),
.Y(n_15)
);

BUFx2_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_L g17 ( 
.A1(n_0),
.A2(n_1),
.B1(n_9),
.B2(n_6),
.Y(n_17)
);

INVx5_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g19 ( 
.A(n_8),
.B(n_6),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_20),
.Y(n_25)
);

OA22x2_ASAP7_75t_L g21 ( 
.A1(n_10),
.A2(n_1),
.B1(n_13),
.B2(n_18),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_L g27 ( 
.A1(n_21),
.A2(n_22),
.B1(n_16),
.B2(n_15),
.Y(n_27)
);

A2O1A1Ixp33_ASAP7_75t_SL g22 ( 
.A1(n_17),
.A2(n_13),
.B(n_16),
.C(n_18),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_14),
.B(n_11),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_23),
.B(n_24),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_14),
.B(n_11),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_27),
.B(n_21),
.Y(n_29)
);

BUFx24_ASAP7_75t_SL g28 ( 
.A(n_26),
.Y(n_28)
);

A2O1A1Ixp33_ASAP7_75t_L g30 ( 
.A1(n_28),
.A2(n_29),
.B(n_23),
.C(n_12),
.Y(n_30)
);

OAI311xp33_ASAP7_75t_L g31 ( 
.A1(n_30),
.A2(n_19),
.A3(n_22),
.B1(n_25),
.C1(n_28),
.Y(n_31)
);


endmodule