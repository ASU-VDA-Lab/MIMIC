module fake_jpeg_19114_n_300 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_300);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_300;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx4f_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

CKINVDCx16_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_13),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx24_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_28),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_39),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_39),
.A2(n_26),
.B1(n_31),
.B2(n_25),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_41),
.A2(n_51),
.B1(n_34),
.B2(n_29),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_33),
.B(n_25),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_44),
.B(n_46),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_33),
.B(n_27),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_39),
.B(n_19),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_50),
.B(n_54),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_39),
.A2(n_26),
.B1(n_31),
.B2(n_29),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_37),
.A2(n_26),
.B1(n_31),
.B2(n_27),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_53),
.A2(n_37),
.B1(n_34),
.B2(n_33),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_33),
.B(n_23),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_55),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_57),
.A2(n_68),
.B1(n_72),
.B2(n_80),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_48),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_58),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_54),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_59),
.B(n_63),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_50),
.A2(n_38),
.B1(n_36),
.B2(n_37),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_60),
.B(n_67),
.Y(n_95)
);

HB1xp67_ASAP7_75t_L g61 ( 
.A(n_50),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_61),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_43),
.A2(n_30),
.B1(n_16),
.B2(n_23),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_62),
.A2(n_32),
.B(n_35),
.Y(n_101)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_47),
.A2(n_16),
.B1(n_30),
.B2(n_36),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_64),
.Y(n_97)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_65),
.B(n_66),
.Y(n_90)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_53),
.A2(n_38),
.B1(n_36),
.B2(n_37),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_41),
.B(n_35),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_47),
.A2(n_30),
.B1(n_16),
.B2(n_36),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_70),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_51),
.A2(n_38),
.B1(n_34),
.B2(n_29),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_71),
.B(n_74),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_47),
.B(n_35),
.Y(n_72)
);

NAND3xp33_ASAP7_75t_L g73 ( 
.A(n_44),
.B(n_19),
.C(n_34),
.Y(n_73)
);

OAI21xp33_ASAP7_75t_L g111 ( 
.A1(n_73),
.A2(n_45),
.B(n_32),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_46),
.A2(n_38),
.B1(n_34),
.B2(n_52),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_49),
.Y(n_75)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_75),
.Y(n_87)
);

OAI22xp33_ASAP7_75t_L g106 ( 
.A1(n_76),
.A2(n_45),
.B1(n_42),
.B2(n_32),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_52),
.A2(n_19),
.B1(n_24),
.B2(n_17),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_77),
.B(n_83),
.Y(n_100)
);

INVx1_ASAP7_75t_SL g78 ( 
.A(n_40),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_78),
.B(n_81),
.Y(n_91)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_79),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_52),
.B(n_35),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_49),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_52),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_82),
.Y(n_107)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_48),
.Y(n_83)
);

OAI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_65),
.A2(n_49),
.B1(n_40),
.B2(n_42),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_86),
.A2(n_98),
.B1(n_106),
.B2(n_60),
.Y(n_123)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_58),
.Y(n_89)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_89),
.Y(n_115)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_58),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_92),
.Y(n_116)
);

A2O1A1Ixp33_ASAP7_75t_L g93 ( 
.A1(n_56),
.A2(n_24),
.B(n_35),
.C(n_32),
.Y(n_93)
);

A2O1A1Ixp33_ASAP7_75t_L g112 ( 
.A1(n_93),
.A2(n_69),
.B(n_62),
.C(n_68),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_59),
.A2(n_42),
.B1(n_45),
.B2(n_40),
.Y(n_94)
);

INVx1_ASAP7_75t_SL g114 ( 
.A(n_94),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_76),
.A2(n_40),
.B1(n_42),
.B2(n_45),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_101),
.A2(n_111),
.B1(n_80),
.B2(n_72),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_56),
.B(n_19),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_102),
.B(n_103),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_55),
.B(n_63),
.Y(n_103)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_72),
.Y(n_105)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_105),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_74),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_110),
.B(n_67),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_112),
.B(n_119),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_113),
.A2(n_104),
.B(n_22),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_117),
.A2(n_22),
.B(n_21),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_103),
.B(n_69),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_90),
.Y(n_120)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_120),
.Y(n_151)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_90),
.Y(n_121)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_121),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_95),
.A2(n_61),
.B1(n_68),
.B2(n_71),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_122),
.A2(n_124),
.B1(n_129),
.B2(n_133),
.Y(n_158)
);

OAI21xp33_ASAP7_75t_SL g154 ( 
.A1(n_123),
.A2(n_104),
.B(n_108),
.Y(n_154)
);

OAI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_97),
.A2(n_79),
.B1(n_66),
.B2(n_83),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_99),
.B(n_82),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_125),
.B(n_137),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_95),
.A2(n_77),
.B1(n_80),
.B2(n_79),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_126),
.A2(n_130),
.B1(n_135),
.B2(n_94),
.Y(n_145)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_91),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_127),
.Y(n_153)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_91),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_128),
.Y(n_165)
);

OAI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_109),
.A2(n_66),
.B1(n_81),
.B2(n_75),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_96),
.A2(n_99),
.B1(n_105),
.B2(n_100),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_84),
.Y(n_131)
);

INVx1_ASAP7_75t_SL g163 ( 
.A(n_131),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_101),
.A2(n_78),
.B1(n_20),
.B2(n_18),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_132),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_96),
.A2(n_85),
.B1(n_100),
.B2(n_102),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_86),
.A2(n_78),
.B1(n_32),
.B2(n_12),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_87),
.A2(n_35),
.B1(n_11),
.B2(n_12),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_136),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_88),
.B(n_20),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_93),
.B(n_18),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_138),
.B(n_35),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_112),
.A2(n_93),
.B(n_88),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_141),
.A2(n_149),
.B(n_150),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_114),
.A2(n_84),
.B1(n_85),
.B2(n_107),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_142),
.Y(n_191)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_115),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_143),
.B(n_166),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_145),
.A2(n_147),
.B1(n_159),
.B2(n_0),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_134),
.B(n_85),
.C(n_107),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_146),
.B(n_156),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_130),
.A2(n_98),
.B1(n_87),
.B2(n_92),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_131),
.Y(n_148)
);

OR2x2_ASAP7_75t_L g170 ( 
.A(n_148),
.B(n_157),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_114),
.A2(n_89),
.B(n_87),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_138),
.A2(n_0),
.B(n_1),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_117),
.A2(n_0),
.B(n_1),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_152),
.A2(n_155),
.B(n_161),
.Y(n_193)
);

OA22x2_ASAP7_75t_L g175 ( 
.A1(n_154),
.A2(n_128),
.B1(n_123),
.B2(n_135),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_118),
.A2(n_18),
.B1(n_20),
.B2(n_17),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_134),
.B(n_35),
.C(n_108),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_126),
.A2(n_108),
.B1(n_104),
.B2(n_22),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_160),
.A2(n_118),
.B1(n_132),
.B2(n_127),
.Y(n_171)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_115),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_120),
.A2(n_22),
.B(n_21),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_167),
.A2(n_161),
.B(n_160),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_119),
.B(n_121),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_168),
.B(n_14),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_133),
.B(n_113),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_169),
.B(n_122),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_171),
.A2(n_183),
.B(n_150),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_151),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_172),
.Y(n_205)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_151),
.Y(n_173)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_173),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_174),
.B(n_181),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_175),
.B(n_177),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_158),
.A2(n_125),
.B1(n_137),
.B2(n_116),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_176),
.A2(n_192),
.B1(n_195),
.B2(n_157),
.Y(n_202)
);

AOI22x1_ASAP7_75t_L g177 ( 
.A1(n_145),
.A2(n_116),
.B1(n_21),
.B2(n_17),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_158),
.A2(n_21),
.B1(n_17),
.B2(n_15),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_178),
.A2(n_186),
.B1(n_188),
.B2(n_189),
.Y(n_204)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_164),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_179),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_180),
.B(n_185),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_146),
.B(n_15),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_164),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_184),
.Y(n_214)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_168),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_144),
.Y(n_186)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_144),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_152),
.A2(n_14),
.B1(n_13),
.B2(n_11),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_190),
.A2(n_194),
.B1(n_196),
.B2(n_198),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_142),
.A2(n_140),
.B1(n_139),
.B2(n_141),
.Y(n_192)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_156),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_140),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_149),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_153),
.B(n_1),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_147),
.A2(n_14),
.B1(n_13),
.B2(n_11),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_199),
.A2(n_163),
.B1(n_143),
.B2(n_10),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_182),
.A2(n_165),
.B1(n_153),
.B2(n_162),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_200),
.B(n_203),
.Y(n_222)
);

CKINVDCx14_ASAP7_75t_R g224 ( 
.A(n_202),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_176),
.A2(n_159),
.B1(n_169),
.B2(n_165),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_206),
.B(n_212),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_182),
.A2(n_148),
.B1(n_163),
.B2(n_167),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_207),
.B(n_171),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_188),
.A2(n_199),
.B1(n_191),
.B2(n_170),
.Y(n_209)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_209),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_191),
.A2(n_163),
.B1(n_155),
.B2(n_166),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_213),
.A2(n_216),
.B1(n_175),
.B2(n_177),
.Y(n_229)
);

INVx3_ASAP7_75t_SL g215 ( 
.A(n_187),
.Y(n_215)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_215),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_192),
.A2(n_175),
.B1(n_177),
.B2(n_197),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_197),
.B(n_2),
.C(n_3),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_217),
.B(n_220),
.C(n_195),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_181),
.B(n_2),
.C(n_4),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_170),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_221),
.B(n_180),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_225),
.B(n_220),
.Y(n_251)
);

CKINVDCx16_ASAP7_75t_R g249 ( 
.A(n_226),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_218),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_227),
.Y(n_254)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_218),
.Y(n_228)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_228),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_229),
.A2(n_238),
.B1(n_201),
.B2(n_207),
.Y(n_241)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_204),
.Y(n_230)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_230),
.Y(n_252)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_210),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_231),
.B(n_211),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_232),
.B(n_222),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_210),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_233),
.B(n_236),
.Y(n_245)
);

NAND3xp33_ASAP7_75t_SL g236 ( 
.A(n_202),
.B(n_193),
.C(n_183),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_219),
.B(n_174),
.C(n_216),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_237),
.B(n_219),
.C(n_203),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_201),
.A2(n_175),
.B1(n_193),
.B2(n_198),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_213),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_239),
.B(n_208),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_240),
.B(n_246),
.Y(n_255)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_241),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_237),
.B(n_206),
.C(n_200),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_243),
.B(n_244),
.C(n_222),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_224),
.B(n_223),
.C(n_231),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_247),
.B(n_248),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_234),
.A2(n_211),
.B1(n_215),
.B2(n_214),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_223),
.B(n_215),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_250),
.B(n_253),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_251),
.B(n_246),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_257),
.B(n_258),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_251),
.B(n_240),
.C(n_244),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_243),
.B(n_232),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_259),
.B(n_264),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_254),
.B(n_214),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_260),
.B(n_265),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_245),
.A2(n_228),
.B(n_205),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_263),
.A2(n_242),
.B1(n_205),
.B2(n_235),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_245),
.B(n_217),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_R g265 ( 
.A(n_253),
.B(n_238),
.C(n_229),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_266),
.B(n_247),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_265),
.A2(n_241),
.B1(n_230),
.B2(n_252),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_267),
.B(n_271),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_270),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_256),
.B(n_249),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_261),
.B(n_252),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_272),
.B(n_273),
.Y(n_279)
);

INVxp67_ASAP7_75t_SL g273 ( 
.A(n_262),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_257),
.A2(n_235),
.B1(n_239),
.B2(n_250),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_274),
.B(n_275),
.Y(n_280)
);

NOR2xp67_ASAP7_75t_SL g281 ( 
.A(n_274),
.B(n_258),
.Y(n_281)
);

AND2x2_ASAP7_75t_L g287 ( 
.A(n_281),
.B(n_269),
.Y(n_287)
);

OR2x2_ASAP7_75t_L g282 ( 
.A(n_276),
.B(n_242),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_282),
.B(n_283),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_268),
.B(n_266),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_276),
.A2(n_255),
.B(n_225),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_284),
.B(n_9),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_SL g285 ( 
.A(n_279),
.B(n_255),
.Y(n_285)
);

INVxp33_ASAP7_75t_L g292 ( 
.A(n_285),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_287),
.B(n_288),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_277),
.B(n_267),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_289),
.A2(n_290),
.B1(n_280),
.B2(n_6),
.Y(n_293)
);

AND2x2_ASAP7_75t_L g290 ( 
.A(n_282),
.B(n_278),
.Y(n_290)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_293),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_291),
.A2(n_286),
.B(n_6),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_294),
.A2(n_4),
.B(n_7),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_296),
.B(n_295),
.C(n_292),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_297),
.B(n_9),
.C(n_7),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_L g299 ( 
.A1(n_298),
.A2(n_8),
.B(n_9),
.Y(n_299)
);

OAI21xp33_ASAP7_75t_L g300 ( 
.A1(n_299),
.A2(n_8),
.B(n_9),
.Y(n_300)
);


endmodule