module fake_jpeg_13895_n_135 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_135);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_135;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_96;

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

INVx2_ASAP7_75t_R g41 ( 
.A(n_36),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_32),
.Y(n_47)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_25),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_18),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_16),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_31),
.B(n_27),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_21),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_2),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_30),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_2),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_4),
.Y(n_57)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_59),
.Y(n_76)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_60),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_41),
.B(n_0),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_61),
.B(n_54),
.Y(n_68)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_62),
.Y(n_73)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_63),
.B(n_65),
.Y(n_72)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

CKINVDCx6p67_ASAP7_75t_R g67 ( 
.A(n_64),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_63),
.B(n_41),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_66),
.B(n_71),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_68),
.B(n_75),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_60),
.A2(n_40),
.B1(n_56),
.B2(n_48),
.Y(n_69)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_69),
.A2(n_48),
.B(n_58),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_59),
.B(n_49),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_70),
.B(n_55),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_64),
.B(n_57),
.Y(n_71)
);

OR2x2_ASAP7_75t_L g75 ( 
.A(n_65),
.B(n_51),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_61),
.B(n_47),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_77),
.B(n_78),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_61),
.B(n_53),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_70),
.A2(n_72),
.B1(n_76),
.B2(n_73),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_79),
.A2(n_90),
.B1(n_8),
.B2(n_9),
.Y(n_97)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_74),
.Y(n_81)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_81),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g98 ( 
.A1(n_82),
.A2(n_87),
.B(n_88),
.Y(n_98)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_74),
.Y(n_84)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_84),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g85 ( 
.A(n_72),
.B(n_52),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_85),
.B(n_94),
.C(n_34),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_69),
.A2(n_55),
.B1(n_43),
.B2(n_42),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_SL g88 ( 
.A1(n_67),
.A2(n_50),
.B(n_1),
.Y(n_88)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_67),
.Y(n_89)
);

NAND2xp33_ASAP7_75t_SL g104 ( 
.A(n_89),
.B(n_92),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_76),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_90)
);

AND2x4_ASAP7_75t_L g92 ( 
.A(n_67),
.B(n_6),
.Y(n_92)
);

OR2x2_ASAP7_75t_L g93 ( 
.A(n_68),
.B(n_6),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_93),
.B(n_95),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_70),
.B(n_20),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_67),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_80),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_96),
.A2(n_15),
.B(n_17),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_97),
.A2(n_24),
.B1(n_26),
.B2(n_28),
.Y(n_118)
);

NOR3xp33_ASAP7_75t_SL g99 ( 
.A(n_91),
.B(n_10),
.C(n_11),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_99),
.B(n_102),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_83),
.B(n_23),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_101),
.B(n_103),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_91),
.B(n_10),
.Y(n_102)
);

BUFx12f_ASAP7_75t_L g105 ( 
.A(n_89),
.Y(n_105)
);

BUFx5_ASAP7_75t_L g119 ( 
.A(n_105),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_95),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_106),
.B(n_110),
.Y(n_114)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_92),
.Y(n_109)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_109),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_86),
.B(n_12),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_84),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_111),
.B(n_33),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_85),
.B(n_13),
.C(n_14),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_112),
.B(n_22),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_113),
.B(n_115),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_117),
.B(n_118),
.C(n_98),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_SL g121 ( 
.A(n_104),
.B(n_29),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_SL g125 ( 
.A(n_121),
.B(n_100),
.Y(n_125)
);

INVx13_ASAP7_75t_L g123 ( 
.A(n_119),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_123),
.B(n_124),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_125),
.B(n_116),
.C(n_102),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g127 ( 
.A(n_122),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_127),
.A2(n_105),
.B1(n_108),
.B2(n_107),
.Y(n_128)
);

FAx1_ASAP7_75t_SL g131 ( 
.A(n_128),
.B(n_130),
.CI(n_120),
.CON(n_131),
.SN(n_131)
);

AOI21x1_ASAP7_75t_L g132 ( 
.A1(n_131),
.A2(n_130),
.B(n_100),
.Y(n_132)
);

NOR3xp33_ASAP7_75t_L g133 ( 
.A(n_132),
.B(n_131),
.C(n_129),
.Y(n_133)
);

AOI322xp5_ASAP7_75t_L g134 ( 
.A1(n_133),
.A2(n_131),
.A3(n_114),
.B1(n_125),
.B2(n_126),
.C1(n_127),
.C2(n_110),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_134),
.B(n_114),
.Y(n_135)
);


endmodule