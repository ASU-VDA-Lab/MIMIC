module fake_netlist_1_10645_n_13 (n_1, n_2, n_0, n_13);
input n_1;
input n_2;
input n_0;
output n_13;
wire n_11;
wire n_12;
wire n_6;
wire n_4;
wire n_3;
wire n_9;
wire n_5;
wire n_7;
wire n_10;
wire n_8;
INVx1_ASAP7_75t_L g3 ( .A(n_2), .Y(n_3) );
BUFx3_ASAP7_75t_L g4 ( .A(n_0), .Y(n_4) );
BUFx6f_ASAP7_75t_L g5 ( .A(n_4), .Y(n_5) );
OA21x2_ASAP7_75t_L g6 ( .A1(n_3), .A2(n_0), .B(n_1), .Y(n_6) );
INVxp67_ASAP7_75t_SL g7 ( .A(n_5), .Y(n_7) );
INVxp67_ASAP7_75t_L g8 ( .A(n_5), .Y(n_8) );
OAI21xp5_ASAP7_75t_L g9 ( .A1(n_7), .A2(n_6), .B(n_4), .Y(n_9) );
AOI222xp33_ASAP7_75t_L g10 ( .A1(n_9), .A2(n_4), .B1(n_3), .B2(n_5), .C1(n_8), .C2(n_1), .Y(n_10) );
NOR3xp33_ASAP7_75t_L g11 ( .A(n_9), .B(n_4), .C(n_8), .Y(n_11) );
OAI22xp5_ASAP7_75t_L g12 ( .A1(n_11), .A2(n_6), .B1(n_1), .B2(n_0), .Y(n_12) );
AOI21xp5_ASAP7_75t_L g13 ( .A1(n_12), .A2(n_10), .B(n_6), .Y(n_13) );
endmodule