module fake_jpeg_3533_n_112 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_112);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_112;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

BUFx4f_ASAP7_75t_SL g33 ( 
.A(n_11),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

INVx11_ASAP7_75t_SL g38 ( 
.A(n_24),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_12),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_23),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_39),
.B(n_0),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_44),
.B(n_40),
.Y(n_51)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_37),
.B(n_1),
.Y(n_49)
);

OR2x2_ASAP7_75t_L g53 ( 
.A(n_49),
.B(n_50),
.Y(n_53)
);

INVx6_ASAP7_75t_SL g50 ( 
.A(n_38),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_51),
.B(n_60),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_49),
.B(n_41),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_54),
.B(n_55),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_50),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_56),
.B(n_33),
.Y(n_64)
);

AOI21xp33_ASAP7_75t_L g60 ( 
.A1(n_47),
.A2(n_38),
.B(n_33),
.Y(n_60)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_58),
.Y(n_63)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_63),
.Y(n_72)
);

INVx1_ASAP7_75t_SL g77 ( 
.A(n_64),
.Y(n_77)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_58),
.Y(n_65)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_65),
.Y(n_76)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_56),
.Y(n_66)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_66),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_53),
.B(n_33),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_67),
.B(n_68),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_53),
.B(n_43),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_57),
.B(n_1),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_69),
.B(n_2),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_59),
.A2(n_48),
.B1(n_46),
.B2(n_36),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_70),
.A2(n_52),
.B1(n_48),
.B2(n_46),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_59),
.B(n_43),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_71),
.B(n_2),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_73),
.B(n_74),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_63),
.A2(n_52),
.B1(n_36),
.B2(n_42),
.Y(n_74)
);

NAND3xp33_ASAP7_75t_L g91 ( 
.A(n_75),
.B(n_3),
.C(n_4),
.Y(n_91)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_65),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_79),
.B(n_3),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_61),
.B(n_69),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_80),
.B(n_62),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_81),
.Y(n_86)
);

AND2x4_ASAP7_75t_SL g82 ( 
.A(n_61),
.B(n_42),
.Y(n_82)
);

CKINVDCx14_ASAP7_75t_R g88 ( 
.A(n_82),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_84),
.B(n_85),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_80),
.B(n_66),
.Y(n_85)
);

XOR2xp5_ASAP7_75t_L g87 ( 
.A(n_83),
.B(n_19),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_87),
.B(n_90),
.C(n_92),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_77),
.B(n_20),
.C(n_31),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_91),
.B(n_9),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_78),
.B(n_18),
.C(n_30),
.Y(n_92)
);

A2O1A1O1Ixp25_ASAP7_75t_L g93 ( 
.A1(n_82),
.A2(n_16),
.B(n_29),
.C(n_28),
.D(n_27),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_93),
.A2(n_14),
.B(n_26),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_94),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_88),
.A2(n_75),
.B1(n_76),
.B2(n_72),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_95),
.A2(n_7),
.B1(n_8),
.B2(n_32),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_98),
.B(n_99),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_89),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_101),
.A2(n_86),
.B1(n_94),
.B2(n_89),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_103),
.B(n_104),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_100),
.B(n_5),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_105),
.B(n_99),
.C(n_96),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_107),
.A2(n_96),
.B(n_102),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_108),
.A2(n_97),
.B(n_106),
.Y(n_109)
);

OAI21xp33_ASAP7_75t_SL g110 ( 
.A1(n_109),
.A2(n_105),
.B(n_21),
.Y(n_110)
);

AOI21x1_ASAP7_75t_SL g111 ( 
.A1(n_110),
.A2(n_22),
.B(n_7),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_111),
.B(n_8),
.Y(n_112)
);


endmodule