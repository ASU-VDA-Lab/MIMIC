module real_jpeg_4878_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_498;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_378;
wire n_98;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_543;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_548;
wire n_319;
wire n_493;
wire n_93;
wire n_242;
wire n_487;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_546;
wire n_531;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_450;
wire n_333;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_343;
wire n_292;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AND2x2_ASAP7_75t_L g147 ( 
.A(n_0),
.B(n_148),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_0),
.B(n_177),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_0),
.B(n_202),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g207 ( 
.A(n_0),
.B(n_208),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g238 ( 
.A(n_0),
.B(n_239),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_0),
.B(n_322),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_0),
.B(n_354),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_0),
.B(n_38),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_1),
.B(n_110),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_1),
.B(n_119),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_1),
.B(n_156),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_1),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_1),
.B(n_129),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_1),
.B(n_246),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_1),
.B(n_259),
.Y(n_258)
);

INVx1_ASAP7_75t_SL g33 ( 
.A(n_2),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_2),
.B(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_2),
.B(n_42),
.Y(n_41)
);

AND2x2_ASAP7_75t_SL g61 ( 
.A(n_2),
.B(n_62),
.Y(n_61)
);

AND2x2_ASAP7_75t_SL g75 ( 
.A(n_2),
.B(n_76),
.Y(n_75)
);

AND2x2_ASAP7_75t_SL g369 ( 
.A(n_2),
.B(n_370),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_2),
.B(n_450),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_3),
.B(n_68),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_3),
.B(n_102),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_3),
.B(n_208),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_3),
.B(n_340),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_3),
.B(n_400),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_3),
.B(n_62),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_3),
.B(n_482),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_3),
.B(n_57),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_4),
.B(n_102),
.Y(n_101)
);

AND2x2_ASAP7_75t_SL g128 ( 
.A(n_4),
.B(n_129),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_4),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_4),
.B(n_307),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_4),
.B(n_357),
.Y(n_356)
);

AND2x2_ASAP7_75t_L g413 ( 
.A(n_4),
.B(n_414),
.Y(n_413)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_5),
.Y(n_104)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_5),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_5),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_5),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g370 ( 
.A(n_5),
.Y(n_370)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_6),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_6),
.Y(n_68)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_6),
.Y(n_74)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_6),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g437 ( 
.A(n_6),
.Y(n_437)
);

BUFx5_ASAP7_75t_L g477 ( 
.A(n_6),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_7),
.B(n_42),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_7),
.B(n_139),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_7),
.B(n_158),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_7),
.B(n_102),
.Y(n_220)
);

AND2x2_ASAP7_75t_L g234 ( 
.A(n_7),
.B(n_235),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_7),
.B(n_202),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_7),
.B(n_316),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_7),
.B(n_68),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_8),
.B(n_47),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_8),
.B(n_55),
.Y(n_54)
);

AND2x2_ASAP7_75t_SL g296 ( 
.A(n_8),
.B(n_206),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_8),
.B(n_366),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_8),
.B(n_402),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_8),
.B(n_461),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_8),
.B(n_480),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_8),
.B(n_507),
.Y(n_506)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_9),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g185 ( 
.A(n_9),
.Y(n_185)
);

INVx3_ASAP7_75t_L g494 ( 
.A(n_9),
.Y(n_494)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_11),
.Y(n_131)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_11),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_11),
.Y(n_202)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_12),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_13),
.B(n_72),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_13),
.B(n_172),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_13),
.B(n_187),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_13),
.B(n_320),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_13),
.B(n_350),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_13),
.B(n_396),
.Y(n_395)
);

AND2x2_ASAP7_75t_L g441 ( 
.A(n_13),
.B(n_442),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_SL g492 ( 
.A(n_13),
.B(n_493),
.Y(n_492)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_14),
.Y(n_99)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_14),
.Y(n_170)
);

BUFx3_ASAP7_75t_L g368 ( 
.A(n_14),
.Y(n_368)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_15),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_16),
.B(n_97),
.Y(n_96)
);

AND2x2_ASAP7_75t_SL g124 ( 
.A(n_16),
.B(n_125),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_16),
.B(n_143),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g204 ( 
.A(n_16),
.B(n_205),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_16),
.B(n_313),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_16),
.B(n_343),
.Y(n_342)
);

CKINVDCx16_ASAP7_75t_R g386 ( 
.A(n_16),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_16),
.B(n_437),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_17),
.B(n_106),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_17),
.B(n_162),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_17),
.B(n_183),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_17),
.B(n_218),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g224 ( 
.A(n_17),
.B(n_225),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_17),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_17),
.B(n_38),
.Y(n_293)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_19),
.A2(n_21),
.B1(n_24),
.B2(n_26),
.Y(n_20)
);

INVx13_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_23),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

O2A1O1Ixp33_ASAP7_75t_SL g26 ( 
.A1(n_27),
.A2(n_36),
.B(n_83),
.C(n_549),
.Y(n_26)
);

CKINVDCx14_ASAP7_75t_R g27 ( 
.A(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_50),
.Y(n_28)
);

OR2x2_ASAP7_75t_L g549 ( 
.A(n_29),
.B(n_50),
.Y(n_549)
);

XNOR2xp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_40),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_31),
.A2(n_32),
.B1(n_36),
.B2(n_37),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_31),
.A2(n_32),
.B1(n_41),
.B2(n_66),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g31 ( 
.A(n_32),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_32),
.B(n_41),
.C(n_46),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_34),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_33),
.B(n_390),
.Y(n_389)
);

INVx6_ASAP7_75t_L g316 ( 
.A(n_34),
.Y(n_316)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_35),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_37),
.Y(n_36)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_41),
.A2(n_60),
.B1(n_61),
.B2(n_66),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_41),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_41),
.B(n_54),
.C(n_61),
.Y(n_80)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_44),
.Y(n_108)
);

BUFx5_ASAP7_75t_L g156 ( 
.A(n_44),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g323 ( 
.A(n_44),
.Y(n_323)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g344 ( 
.A(n_45),
.Y(n_344)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_45),
.Y(n_416)
);

BUFx5_ASAP7_75t_L g446 ( 
.A(n_45),
.Y(n_446)
);

INVx3_ASAP7_75t_L g509 ( 
.A(n_45),
.Y(n_509)
);

XNOR2xp5_ASAP7_75t_L g81 ( 
.A(n_46),
.B(n_82),
.Y(n_81)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_79),
.C(n_81),
.Y(n_50)
);

XNOR2xp5_ASAP7_75t_L g538 ( 
.A(n_51),
.B(n_539),
.Y(n_538)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_67),
.C(n_69),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g534 ( 
.A1(n_52),
.A2(n_53),
.B1(n_535),
.B2(n_536),
.Y(n_534)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

XOR2xp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_59),
.Y(n_53)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_60),
.B(n_70),
.C(n_75),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g498 ( 
.A1(n_60),
.A2(n_61),
.B1(n_75),
.B2(n_495),
.Y(n_498)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_61),
.Y(n_60)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx4_ASAP7_75t_L g314 ( 
.A(n_64),
.Y(n_314)
);

BUFx6f_ASAP7_75t_L g359 ( 
.A(n_64),
.Y(n_359)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_65),
.Y(n_141)
);

BUFx3_ASAP7_75t_L g163 ( 
.A(n_65),
.Y(n_163)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_65),
.Y(n_180)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_65),
.Y(n_259)
);

INVx3_ASAP7_75t_L g398 ( 
.A(n_65),
.Y(n_398)
);

XOR2xp5_ASAP7_75t_L g536 ( 
.A(n_67),
.B(n_69),
.Y(n_536)
);

AOI22xp5_ASAP7_75t_L g496 ( 
.A1(n_70),
.A2(n_71),
.B1(n_497),
.B2(n_498),
.Y(n_496)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g495 ( 
.A(n_75),
.Y(n_495)
);

OAI22xp5_ASAP7_75t_L g513 ( 
.A1(n_75),
.A2(n_448),
.B1(n_449),
.B2(n_495),
.Y(n_513)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx3_ASAP7_75t_L g400 ( 
.A(n_77),
.Y(n_400)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_78),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g151 ( 
.A(n_78),
.Y(n_151)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_78),
.Y(n_159)
);

INVx11_ASAP7_75t_L g231 ( 
.A(n_78),
.Y(n_231)
);

INVx3_ASAP7_75t_L g352 ( 
.A(n_78),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_L g539 ( 
.A1(n_79),
.A2(n_80),
.B1(n_81),
.B2(n_540),
.Y(n_539)
);

CKINVDCx14_ASAP7_75t_R g79 ( 
.A(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_81),
.Y(n_540)
);

AO21x1_ASAP7_75t_SL g83 ( 
.A1(n_84),
.A2(n_467),
.B(n_542),
.Y(n_83)
);

OAI21x1_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_423),
.B(n_466),
.Y(n_84)
);

AOI21x1_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_378),
.B(n_422),
.Y(n_85)
);

OAI21x1_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_327),
.B(n_377),
.Y(n_86)
);

AOI21x1_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_286),
.B(n_326),
.Y(n_87)
);

AO21x1_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_211),
.B(n_285),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_90),
.B(n_195),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_90),
.B(n_195),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_91),
.A2(n_92),
.B1(n_134),
.B2(n_194),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_91),
.B(n_135),
.C(n_174),
.Y(n_325)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_112),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_93),
.B(n_113),
.C(n_133),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_105),
.C(n_109),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_94),
.B(n_210),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_100),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_95),
.A2(n_96),
.B1(n_100),
.B2(n_101),
.Y(n_200)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_97),
.Y(n_219)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_99),
.Y(n_208)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx8_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx3_ASAP7_75t_L g246 ( 
.A(n_104),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_105),
.B(n_109),
.Y(n_210)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_111),
.B(n_386),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_117),
.B1(n_132),
.B2(n_133),
.Y(n_112)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_113),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_114),
.A2(n_115),
.B(n_116),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_114),
.B(n_115),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_SL g299 ( 
.A(n_116),
.B(n_300),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_116),
.B(n_291),
.C(n_300),
.Y(n_334)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_117),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_123),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_118),
.B(n_124),
.C(n_128),
.Y(n_324)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_128),
.Y(n_123)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx8_ASAP7_75t_L g320 ( 
.A(n_130),
.Y(n_320)
);

BUFx5_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g341 ( 
.A(n_131),
.Y(n_341)
);

BUFx3_ASAP7_75t_L g451 ( 
.A(n_131),
.Y(n_451)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_134),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_SL g134 ( 
.A(n_135),
.B(n_174),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_152),
.C(n_164),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_136),
.B(n_197),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_147),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_142),
.Y(n_137)
);

MAJx2_ASAP7_75t_L g193 ( 
.A(n_138),
.B(n_142),
.C(n_147),
.Y(n_193)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_146),
.Y(n_226)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_152),
.A2(n_153),
.B1(n_164),
.B2(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

MAJx2_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_157),
.C(n_160),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_154),
.A2(n_155),
.B1(n_160),
.B2(n_161),
.Y(n_278)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_157),
.B(n_278),
.Y(n_277)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx6_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_164),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_171),
.Y(n_164)
);

AND2x2_ASAP7_75t_L g192 ( 
.A(n_165),
.B(n_171),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_167),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_166),
.B(n_456),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_166),
.B(n_476),
.Y(n_475)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx8_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_170),
.Y(n_188)
);

BUFx3_ASAP7_75t_L g237 ( 
.A(n_170),
.Y(n_237)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

XOR2x1_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_191),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_175),
.B(n_192),
.C(n_193),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_181),
.Y(n_175)
);

MAJx2_ASAP7_75t_L g300 ( 
.A(n_176),
.B(n_186),
.C(n_189),
.Y(n_300)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_179),
.Y(n_480)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_182),
.A2(n_186),
.B1(n_189),
.B2(n_190),
.Y(n_181)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_182),
.Y(n_189)
);

INVx4_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx4_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_185),
.Y(n_355)
);

INVx3_ASAP7_75t_SL g456 ( 
.A(n_185),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_186),
.Y(n_190)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g390 ( 
.A(n_188),
.Y(n_390)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_193),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_199),
.C(n_209),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_196),
.B(n_283),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_199),
.B(n_209),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_201),
.C(n_203),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_200),
.B(n_201),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_203),
.B(n_271),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_204),
.B(n_207),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_204),
.B(n_207),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

OAI21x1_ASAP7_75t_L g211 ( 
.A1(n_212),
.A2(n_280),
.B(n_284),
.Y(n_211)
);

OA21x2_ASAP7_75t_L g212 ( 
.A1(n_213),
.A2(n_265),
.B(n_279),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_214),
.A2(n_249),
.B(n_264),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_215),
.A2(n_240),
.B(n_248),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_221),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_216),
.B(n_221),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_220),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_217),
.B(n_220),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_217),
.B(n_245),
.Y(n_244)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_222),
.A2(n_223),
.B1(n_232),
.B2(n_233),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_227),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_224),
.B(n_227),
.C(n_232),
.Y(n_263)
);

INVx4_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_229),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_229),
.B(n_256),
.Y(n_255)
);

INVx4_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx6_ASAP7_75t_L g310 ( 
.A(n_231),
.Y(n_310)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_SL g233 ( 
.A(n_234),
.B(n_238),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_234),
.B(n_238),
.Y(n_253)
);

INVx4_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_241),
.A2(n_244),
.B(n_247),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_242),
.B(n_243),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_242),
.B(n_243),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_250),
.B(n_263),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_250),
.B(n_263),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_254),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_253),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_252),
.B(n_253),
.C(n_267),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_254),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_SL g254 ( 
.A(n_255),
.B(n_257),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_255),
.B(n_260),
.C(n_262),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_258),
.A2(n_260),
.B1(n_261),
.B2(n_262),
.Y(n_257)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_258),
.Y(n_262)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_268),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_266),
.B(n_268),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_269),
.A2(n_270),
.B1(n_272),
.B2(n_273),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_269),
.B(n_275),
.C(n_276),
.Y(n_281)
);

INVx1_ASAP7_75t_SL g269 ( 
.A(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_274),
.A2(n_275),
.B1(n_276),
.B2(n_277),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx1_ASAP7_75t_SL g276 ( 
.A(n_277),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_282),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_281),
.B(n_282),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_287),
.B(n_325),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_287),
.B(n_325),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_302),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_290),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_289),
.B(n_290),
.C(n_302),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_291),
.A2(n_292),
.B1(n_299),
.B2(n_301),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_SL g292 ( 
.A(n_293),
.B(n_294),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_293),
.B(n_296),
.C(n_297),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_295),
.A2(n_296),
.B1(n_297),
.B2(n_298),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_296),
.Y(n_295)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_299),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_SL g302 ( 
.A(n_303),
.B(n_304),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_303),
.B(n_305),
.C(n_317),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_317),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_311),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_306),
.B(n_312),
.C(n_315),
.Y(n_361)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx6_ASAP7_75t_L g463 ( 
.A(n_310),
.Y(n_463)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_315),
.Y(n_311)
);

INVx6_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_324),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_321),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_319),
.B(n_321),
.C(n_324),
.Y(n_336)
);

BUFx2_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_329),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_328),
.B(n_329),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_331),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_330),
.B(n_347),
.C(n_375),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_332),
.A2(n_347),
.B1(n_375),
.B2(n_376),
.Y(n_331)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_332),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_333),
.A2(n_334),
.B1(n_335),
.B2(n_346),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_333),
.B(n_336),
.C(n_337),
.Y(n_380)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_335),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_SL g335 ( 
.A(n_336),
.B(n_337),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_345),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_339),
.B(n_342),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_339),
.B(n_342),
.C(n_345),
.Y(n_409)
);

INVx3_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

HB1xp67_ASAP7_75t_L g403 ( 
.A(n_341),
.Y(n_403)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_347),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_348),
.B(n_360),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_348),
.B(n_361),
.C(n_362),
.Y(n_407)
);

BUFx24_ASAP7_75t_SL g550 ( 
.A(n_348),
.Y(n_550)
);

FAx1_ASAP7_75t_SL g348 ( 
.A(n_349),
.B(n_353),
.CI(n_356),
.CON(n_348),
.SN(n_348)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_349),
.B(n_353),
.C(n_356),
.Y(n_419)
);

INVx5_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

INVx3_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

INVx5_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

INVx5_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_361),
.B(n_362),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_363),
.A2(n_364),
.B1(n_373),
.B2(n_374),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_365),
.A2(n_369),
.B1(n_371),
.B2(n_372),
.Y(n_364)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_365),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_365),
.B(n_372),
.C(n_373),
.Y(n_392)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_369),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_369),
.A2(n_372),
.B1(n_388),
.B2(n_389),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_372),
.B(n_385),
.C(n_389),
.Y(n_434)
);

CKINVDCx14_ASAP7_75t_R g373 ( 
.A(n_374),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_SL g378 ( 
.A(n_379),
.B(n_421),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_379),
.B(n_421),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_380),
.B(n_381),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_380),
.B(n_382),
.C(n_405),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_382),
.B(n_405),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_383),
.A2(n_384),
.B1(n_391),
.B2(n_404),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_383),
.B(n_392),
.C(n_393),
.Y(n_428)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_SL g384 ( 
.A(n_385),
.B(n_387),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g447 ( 
.A1(n_388),
.A2(n_389),
.B1(n_448),
.B2(n_449),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g514 ( 
.A(n_388),
.B(n_441),
.C(n_448),
.Y(n_514)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_391),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_SL g391 ( 
.A(n_392),
.B(n_393),
.Y(n_391)
);

XOR2xp5_ASAP7_75t_L g393 ( 
.A(n_394),
.B(n_401),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g394 ( 
.A(n_395),
.B(n_399),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_395),
.B(n_399),
.C(n_401),
.Y(n_453)
);

INVx4_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

INVx6_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_406),
.A2(n_407),
.B1(n_408),
.B2(n_420),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_406),
.B(n_409),
.C(n_410),
.Y(n_425)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_408),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_SL g408 ( 
.A(n_409),
.B(n_410),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_L g410 ( 
.A(n_411),
.B(n_419),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_412),
.A2(n_413),
.B1(n_417),
.B2(n_418),
.Y(n_411)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_412),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_413),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_413),
.B(n_417),
.C(n_432),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_L g435 ( 
.A1(n_413),
.A2(n_418),
.B1(n_436),
.B2(n_438),
.Y(n_435)
);

INVx5_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

INVx6_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_418),
.B(n_434),
.C(n_438),
.Y(n_487)
);

INVxp67_ASAP7_75t_L g432 ( 
.A(n_419),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_SL g423 ( 
.A(n_424),
.B(n_465),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_424),
.B(n_465),
.Y(n_466)
);

BUFx24_ASAP7_75t_SL g551 ( 
.A(n_424),
.Y(n_551)
);

FAx1_ASAP7_75t_SL g424 ( 
.A(n_425),
.B(n_426),
.CI(n_439),
.CON(n_424),
.SN(n_424)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_425),
.B(n_426),
.C(n_439),
.Y(n_526)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_427),
.A2(n_428),
.B1(n_429),
.B2(n_430),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_427),
.B(n_431),
.C(n_433),
.Y(n_522)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

XOR2xp5_ASAP7_75t_L g430 ( 
.A(n_431),
.B(n_433),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_L g433 ( 
.A(n_434),
.B(n_435),
.Y(n_433)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_436),
.Y(n_438)
);

XOR2xp5_ASAP7_75t_L g439 ( 
.A(n_440),
.B(n_452),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_440),
.B(n_453),
.C(n_454),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_441),
.B(n_447),
.Y(n_440)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

INVx3_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

BUFx2_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);

INVx6_ASAP7_75t_L g445 ( 
.A(n_446),
.Y(n_445)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_446),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_448),
.B(n_492),
.C(n_495),
.Y(n_491)
);

CKINVDCx16_ASAP7_75t_R g448 ( 
.A(n_449),
.Y(n_448)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_451),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_L g452 ( 
.A(n_453),
.B(n_454),
.Y(n_452)
);

XNOR2xp5_ASAP7_75t_SL g454 ( 
.A(n_455),
.B(n_457),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_455),
.B(n_459),
.C(n_464),
.Y(n_515)
);

AOI22xp5_ASAP7_75t_L g457 ( 
.A1(n_458),
.A2(n_459),
.B1(n_460),
.B2(n_464),
.Y(n_457)
);

CKINVDCx14_ASAP7_75t_R g464 ( 
.A(n_458),
.Y(n_464)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_460),
.Y(n_459)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_462),
.Y(n_461)
);

INVx3_ASAP7_75t_L g462 ( 
.A(n_463),
.Y(n_462)
);

NOR3xp33_ASAP7_75t_L g467 ( 
.A(n_468),
.B(n_527),
.C(n_537),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_469),
.B(n_523),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_470),
.Y(n_469)
);

OAI21xp5_ASAP7_75t_L g545 ( 
.A1(n_470),
.A2(n_546),
.B(n_547),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_SL g470 ( 
.A(n_471),
.B(n_516),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_471),
.B(n_516),
.Y(n_547)
);

XOR2xp5_ASAP7_75t_L g471 ( 
.A(n_472),
.B(n_488),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g529 ( 
.A(n_472),
.B(n_489),
.C(n_511),
.Y(n_529)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_473),
.B(n_474),
.C(n_486),
.Y(n_472)
);

XNOR2xp5_ASAP7_75t_SL g517 ( 
.A(n_473),
.B(n_518),
.Y(n_517)
);

AOI22xp5_ASAP7_75t_L g518 ( 
.A1(n_474),
.A2(n_486),
.B1(n_487),
.B2(n_519),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_474),
.Y(n_519)
);

XNOR2xp5_ASAP7_75t_L g474 ( 
.A(n_475),
.B(n_478),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_475),
.B(n_479),
.C(n_481),
.Y(n_502)
);

INVx3_ASAP7_75t_L g476 ( 
.A(n_477),
.Y(n_476)
);

XNOR2xp5_ASAP7_75t_L g478 ( 
.A(n_479),
.B(n_481),
.Y(n_478)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_483),
.Y(n_482)
);

HB1xp67_ASAP7_75t_L g483 ( 
.A(n_484),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_485),
.Y(n_484)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_487),
.Y(n_486)
);

XOR2xp5_ASAP7_75t_L g488 ( 
.A(n_489),
.B(n_511),
.Y(n_488)
);

XNOR2xp5_ASAP7_75t_L g489 ( 
.A(n_490),
.B(n_501),
.Y(n_489)
);

AOI22xp5_ASAP7_75t_L g490 ( 
.A1(n_491),
.A2(n_496),
.B1(n_499),
.B2(n_500),
.Y(n_490)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_491),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g531 ( 
.A(n_491),
.B(n_500),
.C(n_501),
.Y(n_531)
);

XOR2xp5_ASAP7_75t_L g512 ( 
.A(n_492),
.B(n_513),
.Y(n_512)
);

INVx6_ASAP7_75t_L g493 ( 
.A(n_494),
.Y(n_493)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_496),
.Y(n_500)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_498),
.Y(n_497)
);

XNOR2xp5_ASAP7_75t_SL g501 ( 
.A(n_502),
.B(n_503),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g533 ( 
.A(n_502),
.B(n_505),
.C(n_510),
.Y(n_533)
);

AOI22xp5_ASAP7_75t_L g503 ( 
.A1(n_504),
.A2(n_505),
.B1(n_506),
.B2(n_510),
.Y(n_503)
);

CKINVDCx16_ASAP7_75t_R g510 ( 
.A(n_504),
.Y(n_510)
);

CKINVDCx16_ASAP7_75t_R g505 ( 
.A(n_506),
.Y(n_505)
);

INVx8_ASAP7_75t_L g507 ( 
.A(n_508),
.Y(n_507)
);

INVx4_ASAP7_75t_L g508 ( 
.A(n_509),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_512),
.B(n_514),
.C(n_515),
.Y(n_511)
);

XNOR2xp5_ASAP7_75t_L g520 ( 
.A(n_512),
.B(n_521),
.Y(n_520)
);

XNOR2xp5_ASAP7_75t_L g521 ( 
.A(n_514),
.B(n_515),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_517),
.B(n_520),
.C(n_522),
.Y(n_516)
);

XOR2xp5_ASAP7_75t_L g525 ( 
.A(n_517),
.B(n_520),
.Y(n_525)
);

XNOR2xp5_ASAP7_75t_L g524 ( 
.A(n_522),
.B(n_525),
.Y(n_524)
);

OR2x2_ASAP7_75t_L g523 ( 
.A(n_524),
.B(n_526),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_524),
.B(n_526),
.Y(n_546)
);

INVxp67_ASAP7_75t_L g527 ( 
.A(n_528),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_528),
.B(n_545),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_529),
.B(n_530),
.Y(n_528)
);

OR2x2_ASAP7_75t_L g543 ( 
.A(n_529),
.B(n_530),
.Y(n_543)
);

XNOR2xp5_ASAP7_75t_L g530 ( 
.A(n_531),
.B(n_532),
.Y(n_530)
);

MAJIxp5_ASAP7_75t_L g541 ( 
.A(n_531),
.B(n_533),
.C(n_534),
.Y(n_541)
);

XNOR2xp5_ASAP7_75t_L g532 ( 
.A(n_533),
.B(n_534),
.Y(n_532)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_536),
.Y(n_535)
);

A2O1A1Ixp33_ASAP7_75t_L g542 ( 
.A1(n_537),
.A2(n_543),
.B(n_544),
.C(n_548),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_538),
.B(n_541),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_538),
.B(n_541),
.Y(n_548)
);


endmodule