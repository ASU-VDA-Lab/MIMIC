module fake_jpeg_1025_n_124 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_124);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_124;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_93;
wire n_54;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_10),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_9),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_7),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

BUFx8_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx2_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_25),
.Y(n_27)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_27),
.Y(n_64)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_28),
.Y(n_65)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_29),
.Y(n_60)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_30),
.Y(n_69)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_31),
.B(n_34),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

INVx13_ASAP7_75t_L g62 ( 
.A(n_32),
.Y(n_62)
);

OR2x2_ASAP7_75t_L g33 ( 
.A(n_22),
.B(n_0),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_33),
.B(n_37),
.Y(n_72)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_23),
.A2(n_8),
.B1(n_3),
.B2(n_4),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_35),
.A2(n_5),
.B1(n_16),
.B2(n_42),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_36),
.Y(n_54)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_26),
.B(n_1),
.Y(n_38)
);

NOR2x1_ASAP7_75t_L g67 ( 
.A(n_38),
.B(n_44),
.Y(n_67)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_11),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_39),
.B(n_40),
.Y(n_73)
);

INVx2_ASAP7_75t_SL g40 ( 
.A(n_11),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_12),
.B(n_8),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_41),
.B(n_43),
.Y(n_55)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_42),
.A2(n_48),
.B1(n_50),
.B2(n_17),
.Y(n_58)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_22),
.B(n_3),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_45),
.B(n_46),
.Y(n_59)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_15),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_24),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_47),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_24),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_12),
.B(n_4),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_49),
.B(n_51),
.Y(n_63)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_22),
.Y(n_50)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_19),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_14),
.B(n_4),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_52),
.B(n_41),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_47),
.A2(n_19),
.B1(n_20),
.B2(n_21),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_53),
.A2(n_57),
.B1(n_70),
.B2(n_71),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_45),
.A2(n_21),
.B1(n_20),
.B2(n_15),
.Y(n_57)
);

BUFx2_ASAP7_75t_SL g86 ( 
.A(n_58),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_40),
.B(n_33),
.C(n_52),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_61),
.B(n_66),
.Y(n_82)
);

OA22x2_ASAP7_75t_L g70 ( 
.A1(n_50),
.A2(n_5),
.B1(n_6),
.B2(n_14),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_72),
.B(n_16),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_74),
.B(n_75),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_63),
.B(n_32),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_55),
.B(n_32),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_76),
.B(n_77),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_63),
.B(n_5),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_59),
.B(n_55),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_78),
.B(n_80),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_66),
.B(n_61),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_79),
.B(n_83),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_59),
.B(n_73),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_56),
.Y(n_81)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_81),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_67),
.B(n_57),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_67),
.B(n_60),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_84),
.B(n_87),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_60),
.B(n_64),
.Y(n_87)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_81),
.Y(n_90)
);

HB1xp67_ASAP7_75t_L g99 ( 
.A(n_90),
.Y(n_99)
);

OAI32xp33_ASAP7_75t_L g93 ( 
.A1(n_78),
.A2(n_83),
.A3(n_82),
.B1(n_80),
.B2(n_85),
.Y(n_93)
);

AOI221xp5_ASAP7_75t_L g102 ( 
.A1(n_93),
.A2(n_56),
.B1(n_64),
.B2(n_68),
.C(n_69),
.Y(n_102)
);

CKINVDCx14_ASAP7_75t_R g94 ( 
.A(n_85),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_94),
.B(n_70),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g95 ( 
.A1(n_82),
.A2(n_53),
.B(n_70),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g104 ( 
.A1(n_95),
.A2(n_65),
.B(n_62),
.Y(n_104)
);

INVx1_ASAP7_75t_SL g106 ( 
.A(n_98),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_92),
.A2(n_86),
.B1(n_70),
.B2(n_54),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_100),
.A2(n_101),
.B(n_104),
.Y(n_108)
);

XNOR2x1_ASAP7_75t_SL g101 ( 
.A(n_91),
.B(n_56),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_102),
.B(n_103),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_97),
.B(n_69),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_97),
.B(n_65),
.Y(n_105)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_105),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_101),
.B(n_91),
.C(n_96),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_107),
.B(n_96),
.C(n_109),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_111),
.B(n_113),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_108),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_112),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_107),
.B(n_88),
.C(n_92),
.Y(n_113)
);

A2O1A1Ixp33_ASAP7_75t_SL g114 ( 
.A1(n_110),
.A2(n_104),
.B(n_100),
.C(n_95),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_114),
.A2(n_106),
.B1(n_93),
.B2(n_99),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_116),
.Y(n_119)
);

AOI322xp5_ASAP7_75t_L g118 ( 
.A1(n_117),
.A2(n_62),
.A3(n_88),
.B1(n_89),
.B2(n_90),
.C1(n_106),
.C2(n_115),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_118),
.A2(n_117),
.B(n_115),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_120),
.B(n_121),
.C(n_116),
.Y(n_122)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_119),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_122),
.Y(n_123)
);

OR2x2_ASAP7_75t_L g124 ( 
.A(n_123),
.B(n_89),
.Y(n_124)
);


endmodule