module fake_jpeg_863_n_230 (n_13, n_21, n_53, n_33, n_54, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_230);

input n_13;
input n_21;
input n_53;
input n_33;
input n_54;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_230;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_223;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_12),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

BUFx4f_ASAP7_75t_L g58 ( 
.A(n_32),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_54),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_52),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_53),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_21),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

INVx11_ASAP7_75t_SL g66 ( 
.A(n_5),
.Y(n_66)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_19),
.Y(n_67)
);

INVx1_ASAP7_75t_SL g68 ( 
.A(n_51),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_38),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_18),
.Y(n_70)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_50),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_27),
.Y(n_72)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_20),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_9),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_14),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_5),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_12),
.Y(n_77)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_6),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_31),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_39),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_47),
.Y(n_81)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_66),
.Y(n_82)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_82),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_74),
.B(n_49),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_83),
.B(n_88),
.Y(n_100)
);

BUFx12f_ASAP7_75t_L g84 ( 
.A(n_66),
.Y(n_84)
);

BUFx4f_ASAP7_75t_SL g99 ( 
.A(n_84),
.Y(n_99)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_71),
.Y(n_85)
);

INVx8_ASAP7_75t_L g102 ( 
.A(n_85),
.Y(n_102)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_73),
.Y(n_86)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_86),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_60),
.Y(n_87)
);

CKINVDCx6p67_ASAP7_75t_R g101 ( 
.A(n_87),
.Y(n_101)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_73),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_78),
.A2(n_45),
.B1(n_44),
.B2(n_43),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_89),
.B(n_0),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_67),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_90),
.B(n_69),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_82),
.A2(n_78),
.B1(n_67),
.B2(n_76),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_91),
.A2(n_96),
.B1(n_84),
.B2(n_68),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_94),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_95),
.B(n_97),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_86),
.A2(n_76),
.B1(n_70),
.B2(n_77),
.Y(n_96)
);

OR2x2_ASAP7_75t_L g97 ( 
.A(n_88),
.B(n_75),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_83),
.B(n_56),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_98),
.B(n_58),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_90),
.B(n_55),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_103),
.B(n_80),
.Y(n_122)
);

OR2x2_ASAP7_75t_L g104 ( 
.A(n_100),
.B(n_97),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_104),
.B(n_111),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_105),
.B(n_106),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_98),
.B(n_64),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_100),
.B(n_65),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_107),
.B(n_119),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_95),
.A2(n_87),
.B1(n_89),
.B2(n_85),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_109),
.A2(n_114),
.B1(n_116),
.B2(n_118),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_93),
.B(n_79),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_93),
.B(n_59),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_112),
.B(n_117),
.Y(n_139)
);

INVx13_ASAP7_75t_L g113 ( 
.A(n_99),
.Y(n_113)
);

INVx1_ASAP7_75t_SL g129 ( 
.A(n_113),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_101),
.A2(n_71),
.B1(n_57),
.B2(n_58),
.Y(n_114)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_101),
.Y(n_115)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_115),
.Y(n_124)
);

A2O1A1Ixp33_ASAP7_75t_L g117 ( 
.A1(n_101),
.A2(n_72),
.B(n_68),
.C(n_61),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_101),
.A2(n_57),
.B1(n_81),
.B2(n_62),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_92),
.B(n_60),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_92),
.B(n_63),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_120),
.B(n_121),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_99),
.B(n_63),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_122),
.B(n_99),
.Y(n_140)
);

INVx2_ASAP7_75t_SL g123 ( 
.A(n_102),
.Y(n_123)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_123),
.Y(n_135)
);

INVx13_ASAP7_75t_L g125 ( 
.A(n_113),
.Y(n_125)
);

INVx1_ASAP7_75t_SL g148 ( 
.A(n_125),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_110),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_128),
.B(n_130),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_110),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_119),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_131),
.B(n_136),
.Y(n_169)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_115),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g150 ( 
.A(n_132),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_123),
.Y(n_133)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_133),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_107),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_140),
.B(n_143),
.Y(n_147)
);

INVx13_ASAP7_75t_L g141 ( 
.A(n_123),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_141),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_105),
.B(n_80),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_142),
.B(n_40),
.Y(n_151)
);

AND2x6_ASAP7_75t_L g143 ( 
.A(n_104),
.B(n_42),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_117),
.A2(n_84),
.B(n_102),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_144),
.A2(n_37),
.B(n_36),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_109),
.A2(n_61),
.B1(n_81),
.B2(n_62),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_145),
.B(n_26),
.Y(n_156)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_118),
.Y(n_146)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_146),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_126),
.A2(n_108),
.B1(n_1),
.B2(n_2),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_149),
.A2(n_156),
.B1(n_11),
.B2(n_13),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_151),
.B(n_166),
.Y(n_186)
);

NAND2x1_ASAP7_75t_L g177 ( 
.A(n_152),
.B(n_25),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_126),
.B(n_33),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_153),
.B(n_6),
.C(n_7),
.Y(n_182)
);

AO22x1_ASAP7_75t_SL g154 ( 
.A1(n_134),
.A2(n_30),
.B1(n_29),
.B2(n_28),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_154),
.B(n_158),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_137),
.B(n_0),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_124),
.Y(n_159)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_159),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_144),
.A2(n_1),
.B(n_2),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_160),
.A2(n_3),
.B(n_4),
.Y(n_176)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_124),
.Y(n_162)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_162),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_135),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_163),
.B(n_164),
.Y(n_179)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_135),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_139),
.A2(n_3),
.B(n_4),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_165),
.A2(n_168),
.B(n_170),
.Y(n_172)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_132),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_133),
.Y(n_168)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_129),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_125),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_171),
.A2(n_129),
.B(n_127),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_173),
.B(n_177),
.Y(n_201)
);

OAI32xp33_ASAP7_75t_L g174 ( 
.A1(n_169),
.A2(n_138),
.A3(n_143),
.B1(n_141),
.B2(n_7),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_174),
.B(n_176),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_167),
.B(n_24),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_178),
.B(n_183),
.C(n_188),
.Y(n_193)
);

OR2x6_ASAP7_75t_SL g180 ( 
.A(n_155),
.B(n_23),
.Y(n_180)
);

HB1xp67_ASAP7_75t_SL g192 ( 
.A(n_180),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_182),
.B(n_189),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_163),
.B(n_154),
.C(n_161),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_147),
.A2(n_22),
.B(n_9),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_184),
.A2(n_187),
.B(n_15),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_156),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_185),
.A2(n_191),
.B1(n_13),
.B2(n_14),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_165),
.A2(n_148),
.B(n_154),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_148),
.B(n_20),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_150),
.B(n_8),
.C(n_10),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_183),
.A2(n_168),
.B1(n_157),
.B2(n_150),
.Y(n_195)
);

OAI21xp33_ASAP7_75t_SL g206 ( 
.A1(n_195),
.A2(n_180),
.B(n_188),
.Y(n_206)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_175),
.Y(n_196)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_196),
.Y(n_209)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_181),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_197),
.B(n_199),
.Y(n_205)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_179),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_200),
.B(n_203),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_202),
.Y(n_204)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_172),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_206),
.B(n_211),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_193),
.B(n_186),
.C(n_178),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_207),
.B(n_208),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_193),
.B(n_190),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_201),
.A2(n_198),
.B(n_195),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_194),
.B(n_177),
.Y(n_212)
);

BUFx2_ASAP7_75t_L g216 ( 
.A(n_212),
.Y(n_216)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_205),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g220 ( 
.A(n_213),
.Y(n_220)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_209),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_217),
.A2(n_218),
.B(n_206),
.Y(n_221)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_210),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_214),
.A2(n_204),
.B(n_202),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_219),
.B(n_216),
.Y(n_223)
);

NOR2xp67_ASAP7_75t_L g222 ( 
.A(n_221),
.B(n_214),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_222),
.A2(n_223),
.B(n_192),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_224),
.B(n_220),
.C(n_215),
.Y(n_225)
);

AOI322xp5_ASAP7_75t_L g226 ( 
.A1(n_225),
.A2(n_180),
.A3(n_194),
.B1(n_182),
.B2(n_189),
.C1(n_15),
.C2(n_18),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_226),
.A2(n_16),
.B(n_17),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_227),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_228),
.A2(n_19),
.B(n_16),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_229),
.B(n_17),
.Y(n_230)
);


endmodule