module real_jpeg_32605_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_598, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_598;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_574;
wire n_595;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_578;
wire n_456;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_128;
wire n_202;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_393;
wire n_221;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_214;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_593;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_590;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_592;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_559;
wire n_232;
wire n_582;
wire n_448;
wire n_212;
wire n_284;
wire n_579;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_583;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_589;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_215;
wire n_176;
wire n_166;
wire n_323;
wire n_596;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_594;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_572;
wire n_586;
wire n_548;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_531;
wire n_546;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_18;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_575;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_584;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_585;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_581;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_587;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_588;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_568;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_447;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_591;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

BUFx3_ASAP7_75t_L g135 ( 
.A(n_0),
.Y(n_135)
);

BUFx12f_ASAP7_75t_L g138 ( 
.A(n_0),
.Y(n_138)
);

HB1xp67_ASAP7_75t_L g204 ( 
.A(n_0),
.Y(n_204)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_0),
.Y(n_288)
);

BUFx6f_ASAP7_75t_L g335 ( 
.A(n_0),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_1),
.A2(n_68),
.B1(n_74),
.B2(n_79),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_1),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_1),
.A2(n_79),
.B1(n_207),
.B2(n_211),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_1),
.A2(n_79),
.B1(n_240),
.B2(n_243),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_1),
.A2(n_79),
.B1(n_290),
.B2(n_292),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_2),
.B(n_189),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_2),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_2),
.B(n_367),
.Y(n_375)
);

AOI22xp33_ASAP7_75t_SL g421 ( 
.A1(n_2),
.A2(n_315),
.B1(n_422),
.B2(n_425),
.Y(n_421)
);

OAI21xp33_ASAP7_75t_L g500 ( 
.A1(n_2),
.A2(n_201),
.B(n_447),
.Y(n_500)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_3),
.A2(n_178),
.B1(n_186),
.B2(n_187),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_3),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_3),
.A2(n_186),
.B1(n_216),
.B2(n_220),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_3),
.A2(n_186),
.B1(n_281),
.B2(n_283),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_3),
.A2(n_186),
.B1(n_394),
.B2(n_395),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_4),
.A2(n_109),
.B1(n_272),
.B2(n_273),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_4),
.Y(n_272)
);

AOI22xp33_ASAP7_75t_L g412 ( 
.A1(n_4),
.A2(n_272),
.B1(n_413),
.B2(n_417),
.Y(n_412)
);

AOI22xp33_ASAP7_75t_SL g458 ( 
.A1(n_4),
.A2(n_272),
.B1(n_459),
.B2(n_463),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_L g535 ( 
.A1(n_4),
.A2(n_272),
.B1(n_536),
.B2(n_539),
.Y(n_535)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_5),
.Y(n_166)
);

BUFx3_ASAP7_75t_L g175 ( 
.A(n_5),
.Y(n_175)
);

BUFx3_ASAP7_75t_L g179 ( 
.A(n_5),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_6),
.Y(n_85)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_6),
.Y(n_90)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_7),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_7),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g341 ( 
.A(n_7),
.Y(n_341)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_8),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_8),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g302 ( 
.A(n_8),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_9),
.A2(n_177),
.B1(n_180),
.B2(n_181),
.Y(n_176)
);

INVx1_ASAP7_75t_SL g180 ( 
.A(n_9),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_9),
.A2(n_74),
.B1(n_180),
.B2(n_253),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_9),
.A2(n_180),
.B1(n_308),
.B2(n_311),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_9),
.A2(n_180),
.B1(n_338),
.B2(n_342),
.Y(n_337)
);

AO22x1_ASAP7_75t_L g23 ( 
.A1(n_10),
.A2(n_24),
.B1(n_28),
.B2(n_29),
.Y(n_23)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_10),
.A2(n_28),
.B1(n_250),
.B2(n_252),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_11),
.Y(n_155)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_11),
.Y(n_383)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_12),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_13),
.A2(n_228),
.B1(n_229),
.B2(n_233),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_13),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_SL g297 ( 
.A1(n_13),
.A2(n_228),
.B1(n_298),
.B2(n_303),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g399 ( 
.A1(n_13),
.A2(n_228),
.B1(n_400),
.B2(n_401),
.Y(n_399)
);

AOI22xp33_ASAP7_75t_SL g440 ( 
.A1(n_13),
.A2(n_228),
.B1(n_441),
.B2(n_442),
.Y(n_440)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_14),
.Y(n_73)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_14),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_14),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_14),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_15),
.A2(n_109),
.B1(n_113),
.B2(n_114),
.Y(n_108)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_15),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_15),
.A2(n_61),
.B1(n_113),
.B2(n_127),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g358 ( 
.A1(n_15),
.A2(n_113),
.B1(n_359),
.B2(n_363),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_16),
.A2(n_57),
.B1(n_60),
.B2(n_61),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_16),
.Y(n_60)
);

AO22x1_ASAP7_75t_SL g141 ( 
.A1(n_16),
.A2(n_60),
.B1(n_142),
.B2(n_145),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_261),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_260),
.Y(n_18)
);

OR2x2_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_236),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_20),
.B(n_236),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_122),
.C(n_190),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g554 ( 
.A(n_21),
.B(n_191),
.Y(n_554)
);

OAI21xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_66),
.B(n_121),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_22),
.B(n_66),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_32),
.B1(n_56),
.B2(n_65),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_23),
.B(n_65),
.Y(n_124)
);

INVx1_ASAP7_75t_SL g24 ( 
.A(n_25),
.Y(n_24)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_25),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_26),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g310 ( 
.A(n_27),
.Y(n_310)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_27),
.Y(n_416)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_28),
.A2(n_196),
.B(n_199),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_28),
.B(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_SL g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx2_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_31),
.A2(n_49),
.B1(n_52),
.B2(n_54),
.Y(n_48)
);

OA21x2_ASAP7_75t_L g247 ( 
.A1(n_32),
.A2(n_56),
.B(n_65),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_SL g391 ( 
.A1(n_32),
.A2(n_65),
.B1(n_307),
.B2(n_392),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_32),
.B(n_307),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_32),
.B(n_494),
.Y(n_493)
);

INVx2_ASAP7_75t_SL g32 ( 
.A(n_33),
.Y(n_32)
);

OR2x2_ASAP7_75t_L g125 ( 
.A(n_33),
.B(n_126),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_33),
.A2(n_126),
.B1(n_206),
.B2(n_212),
.Y(n_205)
);

BUFx2_ASAP7_75t_L g296 ( 
.A(n_33),
.Y(n_296)
);

OA22x2_ASAP7_75t_L g528 ( 
.A1(n_33),
.A2(n_206),
.B1(n_212),
.B2(n_393),
.Y(n_528)
);

OR2x2_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_48),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_34),
.Y(n_65)
);

OAI22x1_ASAP7_75t_L g34 ( 
.A1(n_35),
.A2(n_39),
.B1(n_42),
.B2(n_44),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_39),
.Y(n_200)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g285 ( 
.A(n_40),
.Y(n_285)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_41),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_41),
.Y(n_140)
);

INVx3_ASAP7_75t_L g362 ( 
.A(n_41),
.Y(n_362)
);

BUFx6f_ASAP7_75t_L g446 ( 
.A(n_41),
.Y(n_446)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_41),
.Y(n_508)
);

BUFx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx3_ASAP7_75t_L g291 ( 
.A(n_43),
.Y(n_291)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_45),
.Y(n_479)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_50),
.Y(n_59)
);

INVx4_ASAP7_75t_L g305 ( 
.A(n_50),
.Y(n_305)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_51),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_51),
.Y(n_131)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx4_ASAP7_75t_L g311 ( 
.A(n_57),
.Y(n_311)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx4_ASAP7_75t_SL g61 ( 
.A(n_62),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_62),
.B(n_315),
.Y(n_481)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx2_ASAP7_75t_SL g87 ( 
.A(n_64),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g319 ( 
.A(n_64),
.Y(n_319)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_65),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_65),
.B(n_307),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_67),
.A2(n_80),
.B1(n_108),
.B2(n_118),
.Y(n_66)
);

AOI22x1_ASAP7_75t_L g214 ( 
.A1(n_67),
.A2(n_80),
.B1(n_120),
.B2(n_215),
.Y(n_214)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVxp67_ASAP7_75t_SL g69 ( 
.A(n_70),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_72),
.Y(n_107)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_73),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_73),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_73),
.Y(n_222)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_77),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g317 ( 
.A(n_77),
.Y(n_317)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_78),
.Y(n_161)
);

BUFx5_ASAP7_75t_L g428 ( 
.A(n_78),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_80),
.A2(n_108),
.B1(n_118),
.B2(n_249),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_80),
.B(n_276),
.Y(n_275)
);

AOI22x1_ASAP7_75t_L g397 ( 
.A1(n_80),
.A2(n_118),
.B1(n_271),
.B2(n_398),
.Y(n_397)
);

INVx2_ASAP7_75t_SL g420 ( 
.A(n_80),
.Y(n_420)
);

AND2x4_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_94),
.Y(n_80)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_81),
.Y(n_120)
);

AOI22x1_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_86),
.B1(n_88),
.B2(n_91),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_85),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g331 ( 
.A(n_85),
.Y(n_331)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_90),
.Y(n_102)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g418 ( 
.A(n_93),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_95),
.A2(n_99),
.B1(n_103),
.B2(n_107),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

BUFx2_ASAP7_75t_L g402 ( 
.A(n_97),
.Y(n_402)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx3_ASAP7_75t_L g424 ( 
.A(n_98),
.Y(n_424)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_110),
.Y(n_400)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx8_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_112),
.Y(n_274)
);

BUFx6f_ASAP7_75t_L g379 ( 
.A(n_112),
.Y(n_379)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_116),
.Y(n_254)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_117),
.Y(n_327)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_119),
.A2(n_270),
.B(n_275),
.Y(n_269)
);

OR2x2_ASAP7_75t_L g450 ( 
.A(n_119),
.B(n_315),
.Y(n_450)
);

OAI22x1_ASAP7_75t_L g542 ( 
.A1(n_119),
.A2(n_420),
.B1(n_543),
.B2(n_544),
.Y(n_542)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_120),
.B(n_276),
.Y(n_429)
);

HB1xp67_ASAP7_75t_L g257 ( 
.A(n_121),
.Y(n_257)
);

XNOR2x1_ASAP7_75t_L g553 ( 
.A(n_122),
.B(n_554),
.Y(n_553)
);

XOR2x2_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_148),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g256 ( 
.A1(n_123),
.A2(n_132),
.B(n_150),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_124),
.A2(n_125),
.B(n_132),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_124),
.B(n_125),
.Y(n_548)
);

BUFx3_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_131),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_132),
.A2(n_133),
.B1(n_149),
.B2(n_150),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g546 ( 
.A1(n_132),
.A2(n_133),
.B1(n_547),
.B2(n_548),
.Y(n_546)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_133),
.Y(n_132)
);

OA21x2_ASAP7_75t_L g133 ( 
.A1(n_134),
.A2(n_136),
.B(n_141),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx5_ASAP7_75t_L g357 ( 
.A(n_135),
.Y(n_357)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_136),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_136),
.B(n_337),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_136),
.A2(n_355),
.B1(n_356),
.B2(n_358),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g456 ( 
.A1(n_136),
.A2(n_457),
.B1(n_466),
.B2(n_468),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_136),
.B(n_358),
.Y(n_533)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_139),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g467 ( 
.A(n_137),
.Y(n_467)
);

INVx8_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx4_ASAP7_75t_SL g449 ( 
.A(n_138),
.Y(n_449)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx6_ASAP7_75t_L g364 ( 
.A(n_140),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_141),
.B(n_203),
.Y(n_202)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_145),
.Y(n_475)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx4_ASAP7_75t_L g198 ( 
.A(n_146),
.Y(n_198)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

BUFx2_ASAP7_75t_L g282 ( 
.A(n_147),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_147),
.Y(n_293)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_147),
.Y(n_462)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_151),
.B(n_184),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g566 ( 
.A(n_151),
.B(n_567),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_152),
.B(n_176),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_152),
.B(n_227),
.Y(n_226)
);

BUFx2_ASAP7_75t_L g245 ( 
.A(n_152),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g385 ( 
.A1(n_152),
.A2(n_386),
.B(n_389),
.Y(n_385)
);

AO22x1_ASAP7_75t_SL g534 ( 
.A1(n_152),
.A2(n_189),
.B1(n_227),
.B2(n_535),
.Y(n_534)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_162),
.Y(n_152)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_153),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_156),
.B1(n_158),
.B2(n_160),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_155),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_155),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_155),
.Y(n_170)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_159),
.Y(n_371)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_163),
.A2(n_167),
.B1(n_169),
.B2(n_171),
.Y(n_162)
);

BUFx2_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_166),
.Y(n_188)
);

INVx6_ASAP7_75t_L g232 ( 
.A(n_166),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_166),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_166),
.Y(n_242)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx6_ASAP7_75t_L g183 ( 
.A(n_174),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_176),
.B(n_189),
.Y(n_225)
);

INVx2_ASAP7_75t_SL g243 ( 
.A(n_177),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

BUFx3_ASAP7_75t_L g538 ( 
.A(n_179),
.Y(n_538)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_189),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_185),
.A2(n_239),
.B1(n_244),
.B2(n_245),
.Y(n_238)
);

INVx2_ASAP7_75t_SL g187 ( 
.A(n_188),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g387 ( 
.A(n_188),
.Y(n_387)
);

HB1xp67_ASAP7_75t_L g244 ( 
.A(n_189),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_189),
.B(n_535),
.Y(n_567)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_213),
.C(n_223),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g550 ( 
.A(n_193),
.B(n_551),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_205),
.Y(n_193)
);

XOR2x2_ASAP7_75t_L g560 ( 
.A(n_194),
.B(n_561),
.Y(n_560)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_195),
.A2(n_201),
.B(n_202),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g529 ( 
.A1(n_195),
.A2(n_530),
.B(n_533),
.Y(n_529)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_196),
.Y(n_441)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx4_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_201),
.A2(n_280),
.B1(n_286),
.B2(n_289),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_L g439 ( 
.A1(n_201),
.A2(n_440),
.B(n_447),
.Y(n_439)
);

BUFx4f_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

HB1xp67_ASAP7_75t_L g561 ( 
.A(n_205),
.Y(n_561)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

BUFx3_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g411 ( 
.A1(n_212),
.A2(n_296),
.B1(n_297),
.B2(n_412),
.Y(n_411)
);

OAI21xp5_ASAP7_75t_L g452 ( 
.A1(n_212),
.A2(n_412),
.B(n_453),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_SL g497 ( 
.A(n_212),
.B(n_315),
.Y(n_497)
);

INVxp33_ASAP7_75t_SL g213 ( 
.A(n_214),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g551 ( 
.A(n_214),
.B(n_224),
.Y(n_551)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_215),
.Y(n_544)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx2_ASAP7_75t_SL g251 ( 
.A(n_219),
.Y(n_251)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_219),
.Y(n_374)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

HB1xp67_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_226),
.Y(n_224)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_225),
.Y(n_389)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx3_ASAP7_75t_L g368 ( 
.A(n_232),
.Y(n_368)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

BUFx4f_ASAP7_75t_SL g234 ( 
.A(n_235),
.Y(n_234)
);

BUFx12f_ASAP7_75t_L g540 ( 
.A(n_235),
.Y(n_540)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_255),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_246),
.Y(n_237)
);

INVx5_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx4_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_248),
.Y(n_246)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

HB1xp67_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_256),
.A2(n_257),
.B1(n_258),
.B2(n_259),
.Y(n_255)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_256),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_257),
.Y(n_259)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

NAND2x1p5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_588),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_521),
.Y(n_263)
);

OAI21x1_ASAP7_75t_L g264 ( 
.A1(n_265),
.A2(n_403),
.B(n_519),
.Y(n_264)
);

AND2x2_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_345),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_267),
.B(n_520),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_294),
.C(n_312),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_SL g405 ( 
.A(n_268),
.B(n_406),
.Y(n_405)
);

XOR2xp5_ASAP7_75t_SL g268 ( 
.A(n_269),
.B(n_277),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g348 ( 
.A1(n_269),
.A2(n_349),
.B(n_351),
.Y(n_348)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx8_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_276),
.Y(n_543)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_279),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_SL g349 ( 
.A(n_278),
.B(n_350),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_278),
.B(n_350),
.Y(n_351)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_279),
.Y(n_350)
);

OAI21xp5_ASAP7_75t_L g332 ( 
.A1(n_280),
.A2(n_333),
.B(n_336),
.Y(n_332)
);

INVx2_ASAP7_75t_SL g281 ( 
.A(n_282),
.Y(n_281)
);

INVx1_ASAP7_75t_SL g283 ( 
.A(n_284),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx2_ASAP7_75t_SL g505 ( 
.A(n_287),
.Y(n_505)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_289),
.Y(n_355)
);

HB1xp67_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

BUFx2_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g406 ( 
.A1(n_294),
.A2(n_295),
.B1(n_312),
.B2(n_407),
.Y(n_406)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

OAI21xp33_ASAP7_75t_SL g295 ( 
.A1(n_296),
.A2(n_297),
.B(n_306),
.Y(n_295)
);

INVx1_ASAP7_75t_SL g298 ( 
.A(n_299),
.Y(n_298)
);

OAI21xp33_ASAP7_75t_SL g494 ( 
.A1(n_299),
.A2(n_315),
.B(n_481),
.Y(n_494)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx4_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

BUFx6f_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

BUFx6f_ASAP7_75t_L g491 ( 
.A(n_302),
.Y(n_491)
);

INVx3_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

AND2x2_ASAP7_75t_L g492 ( 
.A(n_306),
.B(n_493),
.Y(n_492)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx1_ASAP7_75t_SL g394 ( 
.A(n_310),
.Y(n_394)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_312),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_332),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g409 ( 
.A(n_313),
.B(n_332),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_314),
.A2(n_318),
.B1(n_320),
.B2(n_324),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_316),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_315),
.B(n_321),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_SL g386 ( 
.A1(n_315),
.A2(n_387),
.B(n_388),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_315),
.B(n_503),
.Y(n_502)
);

INVx4_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

BUFx6f_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVx4_ASAP7_75t_L g323 ( 
.A(n_319),
.Y(n_323)
);

INVx5_ASAP7_75t_L g396 ( 
.A(n_319),
.Y(n_396)
);

INVx3_ASAP7_75t_SL g321 ( 
.A(n_322),
.Y(n_321)
);

INVx4_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_328),
.Y(n_324)
);

INVx3_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

BUFx3_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx3_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

INVx8_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

BUFx6f_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

BUFx6f_ASAP7_75t_L g532 ( 
.A(n_335),
.Y(n_532)
);

OAI21xp5_ASAP7_75t_SL g498 ( 
.A1(n_336),
.A2(n_458),
.B(n_467),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_337),
.B(n_448),
.Y(n_447)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx4_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVx3_ASAP7_75t_L g344 ( 
.A(n_340),
.Y(n_344)
);

BUFx6f_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_341),
.Y(n_486)
);

INVx1_ASAP7_75t_SL g342 ( 
.A(n_343),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_345),
.Y(n_520)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_346),
.B(n_384),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_347),
.A2(n_348),
.B1(n_352),
.B2(n_353),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g587 ( 
.A(n_347),
.B(n_353),
.C(n_384),
.Y(n_587)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_354),
.B(n_365),
.Y(n_353)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_354),
.Y(n_569)
);

INVx4_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

INVx3_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

INVx3_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

INVx4_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

BUFx3_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_SL g568 ( 
.A(n_365),
.B(n_569),
.Y(n_568)
);

AO32x1_ASAP7_75t_L g365 ( 
.A1(n_366),
.A2(n_369),
.A3(n_372),
.B1(n_375),
.B2(n_376),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

INVx1_ASAP7_75t_SL g369 ( 
.A(n_370),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_375),
.Y(n_388)
);

NAND2xp33_ASAP7_75t_SL g376 ( 
.A(n_377),
.B(n_380),
.Y(n_376)
);

INVx1_ASAP7_75t_SL g377 ( 
.A(n_378),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

INVx3_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

INVx3_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

XOR2xp5_ASAP7_75t_L g384 ( 
.A(n_385),
.B(n_390),
.Y(n_384)
);

MAJx2_ASAP7_75t_L g583 ( 
.A(n_385),
.B(n_391),
.C(n_397),
.Y(n_583)
);

XNOR2xp5_ASAP7_75t_SL g390 ( 
.A(n_391),
.B(n_397),
.Y(n_390)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

INVx3_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

OAI21xp5_ASAP7_75t_L g564 ( 
.A1(n_399),
.A2(n_420),
.B(n_429),
.Y(n_564)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

AOI21xp5_ASAP7_75t_L g403 ( 
.A1(n_404),
.A2(n_430),
.B(n_518),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_SL g404 ( 
.A(n_405),
.B(n_408),
.Y(n_404)
);

NOR2xp67_ASAP7_75t_L g518 ( 
.A(n_405),
.B(n_408),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_409),
.B(n_410),
.C(n_419),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_409),
.B(n_433),
.Y(n_432)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_409),
.Y(n_436)
);

AOI22xp33_ASAP7_75t_L g517 ( 
.A1(n_409),
.A2(n_433),
.B1(n_434),
.B2(n_436),
.Y(n_517)
);

HB1xp67_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_L g434 ( 
.A(n_411),
.B(n_419),
.Y(n_434)
);

BUFx4f_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

INVx4_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

INVx4_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

INVx4_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

OAI21xp5_ASAP7_75t_SL g419 ( 
.A1(n_420),
.A2(n_421),
.B(n_429),
.Y(n_419)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_427),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

OAI321xp33_ASAP7_75t_L g430 ( 
.A1(n_431),
.A2(n_454),
.A3(n_511),
.B1(n_515),
.B2(n_516),
.C(n_598),
.Y(n_430)
);

AOI21x1_ASAP7_75t_L g431 ( 
.A1(n_432),
.A2(n_435),
.B(n_437),
.Y(n_431)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_434),
.B(n_436),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_437),
.B(n_517),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_438),
.B(n_450),
.C(n_451),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_L g513 ( 
.A(n_439),
.B(n_514),
.Y(n_513)
);

INVxp67_ASAP7_75t_L g468 ( 
.A(n_440),
.Y(n_468)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);

HB1xp67_ASAP7_75t_L g445 ( 
.A(n_446),
.Y(n_445)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_446),
.Y(n_465)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_449),
.Y(n_448)
);

XOR2xp5_ASAP7_75t_L g514 ( 
.A(n_450),
.B(n_452),
.Y(n_514)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_452),
.Y(n_451)
);

AOI21xp5_ASAP7_75t_L g454 ( 
.A1(n_455),
.A2(n_495),
.B(n_510),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_456),
.B(n_469),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_456),
.B(n_469),
.Y(n_510)
);

INVxp67_ASAP7_75t_L g457 ( 
.A(n_458),
.Y(n_457)
);

BUFx2_ASAP7_75t_L g459 ( 
.A(n_460),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_461),
.Y(n_460)
);

INVx4_ASAP7_75t_L g461 ( 
.A(n_462),
.Y(n_461)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_464),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_465),
.Y(n_464)
);

INVx1_ASAP7_75t_SL g466 ( 
.A(n_467),
.Y(n_466)
);

XNOR2xp5_ASAP7_75t_L g469 ( 
.A(n_470),
.B(n_492),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_470),
.B(n_492),
.Y(n_512)
);

AOI22xp5_ASAP7_75t_L g470 ( 
.A1(n_471),
.A2(n_480),
.B1(n_482),
.B2(n_487),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_SL g471 ( 
.A(n_472),
.B(n_476),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_473),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_474),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_475),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_476),
.B(n_488),
.Y(n_487)
);

BUFx2_ASAP7_75t_L g476 ( 
.A(n_477),
.Y(n_476)
);

HB1xp67_ASAP7_75t_L g477 ( 
.A(n_478),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_479),
.Y(n_478)
);

INVxp67_ASAP7_75t_L g480 ( 
.A(n_481),
.Y(n_480)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_483),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_484),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_485),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_486),
.Y(n_485)
);

HB1xp67_ASAP7_75t_L g488 ( 
.A(n_489),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_490),
.Y(n_489)
);

HB1xp67_ASAP7_75t_L g490 ( 
.A(n_491),
.Y(n_490)
);

OAI21xp5_ASAP7_75t_SL g495 ( 
.A1(n_496),
.A2(n_499),
.B(n_509),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_497),
.B(n_498),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_SL g509 ( 
.A(n_497),
.B(n_498),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_SL g499 ( 
.A(n_500),
.B(n_501),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_SL g501 ( 
.A(n_502),
.B(n_506),
.Y(n_501)
);

INVx4_ASAP7_75t_L g503 ( 
.A(n_504),
.Y(n_503)
);

INVx4_ASAP7_75t_L g504 ( 
.A(n_505),
.Y(n_504)
);

INVx5_ASAP7_75t_L g506 ( 
.A(n_507),
.Y(n_506)
);

BUFx6f_ASAP7_75t_L g507 ( 
.A(n_508),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_512),
.B(n_513),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_512),
.B(n_513),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_SL g521 ( 
.A(n_522),
.B(n_573),
.Y(n_521)
);

INVxp67_ASAP7_75t_L g592 ( 
.A(n_522),
.Y(n_592)
);

OAI21xp5_ASAP7_75t_SL g522 ( 
.A1(n_523),
.A2(n_552),
.B(n_555),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_523),
.B(n_552),
.Y(n_596)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_524),
.Y(n_523)
);

AND2x2_ASAP7_75t_L g594 ( 
.A(n_524),
.B(n_553),
.Y(n_594)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_525),
.B(n_545),
.C(n_549),
.Y(n_524)
);

XNOR2xp5_ASAP7_75t_L g570 ( 
.A(n_525),
.B(n_571),
.Y(n_570)
);

MAJx2_ASAP7_75t_L g525 ( 
.A(n_526),
.B(n_534),
.C(n_541),
.Y(n_525)
);

XOR2x1_ASAP7_75t_SL g558 ( 
.A(n_526),
.B(n_559),
.Y(n_558)
);

AND2x2_ASAP7_75t_L g526 ( 
.A(n_527),
.B(n_529),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_528),
.Y(n_527)
);

XOR2xp5_ASAP7_75t_L g581 ( 
.A(n_528),
.B(n_529),
.Y(n_581)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_531),
.Y(n_530)
);

HB1xp67_ASAP7_75t_L g531 ( 
.A(n_532),
.Y(n_531)
);

XNOR2x1_ASAP7_75t_SL g559 ( 
.A(n_534),
.B(n_542),
.Y(n_559)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_537),
.Y(n_536)
);

INVx2_ASAP7_75t_SL g537 ( 
.A(n_538),
.Y(n_537)
);

INVx11_ASAP7_75t_L g539 ( 
.A(n_540),
.Y(n_539)
);

HB1xp67_ASAP7_75t_L g541 ( 
.A(n_542),
.Y(n_541)
);

HB1xp67_ASAP7_75t_L g545 ( 
.A(n_546),
.Y(n_545)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_546),
.Y(n_572)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_548),
.Y(n_547)
);

INVxp67_ASAP7_75t_SL g549 ( 
.A(n_550),
.Y(n_549)
);

XOR2xp5_ASAP7_75t_L g571 ( 
.A(n_550),
.B(n_572),
.Y(n_571)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_553),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_556),
.B(n_570),
.Y(n_555)
);

OR2x2_ASAP7_75t_L g595 ( 
.A(n_556),
.B(n_570),
.Y(n_595)
);

MAJIxp5_ASAP7_75t_L g556 ( 
.A(n_557),
.B(n_560),
.C(n_562),
.Y(n_556)
);

INVxp33_ASAP7_75t_L g557 ( 
.A(n_558),
.Y(n_557)
);

XOR2x1_ASAP7_75t_L g575 ( 
.A(n_558),
.B(n_560),
.Y(n_575)
);

XNOR2x1_ASAP7_75t_L g574 ( 
.A(n_562),
.B(n_575),
.Y(n_574)
);

MAJIxp5_ASAP7_75t_L g562 ( 
.A(n_563),
.B(n_565),
.C(n_568),
.Y(n_562)
);

OAI22xp5_ASAP7_75t_L g579 ( 
.A1(n_563),
.A2(n_564),
.B1(n_565),
.B2(n_566),
.Y(n_579)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_564),
.Y(n_563)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_566),
.Y(n_565)
);

XNOR2xp5_ASAP7_75t_L g578 ( 
.A(n_568),
.B(n_579),
.Y(n_578)
);

OAI21xp5_ASAP7_75t_L g573 ( 
.A1(n_574),
.A2(n_576),
.B(n_584),
.Y(n_573)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_574),
.Y(n_590)
);

INVx1_ASAP7_75t_SL g576 ( 
.A(n_577),
.Y(n_576)
);

MAJIxp5_ASAP7_75t_L g589 ( 
.A(n_577),
.B(n_590),
.C(n_591),
.Y(n_589)
);

MAJx2_ASAP7_75t_L g577 ( 
.A(n_578),
.B(n_580),
.C(n_582),
.Y(n_577)
);

XNOR2xp5_ASAP7_75t_L g585 ( 
.A(n_578),
.B(n_586),
.Y(n_585)
);

HB1xp67_ASAP7_75t_L g580 ( 
.A(n_581),
.Y(n_580)
);

XNOR2xp5_ASAP7_75t_L g586 ( 
.A(n_581),
.B(n_583),
.Y(n_586)
);

HB1xp67_ASAP7_75t_L g582 ( 
.A(n_583),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_585),
.B(n_587),
.Y(n_584)
);

OR2x2_ASAP7_75t_L g591 ( 
.A(n_585),
.B(n_587),
.Y(n_591)
);

AOI21x1_ASAP7_75t_L g588 ( 
.A1(n_589),
.A2(n_592),
.B(n_593),
.Y(n_588)
);

OAI21xp5_ASAP7_75t_L g593 ( 
.A1(n_594),
.A2(n_595),
.B(n_596),
.Y(n_593)
);


endmodule