module fake_ariane_1711_n_770 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_18, n_86, n_75, n_89, n_67, n_34, n_69, n_95, n_92, n_143, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_52, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_136, n_28, n_80, n_97, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_127, n_35, n_54, n_25, n_770);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_34;
input n_69;
input n_95;
input n_92;
input n_143;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_52;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_136;
input n_28;
input n_80;
input n_97;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_127;
input n_35;
input n_54;
input n_25;

output n_770;

wire n_295;
wire n_356;
wire n_556;
wire n_170;
wire n_190;
wire n_698;
wire n_695;
wire n_160;
wire n_180;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_581;
wire n_294;
wire n_646;
wire n_197;
wire n_640;
wire n_463;
wire n_176;
wire n_691;
wire n_404;
wire n_172;
wire n_678;
wire n_651;
wire n_347;
wire n_423;
wire n_183;
wire n_469;
wire n_479;
wire n_726;
wire n_603;
wire n_373;
wire n_299;
wire n_541;
wire n_499;
wire n_564;
wire n_610;
wire n_205;
wire n_752;
wire n_341;
wire n_245;
wire n_421;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_760;
wire n_690;
wire n_416;
wire n_283;
wire n_187;
wire n_525;
wire n_367;
wire n_713;
wire n_649;
wire n_598;
wire n_374;
wire n_345;
wire n_318;
wire n_244;
wire n_643;
wire n_679;
wire n_226;
wire n_261;
wire n_220;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_189;
wire n_717;
wire n_286;
wire n_443;
wire n_586;
wire n_686;
wire n_605;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_524;
wire n_391;
wire n_349;
wire n_634;
wire n_756;
wire n_466;
wire n_346;
wire n_214;
wire n_764;
wire n_348;
wire n_552;
wire n_462;
wire n_607;
wire n_670;
wire n_410;
wire n_379;
wire n_445;
wire n_515;
wire n_162;
wire n_765;
wire n_264;
wire n_737;
wire n_198;
wire n_232;
wire n_441;
wire n_568;
wire n_385;
wire n_637;
wire n_327;
wire n_766;
wire n_372;
wire n_377;
wire n_396;
wire n_631;
wire n_399;
wire n_554;
wire n_520;
wire n_714;
wire n_279;
wire n_702;
wire n_207;
wire n_363;
wire n_720;
wire n_354;
wire n_725;
wire n_419;
wire n_151;
wire n_146;
wire n_230;
wire n_270;
wire n_194;
wire n_633;
wire n_154;
wire n_338;
wire n_285;
wire n_473;
wire n_186;
wire n_202;
wire n_193;
wire n_733;
wire n_761;
wire n_500;
wire n_665;
wire n_336;
wire n_731;
wire n_754;
wire n_315;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_668;
wire n_339;
wire n_738;
wire n_758;
wire n_672;
wire n_487;
wire n_740;
wire n_167;
wire n_422;
wire n_153;
wire n_648;
wire n_269;
wire n_597;
wire n_158;
wire n_259;
wire n_446;
wire n_553;
wire n_753;
wire n_566;
wire n_578;
wire n_701;
wire n_625;
wire n_152;
wire n_405;
wire n_557;
wire n_169;
wire n_173;
wire n_242;
wire n_645;
wire n_331;
wire n_320;
wire n_309;
wire n_559;
wire n_485;
wire n_401;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_344;
wire n_381;
wire n_426;
wire n_433;
wire n_481;
wire n_600;
wire n_721;
wire n_398;
wire n_210;
wire n_200;
wire n_529;
wire n_502;
wire n_166;
wire n_253;
wire n_561;
wire n_218;
wire n_271;
wire n_507;
wire n_465;
wire n_486;
wire n_759;
wire n_247;
wire n_569;
wire n_567;
wire n_732;
wire n_240;
wire n_369;
wire n_224;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_222;
wire n_478;
wire n_703;
wire n_748;
wire n_510;
wire n_256;
wire n_326;
wire n_681;
wire n_227;
wire n_188;
wire n_323;
wire n_550;
wire n_635;
wire n_707;
wire n_330;
wire n_400;
wire n_694;
wire n_689;
wire n_282;
wire n_328;
wire n_368;
wire n_590;
wire n_699;
wire n_727;
wire n_277;
wire n_248;
wire n_301;
wire n_467;
wire n_432;
wire n_545;
wire n_536;
wire n_644;
wire n_293;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_693;
wire n_303;
wire n_671;
wire n_442;
wire n_168;
wire n_206;
wire n_352;
wire n_538;
wire n_576;
wire n_511;
wire n_611;
wire n_238;
wire n_365;
wire n_429;
wire n_455;
wire n_654;
wire n_588;
wire n_638;
wire n_334;
wire n_192;
wire n_729;
wire n_661;
wire n_488;
wire n_667;
wire n_300;
wire n_533;
wire n_505;
wire n_163;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_512;
wire n_715;
wire n_579;
wire n_459;
wire n_685;
wire n_221;
wire n_321;
wire n_361;
wire n_458;
wire n_149;
wire n_383;
wire n_623;
wire n_237;
wire n_175;
wire n_711;
wire n_453;
wire n_734;
wire n_491;
wire n_181;
wire n_723;
wire n_616;
wire n_617;
wire n_658;
wire n_630;
wire n_705;
wire n_570;
wire n_260;
wire n_543;
wire n_362;
wire n_310;
wire n_709;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_281;
wire n_628;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_743;
wire n_225;
wire n_235;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_297;
wire n_662;
wire n_641;
wire n_503;
wire n_700;
wire n_290;
wire n_527;
wire n_741;
wire n_747;
wire n_371;
wire n_199;
wire n_639;
wire n_217;
wire n_452;
wire n_673;
wire n_676;
wire n_178;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_201;
wire n_572;
wire n_343;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_582;
wire n_284;
wire n_448;
wire n_593;
wire n_755;
wire n_710;
wire n_249;
wire n_534;
wire n_212;
wire n_444;
wire n_355;
wire n_609;
wire n_278;
wire n_255;
wire n_560;
wire n_450;
wire n_257;
wire n_148;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_468;
wire n_526;
wire n_716;
wire n_742;
wire n_182;
wire n_696;
wire n_674;
wire n_482;
wire n_316;
wire n_196;
wire n_769;
wire n_577;
wire n_407;
wire n_254;
wire n_596;
wire n_476;
wire n_460;
wire n_219;
wire n_535;
wire n_231;
wire n_366;
wire n_744;
wire n_762;
wire n_656;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_280;
wire n_215;
wire n_252;
wire n_629;
wire n_664;
wire n_161;
wire n_454;
wire n_298;
wire n_532;
wire n_415;
wire n_763;
wire n_655;
wire n_544;
wire n_540;
wire n_216;
wire n_692;
wire n_599;
wire n_768;
wire n_514;
wire n_418;
wire n_537;
wire n_223;
wire n_403;
wire n_750;
wire n_389;
wire n_657;
wire n_513;
wire n_288;
wire n_179;
wire n_395;
wire n_621;
wire n_195;
wire n_606;
wire n_213;
wire n_304;
wire n_659;
wire n_583;
wire n_509;
wire n_724;
wire n_306;
wire n_666;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_203;
wire n_378;
wire n_436;
wire n_150;
wire n_757;
wire n_375;
wire n_324;
wire n_585;
wire n_669;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_622;
wire n_697;
wire n_472;
wire n_296;
wire n_265;
wire n_746;
wire n_208;
wire n_456;
wire n_156;
wire n_292;
wire n_174;
wire n_275;
wire n_704;
wire n_147;
wire n_204;
wire n_751;
wire n_615;
wire n_521;
wire n_496;
wire n_739;
wire n_342;
wire n_246;
wire n_517;
wire n_530;
wire n_428;
wire n_159;
wire n_358;
wire n_580;
wire n_608;
wire n_494;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_563;
wire n_229;
wire n_394;
wire n_250;
wire n_165;
wire n_317;
wire n_243;
wire n_329;
wire n_718;
wire n_185;
wire n_340;
wire n_749;
wire n_289;
wire n_548;
wire n_542;
wire n_523;
wire n_268;
wire n_266;
wire n_470;
wire n_457;
wire n_164;
wire n_157;
wire n_632;
wire n_184;
wire n_177;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_425;
wire n_431;
wire n_508;
wire n_624;
wire n_618;
wire n_484;
wire n_411;
wire n_712;
wire n_353;
wire n_736;
wire n_767;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_191;
wire n_382;
wire n_489;
wire n_480;
wire n_211;
wire n_642;
wire n_408;
wire n_595;
wire n_322;
wire n_251;
wire n_506;
wire n_602;
wire n_558;
wire n_592;
wire n_397;
wire n_471;
wire n_351;
wire n_393;
wire n_474;
wire n_653;
wire n_359;
wire n_155;
wire n_573;
wire n_531;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g146 ( 
.A(n_75),
.Y(n_146)
);

CKINVDCx5p33_ASAP7_75t_R g147 ( 
.A(n_82),
.Y(n_147)
);

CKINVDCx5p33_ASAP7_75t_R g148 ( 
.A(n_143),
.Y(n_148)
);

CKINVDCx5p33_ASAP7_75t_R g149 ( 
.A(n_6),
.Y(n_149)
);

CKINVDCx5p33_ASAP7_75t_R g150 ( 
.A(n_98),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_27),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_10),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_79),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_3),
.Y(n_154)
);

INVxp67_ASAP7_75t_SL g155 ( 
.A(n_123),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_139),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_89),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_19),
.Y(n_158)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_74),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_91),
.Y(n_160)
);

CKINVDCx14_ASAP7_75t_R g161 ( 
.A(n_108),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_6),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_109),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_141),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_81),
.Y(n_165)
);

INVx1_ASAP7_75t_SL g166 ( 
.A(n_96),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_121),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_3),
.Y(n_168)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_56),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_30),
.Y(n_170)
);

BUFx10_ASAP7_75t_L g171 ( 
.A(n_63),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_113),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_101),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_115),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_134),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_18),
.Y(n_176)
);

INVx1_ASAP7_75t_SL g177 ( 
.A(n_43),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_58),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_117),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_100),
.Y(n_180)
);

BUFx3_ASAP7_75t_L g181 ( 
.A(n_105),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_95),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_76),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_77),
.Y(n_184)
);

INVx2_ASAP7_75t_SL g185 ( 
.A(n_53),
.Y(n_185)
);

BUFx2_ASAP7_75t_L g186 ( 
.A(n_10),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_47),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_126),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_64),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_61),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_31),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_51),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_34),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_32),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_102),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_9),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_29),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_142),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_44),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_181),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_181),
.Y(n_201)
);

AND2x4_ASAP7_75t_L g202 ( 
.A(n_185),
.B(n_0),
.Y(n_202)
);

BUFx12f_ASAP7_75t_L g203 ( 
.A(n_171),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_151),
.B(n_164),
.Y(n_204)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_171),
.Y(n_205)
);

INVx5_ASAP7_75t_L g206 ( 
.A(n_185),
.Y(n_206)
);

AND2x2_ASAP7_75t_L g207 ( 
.A(n_186),
.B(n_161),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_159),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_159),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_169),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_179),
.B(n_180),
.Y(n_211)
);

INVx2_ASAP7_75t_SL g212 ( 
.A(n_171),
.Y(n_212)
);

AND2x4_ASAP7_75t_L g213 ( 
.A(n_169),
.B(n_158),
.Y(n_213)
);

INVx5_ASAP7_75t_L g214 ( 
.A(n_156),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_182),
.B(n_0),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_162),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_187),
.B(n_189),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_191),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_155),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_146),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_153),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_195),
.B(n_1),
.Y(n_222)
);

BUFx2_ASAP7_75t_L g223 ( 
.A(n_149),
.Y(n_223)
);

AND2x2_ASAP7_75t_L g224 ( 
.A(n_149),
.B(n_1),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_147),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_152),
.B(n_2),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_147),
.B(n_148),
.Y(n_227)
);

INVx4_ASAP7_75t_L g228 ( 
.A(n_148),
.Y(n_228)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_150),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_150),
.B(n_2),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_199),
.B(n_4),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_157),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_160),
.Y(n_233)
);

INVx2_ASAP7_75t_SL g234 ( 
.A(n_154),
.Y(n_234)
);

BUFx2_ASAP7_75t_L g235 ( 
.A(n_168),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_199),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_172),
.B(n_23),
.Y(n_237)
);

INVx4_ASAP7_75t_L g238 ( 
.A(n_163),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_165),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_200),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_237),
.A2(n_172),
.B1(n_196),
.B2(n_176),
.Y(n_241)
);

OAI22xp33_ASAP7_75t_L g242 ( 
.A1(n_222),
.A2(n_166),
.B1(n_177),
.B2(n_194),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_208),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_200),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_200),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_200),
.Y(n_246)
);

OAI22xp33_ASAP7_75t_SL g247 ( 
.A1(n_219),
.A2(n_198),
.B1(n_197),
.B2(n_193),
.Y(n_247)
);

INVx3_ASAP7_75t_L g248 ( 
.A(n_200),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g249 ( 
.A(n_208),
.Y(n_249)
);

INVx2_ASAP7_75t_SL g250 ( 
.A(n_203),
.Y(n_250)
);

BUFx2_ASAP7_75t_L g251 ( 
.A(n_235),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_207),
.A2(n_192),
.B1(n_190),
.B2(n_188),
.Y(n_252)
);

OAI22xp33_ASAP7_75t_L g253 ( 
.A1(n_212),
.A2(n_184),
.B1(n_183),
.B2(n_178),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_207),
.A2(n_175),
.B1(n_174),
.B2(n_173),
.Y(n_254)
);

OAI22xp33_ASAP7_75t_L g255 ( 
.A1(n_205),
.A2(n_212),
.B1(n_223),
.B2(n_203),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_201),
.Y(n_256)
);

OR2x6_ASAP7_75t_L g257 ( 
.A(n_223),
.B(n_4),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g258 ( 
.A(n_205),
.B(n_167),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g259 ( 
.A(n_205),
.B(n_170),
.Y(n_259)
);

OR2x6_ASAP7_75t_L g260 ( 
.A(n_224),
.B(n_5),
.Y(n_260)
);

INVxp67_ASAP7_75t_SL g261 ( 
.A(n_209),
.Y(n_261)
);

AO22x2_ASAP7_75t_L g262 ( 
.A1(n_202),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_235),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_219),
.B(n_24),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_202),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_265)
);

AND2x2_ASAP7_75t_L g266 ( 
.A(n_214),
.B(n_11),
.Y(n_266)
);

AND2x2_ASAP7_75t_L g267 ( 
.A(n_214),
.B(n_12),
.Y(n_267)
);

INVx1_ASAP7_75t_SL g268 ( 
.A(n_227),
.Y(n_268)
);

OAI22xp33_ASAP7_75t_L g269 ( 
.A1(n_204),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_269)
);

INVx3_ASAP7_75t_L g270 ( 
.A(n_201),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_234),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_201),
.Y(n_272)
);

OAI22xp33_ASAP7_75t_R g273 ( 
.A1(n_234),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_201),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_201),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_208),
.Y(n_276)
);

OAI22xp33_ASAP7_75t_L g277 ( 
.A1(n_211),
.A2(n_17),
.B1(n_19),
.B2(n_20),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_216),
.Y(n_278)
);

OAI22xp33_ASAP7_75t_L g279 ( 
.A1(n_217),
.A2(n_20),
.B1(n_21),
.B2(n_22),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_202),
.A2(n_226),
.B1(n_224),
.B2(n_236),
.Y(n_280)
);

OAI22xp33_ASAP7_75t_SL g281 ( 
.A1(n_202),
.A2(n_21),
.B1(n_22),
.B2(n_25),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_216),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_226),
.A2(n_26),
.B1(n_28),
.B2(n_33),
.Y(n_283)
);

OAI22xp33_ASAP7_75t_L g284 ( 
.A1(n_230),
.A2(n_35),
.B1(n_36),
.B2(n_37),
.Y(n_284)
);

OAI22xp33_ASAP7_75t_L g285 ( 
.A1(n_215),
.A2(n_38),
.B1(n_39),
.B2(n_40),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_213),
.B(n_41),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_250),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_278),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_241),
.B(n_225),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_251),
.B(n_225),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_282),
.Y(n_291)
);

XNOR2x2_ASAP7_75t_L g292 ( 
.A(n_262),
.B(n_231),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_261),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_255),
.B(n_236),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_261),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_248),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_268),
.A2(n_239),
.B(n_229),
.Y(n_297)
);

AND2x2_ASAP7_75t_L g298 ( 
.A(n_268),
.B(n_213),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_248),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_276),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_240),
.Y(n_301)
);

CKINVDCx16_ASAP7_75t_R g302 ( 
.A(n_260),
.Y(n_302)
);

INVxp33_ASAP7_75t_L g303 ( 
.A(n_286),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_258),
.B(n_214),
.Y(n_304)
);

OR2x2_ASAP7_75t_L g305 ( 
.A(n_257),
.B(n_218),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_SL g306 ( 
.A(n_255),
.B(n_214),
.Y(n_306)
);

INVx2_ASAP7_75t_SL g307 ( 
.A(n_259),
.Y(n_307)
);

AND2x2_ASAP7_75t_L g308 ( 
.A(n_280),
.B(n_213),
.Y(n_308)
);

XOR2x2_ASAP7_75t_L g309 ( 
.A(n_247),
.B(n_213),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_270),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_244),
.Y(n_311)
);

INVx3_ASAP7_75t_R g312 ( 
.A(n_245),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_270),
.Y(n_313)
);

INVxp67_ASAP7_75t_SL g314 ( 
.A(n_246),
.Y(n_314)
);

BUFx6f_ASAP7_75t_L g315 ( 
.A(n_243),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_257),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_256),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_272),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_274),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_252),
.B(n_228),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_275),
.Y(n_321)
);

AND2x2_ASAP7_75t_L g322 ( 
.A(n_260),
.B(n_218),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_243),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_264),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_264),
.Y(n_325)
);

BUFx3_ASAP7_75t_L g326 ( 
.A(n_243),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_249),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_249),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_249),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_266),
.Y(n_330)
);

AND2x2_ASAP7_75t_L g331 ( 
.A(n_260),
.B(n_209),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_267),
.Y(n_332)
);

BUFx3_ASAP7_75t_L g333 ( 
.A(n_283),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_265),
.Y(n_334)
);

AND2x2_ASAP7_75t_L g335 ( 
.A(n_257),
.B(n_210),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_254),
.B(n_247),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_262),
.Y(n_337)
);

AND2x2_ASAP7_75t_L g338 ( 
.A(n_262),
.B(n_228),
.Y(n_338)
);

NOR2xp67_ASAP7_75t_L g339 ( 
.A(n_253),
.B(n_214),
.Y(n_339)
);

INVx4_ASAP7_75t_SL g340 ( 
.A(n_271),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_242),
.B(n_239),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_281),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_281),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_277),
.B(n_228),
.Y(n_344)
);

XOR2x2_ASAP7_75t_L g345 ( 
.A(n_263),
.B(n_210),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_279),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_269),
.Y(n_347)
);

INVx1_ASAP7_75t_SL g348 ( 
.A(n_273),
.Y(n_348)
);

BUFx6f_ASAP7_75t_L g349 ( 
.A(n_284),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_269),
.Y(n_350)
);

OR2x6_ASAP7_75t_L g351 ( 
.A(n_337),
.B(n_208),
.Y(n_351)
);

OAI21x1_ASAP7_75t_L g352 ( 
.A1(n_324),
.A2(n_229),
.B(n_285),
.Y(n_352)
);

AND2x2_ASAP7_75t_SL g353 ( 
.A(n_306),
.B(n_285),
.Y(n_353)
);

OAI21xp5_ASAP7_75t_L g354 ( 
.A1(n_325),
.A2(n_229),
.B(n_206),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_300),
.Y(n_355)
);

AND2x2_ASAP7_75t_L g356 ( 
.A(n_298),
.B(n_214),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_300),
.Y(n_357)
);

AND2x2_ASAP7_75t_L g358 ( 
.A(n_298),
.B(n_308),
.Y(n_358)
);

OR2x2_ASAP7_75t_SL g359 ( 
.A(n_302),
.B(n_220),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_307),
.B(n_293),
.Y(n_360)
);

AND2x2_ASAP7_75t_L g361 ( 
.A(n_322),
.B(n_208),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_301),
.Y(n_362)
);

AND2x6_ASAP7_75t_L g363 ( 
.A(n_349),
.B(n_338),
.Y(n_363)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_301),
.Y(n_364)
);

AND2x2_ASAP7_75t_L g365 ( 
.A(n_322),
.B(n_238),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_311),
.Y(n_366)
);

AND2x4_ASAP7_75t_L g367 ( 
.A(n_331),
.B(n_238),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_320),
.B(n_238),
.Y(n_368)
);

AND2x6_ASAP7_75t_L g369 ( 
.A(n_349),
.B(n_220),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_307),
.B(n_220),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_311),
.Y(n_371)
);

AND2x4_ASAP7_75t_L g372 ( 
.A(n_331),
.B(n_220),
.Y(n_372)
);

AND2x4_ASAP7_75t_L g373 ( 
.A(n_335),
.B(n_220),
.Y(n_373)
);

OR2x6_ASAP7_75t_L g374 ( 
.A(n_333),
.B(n_221),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_319),
.Y(n_375)
);

BUFx3_ASAP7_75t_L g376 ( 
.A(n_326),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_295),
.B(n_221),
.Y(n_377)
);

OAI21xp5_ASAP7_75t_L g378 ( 
.A1(n_297),
.A2(n_206),
.B(n_232),
.Y(n_378)
);

BUFx6f_ASAP7_75t_L g379 ( 
.A(n_315),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_321),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_320),
.B(n_221),
.Y(n_381)
);

HB1xp67_ASAP7_75t_L g382 ( 
.A(n_290),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_317),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_318),
.Y(n_384)
);

OAI21xp5_ASAP7_75t_L g385 ( 
.A1(n_304),
.A2(n_206),
.B(n_232),
.Y(n_385)
);

AND2x2_ASAP7_75t_L g386 ( 
.A(n_335),
.B(n_206),
.Y(n_386)
);

AND2x2_ASAP7_75t_L g387 ( 
.A(n_342),
.B(n_206),
.Y(n_387)
);

AND2x2_ASAP7_75t_L g388 ( 
.A(n_343),
.B(n_206),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_344),
.B(n_221),
.Y(n_389)
);

INVx2_ASAP7_75t_SL g390 ( 
.A(n_305),
.Y(n_390)
);

INVx3_ASAP7_75t_L g391 ( 
.A(n_326),
.Y(n_391)
);

HB1xp67_ASAP7_75t_L g392 ( 
.A(n_287),
.Y(n_392)
);

AND2x4_ASAP7_75t_L g393 ( 
.A(n_333),
.B(n_334),
.Y(n_393)
);

OR2x2_ASAP7_75t_L g394 ( 
.A(n_348),
.B(n_294),
.Y(n_394)
);

OR2x2_ASAP7_75t_L g395 ( 
.A(n_347),
.B(n_221),
.Y(n_395)
);

AND2x2_ASAP7_75t_SL g396 ( 
.A(n_349),
.B(n_232),
.Y(n_396)
);

AND2x2_ASAP7_75t_L g397 ( 
.A(n_350),
.B(n_232),
.Y(n_397)
);

AND2x2_ASAP7_75t_L g398 ( 
.A(n_346),
.B(n_288),
.Y(n_398)
);

INVx3_ASAP7_75t_L g399 ( 
.A(n_323),
.Y(n_399)
);

AND2x2_ASAP7_75t_SL g400 ( 
.A(n_349),
.B(n_292),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_296),
.Y(n_401)
);

OAI21x1_ASAP7_75t_L g402 ( 
.A1(n_323),
.A2(n_233),
.B(n_232),
.Y(n_402)
);

INVx3_ASAP7_75t_L g403 ( 
.A(n_315),
.Y(n_403)
);

HB1xp67_ASAP7_75t_L g404 ( 
.A(n_287),
.Y(n_404)
);

HB1xp67_ASAP7_75t_L g405 ( 
.A(n_289),
.Y(n_405)
);

INVx4_ASAP7_75t_L g406 ( 
.A(n_315),
.Y(n_406)
);

INVxp67_ASAP7_75t_L g407 ( 
.A(n_341),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_291),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_344),
.B(n_233),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_299),
.Y(n_410)
);

BUFx6f_ASAP7_75t_L g411 ( 
.A(n_315),
.Y(n_411)
);

AND2x2_ASAP7_75t_L g412 ( 
.A(n_330),
.B(n_233),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_332),
.B(n_339),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_314),
.B(n_310),
.Y(n_414)
);

BUFx6f_ASAP7_75t_L g415 ( 
.A(n_327),
.Y(n_415)
);

OAI21xp5_ASAP7_75t_L g416 ( 
.A1(n_314),
.A2(n_233),
.B(n_45),
.Y(n_416)
);

AND2x2_ASAP7_75t_L g417 ( 
.A(n_309),
.B(n_233),
.Y(n_417)
);

BUFx2_ASAP7_75t_L g418 ( 
.A(n_374),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_408),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_408),
.Y(n_420)
);

BUFx3_ASAP7_75t_L g421 ( 
.A(n_393),
.Y(n_421)
);

BUFx2_ASAP7_75t_SL g422 ( 
.A(n_390),
.Y(n_422)
);

OR2x2_ASAP7_75t_L g423 ( 
.A(n_394),
.B(n_303),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_383),
.Y(n_424)
);

OR2x2_ASAP7_75t_L g425 ( 
.A(n_394),
.B(n_303),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_392),
.B(n_336),
.Y(n_426)
);

BUFx12f_ASAP7_75t_L g427 ( 
.A(n_359),
.Y(n_427)
);

AND2x4_ASAP7_75t_L g428 ( 
.A(n_393),
.B(n_340),
.Y(n_428)
);

INVx6_ASAP7_75t_L g429 ( 
.A(n_376),
.Y(n_429)
);

OR2x6_ASAP7_75t_L g430 ( 
.A(n_393),
.B(n_292),
.Y(n_430)
);

BUFx4f_ASAP7_75t_L g431 ( 
.A(n_363),
.Y(n_431)
);

AND2x2_ASAP7_75t_SL g432 ( 
.A(n_400),
.B(n_316),
.Y(n_432)
);

AND2x4_ASAP7_75t_L g433 ( 
.A(n_358),
.B(n_390),
.Y(n_433)
);

BUFx12f_ASAP7_75t_L g434 ( 
.A(n_359),
.Y(n_434)
);

BUFx12f_ASAP7_75t_L g435 ( 
.A(n_367),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_358),
.B(n_309),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_364),
.Y(n_437)
);

INVx4_ASAP7_75t_L g438 ( 
.A(n_376),
.Y(n_438)
);

AND2x4_ASAP7_75t_L g439 ( 
.A(n_367),
.B(n_340),
.Y(n_439)
);

OR2x2_ASAP7_75t_L g440 ( 
.A(n_382),
.B(n_345),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_368),
.B(n_313),
.Y(n_441)
);

BUFx3_ASAP7_75t_L g442 ( 
.A(n_404),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_397),
.B(n_353),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_364),
.Y(n_444)
);

INVxp67_ASAP7_75t_L g445 ( 
.A(n_365),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_397),
.B(n_328),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_353),
.B(n_329),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_383),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_384),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_353),
.B(n_345),
.Y(n_450)
);

AND2x2_ASAP7_75t_L g451 ( 
.A(n_417),
.B(n_340),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_396),
.B(n_316),
.Y(n_452)
);

OR2x2_ASAP7_75t_L g453 ( 
.A(n_405),
.B(n_417),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_396),
.B(n_42),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_384),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_396),
.B(n_46),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_398),
.B(n_48),
.Y(n_457)
);

OR2x6_ASAP7_75t_L g458 ( 
.A(n_374),
.B(n_312),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_371),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_367),
.B(n_400),
.Y(n_460)
);

AND2x4_ASAP7_75t_L g461 ( 
.A(n_398),
.B(n_49),
.Y(n_461)
);

INVx4_ASAP7_75t_L g462 ( 
.A(n_363),
.Y(n_462)
);

AO21x2_ASAP7_75t_L g463 ( 
.A1(n_416),
.A2(n_50),
.B(n_52),
.Y(n_463)
);

AND2x2_ASAP7_75t_L g464 ( 
.A(n_365),
.B(n_54),
.Y(n_464)
);

BUFx2_ASAP7_75t_L g465 ( 
.A(n_374),
.Y(n_465)
);

BUFx8_ASAP7_75t_L g466 ( 
.A(n_373),
.Y(n_466)
);

AND2x4_ASAP7_75t_L g467 ( 
.A(n_372),
.B(n_55),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_412),
.Y(n_468)
);

AND2x2_ASAP7_75t_L g469 ( 
.A(n_407),
.B(n_361),
.Y(n_469)
);

INVx2_ASAP7_75t_SL g470 ( 
.A(n_373),
.Y(n_470)
);

HB1xp67_ASAP7_75t_L g471 ( 
.A(n_361),
.Y(n_471)
);

NOR2xp67_ASAP7_75t_L g472 ( 
.A(n_370),
.B(n_57),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_400),
.B(n_145),
.Y(n_473)
);

BUFx6f_ASAP7_75t_L g474 ( 
.A(n_379),
.Y(n_474)
);

HB1xp67_ASAP7_75t_L g475 ( 
.A(n_442),
.Y(n_475)
);

CKINVDCx20_ASAP7_75t_R g476 ( 
.A(n_422),
.Y(n_476)
);

INVx4_ASAP7_75t_L g477 ( 
.A(n_431),
.Y(n_477)
);

BUFx3_ASAP7_75t_L g478 ( 
.A(n_431),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_427),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_437),
.Y(n_480)
);

INVx2_ASAP7_75t_SL g481 ( 
.A(n_429),
.Y(n_481)
);

INVx1_ASAP7_75t_SL g482 ( 
.A(n_423),
.Y(n_482)
);

BUFx2_ASAP7_75t_L g483 ( 
.A(n_435),
.Y(n_483)
);

INVx3_ASAP7_75t_L g484 ( 
.A(n_462),
.Y(n_484)
);

BUFx12f_ASAP7_75t_L g485 ( 
.A(n_425),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_444),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_459),
.Y(n_487)
);

BUFx3_ASAP7_75t_L g488 ( 
.A(n_462),
.Y(n_488)
);

AND2x2_ASAP7_75t_L g489 ( 
.A(n_450),
.B(n_356),
.Y(n_489)
);

NAND2x1p5_ASAP7_75t_L g490 ( 
.A(n_467),
.B(n_406),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_450),
.B(n_360),
.Y(n_491)
);

AOI22xp33_ASAP7_75t_L g492 ( 
.A1(n_430),
.A2(n_363),
.B1(n_356),
.B2(n_372),
.Y(n_492)
);

INVx3_ASAP7_75t_SL g493 ( 
.A(n_439),
.Y(n_493)
);

INVx2_ASAP7_75t_SL g494 ( 
.A(n_429),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_424),
.Y(n_495)
);

AND2x2_ASAP7_75t_L g496 ( 
.A(n_460),
.B(n_363),
.Y(n_496)
);

BUFx3_ASAP7_75t_L g497 ( 
.A(n_466),
.Y(n_497)
);

INVx6_ASAP7_75t_SL g498 ( 
.A(n_458),
.Y(n_498)
);

BUFx12f_ASAP7_75t_L g499 ( 
.A(n_428),
.Y(n_499)
);

BUFx12f_ASAP7_75t_L g500 ( 
.A(n_428),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_419),
.Y(n_501)
);

BUFx3_ASAP7_75t_L g502 ( 
.A(n_466),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_420),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_448),
.Y(n_504)
);

INVx2_ASAP7_75t_SL g505 ( 
.A(n_429),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_449),
.Y(n_506)
);

BUFx8_ASAP7_75t_L g507 ( 
.A(n_439),
.Y(n_507)
);

OR2x2_ASAP7_75t_L g508 ( 
.A(n_436),
.B(n_452),
.Y(n_508)
);

INVx1_ASAP7_75t_SL g509 ( 
.A(n_453),
.Y(n_509)
);

AND2x4_ASAP7_75t_L g510 ( 
.A(n_421),
.B(n_363),
.Y(n_510)
);

NAND2x1p5_ASAP7_75t_L g511 ( 
.A(n_467),
.B(n_406),
.Y(n_511)
);

BUFx2_ASAP7_75t_SL g512 ( 
.A(n_474),
.Y(n_512)
);

HB1xp67_ASAP7_75t_L g513 ( 
.A(n_433),
.Y(n_513)
);

AOI22xp5_ASAP7_75t_SL g514 ( 
.A1(n_426),
.A2(n_363),
.B1(n_369),
.B2(n_381),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_455),
.Y(n_515)
);

INVx4_ASAP7_75t_L g516 ( 
.A(n_474),
.Y(n_516)
);

BUFx3_ASAP7_75t_L g517 ( 
.A(n_474),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_446),
.Y(n_518)
);

INVx5_ASAP7_75t_L g519 ( 
.A(n_458),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_445),
.B(n_363),
.Y(n_520)
);

CKINVDCx11_ASAP7_75t_R g521 ( 
.A(n_476),
.Y(n_521)
);

AOI22xp33_ASAP7_75t_L g522 ( 
.A1(n_491),
.A2(n_430),
.B1(n_436),
.B2(n_440),
.Y(n_522)
);

INVx6_ASAP7_75t_L g523 ( 
.A(n_507),
.Y(n_523)
);

AOI22xp33_ASAP7_75t_L g524 ( 
.A1(n_489),
.A2(n_430),
.B1(n_432),
.B2(n_473),
.Y(n_524)
);

CKINVDCx20_ASAP7_75t_R g525 ( 
.A(n_497),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_501),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_495),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_485),
.Y(n_528)
);

HB1xp67_ASAP7_75t_SL g529 ( 
.A(n_507),
.Y(n_529)
);

AOI22xp33_ASAP7_75t_L g530 ( 
.A1(n_489),
.A2(n_469),
.B1(n_451),
.B2(n_492),
.Y(n_530)
);

AOI22xp33_ASAP7_75t_L g531 ( 
.A1(n_508),
.A2(n_433),
.B1(n_443),
.B2(n_452),
.Y(n_531)
);

AOI22xp33_ASAP7_75t_SL g532 ( 
.A1(n_514),
.A2(n_461),
.B1(n_434),
.B2(n_374),
.Y(n_532)
);

AOI22xp33_ASAP7_75t_SL g533 ( 
.A1(n_514),
.A2(n_461),
.B1(n_454),
.B2(n_456),
.Y(n_533)
);

CKINVDCx11_ASAP7_75t_R g534 ( 
.A(n_485),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_501),
.Y(n_535)
);

BUFx8_ASAP7_75t_L g536 ( 
.A(n_483),
.Y(n_536)
);

INVx2_ASAP7_75t_R g537 ( 
.A(n_488),
.Y(n_537)
);

BUFx2_ASAP7_75t_L g538 ( 
.A(n_475),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_479),
.Y(n_539)
);

OAI22xp5_ASAP7_75t_L g540 ( 
.A1(n_490),
.A2(n_445),
.B1(n_471),
.B2(n_464),
.Y(n_540)
);

AOI22xp33_ASAP7_75t_L g541 ( 
.A1(n_508),
.A2(n_509),
.B1(n_482),
.B2(n_443),
.Y(n_541)
);

AOI22xp33_ASAP7_75t_L g542 ( 
.A1(n_513),
.A2(n_372),
.B1(n_373),
.B2(n_470),
.Y(n_542)
);

AOI22xp33_ASAP7_75t_SL g543 ( 
.A1(n_496),
.A2(n_369),
.B1(n_456),
.B2(n_454),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_503),
.Y(n_544)
);

OAI22xp5_ASAP7_75t_L g545 ( 
.A1(n_490),
.A2(n_471),
.B1(n_441),
.B2(n_457),
.Y(n_545)
);

AOI22xp33_ASAP7_75t_SL g546 ( 
.A1(n_496),
.A2(n_369),
.B1(n_457),
.B2(n_409),
.Y(n_546)
);

CKINVDCx8_ASAP7_75t_R g547 ( 
.A(n_483),
.Y(n_547)
);

CKINVDCx11_ASAP7_75t_R g548 ( 
.A(n_497),
.Y(n_548)
);

AOI22xp33_ASAP7_75t_L g549 ( 
.A1(n_495),
.A2(n_418),
.B1(n_465),
.B2(n_468),
.Y(n_549)
);

OAI21xp33_ASAP7_75t_L g550 ( 
.A1(n_518),
.A2(n_389),
.B(n_412),
.Y(n_550)
);

AOI21xp5_ASAP7_75t_L g551 ( 
.A1(n_490),
.A2(n_354),
.B(n_441),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_503),
.Y(n_552)
);

AOI21xp5_ASAP7_75t_L g553 ( 
.A1(n_511),
.A2(n_352),
.B(n_463),
.Y(n_553)
);

AOI22xp33_ASAP7_75t_SL g554 ( 
.A1(n_507),
.A2(n_369),
.B1(n_463),
.B2(n_352),
.Y(n_554)
);

AOI22xp33_ASAP7_75t_L g555 ( 
.A1(n_504),
.A2(n_458),
.B1(n_375),
.B2(n_380),
.Y(n_555)
);

INVx6_ASAP7_75t_L g556 ( 
.A(n_507),
.Y(n_556)
);

BUFx6f_ASAP7_75t_L g557 ( 
.A(n_519),
.Y(n_557)
);

BUFx3_ASAP7_75t_L g558 ( 
.A(n_497),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_504),
.Y(n_559)
);

AOI22xp33_ASAP7_75t_L g560 ( 
.A1(n_515),
.A2(n_518),
.B1(n_510),
.B2(n_487),
.Y(n_560)
);

HB1xp67_ASAP7_75t_L g561 ( 
.A(n_481),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_527),
.Y(n_562)
);

OAI22xp33_ASAP7_75t_L g563 ( 
.A1(n_525),
.A2(n_502),
.B1(n_519),
.B2(n_520),
.Y(n_563)
);

AOI22xp33_ASAP7_75t_L g564 ( 
.A1(n_522),
.A2(n_515),
.B1(n_487),
.B2(n_510),
.Y(n_564)
);

AOI22xp33_ASAP7_75t_SL g565 ( 
.A1(n_540),
.A2(n_369),
.B1(n_519),
.B2(n_510),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_526),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_535),
.Y(n_567)
);

AOI22xp33_ASAP7_75t_L g568 ( 
.A1(n_524),
.A2(n_510),
.B1(n_375),
.B2(n_380),
.Y(n_568)
);

INVx3_ASAP7_75t_L g569 ( 
.A(n_557),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_559),
.Y(n_570)
);

CKINVDCx11_ASAP7_75t_R g571 ( 
.A(n_548),
.Y(n_571)
);

OAI22xp5_ASAP7_75t_L g572 ( 
.A1(n_533),
.A2(n_511),
.B1(n_519),
.B2(n_413),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_544),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_552),
.Y(n_574)
);

AOI22xp33_ASAP7_75t_L g575 ( 
.A1(n_532),
.A2(n_486),
.B1(n_480),
.B2(n_369),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_561),
.Y(n_576)
);

BUFx2_ASAP7_75t_L g577 ( 
.A(n_538),
.Y(n_577)
);

BUFx6f_ASAP7_75t_L g578 ( 
.A(n_557),
.Y(n_578)
);

AND2x2_ASAP7_75t_L g579 ( 
.A(n_531),
.B(n_506),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_541),
.Y(n_580)
);

AOI21xp5_ASAP7_75t_L g581 ( 
.A1(n_551),
.A2(n_511),
.B(n_484),
.Y(n_581)
);

NAND3xp33_ASAP7_75t_L g582 ( 
.A(n_554),
.B(n_395),
.C(n_506),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_560),
.Y(n_583)
);

AOI22xp33_ASAP7_75t_L g584 ( 
.A1(n_530),
.A2(n_486),
.B1(n_480),
.B2(n_369),
.Y(n_584)
);

BUFx6f_ASAP7_75t_L g585 ( 
.A(n_557),
.Y(n_585)
);

INVx3_ASAP7_75t_L g586 ( 
.A(n_523),
.Y(n_586)
);

AOI22xp33_ASAP7_75t_L g587 ( 
.A1(n_543),
.A2(n_499),
.B1(n_500),
.B2(n_502),
.Y(n_587)
);

INVx2_ASAP7_75t_SL g588 ( 
.A(n_523),
.Y(n_588)
);

AOI22xp33_ASAP7_75t_L g589 ( 
.A1(n_543),
.A2(n_499),
.B1(n_500),
.B2(n_502),
.Y(n_589)
);

OAI22xp5_ASAP7_75t_L g590 ( 
.A1(n_545),
.A2(n_519),
.B1(n_447),
.B2(n_395),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_550),
.Y(n_591)
);

AOI22xp33_ASAP7_75t_L g592 ( 
.A1(n_534),
.A2(n_447),
.B1(n_519),
.B2(n_498),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_549),
.Y(n_593)
);

AOI22xp33_ASAP7_75t_L g594 ( 
.A1(n_546),
.A2(n_498),
.B1(n_386),
.B2(n_446),
.Y(n_594)
);

AND2x4_ASAP7_75t_L g595 ( 
.A(n_558),
.B(n_517),
.Y(n_595)
);

AOI22xp33_ASAP7_75t_L g596 ( 
.A1(n_546),
.A2(n_498),
.B1(n_386),
.B2(n_401),
.Y(n_596)
);

AOI22xp33_ASAP7_75t_SL g597 ( 
.A1(n_523),
.A2(n_556),
.B1(n_536),
.B2(n_528),
.Y(n_597)
);

OAI22xp5_ASAP7_75t_L g598 ( 
.A1(n_547),
.A2(n_529),
.B1(n_555),
.B2(n_556),
.Y(n_598)
);

BUFx6f_ASAP7_75t_L g599 ( 
.A(n_556),
.Y(n_599)
);

AOI22xp5_ASAP7_75t_L g600 ( 
.A1(n_542),
.A2(n_493),
.B1(n_505),
.B2(n_481),
.Y(n_600)
);

AND2x2_ASAP7_75t_L g601 ( 
.A(n_537),
.B(n_554),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_529),
.Y(n_602)
);

BUFx12f_ASAP7_75t_L g603 ( 
.A(n_521),
.Y(n_603)
);

AND2x2_ASAP7_75t_L g604 ( 
.A(n_537),
.B(n_517),
.Y(n_604)
);

BUFx3_ASAP7_75t_L g605 ( 
.A(n_536),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_553),
.Y(n_606)
);

AOI22xp33_ASAP7_75t_L g607 ( 
.A1(n_539),
.A2(n_498),
.B1(n_401),
.B2(n_357),
.Y(n_607)
);

HB1xp67_ASAP7_75t_L g608 ( 
.A(n_538),
.Y(n_608)
);

BUFx4f_ASAP7_75t_SL g609 ( 
.A(n_525),
.Y(n_609)
);

AOI22xp33_ASAP7_75t_L g610 ( 
.A1(n_522),
.A2(n_362),
.B1(n_355),
.B2(n_357),
.Y(n_610)
);

AOI22xp33_ASAP7_75t_L g611 ( 
.A1(n_580),
.A2(n_377),
.B1(n_355),
.B2(n_362),
.Y(n_611)
);

AOI22xp33_ASAP7_75t_SL g612 ( 
.A1(n_582),
.A2(n_478),
.B1(n_488),
.B2(n_477),
.Y(n_612)
);

AOI22xp33_ASAP7_75t_SL g613 ( 
.A1(n_601),
.A2(n_572),
.B1(n_590),
.B2(n_593),
.Y(n_613)
);

OAI21xp5_ASAP7_75t_SL g614 ( 
.A1(n_597),
.A2(n_505),
.B(n_494),
.Y(n_614)
);

AOI22xp33_ASAP7_75t_L g615 ( 
.A1(n_583),
.A2(n_366),
.B1(n_371),
.B2(n_415),
.Y(n_615)
);

AOI22xp33_ASAP7_75t_SL g616 ( 
.A1(n_601),
.A2(n_478),
.B1(n_488),
.B2(n_477),
.Y(n_616)
);

AOI22xp33_ASAP7_75t_L g617 ( 
.A1(n_579),
.A2(n_366),
.B1(n_415),
.B2(n_410),
.Y(n_617)
);

AOI22xp33_ASAP7_75t_SL g618 ( 
.A1(n_579),
.A2(n_478),
.B1(n_477),
.B2(n_438),
.Y(n_618)
);

AND2x2_ASAP7_75t_L g619 ( 
.A(n_566),
.B(n_517),
.Y(n_619)
);

AOI22xp33_ASAP7_75t_L g620 ( 
.A1(n_568),
.A2(n_415),
.B1(n_410),
.B2(n_388),
.Y(n_620)
);

AOI222xp33_ASAP7_75t_L g621 ( 
.A1(n_591),
.A2(n_493),
.B1(n_387),
.B2(n_388),
.C1(n_414),
.C2(n_438),
.Y(n_621)
);

AOI221xp5_ASAP7_75t_L g622 ( 
.A1(n_567),
.A2(n_494),
.B1(n_493),
.B2(n_387),
.C(n_378),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_562),
.Y(n_623)
);

AND2x2_ASAP7_75t_L g624 ( 
.A(n_573),
.B(n_516),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_608),
.B(n_516),
.Y(n_625)
);

AOI22xp5_ASAP7_75t_L g626 ( 
.A1(n_598),
.A2(n_477),
.B1(n_351),
.B2(n_484),
.Y(n_626)
);

OA21x2_ASAP7_75t_L g627 ( 
.A1(n_606),
.A2(n_402),
.B(n_385),
.Y(n_627)
);

AOI221xp5_ASAP7_75t_L g628 ( 
.A1(n_574),
.A2(n_399),
.B1(n_415),
.B2(n_391),
.C(n_516),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_562),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_570),
.Y(n_630)
);

OAI22xp5_ASAP7_75t_L g631 ( 
.A1(n_594),
.A2(n_484),
.B1(n_516),
.B2(n_512),
.Y(n_631)
);

AOI22xp33_ASAP7_75t_L g632 ( 
.A1(n_564),
.A2(n_415),
.B1(n_351),
.B2(n_472),
.Y(n_632)
);

AOI22xp33_ASAP7_75t_L g633 ( 
.A1(n_584),
.A2(n_351),
.B1(n_399),
.B2(n_391),
.Y(n_633)
);

AOI22xp33_ASAP7_75t_SL g634 ( 
.A1(n_599),
.A2(n_512),
.B1(n_484),
.B2(n_351),
.Y(n_634)
);

OAI22xp5_ASAP7_75t_L g635 ( 
.A1(n_596),
.A2(n_391),
.B1(n_403),
.B2(n_406),
.Y(n_635)
);

AOI22xp33_ASAP7_75t_L g636 ( 
.A1(n_610),
.A2(n_399),
.B1(n_403),
.B2(n_411),
.Y(n_636)
);

AOI22xp33_ASAP7_75t_L g637 ( 
.A1(n_565),
.A2(n_403),
.B1(n_411),
.B2(n_379),
.Y(n_637)
);

AND2x2_ASAP7_75t_L g638 ( 
.A(n_577),
.B(n_604),
.Y(n_638)
);

OAI22xp5_ASAP7_75t_L g639 ( 
.A1(n_577),
.A2(n_411),
.B1(n_379),
.B2(n_402),
.Y(n_639)
);

AOI22xp5_ASAP7_75t_L g640 ( 
.A1(n_600),
.A2(n_411),
.B1(n_379),
.B2(n_62),
.Y(n_640)
);

AOI22xp33_ASAP7_75t_L g641 ( 
.A1(n_587),
.A2(n_411),
.B1(n_379),
.B2(n_65),
.Y(n_641)
);

AOI22xp33_ASAP7_75t_L g642 ( 
.A1(n_589),
.A2(n_59),
.B1(n_60),
.B2(n_66),
.Y(n_642)
);

AOI22xp5_ASAP7_75t_L g643 ( 
.A1(n_563),
.A2(n_67),
.B1(n_68),
.B2(n_69),
.Y(n_643)
);

AND2x2_ASAP7_75t_L g644 ( 
.A(n_604),
.B(n_70),
.Y(n_644)
);

AND2x2_ASAP7_75t_L g645 ( 
.A(n_576),
.B(n_71),
.Y(n_645)
);

OAI222xp33_ASAP7_75t_L g646 ( 
.A1(n_592),
.A2(n_575),
.B1(n_607),
.B2(n_570),
.C1(n_588),
.C2(n_602),
.Y(n_646)
);

AOI22xp33_ASAP7_75t_L g647 ( 
.A1(n_599),
.A2(n_72),
.B1(n_73),
.B2(n_78),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_606),
.Y(n_648)
);

AND2x2_ASAP7_75t_L g649 ( 
.A(n_638),
.B(n_605),
.Y(n_649)
);

NAND3xp33_ASAP7_75t_L g650 ( 
.A(n_613),
.B(n_581),
.C(n_599),
.Y(n_650)
);

AND2x2_ASAP7_75t_L g651 ( 
.A(n_638),
.B(n_605),
.Y(n_651)
);

AND2x2_ASAP7_75t_L g652 ( 
.A(n_619),
.B(n_595),
.Y(n_652)
);

AOI221xp5_ASAP7_75t_L g653 ( 
.A1(n_619),
.A2(n_595),
.B1(n_588),
.B2(n_586),
.C(n_599),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_625),
.B(n_595),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_SL g655 ( 
.A(n_612),
.B(n_585),
.Y(n_655)
);

NAND3xp33_ASAP7_75t_L g656 ( 
.A(n_645),
.B(n_599),
.C(n_578),
.Y(n_656)
);

AOI22xp33_ASAP7_75t_L g657 ( 
.A1(n_621),
.A2(n_586),
.B1(n_603),
.B2(n_609),
.Y(n_657)
);

NAND3xp33_ASAP7_75t_L g658 ( 
.A(n_645),
.B(n_585),
.C(n_578),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_624),
.B(n_586),
.Y(n_659)
);

AND2x2_ASAP7_75t_L g660 ( 
.A(n_624),
.B(n_569),
.Y(n_660)
);

OAI22xp5_ASAP7_75t_SL g661 ( 
.A1(n_640),
.A2(n_603),
.B1(n_571),
.B2(n_578),
.Y(n_661)
);

NOR2xp33_ASAP7_75t_L g662 ( 
.A(n_614),
.B(n_571),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_644),
.B(n_569),
.Y(n_663)
);

OAI22xp5_ASAP7_75t_L g664 ( 
.A1(n_641),
.A2(n_569),
.B1(n_585),
.B2(n_578),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_644),
.B(n_578),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_SL g666 ( 
.A(n_618),
.B(n_585),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_SL g667 ( 
.A(n_616),
.B(n_585),
.Y(n_667)
);

NAND3xp33_ASAP7_75t_L g668 ( 
.A(n_622),
.B(n_80),
.C(n_83),
.Y(n_668)
);

NAND3xp33_ASAP7_75t_L g669 ( 
.A(n_628),
.B(n_84),
.C(n_85),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_629),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_617),
.B(n_629),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_623),
.B(n_144),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_623),
.B(n_86),
.Y(n_673)
);

NAND3xp33_ASAP7_75t_L g674 ( 
.A(n_643),
.B(n_642),
.C(n_626),
.Y(n_674)
);

NAND2xp33_ASAP7_75t_SL g675 ( 
.A(n_631),
.B(n_87),
.Y(n_675)
);

AOI21xp5_ASAP7_75t_SL g676 ( 
.A1(n_635),
.A2(n_88),
.B(n_90),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_670),
.Y(n_677)
);

NOR3xp33_ASAP7_75t_SL g678 ( 
.A(n_662),
.B(n_646),
.C(n_639),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_654),
.B(n_648),
.Y(n_679)
);

AND2x2_ASAP7_75t_L g680 ( 
.A(n_652),
.B(n_648),
.Y(n_680)
);

OAI21xp5_ASAP7_75t_L g681 ( 
.A1(n_668),
.A2(n_647),
.B(n_634),
.Y(n_681)
);

NAND4xp75_ASAP7_75t_L g682 ( 
.A(n_662),
.B(n_630),
.C(n_627),
.D(n_637),
.Y(n_682)
);

NAND3xp33_ASAP7_75t_L g683 ( 
.A(n_650),
.B(n_611),
.C(n_636),
.Y(n_683)
);

OR2x2_ASAP7_75t_L g684 ( 
.A(n_659),
.B(n_630),
.Y(n_684)
);

AND2x4_ASAP7_75t_L g685 ( 
.A(n_660),
.B(n_649),
.Y(n_685)
);

NOR2x1_ASAP7_75t_R g686 ( 
.A(n_651),
.B(n_632),
.Y(n_686)
);

NOR2xp33_ASAP7_75t_L g687 ( 
.A(n_663),
.B(n_92),
.Y(n_687)
);

AOI22xp33_ASAP7_75t_L g688 ( 
.A1(n_674),
.A2(n_675),
.B1(n_657),
.B2(n_661),
.Y(n_688)
);

AOI22xp33_ASAP7_75t_L g689 ( 
.A1(n_675),
.A2(n_615),
.B1(n_620),
.B2(n_633),
.Y(n_689)
);

AOI22xp33_ASAP7_75t_L g690 ( 
.A1(n_671),
.A2(n_627),
.B1(n_94),
.B2(n_97),
.Y(n_690)
);

AND2x2_ASAP7_75t_L g691 ( 
.A(n_665),
.B(n_627),
.Y(n_691)
);

AND2x2_ASAP7_75t_L g692 ( 
.A(n_658),
.B(n_93),
.Y(n_692)
);

AOI22xp33_ASAP7_75t_L g693 ( 
.A1(n_667),
.A2(n_99),
.B1(n_103),
.B2(n_104),
.Y(n_693)
);

INVxp67_ASAP7_75t_L g694 ( 
.A(n_656),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_677),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_691),
.Y(n_696)
);

AOI21xp5_ASAP7_75t_L g697 ( 
.A1(n_688),
.A2(n_655),
.B(n_667),
.Y(n_697)
);

BUFx3_ASAP7_75t_L g698 ( 
.A(n_692),
.Y(n_698)
);

XOR2x2_ASAP7_75t_L g699 ( 
.A(n_682),
.B(n_655),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_684),
.Y(n_700)
);

OR2x2_ASAP7_75t_L g701 ( 
.A(n_684),
.B(n_666),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_679),
.Y(n_702)
);

AND2x2_ASAP7_75t_L g703 ( 
.A(n_685),
.B(n_666),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_694),
.B(n_653),
.Y(n_704)
);

HB1xp67_ASAP7_75t_L g705 ( 
.A(n_691),
.Y(n_705)
);

XNOR2xp5_ASAP7_75t_L g706 ( 
.A(n_699),
.B(n_685),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_695),
.Y(n_707)
);

AND2x2_ASAP7_75t_L g708 ( 
.A(n_705),
.B(n_685),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_701),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_702),
.Y(n_710)
);

OA22x2_ASAP7_75t_L g711 ( 
.A1(n_706),
.A2(n_709),
.B1(n_704),
.B2(n_703),
.Y(n_711)
);

OA22x2_ASAP7_75t_L g712 ( 
.A1(n_709),
.A2(n_703),
.B1(n_696),
.B2(n_699),
.Y(n_712)
);

AOI22x1_ASAP7_75t_L g713 ( 
.A1(n_708),
.A2(n_697),
.B1(n_707),
.B2(n_710),
.Y(n_713)
);

CKINVDCx20_ASAP7_75t_R g714 ( 
.A(n_708),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_707),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_715),
.Y(n_716)
);

INVxp67_ASAP7_75t_L g717 ( 
.A(n_713),
.Y(n_717)
);

INVxp67_ASAP7_75t_L g718 ( 
.A(n_711),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_714),
.Y(n_719)
);

AOI22xp5_ASAP7_75t_L g720 ( 
.A1(n_718),
.A2(n_712),
.B1(n_682),
.B2(n_698),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_716),
.Y(n_721)
);

AOI22xp5_ASAP7_75t_L g722 ( 
.A1(n_717),
.A2(n_698),
.B1(n_678),
.B2(n_683),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_721),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_722),
.Y(n_724)
);

A2O1A1Ixp33_ASAP7_75t_L g725 ( 
.A1(n_720),
.A2(n_719),
.B(n_681),
.C(n_687),
.Y(n_725)
);

BUFx2_ASAP7_75t_L g726 ( 
.A(n_721),
.Y(n_726)
);

AOI22xp5_ASAP7_75t_L g727 ( 
.A1(n_725),
.A2(n_696),
.B1(n_692),
.B2(n_701),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_SL g728 ( 
.A(n_724),
.B(n_700),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_726),
.Y(n_729)
);

AOI22xp5_ASAP7_75t_L g730 ( 
.A1(n_725),
.A2(n_689),
.B1(n_693),
.B2(n_690),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_723),
.B(n_680),
.Y(n_731)
);

AOI221xp5_ASAP7_75t_L g732 ( 
.A1(n_725),
.A2(n_676),
.B1(n_664),
.B2(n_669),
.C(n_673),
.Y(n_732)
);

AOI221xp5_ASAP7_75t_L g733 ( 
.A1(n_725),
.A2(n_672),
.B1(n_680),
.B2(n_686),
.C(n_111),
.Y(n_733)
);

INVx1_ASAP7_75t_SL g734 ( 
.A(n_729),
.Y(n_734)
);

AOI22xp5_ASAP7_75t_L g735 ( 
.A1(n_733),
.A2(n_106),
.B1(n_107),
.B2(n_110),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_728),
.B(n_731),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_727),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_730),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_732),
.Y(n_739)
);

AOI22xp5_ASAP7_75t_L g740 ( 
.A1(n_733),
.A2(n_112),
.B1(n_114),
.B2(n_116),
.Y(n_740)
);

BUFx6f_ASAP7_75t_L g741 ( 
.A(n_736),
.Y(n_741)
);

NOR2x1_ASAP7_75t_L g742 ( 
.A(n_734),
.B(n_118),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_739),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_738),
.Y(n_744)
);

AND2x4_ASAP7_75t_L g745 ( 
.A(n_737),
.B(n_119),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_735),
.Y(n_746)
);

BUFx2_ASAP7_75t_L g747 ( 
.A(n_740),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_741),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_741),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_744),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_742),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_743),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_747),
.Y(n_753)
);

AOI22xp5_ASAP7_75t_L g754 ( 
.A1(n_751),
.A2(n_746),
.B1(n_747),
.B2(n_745),
.Y(n_754)
);

AO22x1_ASAP7_75t_L g755 ( 
.A1(n_748),
.A2(n_120),
.B1(n_122),
.B2(n_124),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_753),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_748),
.Y(n_757)
);

HB1xp67_ASAP7_75t_L g758 ( 
.A(n_750),
.Y(n_758)
);

NAND4xp25_ASAP7_75t_L g759 ( 
.A(n_749),
.B(n_125),
.C(n_127),
.D(n_128),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_758),
.Y(n_760)
);

INVx4_ASAP7_75t_L g761 ( 
.A(n_756),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_757),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_754),
.Y(n_763)
);

AOI22xp33_ASAP7_75t_L g764 ( 
.A1(n_760),
.A2(n_752),
.B1(n_759),
.B2(n_755),
.Y(n_764)
);

AOI22xp5_ASAP7_75t_L g765 ( 
.A1(n_761),
.A2(n_129),
.B1(n_130),
.B2(n_131),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_764),
.Y(n_766)
);

AOI22xp5_ASAP7_75t_L g767 ( 
.A1(n_766),
.A2(n_762),
.B1(n_763),
.B2(n_765),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_767),
.Y(n_768)
);

AOI221xp5_ASAP7_75t_L g769 ( 
.A1(n_768),
.A2(n_132),
.B1(n_133),
.B2(n_135),
.C(n_136),
.Y(n_769)
);

AOI22xp33_ASAP7_75t_L g770 ( 
.A1(n_769),
.A2(n_137),
.B1(n_138),
.B2(n_140),
.Y(n_770)
);


endmodule