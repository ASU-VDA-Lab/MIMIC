module fake_jpeg_11802_n_340 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_340);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_340;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_260;
wire n_199;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_3),
.B(n_9),
.Y(n_18)
);

INVx8_ASAP7_75t_SL g19 ( 
.A(n_1),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx11_ASAP7_75t_SL g29 ( 
.A(n_12),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_10),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_12),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_7),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

AOI21xp33_ASAP7_75t_L g37 ( 
.A1(n_18),
.A2(n_0),
.B(n_2),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_0),
.Y(n_50)
);

INVx3_ASAP7_75t_SL g38 ( 
.A(n_19),
.Y(n_38)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVx2_ASAP7_75t_SL g59 ( 
.A(n_39),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

INVx1_ASAP7_75t_SL g60 ( 
.A(n_40),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_21),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_41),
.A2(n_35),
.B1(n_26),
.B2(n_30),
.Y(n_70)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_41),
.B(n_18),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_48),
.B(n_56),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_49),
.B(n_50),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_37),
.B(n_35),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_53),
.B(n_54),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_38),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_36),
.B(n_32),
.Y(n_56)
);

BUFx2_ASAP7_75t_R g57 ( 
.A(n_38),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_57),
.B(n_42),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_43),
.A2(n_20),
.B1(n_23),
.B2(n_33),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_61),
.A2(n_71),
.B1(n_23),
.B2(n_20),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_40),
.B(n_31),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_63),
.B(n_66),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_40),
.B(n_31),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_40),
.B(n_31),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_68),
.B(n_69),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_40),
.B(n_35),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_70),
.A2(n_26),
.B1(n_30),
.B2(n_34),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_43),
.A2(n_20),
.B1(n_23),
.B2(n_22),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_38),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_72),
.B(n_17),
.Y(n_101)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_65),
.Y(n_73)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_73),
.Y(n_129)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_65),
.Y(n_74)
);

BUFx5_ASAP7_75t_L g122 ( 
.A(n_74),
.Y(n_122)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_65),
.Y(n_75)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_75),
.Y(n_108)
);

INVx2_ASAP7_75t_SL g76 ( 
.A(n_55),
.Y(n_76)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_76),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_61),
.A2(n_46),
.B1(n_47),
.B2(n_45),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_77),
.A2(n_81),
.B1(n_59),
.B2(n_60),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_78),
.A2(n_87),
.B1(n_91),
.B2(n_103),
.Y(n_114)
);

AO22x1_ASAP7_75t_SL g79 ( 
.A1(n_48),
.A2(n_44),
.B1(n_19),
.B2(n_34),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_79),
.B(n_72),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_63),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_80),
.B(n_92),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_53),
.A2(n_42),
.B1(n_39),
.B2(n_30),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_82),
.Y(n_111)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_51),
.Y(n_83)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_83),
.Y(n_112)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_55),
.Y(n_85)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_85),
.Y(n_118)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_51),
.Y(n_86)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_86),
.Y(n_123)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_65),
.Y(n_88)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_88),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_56),
.B(n_39),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_89),
.B(n_95),
.C(n_58),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_60),
.A2(n_24),
.B1(n_25),
.B2(n_27),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_90),
.A2(n_57),
.B1(n_59),
.B2(n_17),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_48),
.A2(n_46),
.B1(n_22),
.B2(n_33),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_55),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_66),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_94),
.B(n_98),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_52),
.B(n_46),
.C(n_33),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_68),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_52),
.A2(n_17),
.B1(n_29),
.B2(n_33),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_100),
.A2(n_102),
.B1(n_26),
.B2(n_34),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_101),
.B(n_54),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_64),
.A2(n_17),
.B1(n_29),
.B2(n_27),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_70),
.A2(n_50),
.B1(n_71),
.B2(n_69),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_105),
.B(n_119),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_106),
.B(n_113),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_96),
.B(n_70),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_107),
.B(n_116),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_96),
.B(n_80),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_103),
.A2(n_64),
.B1(n_51),
.B2(n_62),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_115),
.A2(n_121),
.B1(n_77),
.B2(n_76),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_98),
.B(n_62),
.Y(n_116)
);

NOR2xp67_ASAP7_75t_SL g117 ( 
.A(n_93),
.B(n_57),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_117),
.A2(n_128),
.B(n_82),
.Y(n_144)
);

MAJx2_ASAP7_75t_L g120 ( 
.A(n_93),
.B(n_60),
.C(n_59),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_120),
.B(n_92),
.C(n_85),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_91),
.A2(n_62),
.B1(n_59),
.B2(n_58),
.Y(n_121)
);

OAI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_125),
.A2(n_75),
.B1(n_88),
.B2(n_74),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_126),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_101),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_127),
.B(n_131),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_89),
.A2(n_58),
.B1(n_27),
.B2(n_65),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_130),
.B(n_67),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_87),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_97),
.B(n_67),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_132),
.B(n_76),
.Y(n_154)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_118),
.Y(n_135)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_135),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_104),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_136),
.B(n_141),
.Y(n_167)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_118),
.Y(n_138)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_138),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_105),
.A2(n_84),
.B(n_82),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_139),
.A2(n_140),
.B(n_150),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_117),
.A2(n_84),
.B(n_99),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_104),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_109),
.B(n_99),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_142),
.B(n_145),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_144),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_109),
.B(n_97),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_146),
.A2(n_157),
.B1(n_159),
.B2(n_119),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_113),
.B(n_89),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_147),
.B(n_156),
.Y(n_182)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_112),
.Y(n_148)
);

INVx1_ASAP7_75t_SL g184 ( 
.A(n_148),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_116),
.B(n_79),
.Y(n_149)
);

NAND3xp33_ASAP7_75t_L g195 ( 
.A(n_149),
.B(n_161),
.C(n_163),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_111),
.A2(n_89),
.B(n_82),
.Y(n_150)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_110),
.Y(n_152)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_152),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_131),
.A2(n_78),
.B1(n_95),
.B2(n_79),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_153),
.A2(n_121),
.B1(n_128),
.B2(n_125),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_154),
.B(n_123),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_132),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_155),
.B(n_110),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_127),
.B(n_79),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_114),
.A2(n_100),
.B1(n_102),
.B2(n_76),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_158),
.B(n_67),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_114),
.A2(n_86),
.B1(n_83),
.B2(n_25),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_160),
.A2(n_124),
.B1(n_108),
.B2(n_128),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_106),
.B(n_74),
.Y(n_161)
);

INVx6_ASAP7_75t_L g162 ( 
.A(n_122),
.Y(n_162)
);

INVx5_ASAP7_75t_L g177 ( 
.A(n_162),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_107),
.B(n_73),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_164),
.B(n_120),
.C(n_108),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_166),
.A2(n_168),
.B1(n_186),
.B2(n_187),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_134),
.A2(n_130),
.B1(n_115),
.B2(n_120),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_140),
.A2(n_130),
.B(n_126),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_169),
.A2(n_0),
.B(n_4),
.Y(n_226)
);

CKINVDCx14_ASAP7_75t_R g224 ( 
.A(n_170),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_172),
.A2(n_191),
.B1(n_194),
.B2(n_157),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_136),
.B(n_123),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_173),
.B(n_179),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_174),
.B(n_188),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_176),
.A2(n_139),
.B(n_149),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_178),
.B(n_189),
.C(n_164),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_141),
.B(n_112),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_162),
.A2(n_129),
.B1(n_124),
.B2(n_126),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_181),
.A2(n_162),
.B1(n_152),
.B2(n_148),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_134),
.A2(n_129),
.B1(n_73),
.B2(n_75),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_134),
.A2(n_88),
.B1(n_25),
.B2(n_122),
.Y(n_187)
);

A2O1A1Ixp33_ASAP7_75t_L g188 ( 
.A1(n_151),
.A2(n_16),
.B(n_15),
.C(n_14),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_133),
.B(n_67),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_190),
.B(n_193),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_153),
.A2(n_67),
.B1(n_25),
.B2(n_122),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_142),
.B(n_16),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_192),
.B(n_196),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_133),
.B(n_16),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_153),
.A2(n_15),
.B1(n_14),
.B2(n_13),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_137),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_135),
.Y(n_197)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_197),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_137),
.B(n_145),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_198),
.B(n_147),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_200),
.B(n_225),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_183),
.A2(n_143),
.B1(n_134),
.B2(n_160),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_201),
.A2(n_184),
.B(n_177),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_172),
.A2(n_143),
.B1(n_159),
.B2(n_155),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_204),
.B(n_206),
.Y(n_242)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_180),
.Y(n_205)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_205),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_196),
.A2(n_151),
.B1(n_156),
.B2(n_146),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_170),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_207),
.B(n_179),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_208),
.B(n_223),
.C(n_165),
.Y(n_228)
);

AO22x1_ASAP7_75t_SL g209 ( 
.A1(n_182),
.A2(n_166),
.B1(n_168),
.B2(n_195),
.Y(n_209)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_209),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_210),
.A2(n_220),
.B(n_187),
.Y(n_237)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_180),
.Y(n_211)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_211),
.Y(n_245)
);

OAI21xp33_ASAP7_75t_SL g212 ( 
.A1(n_165),
.A2(n_139),
.B(n_154),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_212),
.B(n_226),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_191),
.A2(n_158),
.B1(n_164),
.B2(n_138),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_213),
.B(n_219),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_214),
.B(n_173),
.Y(n_241)
);

AOI322xp5_ASAP7_75t_L g218 ( 
.A1(n_185),
.A2(n_163),
.A3(n_144),
.B1(n_161),
.B2(n_150),
.C1(n_158),
.C2(n_164),
.Y(n_218)
);

NOR4xp25_ASAP7_75t_L g243 ( 
.A(n_218),
.B(n_174),
.C(n_188),
.D(n_194),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_167),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_176),
.A2(n_14),
.B1(n_13),
.B2(n_4),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_221),
.B(n_222),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_169),
.A2(n_28),
.B1(n_3),
.B2(n_4),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_189),
.B(n_28),
.C(n_3),
.Y(n_223)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_171),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_167),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_227),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_228),
.B(n_230),
.C(n_232),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_208),
.B(n_178),
.C(n_182),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_210),
.A2(n_198),
.B(n_185),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_231),
.B(n_247),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_214),
.B(n_213),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_219),
.Y(n_235)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_235),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_237),
.A2(n_200),
.B1(n_204),
.B2(n_222),
.Y(n_259)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_238),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_227),
.B(n_193),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_239),
.B(n_240),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_215),
.B(n_190),
.Y(n_240)
);

CKINVDCx14_ASAP7_75t_R g265 ( 
.A(n_241),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_SL g254 ( 
.A(n_243),
.B(n_209),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_209),
.B(n_197),
.C(n_175),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_246),
.B(n_253),
.C(n_223),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_207),
.B(n_175),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_201),
.A2(n_186),
.B(n_171),
.Y(n_250)
);

INVxp33_ASAP7_75t_L g266 ( 
.A(n_250),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_251),
.B(n_226),
.Y(n_260)
);

BUFx5_ASAP7_75t_L g252 ( 
.A(n_202),
.Y(n_252)
);

INVx1_ASAP7_75t_SL g261 ( 
.A(n_252),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_206),
.B(n_184),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_254),
.B(n_233),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_242),
.A2(n_216),
.B1(n_236),
.B2(n_244),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_255),
.A2(n_256),
.B1(n_234),
.B2(n_241),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_242),
.A2(n_216),
.B1(n_224),
.B2(n_209),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_259),
.A2(n_229),
.B1(n_235),
.B2(n_237),
.Y(n_277)
);

AND2x2_ASAP7_75t_SL g284 ( 
.A(n_260),
.B(n_263),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_262),
.B(n_231),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_229),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_230),
.B(n_203),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_264),
.B(n_267),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_232),
.B(n_203),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_249),
.A2(n_199),
.B1(n_217),
.B2(n_211),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_268),
.A2(n_272),
.B1(n_245),
.B2(n_248),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_228),
.B(n_225),
.C(n_202),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_270),
.B(n_273),
.C(n_247),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_249),
.A2(n_199),
.B1(n_217),
.B2(n_205),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_244),
.B(n_221),
.C(n_177),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_SL g275 ( 
.A1(n_263),
.A2(n_246),
.B(n_236),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_275),
.B(n_277),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_276),
.B(n_278),
.C(n_286),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_262),
.B(n_253),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_279),
.A2(n_258),
.B(n_270),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_280),
.B(n_255),
.C(n_267),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_256),
.A2(n_271),
.B1(n_273),
.B2(n_274),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_281),
.A2(n_289),
.B1(n_265),
.B2(n_284),
.Y(n_294)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_269),
.Y(n_283)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_283),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_257),
.B(n_235),
.C(n_250),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_285),
.B(n_287),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_264),
.B(n_233),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_261),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_261),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_288),
.B(n_290),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_257),
.B(n_251),
.C(n_234),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_291),
.B(n_5),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_292),
.B(n_282),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_293),
.B(n_294),
.Y(n_310)
);

O2A1O1Ixp33_ASAP7_75t_L g295 ( 
.A1(n_284),
.A2(n_266),
.B(n_260),
.C(n_254),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_295),
.A2(n_286),
.B(n_278),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_285),
.B(n_266),
.C(n_248),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_297),
.B(n_305),
.Y(n_315)
);

A2O1A1Ixp33_ASAP7_75t_SL g300 ( 
.A1(n_275),
.A2(n_245),
.B(n_252),
.C(n_243),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_300),
.B(n_6),
.C(n_7),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_276),
.B(n_5),
.C(n_6),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_301),
.B(n_5),
.Y(n_313)
);

BUFx24_ASAP7_75t_SL g303 ( 
.A(n_282),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_303),
.B(n_306),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_291),
.A2(n_5),
.B(n_6),
.Y(n_305)
);

NAND2xp33_ASAP7_75t_SL g307 ( 
.A(n_296),
.B(n_284),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_307),
.B(n_308),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_SL g308 ( 
.A1(n_302),
.A2(n_277),
.B(n_280),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_304),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_309),
.B(n_312),
.Y(n_326)
);

CKINVDCx16_ASAP7_75t_R g322 ( 
.A(n_311),
.Y(n_322)
);

NOR4xp25_ASAP7_75t_L g327 ( 
.A(n_313),
.B(n_8),
.C(n_318),
.D(n_310),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_314),
.A2(n_316),
.B1(n_298),
.B2(n_300),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_296),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_293),
.B(n_299),
.C(n_297),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_SL g325 ( 
.A1(n_317),
.A2(n_8),
.B(n_11),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_319),
.B(n_324),
.Y(n_331)
);

AOI322xp5_ASAP7_75t_L g320 ( 
.A1(n_315),
.A2(n_300),
.A3(n_295),
.B1(n_10),
.B2(n_11),
.C1(n_12),
.C2(n_9),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g333 ( 
.A(n_320),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_314),
.A2(n_300),
.B1(n_9),
.B2(n_11),
.Y(n_323)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_323),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_SL g324 ( 
.A1(n_307),
.A2(n_8),
.B(n_11),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_325),
.B(n_324),
.C(n_323),
.Y(n_330)
);

NOR2xp67_ASAP7_75t_L g328 ( 
.A(n_327),
.B(n_316),
.Y(n_328)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_328),
.Y(n_336)
);

INVxp67_ASAP7_75t_SL g329 ( 
.A(n_321),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_329),
.B(n_330),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_SL g334 ( 
.A1(n_329),
.A2(n_322),
.B(n_317),
.Y(n_334)
);

OAI21x1_ASAP7_75t_L g337 ( 
.A1(n_334),
.A2(n_326),
.B(n_331),
.Y(n_337)
);

AOI321xp33_ASAP7_75t_L g338 ( 
.A1(n_337),
.A2(n_336),
.A3(n_335),
.B1(n_332),
.B2(n_312),
.C(n_311),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_338),
.B(n_319),
.C(n_333),
.Y(n_339)
);

HB1xp67_ASAP7_75t_L g340 ( 
.A(n_339),
.Y(n_340)
);


endmodule