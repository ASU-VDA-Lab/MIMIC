module fake_jpeg_23083_n_280 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_280);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_280;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_240;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

BUFx5_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_2),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx3_ASAP7_75t_SL g22 ( 
.A(n_14),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx10_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_35),
.B(n_24),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_29),
.B(n_0),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_36),
.B(n_40),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_18),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_37),
.B(n_38),
.Y(n_62)
);

INVx2_ASAP7_75t_SL g38 ( 
.A(n_22),
.Y(n_38)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_29),
.B(n_1),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_24),
.B(n_30),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_43),
.B(n_35),
.C(n_20),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_44),
.Y(n_89)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

INVx11_ASAP7_75t_L g101 ( 
.A(n_45),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_43),
.A2(n_29),
.B1(n_28),
.B2(n_20),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_47),
.A2(n_48),
.B1(n_20),
.B2(n_21),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_43),
.A2(n_28),
.B1(n_21),
.B2(n_20),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_49),
.B(n_56),
.Y(n_79)
);

AOI21xp33_ASAP7_75t_L g51 ( 
.A1(n_36),
.A2(n_40),
.B(n_37),
.Y(n_51)
);

A2O1A1Ixp33_ASAP7_75t_L g75 ( 
.A1(n_51),
.A2(n_18),
.B(n_24),
.C(n_17),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_52),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_39),
.A2(n_28),
.B1(n_31),
.B2(n_19),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_53),
.A2(n_59),
.B1(n_31),
.B2(n_21),
.Y(n_71)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_57),
.B(n_60),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_43),
.B(n_34),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_58),
.B(n_31),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_39),
.A2(n_31),
.B1(n_17),
.B2(n_21),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_61),
.B(n_33),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_63),
.B(n_22),
.C(n_25),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_35),
.B(n_33),
.Y(n_64)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_64),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_65),
.B(n_100),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_67),
.A2(n_78),
.B1(n_50),
.B2(n_22),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_63),
.A2(n_42),
.B1(n_21),
.B2(n_17),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_68),
.A2(n_71),
.B1(n_76),
.B2(n_84),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

BUFx2_ASAP7_75t_SL g118 ( 
.A(n_69),
.Y(n_118)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

INVx11_ASAP7_75t_L g108 ( 
.A(n_70),
.Y(n_108)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_72),
.B(n_73),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_61),
.B(n_19),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_74),
.B(n_75),
.Y(n_102)
);

OA22x2_ASAP7_75t_L g76 ( 
.A1(n_48),
.A2(n_38),
.B1(n_41),
.B2(n_42),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_49),
.A2(n_42),
.B1(n_34),
.B2(n_32),
.Y(n_78)
);

OAI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_56),
.A2(n_42),
.B1(n_27),
.B2(n_26),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g122 ( 
.A1(n_81),
.A2(n_90),
.B1(n_22),
.B2(n_5),
.Y(n_122)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_46),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_82),
.B(n_85),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_58),
.B(n_1),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_83),
.B(n_4),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_62),
.A2(n_26),
.B1(n_23),
.B2(n_32),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_44),
.Y(n_85)
);

CKINVDCx9p33_ASAP7_75t_R g86 ( 
.A(n_57),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_86),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_62),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_87),
.B(n_88),
.Y(n_107)
);

OR2x2_ASAP7_75t_L g88 ( 
.A(n_54),
.B(n_41),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_54),
.A2(n_27),
.B1(n_25),
.B2(n_23),
.Y(n_90)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_55),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_91),
.B(n_92),
.Y(n_114)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_46),
.Y(n_92)
);

BUFx12_ASAP7_75t_L g93 ( 
.A(n_45),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_93),
.B(n_94),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_50),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_60),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_95),
.B(n_97),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_96),
.B(n_22),
.C(n_38),
.Y(n_117)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_52),
.Y(n_97)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_52),
.Y(n_98)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_98),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_55),
.B(n_3),
.Y(n_99)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_99),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_50),
.B(n_3),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_96),
.B(n_41),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_106),
.B(n_117),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_110),
.A2(n_115),
.B1(n_120),
.B2(n_98),
.Y(n_146)
);

NOR2x1_ASAP7_75t_L g112 ( 
.A(n_88),
.B(n_41),
.Y(n_112)
);

NOR2x1_ASAP7_75t_L g154 ( 
.A(n_112),
.B(n_101),
.Y(n_154)
);

AOI21xp33_ASAP7_75t_L g113 ( 
.A1(n_79),
.A2(n_24),
.B(n_16),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_SL g138 ( 
.A(n_113),
.B(n_121),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_70),
.A2(n_38),
.B1(n_30),
.B2(n_22),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_83),
.B(n_65),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_116),
.B(n_128),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_67),
.A2(n_75),
.B1(n_76),
.B2(n_68),
.Y(n_120)
);

MAJx2_ASAP7_75t_L g121 ( 
.A(n_65),
.B(n_22),
.C(n_5),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_122),
.B(n_127),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_SL g155 ( 
.A(n_123),
.B(n_6),
.Y(n_155)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_69),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_83),
.B(n_77),
.Y(n_128)
);

AO22x2_ASAP7_75t_L g129 ( 
.A1(n_76),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_129),
.A2(n_91),
.B1(n_94),
.B2(n_92),
.Y(n_134)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_126),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_130),
.B(n_131),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_118),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_104),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_132),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_103),
.B(n_84),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_133),
.B(n_135),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_134),
.A2(n_148),
.B1(n_89),
.B2(n_80),
.Y(n_170)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_114),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_112),
.A2(n_76),
.B(n_86),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_136),
.A2(n_123),
.B(n_7),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_107),
.B(n_66),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_137),
.B(n_139),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_119),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_115),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_140),
.B(n_144),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_105),
.B(n_93),
.Y(n_143)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_143),
.Y(n_168)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_129),
.Y(n_144)
);

BUFx2_ASAP7_75t_L g145 ( 
.A(n_111),
.Y(n_145)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_145),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_146),
.A2(n_108),
.B1(n_124),
.B2(n_117),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_102),
.B(n_93),
.Y(n_147)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_147),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_108),
.A2(n_101),
.B1(n_97),
.B2(n_80),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_111),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_149),
.A2(n_150),
.B1(n_152),
.B2(n_156),
.Y(n_167)
);

INVx3_ASAP7_75t_SL g150 ( 
.A(n_127),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_129),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_151),
.B(n_153),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_129),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_106),
.B(n_102),
.Y(n_153)
);

NAND2xp33_ASAP7_75t_SL g162 ( 
.A(n_154),
.B(n_125),
.Y(n_162)
);

OA21x2_ASAP7_75t_SL g185 ( 
.A1(n_155),
.A2(n_9),
.B(n_10),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_129),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_105),
.B(n_125),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_158),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_157),
.B(n_120),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_160),
.B(n_172),
.Y(n_198)
);

OAI21xp33_ASAP7_75t_SL g207 ( 
.A1(n_162),
.A2(n_170),
.B(n_171),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_153),
.B(n_116),
.Y(n_166)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_166),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_169),
.A2(n_174),
.B1(n_178),
.B2(n_150),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_SL g171 ( 
.A(n_157),
.B(n_124),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_142),
.B(n_109),
.C(n_128),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_142),
.B(n_138),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_173),
.B(n_182),
.Y(n_203)
);

OAI22x1_ASAP7_75t_L g174 ( 
.A1(n_154),
.A2(n_121),
.B1(n_110),
.B2(n_109),
.Y(n_174)
);

NAND3xp33_ASAP7_75t_L g175 ( 
.A(n_130),
.B(n_123),
.C(n_15),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_175),
.B(n_9),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_148),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_177),
.B(n_134),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_146),
.A2(n_89),
.B1(n_85),
.B2(n_72),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_179),
.A2(n_183),
.B(n_182),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_138),
.B(n_6),
.C(n_7),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_136),
.B(n_7),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_139),
.B(n_8),
.Y(n_184)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_184),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_185),
.A2(n_155),
.B(n_141),
.Y(n_191)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_187),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_180),
.B(n_132),
.Y(n_188)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_188),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_167),
.A2(n_151),
.B(n_144),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_189),
.B(n_193),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_184),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_190),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_191),
.B(n_195),
.Y(n_218)
);

XOR2x1_ASAP7_75t_SL g211 ( 
.A(n_192),
.B(n_204),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_181),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_186),
.B(n_156),
.Y(n_195)
);

BUFx12f_ASAP7_75t_L g196 ( 
.A(n_176),
.Y(n_196)
);

INVx6_ASAP7_75t_L g217 ( 
.A(n_196),
.Y(n_217)
);

INVx13_ASAP7_75t_L g197 ( 
.A(n_176),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_197),
.B(n_200),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_163),
.A2(n_177),
.B1(n_140),
.B2(n_152),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_199),
.A2(n_208),
.B1(n_178),
.B2(n_164),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_163),
.A2(n_131),
.B(n_135),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g212 ( 
.A(n_201),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_186),
.B(n_9),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g221 ( 
.A(n_202),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_161),
.B(n_11),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_205),
.B(n_170),
.Y(n_222)
);

OR2x2_ASAP7_75t_L g208 ( 
.A(n_174),
.B(n_150),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_209),
.A2(n_210),
.B1(n_194),
.B2(n_208),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_199),
.A2(n_164),
.B1(n_171),
.B2(n_160),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_198),
.B(n_173),
.C(n_166),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_215),
.B(n_219),
.C(n_224),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_198),
.B(n_172),
.C(n_183),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_222),
.B(n_189),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_203),
.B(n_179),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_223),
.B(n_225),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_203),
.B(n_168),
.C(n_159),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_194),
.B(n_165),
.C(n_145),
.Y(n_225)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_225),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_227),
.B(n_234),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_228),
.B(n_231),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_226),
.A2(n_200),
.B(n_187),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g249 ( 
.A1(n_230),
.A2(n_236),
.B(n_204),
.Y(n_249)
);

AOI221xp5_ASAP7_75t_L g231 ( 
.A1(n_218),
.A2(n_211),
.B1(n_213),
.B2(n_214),
.C(n_207),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_222),
.A2(n_195),
.B1(n_208),
.B2(n_205),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_232),
.A2(n_241),
.B1(n_192),
.B2(n_219),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_216),
.Y(n_234)
);

BUFx12_ASAP7_75t_L g235 ( 
.A(n_211),
.Y(n_235)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_235),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_220),
.B(n_190),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_SL g242 ( 
.A(n_237),
.B(n_223),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_209),
.A2(n_188),
.B1(n_196),
.B2(n_197),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_238),
.A2(n_239),
.B1(n_240),
.B2(n_206),
.Y(n_243)
);

CKINVDCx14_ASAP7_75t_R g239 ( 
.A(n_224),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_217),
.B(n_193),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_217),
.A2(n_210),
.B1(n_206),
.B2(n_196),
.Y(n_241)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_242),
.Y(n_255)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_243),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_SL g261 ( 
.A(n_244),
.B(n_238),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_232),
.A2(n_215),
.B1(n_221),
.B2(n_165),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_245),
.B(n_249),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_229),
.B(n_196),
.C(n_197),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_246),
.B(n_248),
.C(n_230),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_229),
.B(n_191),
.C(n_202),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_233),
.B(n_212),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_251),
.B(n_233),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_249),
.B(n_234),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_253),
.B(n_257),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_254),
.B(n_259),
.C(n_261),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_242),
.B(n_241),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_256),
.B(n_252),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_247),
.B(n_236),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_L g263 ( 
.A1(n_260),
.A2(n_246),
.B(n_248),
.Y(n_263)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_263),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_SL g264 ( 
.A1(n_259),
.A2(n_227),
.B(n_250),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_264),
.B(n_255),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_258),
.B(n_251),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_265),
.B(n_266),
.Y(n_269)
);

AOI322xp5_ASAP7_75t_L g273 ( 
.A1(n_268),
.A2(n_261),
.A3(n_235),
.B1(n_13),
.B2(n_14),
.C1(n_12),
.C2(n_11),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_267),
.B(n_252),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_271),
.B(n_272),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_262),
.B(n_254),
.Y(n_272)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_273),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_270),
.A2(n_269),
.B1(n_235),
.B2(n_13),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_275),
.A2(n_12),
.B(n_274),
.Y(n_276)
);

BUFx24_ASAP7_75t_SL g278 ( 
.A(n_276),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_278),
.B(n_277),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_279),
.B(n_12),
.Y(n_280)
);


endmodule