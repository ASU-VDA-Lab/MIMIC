module fake_jpeg_3806_n_313 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_313);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_313;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx6_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_11),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_14),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_5),
.Y(n_31)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_1),
.B(n_14),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_32),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_34),
.B(n_35),
.Y(n_52)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_32),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_37),
.B(n_39),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_19),
.B(n_0),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_38),
.B(n_21),
.Y(n_48)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_40),
.B(n_16),
.Y(n_60)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_41),
.B(n_24),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

BUFx12_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_43),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_42),
.Y(n_45)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_45),
.Y(n_75)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_46),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_48),
.B(n_49),
.Y(n_76)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_37),
.A2(n_16),
.B1(n_34),
.B2(n_35),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_50),
.A2(n_27),
.B1(n_39),
.B2(n_17),
.Y(n_73)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_53),
.Y(n_77)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_55),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_37),
.A2(n_16),
.B1(n_27),
.B2(n_29),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_56),
.A2(n_62),
.B1(n_30),
.B2(n_20),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_57),
.B(n_60),
.Y(n_81)
);

A2O1A1Ixp33_ASAP7_75t_L g58 ( 
.A1(n_43),
.A2(n_33),
.B(n_17),
.C(n_18),
.Y(n_58)
);

A2O1A1Ixp33_ASAP7_75t_L g78 ( 
.A1(n_58),
.A2(n_66),
.B(n_17),
.C(n_18),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_41),
.B(n_23),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_59),
.B(n_64),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_40),
.A2(n_16),
.B1(n_27),
.B2(n_29),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_63),
.B(n_69),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_36),
.B(n_21),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_36),
.B(n_21),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_65),
.B(n_71),
.Y(n_86)
);

INVx2_ASAP7_75t_R g66 ( 
.A(n_43),
.Y(n_66)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

BUFx2_ASAP7_75t_L g97 ( 
.A(n_67),
.Y(n_97)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_68),
.Y(n_79)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_44),
.B(n_20),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_49),
.A2(n_27),
.B1(n_24),
.B2(n_39),
.Y(n_72)
);

OAI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_72),
.A2(n_94),
.B1(n_23),
.B2(n_19),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_73),
.A2(n_90),
.B1(n_62),
.B2(n_56),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_78),
.B(n_89),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_80),
.A2(n_25),
.B1(n_31),
.B2(n_28),
.Y(n_103)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_66),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_82),
.B(n_83),
.Y(n_102)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_66),
.Y(n_83)
);

INVx13_ASAP7_75t_L g87 ( 
.A(n_63),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_87),
.B(n_93),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_61),
.B(n_33),
.C(n_24),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_88),
.B(n_91),
.C(n_65),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_59),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_58),
.A2(n_24),
.B1(n_18),
.B2(n_28),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_61),
.B(n_20),
.C(n_30),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_54),
.Y(n_92)
);

INVx1_ASAP7_75t_SL g124 ( 
.A(n_92),
.Y(n_124)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_67),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_68),
.A2(n_30),
.B1(n_23),
.B2(n_28),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_47),
.Y(n_96)
);

BUFx24_ASAP7_75t_L g107 ( 
.A(n_96),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_80),
.A2(n_86),
.B1(n_50),
.B2(n_76),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_98),
.A2(n_99),
.B1(n_103),
.B2(n_115),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_86),
.A2(n_53),
.B1(n_54),
.B2(n_55),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_74),
.B(n_71),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_100),
.A2(n_77),
.B(n_91),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_101),
.B(n_70),
.Y(n_139)
);

INVx2_ASAP7_75t_SL g104 ( 
.A(n_85),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_104),
.B(n_106),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_74),
.B(n_48),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_105),
.B(n_108),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_95),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_89),
.B(n_64),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_109),
.A2(n_112),
.B1(n_88),
.B2(n_83),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_95),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_110),
.B(n_113),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g145 ( 
.A1(n_111),
.A2(n_116),
.B1(n_79),
.B2(n_75),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_90),
.A2(n_52),
.B1(n_57),
.B2(n_45),
.Y(n_112)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_97),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_76),
.B(n_69),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_114),
.B(n_117),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_81),
.A2(n_47),
.B1(n_19),
.B2(n_31),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g116 ( 
.A1(n_73),
.A2(n_46),
.B1(n_31),
.B2(n_25),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_81),
.B(n_25),
.Y(n_117)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_97),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_119),
.B(n_121),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_78),
.B(n_0),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_120),
.B(n_0),
.Y(n_141)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_97),
.Y(n_121)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_85),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_123),
.A2(n_79),
.B1(n_96),
.B2(n_70),
.Y(n_150)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_114),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_126),
.B(n_133),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_101),
.B(n_105),
.C(n_98),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_128),
.B(n_139),
.C(n_70),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_129),
.A2(n_140),
.B1(n_143),
.B2(n_99),
.Y(n_160)
);

OA22x2_ASAP7_75t_L g132 ( 
.A1(n_109),
.A2(n_82),
.B1(n_47),
.B2(n_51),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_132),
.A2(n_140),
.B1(n_148),
.B2(n_144),
.Y(n_155)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_121),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_107),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g163 ( 
.A(n_134),
.Y(n_163)
);

INVx13_ASAP7_75t_L g135 ( 
.A(n_104),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_135),
.B(n_136),
.Y(n_162)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_113),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_137),
.A2(n_117),
.B(n_118),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_122),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_138),
.B(n_141),
.Y(n_156)
);

AO21x2_ASAP7_75t_L g140 ( 
.A1(n_124),
.A2(n_51),
.B(n_75),
.Y(n_140)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_115),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_142),
.B(n_110),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_112),
.A2(n_84),
.B1(n_75),
.B2(n_77),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_100),
.B(n_84),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_144),
.B(n_148),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_145),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_118),
.A2(n_87),
.B(n_26),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_147),
.A2(n_151),
.B(n_26),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_100),
.B(n_93),
.Y(n_148)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_119),
.Y(n_149)
);

HB1xp67_ASAP7_75t_L g174 ( 
.A(n_149),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_150),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_108),
.A2(n_26),
.B(n_70),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_154),
.B(n_171),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_155),
.A2(n_161),
.B1(n_170),
.B2(n_51),
.Y(n_196)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_131),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_157),
.B(n_166),
.Y(n_205)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_158),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_130),
.B(n_106),
.Y(n_159)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_159),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_160),
.A2(n_132),
.B1(n_152),
.B2(n_166),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_132),
.A2(n_120),
.B1(n_124),
.B2(n_102),
.Y(n_161)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_140),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_130),
.B(n_102),
.Y(n_167)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_167),
.Y(n_184)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_125),
.Y(n_168)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_168),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_146),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_169),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_132),
.A2(n_152),
.B1(n_142),
.B2(n_129),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_127),
.A2(n_122),
.B(n_3),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_172),
.B(n_179),
.C(n_176),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_143),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_173),
.Y(n_188)
);

CKINVDCx14_ASAP7_75t_R g175 ( 
.A(n_140),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_175),
.B(n_140),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_127),
.A2(n_1),
.B(n_3),
.Y(n_177)
);

MAJx2_ASAP7_75t_L g186 ( 
.A(n_177),
.B(n_147),
.C(n_141),
.Y(n_186)
);

CKINVDCx14_ASAP7_75t_R g197 ( 
.A(n_178),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_128),
.B(n_87),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_182),
.B(n_185),
.C(n_189),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_179),
.B(n_139),
.Y(n_185)
);

OAI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_186),
.A2(n_156),
.B1(n_11),
.B2(n_15),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_172),
.B(n_139),
.C(n_137),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_190),
.B(n_206),
.Y(n_213)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_191),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_160),
.A2(n_126),
.B1(n_138),
.B2(n_151),
.Y(n_192)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_192),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_176),
.B(n_133),
.C(n_136),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_193),
.B(n_163),
.C(n_107),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_173),
.A2(n_165),
.B1(n_154),
.B2(n_155),
.Y(n_194)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_194),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_L g195 ( 
.A1(n_164),
.A2(n_123),
.B1(n_149),
.B2(n_104),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_L g208 ( 
.A1(n_195),
.A2(n_157),
.B1(n_171),
.B2(n_174),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_196),
.A2(n_156),
.B1(n_159),
.B2(n_177),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_165),
.A2(n_135),
.B1(n_26),
.B2(n_96),
.Y(n_198)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_198),
.Y(n_221)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_153),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_199),
.B(n_203),
.Y(n_228)
);

NAND3xp33_ASAP7_75t_L g201 ( 
.A(n_164),
.B(n_169),
.C(n_168),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_201),
.B(n_204),
.Y(n_218)
);

INVx5_ASAP7_75t_L g202 ( 
.A(n_163),
.Y(n_202)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_202),
.Y(n_222)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_153),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_162),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_162),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_183),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_207),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_208),
.B(n_227),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_185),
.B(n_170),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_209),
.B(n_224),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_180),
.B(n_167),
.Y(n_210)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_210),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_202),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_214),
.B(n_229),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_197),
.A2(n_178),
.B1(n_161),
.B2(n_158),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_215),
.A2(n_216),
.B1(n_219),
.B2(n_220),
.Y(n_240)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_217),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_223),
.B(n_230),
.C(n_231),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_SL g224 ( 
.A(n_192),
.B(n_194),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_188),
.A2(n_163),
.B(n_4),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_SL g244 ( 
.A1(n_225),
.A2(n_203),
.B(n_199),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_187),
.B(n_10),
.Y(n_226)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_226),
.Y(n_242)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_205),
.Y(n_227)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_193),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_182),
.B(n_134),
.C(n_107),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_189),
.B(n_107),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_200),
.B(n_15),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_232),
.B(n_200),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_211),
.B(n_184),
.C(n_196),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_237),
.B(n_231),
.C(n_221),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_212),
.A2(n_180),
.B1(n_181),
.B2(n_184),
.Y(n_238)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_238),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_210),
.B(n_181),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_240),
.A2(n_253),
.B1(n_249),
.B2(n_239),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_241),
.B(n_243),
.Y(n_259)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_228),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_244),
.A2(n_251),
.B(n_254),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_209),
.B(n_191),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_245),
.B(n_252),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_213),
.B(n_187),
.Y(n_247)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_247),
.Y(n_270)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_225),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_248),
.B(n_250),
.Y(n_258)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_216),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_223),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_224),
.B(n_186),
.Y(n_252)
);

XOR2x2_ASAP7_75t_L g254 ( 
.A(n_220),
.B(n_215),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_252),
.B(n_211),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_256),
.B(n_268),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_240),
.A2(n_212),
.B1(n_219),
.B2(n_221),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_233),
.B(n_230),
.Y(n_260)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_260),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_246),
.Y(n_261)
);

HB1xp67_ASAP7_75t_L g262 ( 
.A(n_254),
.Y(n_262)
);

CKINVDCx16_ASAP7_75t_R g283 ( 
.A(n_262),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_263),
.B(n_267),
.C(n_271),
.Y(n_274)
);

HB1xp67_ASAP7_75t_L g264 ( 
.A(n_238),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_264),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_235),
.B(n_222),
.C(n_218),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_234),
.B(n_232),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g273 ( 
.A1(n_269),
.A2(n_237),
.B(n_236),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_235),
.B(n_222),
.C(n_198),
.Y(n_271)
);

XNOR2x2_ASAP7_75t_SL g275 ( 
.A(n_265),
.B(n_245),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_259),
.B(n_234),
.C(n_241),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_276),
.B(n_277),
.C(n_281),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_263),
.B(n_242),
.C(n_134),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_261),
.A2(n_255),
.B1(n_258),
.B2(n_270),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_279),
.A2(n_272),
.B1(n_281),
.B2(n_277),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_266),
.B(n_1),
.C(n_4),
.Y(n_281)
);

INVx1_ASAP7_75t_SL g282 ( 
.A(n_257),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_282),
.B(n_266),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_273),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_284),
.B(n_287),
.Y(n_300)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_285),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_280),
.B(n_268),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_286),
.B(n_291),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_SL g287 ( 
.A(n_283),
.B(n_256),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_275),
.A2(n_13),
.B(n_12),
.Y(n_289)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_289),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_278),
.B(n_12),
.Y(n_290)
);

AND2x2_ASAP7_75t_L g292 ( 
.A(n_274),
.B(n_10),
.Y(n_292)
);

AND2x2_ASAP7_75t_L g298 ( 
.A(n_292),
.B(n_293),
.Y(n_298)
);

NOR2xp67_ASAP7_75t_L g293 ( 
.A(n_274),
.B(n_10),
.Y(n_293)
);

OAI21x1_ASAP7_75t_L g294 ( 
.A1(n_292),
.A2(n_280),
.B(n_276),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_294),
.A2(n_299),
.B(n_296),
.Y(n_301)
);

OAI21x1_ASAP7_75t_L g299 ( 
.A1(n_288),
.A2(n_4),
.B(n_5),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_301),
.B(n_304),
.Y(n_308)
);

AOI21xp33_ASAP7_75t_L g302 ( 
.A1(n_297),
.A2(n_284),
.B(n_7),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_302),
.B(n_305),
.C(n_306),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_298),
.B(n_6),
.Y(n_303)
);

OA21x2_ASAP7_75t_L g309 ( 
.A1(n_303),
.A2(n_290),
.B(n_120),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_SL g304 ( 
.A1(n_300),
.A2(n_6),
.B(n_8),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_300),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_295),
.A2(n_6),
.B(n_8),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_309),
.B(n_307),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_310),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_311),
.B(n_308),
.Y(n_312)
);

BUFx24_ASAP7_75t_SL g313 ( 
.A(n_312),
.Y(n_313)
);


endmodule