module fake_netlist_1_1757_n_20 (n_1, n_2, n_4, n_3, n_5, n_0, n_20);
input n_1;
input n_2;
input n_4;
input n_3;
input n_5;
input n_0;
output n_20;
wire n_8;
wire n_11;
wire n_16;
wire n_13;
wire n_18;
wire n_12;
wire n_9;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_19;
wire n_6;
wire n_7;
INVx2_ASAP7_75t_L g6 ( .A(n_4), .Y(n_6) );
HB1xp67_ASAP7_75t_L g7 ( .A(n_5), .Y(n_7) );
INVx2_ASAP7_75t_L g8 ( .A(n_0), .Y(n_8) );
INVx1_ASAP7_75t_L g9 ( .A(n_6), .Y(n_9) );
BUFx6f_ASAP7_75t_L g10 ( .A(n_6), .Y(n_10) );
CKINVDCx5p33_ASAP7_75t_R g11 ( .A(n_7), .Y(n_11) );
AND2x4_ASAP7_75t_L g12 ( .A(n_11), .B(n_8), .Y(n_12) );
OAI22xp5_ASAP7_75t_L g13 ( .A1(n_9), .A2(n_1), .B1(n_2), .B2(n_3), .Y(n_13) );
HB1xp67_ASAP7_75t_L g14 ( .A(n_12), .Y(n_14) );
OR2x6_ASAP7_75t_L g15 ( .A(n_14), .B(n_13), .Y(n_15) );
NAND2xp5_ASAP7_75t_L g16 ( .A(n_15), .B(n_10), .Y(n_16) );
XNOR2xp5_ASAP7_75t_L g17 ( .A(n_16), .B(n_10), .Y(n_17) );
AND2x2_ASAP7_75t_L g18 ( .A(n_17), .B(n_15), .Y(n_18) );
INVxp33_ASAP7_75t_SL g19 ( .A(n_18), .Y(n_19) );
INVx1_ASAP7_75t_L g20 ( .A(n_19), .Y(n_20) );
endmodule