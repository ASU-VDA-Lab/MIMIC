module real_jpeg_8951_n_18 (n_17, n_8, n_0, n_2, n_10, n_9, n_333, n_12, n_6, n_11, n_14, n_7, n_3, n_5, n_4, n_1, n_332, n_16, n_15, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_333;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_332;
input n_16;
input n_15;
input n_13;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_1),
.A2(n_45),
.B(n_96),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_1),
.B(n_45),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_1),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_1),
.A2(n_107),
.B1(n_108),
.B2(n_109),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_1),
.A2(n_32),
.B(n_136),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_1),
.B(n_32),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_1),
.B(n_36),
.Y(n_157)
);

AOI21xp33_ASAP7_75t_L g176 ( 
.A1(n_1),
.A2(n_3),
.B(n_33),
.Y(n_176)
);

OAI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_1),
.A2(n_25),
.B1(n_26),
.B2(n_111),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_2),
.A2(n_45),
.B1(n_46),
.B2(n_98),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_2),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_2),
.A2(n_61),
.B1(n_62),
.B2(n_98),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g137 ( 
.A1(n_2),
.A2(n_32),
.B1(n_33),
.B2(n_98),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_2),
.A2(n_25),
.B1(n_26),
.B2(n_98),
.Y(n_197)
);

INVx2_ASAP7_75t_SL g29 ( 
.A(n_3),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_3),
.A2(n_29),
.B1(n_32),
.B2(n_33),
.Y(n_31)
);

BUFx10_ASAP7_75t_L g88 ( 
.A(n_4),
.Y(n_88)
);

BUFx4f_ASAP7_75t_L g62 ( 
.A(n_5),
.Y(n_62)
);

BUFx10_ASAP7_75t_L g58 ( 
.A(n_6),
.Y(n_58)
);

A2O1A1Ixp33_ASAP7_75t_L g42 ( 
.A1(n_7),
.A2(n_32),
.B(n_43),
.C(n_44),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_7),
.B(n_32),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_7),
.A2(n_45),
.B1(n_46),
.B2(n_47),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_7),
.Y(n_47)
);

BUFx4f_ASAP7_75t_L g46 ( 
.A(n_8),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g23 ( 
.A1(n_9),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_9),
.A2(n_24),
.B1(n_32),
.B2(n_33),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_9),
.A2(n_24),
.B1(n_61),
.B2(n_62),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g258 ( 
.A1(n_9),
.A2(n_24),
.B1(n_45),
.B2(n_46),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_10),
.A2(n_61),
.B1(n_62),
.B2(n_127),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_10),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_10),
.A2(n_45),
.B1(n_46),
.B2(n_127),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_10),
.A2(n_32),
.B1(n_33),
.B2(n_127),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_SL g252 ( 
.A1(n_10),
.A2(n_25),
.B1(n_26),
.B2(n_127),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_11),
.A2(n_61),
.B1(n_62),
.B2(n_146),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_11),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_11),
.A2(n_45),
.B1(n_46),
.B2(n_146),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_11),
.A2(n_32),
.B1(n_33),
.B2(n_146),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_SL g278 ( 
.A1(n_11),
.A2(n_25),
.B1(n_26),
.B2(n_146),
.Y(n_278)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_12),
.A2(n_61),
.B1(n_62),
.B2(n_86),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_12),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_12),
.A2(n_45),
.B1(n_46),
.B2(n_86),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_12),
.A2(n_32),
.B1(n_33),
.B2(n_86),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_12),
.A2(n_25),
.B1(n_26),
.B2(n_86),
.Y(n_209)
);

BUFx2_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_14),
.A2(n_25),
.B1(n_26),
.B2(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_14),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_14),
.A2(n_32),
.B1(n_33),
.B2(n_35),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_14),
.A2(n_35),
.B1(n_45),
.B2(n_46),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g224 ( 
.A1(n_14),
.A2(n_35),
.B1(n_61),
.B2(n_62),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_15),
.A2(n_25),
.B1(n_26),
.B2(n_53),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_15),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_15),
.A2(n_53),
.B1(n_61),
.B2(n_62),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_15),
.A2(n_45),
.B1(n_46),
.B2(n_53),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_SL g249 ( 
.A1(n_15),
.A2(n_32),
.B1(n_33),
.B2(n_53),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_16),
.A2(n_25),
.B1(n_26),
.B2(n_55),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_16),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_16),
.A2(n_55),
.B1(n_61),
.B2(n_62),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_L g226 ( 
.A1(n_16),
.A2(n_45),
.B1(n_46),
.B2(n_55),
.Y(n_226)
);

OAI22xp33_ASAP7_75t_SL g271 ( 
.A1(n_16),
.A2(n_32),
.B1(n_33),
.B2(n_55),
.Y(n_271)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_17),
.A2(n_61),
.B1(n_62),
.B2(n_91),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_17),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g133 ( 
.A1(n_17),
.A2(n_45),
.B1(n_46),
.B2(n_91),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_17),
.A2(n_32),
.B1(n_33),
.B2(n_91),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_17),
.A2(n_25),
.B1(n_26),
.B2(n_91),
.Y(n_234)
);

HAxp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_73),
.CON(n_18),
.SN(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_72),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_37),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_22),
.B(n_37),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_27),
.B1(n_34),
.B2(n_36),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_23),
.A2(n_27),
.B1(n_36),
.B2(n_66),
.Y(n_65)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_25),
.Y(n_26)
);

A2O1A1Ixp33_ASAP7_75t_L g28 ( 
.A1(n_25),
.A2(n_29),
.B(n_30),
.C(n_31),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_25),
.B(n_29),
.Y(n_30)
);

A2O1A1Ixp33_ASAP7_75t_L g175 ( 
.A1(n_25),
.A2(n_29),
.B(n_111),
.C(n_176),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_27),
.A2(n_36),
.B1(n_196),
.B2(n_197),
.Y(n_195)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_28),
.A2(n_31),
.B1(n_52),
.B2(n_54),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_28),
.A2(n_31),
.B1(n_208),
.B2(n_209),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_28),
.A2(n_31),
.B1(n_209),
.B2(n_234),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_28),
.A2(n_31),
.B1(n_234),
.B2(n_252),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_28),
.A2(n_31),
.B1(n_252),
.B2(n_278),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_28),
.A2(n_31),
.B1(n_52),
.B2(n_278),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_31),
.Y(n_36)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_65),
.C(n_67),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_38),
.A2(n_39),
.B1(n_325),
.B2(n_327),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_50),
.C(n_56),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g314 ( 
.A1(n_40),
.A2(n_41),
.B1(n_56),
.B2(n_305),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_41),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_42),
.A2(n_44),
.B1(n_48),
.B2(n_49),
.Y(n_41)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_42),
.A2(n_44),
.B1(n_135),
.B2(n_137),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_42),
.A2(n_44),
.B1(n_137),
.B2(n_154),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_42),
.A2(n_44),
.B1(n_154),
.B2(n_194),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_42),
.A2(n_44),
.B1(n_194),
.B2(n_205),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_42),
.A2(n_44),
.B1(n_205),
.B2(n_231),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_42),
.A2(n_44),
.B1(n_231),
.B2(n_249),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_42),
.A2(n_44),
.B1(n_48),
.B2(n_304),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_43),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_44),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_44),
.B(n_111),
.Y(n_122)
);

A2O1A1Ixp33_ASAP7_75t_SL g57 ( 
.A1(n_45),
.A2(n_58),
.B(n_59),
.C(n_60),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_45),
.B(n_58),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_45),
.B(n_47),
.Y(n_141)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_46),
.A2(n_140),
.B1(n_141),
.B2(n_142),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_49),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_50),
.A2(n_51),
.B1(n_313),
.B2(n_314),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_51),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_54),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_56),
.A2(n_303),
.B1(n_305),
.B2(n_306),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_56),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_SL g56 ( 
.A1(n_57),
.A2(n_60),
.B(n_64),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_57),
.A2(n_60),
.B1(n_95),
.B2(n_97),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_57),
.A2(n_60),
.B1(n_97),
.B2(n_124),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_57),
.A2(n_60),
.B1(n_124),
.B2(n_133),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_57),
.A2(n_60),
.B1(n_133),
.B2(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_57),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_57),
.A2(n_60),
.B1(n_216),
.B2(n_217),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_57),
.A2(n_60),
.B1(n_217),
.B2(n_226),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_57),
.A2(n_60),
.B1(n_226),
.B2(n_258),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_58),
.A2(n_61),
.B1(n_62),
.B2(n_63),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_58),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_59),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_60),
.B(n_111),
.Y(n_110)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_60),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_61),
.B(n_88),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_61),
.B(n_63),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_61),
.B(n_115),
.Y(n_114)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_62),
.A2(n_100),
.B1(n_101),
.B2(n_102),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_64),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_65),
.A2(n_67),
.B1(n_68),
.B2(n_326),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_65),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_68),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_SL g68 ( 
.A1(n_69),
.A2(n_70),
.B(n_71),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_69),
.A2(n_70),
.B1(n_270),
.B2(n_271),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_SL g73 ( 
.A1(n_74),
.A2(n_323),
.B(n_329),
.Y(n_73)
);

OAI321xp33_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_296),
.A3(n_316),
.B1(n_321),
.B2(n_322),
.C(n_332),
.Y(n_74)
);

AOI321xp33_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_242),
.A3(n_284),
.B1(n_290),
.B2(n_295),
.C(n_333),
.Y(n_75)
);

NOR3xp33_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_199),
.C(n_238),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_169),
.B(n_198),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_SL g78 ( 
.A1(n_79),
.A2(n_148),
.B(n_168),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_129),
.B(n_147),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_SL g80 ( 
.A1(n_81),
.A2(n_118),
.B(n_128),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_104),
.B(n_117),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_92),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_83),
.B(n_92),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_84),
.A2(n_87),
.B1(n_88),
.B2(n_89),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_85),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_85),
.A2(n_107),
.B1(n_108),
.B2(n_109),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_87),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_87),
.A2(n_88),
.B1(n_145),
.B2(n_159),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_88),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_90),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_90),
.A2(n_108),
.B1(n_109),
.B2(n_126),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_93),
.A2(n_94),
.B1(n_99),
.B2(n_103),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_93),
.B(n_103),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_94),
.Y(n_93)
);

CKINVDCx14_ASAP7_75t_R g101 ( 
.A(n_96),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_99),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g104 ( 
.A1(n_105),
.A2(n_112),
.B(n_116),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_110),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_106),
.B(n_110),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_108),
.A2(n_109),
.B1(n_126),
.B2(n_144),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_108),
.A2(n_109),
.B1(n_179),
.B2(n_180),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_108),
.A2(n_109),
.B1(n_180),
.B2(n_214),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_108),
.A2(n_109),
.B1(n_214),
.B2(n_224),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_108),
.A2(n_109),
.B(n_224),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_109),
.B(n_111),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_113),
.B(n_114),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_120),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_119),
.B(n_120),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_125),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_123),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_122),
.B(n_123),
.C(n_125),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_131),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_130),
.B(n_131),
.Y(n_147)
);

CKINVDCx5p33_ASAP7_75t_R g149 ( 
.A(n_131),
.Y(n_149)
);

FAx1_ASAP7_75t_SL g131 ( 
.A(n_132),
.B(n_134),
.CI(n_138),
.CON(n_131),
.SN(n_131)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_136),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_143),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_139),
.B(n_143),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_145),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_150),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_149),
.B(n_150),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_151),
.A2(n_152),
.B1(n_161),
.B2(n_162),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_151),
.B(n_164),
.C(n_166),
.Y(n_170)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_153),
.A2(n_155),
.B1(n_156),
.B2(n_160),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_153),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_156),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_158),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_157),
.B(n_158),
.C(n_160),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_159),
.Y(n_179)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_163),
.A2(n_164),
.B1(n_166),
.B2(n_167),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_163),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_164),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_165),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_171),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_170),
.B(n_171),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_184),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_173),
.A2(n_181),
.B1(n_182),
.B2(n_183),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_173),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_173),
.B(n_183),
.C(n_184),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_174),
.A2(n_175),
.B1(n_177),
.B2(n_178),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_174),
.B(n_178),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_175),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_181),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_195),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_186),
.A2(n_187),
.B1(n_192),
.B2(n_193),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_187),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_187),
.B(n_192),
.C(n_195),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_188),
.A2(n_189),
.B1(n_190),
.B2(n_191),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_189),
.A2(n_191),
.B1(n_267),
.B2(n_268),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_190),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_193),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_197),
.Y(n_208)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

AOI21xp33_ASAP7_75t_L g291 ( 
.A1(n_200),
.A2(n_292),
.B(n_293),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_219),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_201),
.B(n_219),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_212),
.C(n_218),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_202),
.B(n_241),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_SL g202 ( 
.A(n_203),
.B(n_211),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_204),
.A2(n_206),
.B1(n_207),
.B2(n_210),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_204),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_SL g236 ( 
.A(n_206),
.B(n_210),
.C(n_211),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_207),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_212),
.B(n_218),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_215),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_213),
.B(n_215),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_220),
.A2(n_221),
.B1(n_236),
.B2(n_237),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_227),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_222),
.B(n_227),
.C(n_237),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_225),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_223),
.B(n_225),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_229),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_228),
.B(n_232),
.C(n_235),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_230),
.A2(n_232),
.B1(n_233),
.B2(n_235),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_230),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_233),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g237 ( 
.A(n_236),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_240),
.Y(n_238)
);

AND2x2_ASAP7_75t_L g292 ( 
.A(n_239),
.B(n_240),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_261),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g295 ( 
.A(n_243),
.B(n_261),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_254),
.C(n_260),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_244),
.A2(n_245),
.B1(n_254),
.B2(n_289),
.Y(n_288)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_247),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_246),
.B(n_250),
.C(n_253),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_248),
.A2(n_250),
.B1(n_251),
.B2(n_253),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_248),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_249),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_251),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g289 ( 
.A(n_254),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_255),
.A2(n_256),
.B1(n_257),
.B2(n_259),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_255),
.A2(n_256),
.B1(n_277),
.B2(n_279),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_L g308 ( 
.A1(n_255),
.A2(n_277),
.B(n_280),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_256),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_256),
.B(n_257),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_257),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_258),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_260),
.B(n_288),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_262),
.A2(n_263),
.B1(n_282),
.B2(n_283),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_264),
.A2(n_265),
.B1(n_273),
.B2(n_274),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_264),
.B(n_274),
.C(n_283),
.Y(n_317)
);

CKINVDCx16_ASAP7_75t_R g264 ( 
.A(n_265),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_L g265 ( 
.A1(n_266),
.A2(n_269),
.B(n_272),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_266),
.B(n_269),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_271),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_272),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_272),
.A2(n_298),
.B1(n_307),
.B2(n_320),
.Y(n_319)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_275),
.A2(n_276),
.B1(n_280),
.B2(n_281),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_277),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_281),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_282),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_L g290 ( 
.A1(n_285),
.A2(n_291),
.B(n_294),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_287),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_286),
.B(n_287),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_309),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_297),
.B(n_309),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_307),
.C(n_308),
.Y(n_297)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_298),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_299),
.A2(n_300),
.B1(n_301),
.B2(n_302),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_299),
.A2(n_300),
.B1(n_311),
.B2(n_312),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_300),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_300),
.B(n_305),
.C(n_306),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_300),
.B(n_311),
.C(n_315),
.Y(n_328)
);

CKINVDCx14_ASAP7_75t_R g301 ( 
.A(n_302),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_303),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_308),
.B(n_319),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_315),
.Y(n_309)
);

CKINVDCx14_ASAP7_75t_R g311 ( 
.A(n_312),
.Y(n_311)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_318),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_317),
.B(n_318),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_328),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_324),
.B(n_328),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_325),
.Y(n_327)
);


endmodule