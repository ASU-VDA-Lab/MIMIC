module fake_jpeg_31204_n_508 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_508);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_508;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx2_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_13),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_16),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_16),
.B(n_6),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_9),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_5),
.Y(n_35)
);

BUFx4f_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_10),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_2),
.B(n_5),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_10),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_3),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_1),
.B(n_15),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_1),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_9),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_9),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_7),
.Y(n_49)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_2),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_0),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_26),
.Y(n_52)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_52),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_20),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_53),
.Y(n_103)
);

INVx13_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g136 ( 
.A(n_54),
.Y(n_136)
);

INVx13_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g138 ( 
.A(n_55),
.Y(n_138)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_56),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g57 ( 
.A(n_27),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_57),
.B(n_58),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_32),
.B(n_17),
.Y(n_58)
);

INVx6_ASAP7_75t_SL g59 ( 
.A(n_36),
.Y(n_59)
);

INVx6_ASAP7_75t_SL g133 ( 
.A(n_59),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_20),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_60),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_30),
.Y(n_61)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_61),
.Y(n_129)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_30),
.Y(n_62)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_62),
.Y(n_112)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_20),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_63),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_30),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g121 ( 
.A(n_64),
.Y(n_121)
);

AND2x2_ASAP7_75t_SL g65 ( 
.A(n_26),
.B(n_0),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_65),
.B(n_66),
.Y(n_127)
);

BUFx12_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_67),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_32),
.B(n_45),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_68),
.B(n_86),
.Y(n_117)
);

BUFx12_ASAP7_75t_L g69 ( 
.A(n_36),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_69),
.B(n_72),
.Y(n_130)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

INVx11_ASAP7_75t_L g144 ( 
.A(n_70),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_20),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_71),
.Y(n_123)
);

CKINVDCx14_ASAP7_75t_R g72 ( 
.A(n_26),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_22),
.Y(n_73)
);

BUFx2_ASAP7_75t_SL g114 ( 
.A(n_73),
.Y(n_114)
);

BUFx4f_ASAP7_75t_SL g74 ( 
.A(n_36),
.Y(n_74)
);

INVx2_ASAP7_75t_SL g147 ( 
.A(n_74),
.Y(n_147)
);

INVx1_ASAP7_75t_SL g75 ( 
.A(n_40),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_75),
.B(n_77),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_22),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_76),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_47),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_47),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_78),
.B(n_79),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_18),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_22),
.Y(n_80)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_80),
.Y(n_102)
);

HB1xp67_ASAP7_75t_L g81 ( 
.A(n_48),
.Y(n_81)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_81),
.Y(n_125)
);

BUFx12_ASAP7_75t_L g82 ( 
.A(n_36),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_82),
.B(n_85),
.Y(n_151)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_27),
.Y(n_83)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_83),
.Y(n_142)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_18),
.Y(n_84)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_84),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_45),
.B(n_19),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_42),
.B(n_17),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_34),
.Y(n_87)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_87),
.Y(n_145)
);

BUFx2_ASAP7_75t_R g88 ( 
.A(n_19),
.Y(n_88)
);

BUFx16f_ASAP7_75t_L g122 ( 
.A(n_88),
.Y(n_122)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_34),
.Y(n_89)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_89),
.Y(n_158)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_28),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_90),
.B(n_101),
.Y(n_153)
);

BUFx5_ASAP7_75t_L g91 ( 
.A(n_29),
.Y(n_91)
);

INVx8_ASAP7_75t_L g139 ( 
.A(n_91),
.Y(n_139)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_18),
.Y(n_92)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_92),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_48),
.Y(n_93)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_93),
.Y(n_135)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_29),
.Y(n_94)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_94),
.Y(n_152)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_29),
.Y(n_95)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_95),
.Y(n_156)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_50),
.Y(n_96)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_96),
.Y(n_105)
);

INVx11_ASAP7_75t_L g97 ( 
.A(n_50),
.Y(n_97)
);

INVx6_ASAP7_75t_L g143 ( 
.A(n_97),
.Y(n_143)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_18),
.Y(n_98)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_98),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_22),
.Y(n_99)
);

INVx6_ASAP7_75t_L g150 ( 
.A(n_99),
.Y(n_150)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_29),
.Y(n_100)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_100),
.Y(n_116)
);

BUFx12f_ASAP7_75t_L g101 ( 
.A(n_38),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_65),
.A2(n_42),
.B1(n_23),
.B2(n_44),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_111),
.A2(n_115),
.B1(n_132),
.B2(n_21),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_53),
.A2(n_23),
.B1(n_46),
.B2(n_44),
.Y(n_115)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_95),
.Y(n_118)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_118),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_88),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_119),
.B(n_141),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_75),
.B(n_49),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_124),
.B(n_157),
.Y(n_162)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_100),
.Y(n_128)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_128),
.Y(n_199)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_56),
.Y(n_131)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_131),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_63),
.A2(n_28),
.B1(n_46),
.B2(n_43),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_61),
.A2(n_29),
.B1(n_50),
.B2(n_38),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_134),
.A2(n_101),
.B1(n_73),
.B2(n_40),
.Y(n_187)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_67),
.Y(n_137)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_137),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_96),
.Y(n_141)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_60),
.Y(n_146)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_146),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_64),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_154),
.B(n_70),
.Y(n_173)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_71),
.Y(n_155)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_155),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_54),
.B(n_21),
.Y(n_157)
);

INVx5_ASAP7_75t_L g159 ( 
.A(n_129),
.Y(n_159)
);

INVx11_ASAP7_75t_L g225 ( 
.A(n_159),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_103),
.Y(n_160)
);

BUFx2_ASAP7_75t_L g226 ( 
.A(n_160),
.Y(n_226)
);

FAx1_ASAP7_75t_SL g161 ( 
.A(n_117),
.B(n_74),
.CI(n_55),
.CON(n_161),
.SN(n_161)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_161),
.B(n_163),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_120),
.B(n_28),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_103),
.Y(n_164)
);

BUFx2_ASAP7_75t_L g240 ( 
.A(n_164),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_142),
.B(n_62),
.C(n_93),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_166),
.B(n_195),
.C(n_39),
.Y(n_233)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_156),
.Y(n_167)
);

INVx3_ASAP7_75t_L g231 ( 
.A(n_167),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_L g169 ( 
.A1(n_102),
.A2(n_99),
.B1(n_80),
.B2(n_76),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_169),
.A2(n_202),
.B1(n_134),
.B2(n_143),
.Y(n_219)
);

BUFx2_ASAP7_75t_L g170 ( 
.A(n_129),
.Y(n_170)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_170),
.Y(n_235)
);

BUFx5_ASAP7_75t_L g171 ( 
.A(n_136),
.Y(n_171)
);

INVx5_ASAP7_75t_L g229 ( 
.A(n_171),
.Y(n_229)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_116),
.Y(n_172)
);

INVx8_ASAP7_75t_L g244 ( 
.A(n_172),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_173),
.B(n_179),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_174),
.B(n_192),
.Y(n_253)
);

INVx6_ASAP7_75t_L g175 ( 
.A(n_104),
.Y(n_175)
);

INVx2_ASAP7_75t_SL g230 ( 
.A(n_175),
.Y(n_230)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_156),
.Y(n_176)
);

HB1xp67_ASAP7_75t_L g218 ( 
.A(n_176),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_127),
.B(n_33),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_177),
.B(n_194),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_104),
.Y(n_178)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_178),
.Y(n_238)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_122),
.Y(n_179)
);

INVx4_ASAP7_75t_SL g180 ( 
.A(n_122),
.Y(n_180)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_180),
.Y(n_213)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_112),
.Y(n_181)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_181),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_123),
.Y(n_182)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_182),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_149),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_183),
.B(n_191),
.Y(n_236)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_112),
.Y(n_184)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_184),
.Y(n_221)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_135),
.Y(n_185)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_185),
.Y(n_224)
);

OAI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_110),
.A2(n_109),
.B1(n_102),
.B2(n_150),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_186),
.A2(n_143),
.B1(n_107),
.B2(n_130),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_187),
.A2(n_193),
.B1(n_197),
.B2(n_209),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_123),
.Y(n_188)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_188),
.Y(n_241)
);

BUFx3_ASAP7_75t_L g189 ( 
.A(n_139),
.Y(n_189)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_189),
.Y(n_250)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_148),
.Y(n_190)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_190),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_153),
.Y(n_191)
);

NAND2xp33_ASAP7_75t_R g192 ( 
.A(n_114),
.B(n_133),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_135),
.A2(n_121),
.B1(n_101),
.B2(n_73),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_145),
.B(n_33),
.Y(n_194)
);

MAJx2_ASAP7_75t_L g195 ( 
.A(n_151),
.B(n_25),
.C(n_24),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_158),
.B(n_35),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_196),
.B(n_198),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_121),
.A2(n_25),
.B1(n_31),
.B2(n_51),
.Y(n_197)
);

BUFx12_ASAP7_75t_L g198 ( 
.A(n_147),
.Y(n_198)
);

A2O1A1Ixp33_ASAP7_75t_L g200 ( 
.A1(n_140),
.A2(n_24),
.B(n_37),
.C(n_31),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_200),
.B(n_204),
.Y(n_256)
);

INVx4_ASAP7_75t_SL g201 ( 
.A(n_107),
.Y(n_201)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_201),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_L g202 ( 
.A1(n_150),
.A2(n_38),
.B1(n_97),
.B2(n_40),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_126),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_203),
.A2(n_208),
.B1(n_212),
.B2(n_138),
.Y(n_215)
);

INVx4_ASAP7_75t_L g204 ( 
.A(n_148),
.Y(n_204)
);

INVx4_ASAP7_75t_L g206 ( 
.A(n_152),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g255 ( 
.A(n_206),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_126),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_109),
.A2(n_39),
.B1(n_35),
.B2(n_49),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_105),
.A2(n_37),
.B1(n_51),
.B2(n_38),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_214),
.A2(n_210),
.B1(n_175),
.B2(n_211),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_215),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_186),
.A2(n_161),
.B1(n_187),
.B2(n_108),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_216),
.A2(n_232),
.B1(n_239),
.B2(n_201),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_219),
.A2(n_254),
.B1(n_164),
.B2(n_4),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_168),
.A2(n_147),
.B(n_125),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_223),
.A2(n_243),
.B(n_167),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_162),
.B(n_113),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_227),
.B(n_237),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_L g232 ( 
.A1(n_202),
.A2(n_105),
.B1(n_152),
.B2(n_106),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_233),
.B(n_198),
.Y(n_281)
);

AOI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_180),
.A2(n_138),
.B1(n_136),
.B2(n_139),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g265 ( 
.A(n_234),
.Y(n_265)
);

AO22x1_ASAP7_75t_SL g237 ( 
.A1(n_195),
.A2(n_74),
.B1(n_82),
.B2(n_69),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_169),
.A2(n_144),
.B1(n_43),
.B2(n_69),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_197),
.A2(n_138),
.B(n_136),
.Y(n_243)
);

OAI22x1_ASAP7_75t_L g245 ( 
.A1(n_212),
.A2(n_193),
.B1(n_189),
.B2(n_144),
.Y(n_245)
);

OA21x2_ASAP7_75t_L g297 ( 
.A1(n_245),
.A2(n_6),
.B(n_7),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_207),
.B(n_1),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_246),
.B(n_247),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_205),
.B(n_1),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_165),
.B(n_2),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_249),
.B(n_247),
.Y(n_294)
);

OAI22xp33_ASAP7_75t_SL g254 ( 
.A1(n_190),
.A2(n_82),
.B1(n_66),
.B2(n_17),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_217),
.B(n_15),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_258),
.B(n_267),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_259),
.A2(n_268),
.B1(n_279),
.B2(n_282),
.Y(n_312)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_257),
.Y(n_260)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_260),
.Y(n_298)
);

BUFx3_ASAP7_75t_L g262 ( 
.A(n_229),
.Y(n_262)
);

BUFx8_ASAP7_75t_L g323 ( 
.A(n_262),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_L g300 ( 
.A1(n_263),
.A2(n_223),
.B(n_250),
.Y(n_300)
);

AOI22xp33_ASAP7_75t_L g334 ( 
.A1(n_266),
.A2(n_297),
.B1(n_240),
.B2(n_220),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_236),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_216),
.A2(n_208),
.B1(n_203),
.B2(n_160),
.Y(n_268)
);

A2O1A1Ixp33_ASAP7_75t_L g269 ( 
.A1(n_228),
.A2(n_198),
.B(n_14),
.C(n_199),
.Y(n_269)
);

NAND2xp33_ASAP7_75t_R g319 ( 
.A(n_269),
.B(n_277),
.Y(n_319)
);

CKINVDCx14_ASAP7_75t_R g270 ( 
.A(n_253),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_270),
.B(n_272),
.Y(n_321)
);

NAND3xp33_ASAP7_75t_L g272 ( 
.A(n_217),
.B(n_14),
.C(n_4),
.Y(n_272)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_222),
.Y(n_273)
);

CKINVDCx14_ASAP7_75t_R g305 ( 
.A(n_273),
.Y(n_305)
);

BUFx2_ASAP7_75t_L g274 ( 
.A(n_238),
.Y(n_274)
);

BUFx2_ASAP7_75t_L g317 ( 
.A(n_274),
.Y(n_317)
);

INVx13_ASAP7_75t_L g275 ( 
.A(n_231),
.Y(n_275)
);

INVxp67_ASAP7_75t_L g302 ( 
.A(n_275),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_SL g276 ( 
.A(n_256),
.B(n_14),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_276),
.B(n_291),
.Y(n_303)
);

OR2x2_ASAP7_75t_SL g277 ( 
.A(n_237),
.B(n_188),
.Y(n_277)
);

INVx13_ASAP7_75t_L g278 ( 
.A(n_231),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_278),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_214),
.A2(n_253),
.B1(n_245),
.B2(n_239),
.Y(n_279)
);

BUFx3_ASAP7_75t_L g280 ( 
.A(n_229),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_280),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_281),
.B(n_285),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_253),
.A2(n_227),
.B1(n_219),
.B2(n_251),
.Y(n_282)
);

O2A1O1Ixp33_ASAP7_75t_SL g283 ( 
.A1(n_243),
.A2(n_170),
.B(n_178),
.C(n_182),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_283),
.A2(n_250),
.B(n_230),
.Y(n_308)
);

INVx3_ASAP7_75t_L g284 ( 
.A(n_226),
.Y(n_284)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_284),
.Y(n_299)
);

NOR2xp67_ASAP7_75t_L g285 ( 
.A(n_237),
.B(n_66),
.Y(n_285)
);

INVx13_ASAP7_75t_L g286 ( 
.A(n_244),
.Y(n_286)
);

CKINVDCx16_ASAP7_75t_R g315 ( 
.A(n_286),
.Y(n_315)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_244),
.Y(n_287)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_287),
.Y(n_306)
);

INVx5_ASAP7_75t_L g288 ( 
.A(n_225),
.Y(n_288)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_288),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_289),
.A2(n_293),
.B1(n_230),
.B2(n_240),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_248),
.B(n_3),
.Y(n_290)
);

CKINVDCx16_ASAP7_75t_R g325 ( 
.A(n_290),
.Y(n_325)
);

INVxp67_ASAP7_75t_L g291 ( 
.A(n_213),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_226),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_292),
.Y(n_320)
);

AOI22xp33_ASAP7_75t_SL g293 ( 
.A1(n_213),
.A2(n_3),
.B1(n_6),
.B2(n_7),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_294),
.B(n_252),
.Y(n_314)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_257),
.Y(n_295)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_295),
.Y(n_310)
);

BUFx2_ASAP7_75t_L g296 ( 
.A(n_238),
.Y(n_296)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_296),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_L g355 ( 
.A1(n_300),
.A2(n_297),
.B(n_265),
.Y(n_355)
);

MAJx2_ASAP7_75t_L g304 ( 
.A(n_264),
.B(n_233),
.C(n_249),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_304),
.B(n_313),
.Y(n_347)
);

OAI21xp5_ASAP7_75t_SL g358 ( 
.A1(n_308),
.A2(n_261),
.B(n_265),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_264),
.B(n_221),
.C(n_224),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_309),
.B(n_327),
.C(n_277),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_271),
.B(n_246),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_314),
.B(n_258),
.Y(n_340)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_260),
.Y(n_316)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_316),
.Y(n_342)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_295),
.Y(n_318)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_318),
.Y(n_350)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_287),
.Y(n_324)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_324),
.Y(n_360)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_271),
.B(n_294),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_274),
.Y(n_328)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_328),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g353 ( 
.A1(n_329),
.A2(n_283),
.B1(n_266),
.B2(n_268),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_282),
.A2(n_230),
.B1(n_220),
.B2(n_241),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_330),
.A2(n_334),
.B1(n_289),
.B2(n_291),
.Y(n_345)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_274),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_332),
.B(n_333),
.Y(n_352)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_296),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_314),
.B(n_273),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_335),
.B(n_344),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_325),
.B(n_267),
.Y(n_336)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_336),
.Y(n_369)
);

INVx4_ASAP7_75t_L g337 ( 
.A(n_323),
.Y(n_337)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_337),
.Y(n_373)
);

INVx13_ASAP7_75t_L g338 ( 
.A(n_302),
.Y(n_338)
);

INVxp67_ASAP7_75t_L g371 ( 
.A(n_338),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_303),
.B(n_276),
.Y(n_339)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_339),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_340),
.B(n_346),
.Y(n_380)
);

XOR2xp5_ASAP7_75t_L g396 ( 
.A(n_341),
.B(n_311),
.Y(n_396)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_327),
.B(n_263),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_343),
.B(n_348),
.C(n_365),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_313),
.B(n_279),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_345),
.A2(n_354),
.B1(n_307),
.B2(n_299),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_SL g346 ( 
.A(n_309),
.B(n_303),
.Y(n_346)
);

XOR2xp5_ASAP7_75t_L g348 ( 
.A(n_304),
.B(n_259),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_SL g349 ( 
.A(n_322),
.B(n_269),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_SL g378 ( 
.A(n_349),
.B(n_351),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_SL g351 ( 
.A(n_305),
.B(n_297),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_353),
.A2(n_307),
.B1(n_306),
.B2(n_324),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_312),
.A2(n_261),
.B1(n_285),
.B2(n_283),
.Y(n_354)
);

INVxp67_ASAP7_75t_L g394 ( 
.A(n_355),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_301),
.B(n_255),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_356),
.B(n_357),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_331),
.B(n_262),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_358),
.Y(n_377)
);

OAI21xp5_ASAP7_75t_L g359 ( 
.A1(n_308),
.A2(n_297),
.B(n_280),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_359),
.B(n_361),
.Y(n_381)
);

INVxp67_ASAP7_75t_L g361 ( 
.A(n_300),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_312),
.B(n_218),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_362),
.B(n_299),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_315),
.B(n_224),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_363),
.B(n_366),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_330),
.B(n_221),
.C(n_252),
.Y(n_365)
);

INVxp67_ASAP7_75t_L g366 ( 
.A(n_319),
.Y(n_366)
);

OAI21xp5_ASAP7_75t_SL g367 ( 
.A1(n_321),
.A2(n_298),
.B(n_310),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_367),
.B(n_292),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_L g370 ( 
.A1(n_349),
.A2(n_320),
.B1(n_329),
.B2(n_316),
.Y(n_370)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_370),
.Y(n_400)
);

OAI32xp33_ASAP7_75t_L g375 ( 
.A1(n_344),
.A2(n_310),
.A3(n_318),
.B1(n_298),
.B2(n_306),
.Y(n_375)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_375),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_376),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_352),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_379),
.B(n_384),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_382),
.A2(n_365),
.B1(n_335),
.B2(n_361),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_SL g412 ( 
.A(n_383),
.B(n_396),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_348),
.B(n_326),
.C(n_302),
.Y(n_384)
);

CKINVDCx14_ASAP7_75t_R g407 ( 
.A(n_386),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_L g387 ( 
.A(n_347),
.B(n_333),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_387),
.B(n_388),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_L g388 ( 
.A(n_347),
.B(n_332),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_353),
.A2(n_328),
.B1(n_311),
.B2(n_317),
.Y(n_389)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_389),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_367),
.B(n_323),
.Y(n_390)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_390),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_340),
.B(n_323),
.Y(n_391)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_391),
.Y(n_415)
);

INVx4_ASAP7_75t_L g392 ( 
.A(n_337),
.Y(n_392)
);

INVx1_ASAP7_75t_SL g398 ( 
.A(n_392),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_341),
.B(n_326),
.C(n_242),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g421 ( 
.A(n_393),
.B(n_397),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_343),
.B(n_286),
.Y(n_397)
);

AOI22xp33_ASAP7_75t_SL g399 ( 
.A1(n_377),
.A2(n_358),
.B1(n_359),
.B2(n_355),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_L g436 ( 
.A1(n_399),
.A2(n_409),
.B1(n_383),
.B2(n_371),
.Y(n_436)
);

INVxp67_ASAP7_75t_L g403 ( 
.A(n_374),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_403),
.B(n_406),
.Y(n_425)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_375),
.Y(n_405)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_405),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_L g408 ( 
.A1(n_372),
.A2(n_378),
.B1(n_369),
.B2(n_382),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_408),
.B(n_410),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_SL g409 ( 
.A1(n_394),
.A2(n_366),
.B1(n_346),
.B2(n_362),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_SL g410 ( 
.A(n_380),
.B(n_350),
.Y(n_410)
);

XOR2xp5_ASAP7_75t_L g411 ( 
.A(n_368),
.B(n_354),
.Y(n_411)
);

XOR2xp5_ASAP7_75t_L g426 ( 
.A(n_411),
.B(n_418),
.Y(n_426)
);

AO21x1_ASAP7_75t_L g413 ( 
.A1(n_381),
.A2(n_351),
.B(n_352),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_413),
.B(n_385),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_371),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_416),
.Y(n_430)
);

XOR2xp5_ASAP7_75t_L g418 ( 
.A(n_368),
.B(n_345),
.Y(n_418)
);

AOI21xp5_ASAP7_75t_L g420 ( 
.A1(n_394),
.A2(n_389),
.B(n_376),
.Y(n_420)
);

INVxp33_ASAP7_75t_L g424 ( 
.A(n_420),
.Y(n_424)
);

XOR2xp5_ASAP7_75t_L g422 ( 
.A(n_396),
.B(n_350),
.Y(n_422)
);

XOR2xp5_ASAP7_75t_L g435 ( 
.A(n_422),
.B(n_412),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_SL g445 ( 
.A(n_427),
.B(n_429),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g428 ( 
.A(n_418),
.B(n_387),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_428),
.B(n_419),
.Y(n_447)
);

CKINVDCx16_ASAP7_75t_R g429 ( 
.A(n_415),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_SL g431 ( 
.A1(n_400),
.A2(n_395),
.B1(n_380),
.B2(n_384),
.Y(n_431)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_431),
.Y(n_456)
);

XOR2x2_ASAP7_75t_SL g432 ( 
.A(n_411),
.B(n_397),
.Y(n_432)
);

BUFx12_ASAP7_75t_L g451 ( 
.A(n_432),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_421),
.B(n_393),
.C(n_388),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_433),
.B(n_437),
.C(n_438),
.Y(n_450)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_414),
.Y(n_434)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_434),
.Y(n_455)
);

XOR2xp5_ASAP7_75t_L g448 ( 
.A(n_435),
.B(n_436),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_421),
.B(n_360),
.C(n_364),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_422),
.B(n_360),
.C(n_364),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_404),
.A2(n_342),
.B1(n_373),
.B2(n_392),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_439),
.B(n_442),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_417),
.B(n_342),
.C(n_373),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_440),
.B(n_406),
.C(n_409),
.Y(n_453)
);

OAI22xp5_ASAP7_75t_SL g442 ( 
.A1(n_404),
.A2(n_317),
.B1(n_241),
.B2(n_284),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_SL g443 ( 
.A1(n_423),
.A2(n_401),
.B1(n_405),
.B2(n_402),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_L g473 ( 
.A1(n_443),
.A2(n_338),
.B1(n_288),
.B2(n_296),
.Y(n_473)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_441),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_444),
.B(n_454),
.Y(n_463)
);

XNOR2xp5_ASAP7_75t_L g466 ( 
.A(n_447),
.B(n_449),
.Y(n_466)
);

XOR2xp5_ASAP7_75t_L g449 ( 
.A(n_426),
.B(n_419),
.Y(n_449)
);

AOI21xp5_ASAP7_75t_L g452 ( 
.A1(n_427),
.A2(n_413),
.B(n_420),
.Y(n_452)
);

AOI21xp5_ASAP7_75t_L g470 ( 
.A1(n_452),
.A2(n_433),
.B(n_426),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_453),
.B(n_458),
.C(n_438),
.Y(n_459)
);

INVxp67_ASAP7_75t_L g454 ( 
.A(n_440),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_430),
.B(n_403),
.Y(n_457)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_457),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_437),
.B(n_412),
.C(n_402),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g480 ( 
.A(n_459),
.B(n_472),
.Y(n_480)
);

OAI22xp5_ASAP7_75t_L g460 ( 
.A1(n_456),
.A2(n_407),
.B1(n_401),
.B2(n_425),
.Y(n_460)
);

AOI22xp5_ASAP7_75t_L g481 ( 
.A1(n_460),
.A2(n_462),
.B1(n_465),
.B2(n_448),
.Y(n_481)
);

OAI22xp5_ASAP7_75t_L g462 ( 
.A1(n_456),
.A2(n_424),
.B1(n_398),
.B2(n_439),
.Y(n_462)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_457),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_464),
.B(n_467),
.Y(n_474)
);

OAI22xp5_ASAP7_75t_SL g465 ( 
.A1(n_446),
.A2(n_424),
.B1(n_432),
.B2(n_431),
.Y(n_465)
);

FAx1_ASAP7_75t_SL g467 ( 
.A(n_443),
.B(n_428),
.CI(n_435),
.CON(n_467),
.SN(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_455),
.B(n_398),
.Y(n_468)
);

CKINVDCx14_ASAP7_75t_R g475 ( 
.A(n_468),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_452),
.B(n_442),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_469),
.B(n_471),
.Y(n_479)
);

XOR2xp5_ASAP7_75t_L g483 ( 
.A(n_470),
.B(n_473),
.Y(n_483)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_445),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_446),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_463),
.B(n_454),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_476),
.B(n_477),
.Y(n_487)
);

OAI22xp5_ASAP7_75t_SL g477 ( 
.A1(n_461),
.A2(n_453),
.B1(n_458),
.B2(n_450),
.Y(n_477)
);

XOR2x2_ASAP7_75t_L g478 ( 
.A(n_463),
.B(n_448),
.Y(n_478)
);

OAI21x1_ASAP7_75t_L g492 ( 
.A1(n_478),
.A2(n_278),
.B(n_275),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_481),
.B(n_482),
.Y(n_491)
);

XNOR2xp5_ASAP7_75t_L g482 ( 
.A(n_459),
.B(n_450),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_L g484 ( 
.A(n_466),
.B(n_449),
.Y(n_484)
);

XOR2xp5_ASAP7_75t_L g490 ( 
.A(n_484),
.B(n_451),
.Y(n_490)
);

OAI21xp5_ASAP7_75t_L g485 ( 
.A1(n_470),
.A2(n_451),
.B(n_338),
.Y(n_485)
);

AOI21xp5_ASAP7_75t_L g488 ( 
.A1(n_485),
.A2(n_468),
.B(n_467),
.Y(n_488)
);

AOI22xp5_ASAP7_75t_L g486 ( 
.A1(n_475),
.A2(n_465),
.B1(n_473),
.B2(n_467),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_486),
.B(n_488),
.Y(n_494)
);

OAI21xp5_ASAP7_75t_SL g489 ( 
.A1(n_480),
.A2(n_466),
.B(n_451),
.Y(n_489)
);

AOI21xp5_ASAP7_75t_L g498 ( 
.A1(n_489),
.A2(n_483),
.B(n_235),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_490),
.B(n_483),
.C(n_484),
.Y(n_497)
);

AOI22xp33_ASAP7_75t_SL g496 ( 
.A1(n_492),
.A2(n_493),
.B1(n_478),
.B2(n_242),
.Y(n_496)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_479),
.Y(n_493)
);

NOR3xp33_ASAP7_75t_SL g495 ( 
.A(n_487),
.B(n_474),
.C(n_482),
.Y(n_495)
);

CKINVDCx20_ASAP7_75t_R g501 ( 
.A(n_495),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_496),
.B(n_497),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_498),
.B(n_486),
.C(n_491),
.Y(n_499)
);

OAI22xp5_ASAP7_75t_L g502 ( 
.A1(n_499),
.A2(n_494),
.B1(n_490),
.B2(n_235),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_SL g504 ( 
.A(n_502),
.B(n_503),
.Y(n_504)
);

AOI322xp5_ASAP7_75t_L g503 ( 
.A1(n_501),
.A2(n_225),
.A3(n_8),
.B1(n_9),
.B2(n_10),
.C1(n_11),
.C2(n_12),
.Y(n_503)
);

A2O1A1Ixp33_ASAP7_75t_SL g505 ( 
.A1(n_504),
.A2(n_500),
.B(n_8),
.C(n_10),
.Y(n_505)
);

O2A1O1Ixp33_ASAP7_75t_SL g506 ( 
.A1(n_505),
.A2(n_6),
.B(n_11),
.C(n_12),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_506),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_507),
.B(n_11),
.Y(n_508)
);


endmodule