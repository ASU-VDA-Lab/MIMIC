module fake_jpeg_4318_n_279 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_279);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_279;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_155;
wire n_118;
wire n_258;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

INVx8_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_12),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_5),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

INVx13_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_30),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_24),
.B(n_0),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_34),
.B(n_16),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_35),
.Y(n_48)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_36),
.B(n_38),
.Y(n_42)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_37),
.B(n_39),
.Y(n_59)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_L g43 ( 
.A1(n_37),
.A2(n_21),
.B1(n_23),
.B2(n_29),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_43),
.A2(n_27),
.B1(n_28),
.B2(n_24),
.Y(n_88)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_44),
.B(n_47),
.Y(n_67)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVx1_ASAP7_75t_SL g80 ( 
.A(n_45),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_46),
.B(n_51),
.Y(n_83)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_50),
.B(n_18),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_16),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_16),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_52),
.B(n_57),
.Y(n_74)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_53),
.Y(n_61)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_54),
.B(n_56),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_55),
.Y(n_72)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_35),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_58),
.Y(n_73)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_60),
.Y(n_65)
);

OAI22xp33_ASAP7_75t_L g62 ( 
.A1(n_49),
.A2(n_36),
.B1(n_35),
.B2(n_26),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_62),
.A2(n_68),
.B1(n_78),
.B2(n_85),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_51),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_63),
.B(n_81),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_50),
.A2(n_21),
.B1(n_23),
.B2(n_29),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_64),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_54),
.A2(n_21),
.B1(n_29),
.B2(n_17),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_66),
.Y(n_96)
);

OAI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_58),
.A2(n_19),
.B1(n_21),
.B2(n_17),
.Y(n_68)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_49),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_69),
.B(n_70),
.Y(n_104)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_60),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_56),
.A2(n_17),
.B1(n_29),
.B2(n_19),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_75),
.B(n_77),
.Y(n_110)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_76),
.Y(n_93)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_45),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_44),
.A2(n_17),
.B1(n_19),
.B2(n_27),
.Y(n_78)
);

AOI32xp33_ASAP7_75t_L g79 ( 
.A1(n_59),
.A2(n_35),
.A3(n_20),
.B1(n_31),
.B2(n_22),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_79),
.B(n_84),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_52),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_47),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_82),
.B(n_41),
.Y(n_109)
);

FAx1_ASAP7_75t_SL g84 ( 
.A(n_46),
.B(n_35),
.CI(n_25),
.CON(n_84),
.SN(n_84)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_53),
.A2(n_18),
.B1(n_27),
.B2(n_28),
.Y(n_85)
);

OA22x2_ASAP7_75t_L g86 ( 
.A1(n_59),
.A2(n_25),
.B1(n_26),
.B2(n_31),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_86),
.A2(n_87),
.B1(n_88),
.B2(n_20),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_42),
.A2(n_24),
.B1(n_28),
.B2(n_18),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_81),
.B(n_57),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_89),
.B(n_100),
.Y(n_127)
);

BUFx24_ASAP7_75t_SL g91 ( 
.A(n_83),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_91),
.B(n_94),
.Y(n_137)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_86),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_67),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_95),
.B(n_97),
.Y(n_140)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_87),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_63),
.B(n_48),
.Y(n_98)
);

OR2x4_ASAP7_75t_L g122 ( 
.A(n_98),
.B(n_25),
.Y(n_122)
);

HB1xp67_ASAP7_75t_L g99 ( 
.A(n_86),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_99),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_83),
.B(n_48),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_71),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_101),
.B(n_103),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_83),
.B(n_25),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_102),
.B(n_114),
.Y(n_129)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_71),
.Y(n_103)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_76),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_105),
.B(n_112),
.Y(n_126)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_74),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_106),
.Y(n_120)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_109),
.Y(n_128)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_111),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_74),
.B(n_84),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_88),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_113),
.B(n_12),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_84),
.B(n_25),
.Y(n_114)
);

AO21x2_ASAP7_75t_L g115 ( 
.A1(n_98),
.A2(n_86),
.B(n_62),
.Y(n_115)
);

AO22x1_ASAP7_75t_SL g143 ( 
.A1(n_115),
.A2(n_98),
.B1(n_89),
.B2(n_108),
.Y(n_143)
);

HB1xp67_ASAP7_75t_SL g116 ( 
.A(n_110),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_116),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_92),
.B(n_64),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_117),
.B(n_107),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_113),
.A2(n_92),
.B1(n_90),
.B2(n_97),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_119),
.A2(n_133),
.B1(n_138),
.B2(n_141),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_111),
.A2(n_79),
.B1(n_70),
.B2(n_69),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_121),
.A2(n_125),
.B1(n_132),
.B2(n_115),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_122),
.A2(n_136),
.B(n_2),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_93),
.B(n_61),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_124),
.B(n_134),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_114),
.A2(n_65),
.B1(n_82),
.B2(n_61),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_112),
.A2(n_25),
.B(n_55),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_131),
.A2(n_32),
.B(n_80),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_108),
.A2(n_65),
.B1(n_73),
.B2(n_41),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_94),
.A2(n_41),
.B1(n_55),
.B2(n_77),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_106),
.B(n_0),
.Y(n_134)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_104),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_135),
.B(n_142),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_96),
.A2(n_73),
.B1(n_31),
.B2(n_22),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_102),
.A2(n_26),
.B1(n_31),
.B2(n_22),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_139),
.B(n_10),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_100),
.A2(n_26),
.B1(n_22),
.B2(n_20),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_107),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_143),
.A2(n_148),
.B1(n_130),
.B2(n_138),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_145),
.B(n_6),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_115),
.A2(n_105),
.B1(n_93),
.B2(n_103),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_147),
.A2(n_149),
.B1(n_158),
.B2(n_132),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_115),
.A2(n_101),
.B1(n_95),
.B2(n_109),
.Y(n_149)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_151),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_123),
.B(n_72),
.Y(n_152)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_152),
.Y(n_175)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_124),
.Y(n_153)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_153),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_123),
.B(n_72),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_154),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_127),
.B(n_1),
.Y(n_155)
);

FAx1_ASAP7_75t_SL g184 ( 
.A(n_155),
.B(n_156),
.CI(n_157),
.CON(n_184),
.SN(n_184)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_127),
.B(n_1),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_142),
.B(n_120),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_115),
.A2(n_72),
.B1(n_32),
.B2(n_4),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_117),
.B(n_80),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_159),
.B(n_163),
.C(n_134),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_140),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_160),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_161),
.A2(n_162),
.B(n_165),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_128),
.B(n_32),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_129),
.B(n_32),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_120),
.B(n_2),
.Y(n_164)
);

OAI21xp33_ASAP7_75t_L g188 ( 
.A1(n_164),
.A2(n_3),
.B(n_4),
.Y(n_188)
);

AND2x6_ASAP7_75t_L g166 ( 
.A(n_122),
.B(n_9),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_166),
.B(n_119),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_128),
.B(n_2),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_167),
.A2(n_168),
.B(n_169),
.Y(n_176)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_125),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_118),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_126),
.B(n_10),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_170),
.A2(n_130),
.B1(n_133),
.B2(n_137),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_173),
.B(n_186),
.Y(n_203)
);

OA21x2_ASAP7_75t_L g177 ( 
.A1(n_143),
.A2(n_166),
.B(n_158),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_177),
.A2(n_189),
.B(n_191),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_145),
.B(n_129),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_178),
.B(n_179),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_159),
.B(n_131),
.Y(n_179)
);

CKINVDCx14_ASAP7_75t_R g197 ( 
.A(n_180),
.Y(n_197)
);

AOI22x1_ASAP7_75t_L g182 ( 
.A1(n_143),
.A2(n_135),
.B1(n_136),
.B2(n_141),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_182),
.A2(n_180),
.B1(n_181),
.B2(n_147),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_183),
.B(n_193),
.C(n_169),
.Y(n_205)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_187),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_SL g210 ( 
.A(n_188),
.B(n_165),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_168),
.A2(n_121),
.B(n_3),
.Y(n_189)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_157),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_190),
.B(n_194),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g191 ( 
.A(n_149),
.B(n_11),
.Y(n_191)
);

OAI21xp33_ASAP7_75t_L g192 ( 
.A1(n_153),
.A2(n_3),
.B(n_5),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_192),
.A2(n_164),
.B(n_151),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_163),
.B(n_6),
.C(n_8),
.Y(n_193)
);

INVx2_ASAP7_75t_SL g194 ( 
.A(n_150),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_195),
.B(n_156),
.Y(n_212)
);

XOR2x2_ASAP7_75t_L g198 ( 
.A(n_182),
.B(n_161),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_SL g226 ( 
.A(n_198),
.B(n_177),
.Y(n_226)
);

BUFx5_ASAP7_75t_L g200 ( 
.A(n_194),
.Y(n_200)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_200),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_184),
.B(n_146),
.Y(n_202)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_202),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_205),
.B(n_212),
.C(n_195),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_172),
.A2(n_148),
.B(n_144),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_206),
.B(n_209),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_207),
.A2(n_171),
.B1(n_175),
.B2(n_196),
.Y(n_229)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_176),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_208),
.B(n_213),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_178),
.B(n_146),
.Y(n_209)
);

NAND3xp33_ASAP7_75t_L g221 ( 
.A(n_210),
.B(n_184),
.C(n_191),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_185),
.Y(n_214)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_214),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_184),
.B(n_155),
.Y(n_215)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_215),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_179),
.B(n_183),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_216),
.B(n_217),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_177),
.A2(n_144),
.B(n_160),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_218),
.B(n_230),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_204),
.B(n_189),
.C(n_193),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_219),
.B(n_220),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_204),
.B(n_174),
.C(n_171),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_SL g242 ( 
.A(n_221),
.B(n_226),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_197),
.A2(n_201),
.B1(n_198),
.B2(n_173),
.Y(n_223)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_223),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_229),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_216),
.B(n_192),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_209),
.B(n_188),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_232),
.B(n_202),
.Y(n_244)
);

INVx1_ASAP7_75t_SL g235 ( 
.A(n_228),
.Y(n_235)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_235),
.Y(n_248)
);

INVx13_ASAP7_75t_L g236 ( 
.A(n_224),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_236),
.B(n_245),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_SL g237 ( 
.A1(n_233),
.A2(n_200),
.B1(n_210),
.B2(n_206),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_237),
.A2(n_207),
.B1(n_217),
.B2(n_211),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_220),
.B(n_212),
.Y(n_238)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_238),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_231),
.A2(n_203),
.B(n_199),
.Y(n_239)
);

AO21x1_ASAP7_75t_L g255 ( 
.A1(n_239),
.A2(n_242),
.B(n_241),
.Y(n_255)
);

MAJx2_ASAP7_75t_L g251 ( 
.A(n_244),
.B(n_225),
.C(n_232),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_222),
.B(n_215),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_234),
.B(n_225),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_246),
.B(n_251),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_243),
.B(n_227),
.C(n_218),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_247),
.B(n_249),
.C(n_244),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_243),
.B(n_227),
.C(n_219),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_234),
.B(n_226),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_252),
.B(n_254),
.C(n_239),
.Y(n_261)
);

AND2x2_ASAP7_75t_L g258 ( 
.A(n_255),
.B(n_242),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_256),
.B(n_261),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_248),
.B(n_235),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_257),
.B(n_258),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_250),
.B(n_236),
.Y(n_259)
);

AOI221xp5_ASAP7_75t_L g269 ( 
.A1(n_259),
.A2(n_251),
.B1(n_247),
.B2(n_10),
.C(n_11),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_253),
.B(n_213),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_260),
.B(n_262),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_255),
.A2(n_240),
.B1(n_199),
.B2(n_230),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_258),
.B(n_205),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_267),
.A2(n_6),
.B(n_8),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_263),
.B(n_249),
.Y(n_268)
);

AO21x1_ASAP7_75t_L g272 ( 
.A1(n_268),
.A2(n_269),
.B(n_15),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_265),
.A2(n_256),
.B1(n_263),
.B2(n_11),
.Y(n_270)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_270),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_271),
.B(n_272),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_SL g273 ( 
.A1(n_266),
.A2(n_8),
.B(n_12),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_275),
.B(n_264),
.C(n_273),
.Y(n_276)
);

AOI322xp5_ASAP7_75t_L g277 ( 
.A1(n_276),
.A2(n_13),
.A3(n_14),
.B1(n_15),
.B2(n_274),
.C1(n_266),
.C2(n_259),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_277),
.B(n_15),
.Y(n_278)
);

OR2x2_ASAP7_75t_L g279 ( 
.A(n_278),
.B(n_13),
.Y(n_279)
);


endmodule