module real_aes_6212_n_105 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_104, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_105);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_104;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_105;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_766;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_565;
wire n_443;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_754;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_505;
wire n_434;
wire n_769;
wire n_502;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_756;
wire n_147;
wire n_288;
wire n_404;
wire n_713;
wire n_598;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_765;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_633;
wire n_520;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_753;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_762;
wire n_212;
wire n_210;
wire n_325;
wire n_575;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g561 ( .A1(n_0), .A2(n_199), .B(n_562), .C(n_565), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_1), .B(n_550), .Y(n_566) );
NAND3xp33_ASAP7_75t_SL g111 ( .A(n_2), .B(n_92), .C(n_112), .Y(n_111) );
INVx1_ASAP7_75t_L g125 ( .A(n_2), .Y(n_125) );
AOI22xp5_ASAP7_75t_L g127 ( .A1(n_3), .A2(n_128), .B1(n_129), .B2(n_132), .Y(n_127) );
INVx1_ASAP7_75t_L g132 ( .A(n_3), .Y(n_132) );
INVx1_ASAP7_75t_L g217 ( .A(n_4), .Y(n_217) );
NAND2xp5_ASAP7_75t_SL g487 ( .A(n_5), .B(n_188), .Y(n_487) );
AOI21xp5_ASAP7_75t_L g543 ( .A1(n_6), .A2(n_465), .B(n_544), .Y(n_543) );
AO21x2_ASAP7_75t_L g511 ( .A1(n_7), .A2(n_164), .B(n_512), .Y(n_511) );
AOI22xp33_ASAP7_75t_L g198 ( .A1(n_8), .A2(n_39), .B1(n_144), .B2(n_153), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_9), .B(n_164), .Y(n_228) );
AND2x6_ASAP7_75t_L g162 ( .A(n_10), .B(n_163), .Y(n_162) );
A2O1A1Ixp33_ASAP7_75t_L g524 ( .A1(n_11), .A2(n_162), .B(n_468), .C(n_525), .Y(n_524) );
NOR2xp33_ASAP7_75t_L g109 ( .A(n_12), .B(n_40), .Y(n_109) );
AOI22xp33_ASAP7_75t_L g105 ( .A1(n_13), .A2(n_106), .B1(n_115), .B2(n_771), .Y(n_105) );
INVx1_ASAP7_75t_L g160 ( .A(n_14), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_15), .B(n_151), .Y(n_171) );
INVx1_ASAP7_75t_L g209 ( .A(n_16), .Y(n_209) );
NAND2xp5_ASAP7_75t_SL g517 ( .A(n_17), .B(n_188), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_18), .B(n_165), .Y(n_233) );
AO32x2_ASAP7_75t_L g196 ( .A1(n_19), .A2(n_161), .A3(n_164), .B1(n_197), .B2(n_201), .Y(n_196) );
NAND2xp5_ASAP7_75t_SL g175 ( .A(n_20), .B(n_153), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_21), .B(n_165), .Y(n_219) );
AOI22xp33_ASAP7_75t_L g200 ( .A1(n_22), .A2(n_56), .B1(n_144), .B2(n_153), .Y(n_200) );
AOI22xp33_ASAP7_75t_SL g150 ( .A1(n_23), .A2(n_83), .B1(n_151), .B2(n_153), .Y(n_150) );
NAND2xp5_ASAP7_75t_SL g190 ( .A(n_24), .B(n_153), .Y(n_190) );
A2O1A1Ixp33_ASAP7_75t_L g467 ( .A1(n_25), .A2(n_161), .B(n_468), .C(n_470), .Y(n_467) );
AOI222xp33_ASAP7_75t_L g446 ( .A1(n_26), .A2(n_447), .B1(n_752), .B2(n_753), .C1(n_762), .C2(n_766), .Y(n_446) );
A2O1A1Ixp33_ASAP7_75t_L g514 ( .A1(n_27), .A2(n_161), .B(n_468), .C(n_515), .Y(n_514) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_28), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_29), .B(n_156), .Y(n_253) );
OAI22xp5_ASAP7_75t_SL g756 ( .A1(n_30), .A2(n_757), .B1(n_760), .B2(n_761), .Y(n_756) );
CKINVDCx20_ASAP7_75t_R g761 ( .A(n_30), .Y(n_761) );
AOI21xp5_ASAP7_75t_L g558 ( .A1(n_31), .A2(n_465), .B(n_559), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_32), .B(n_156), .Y(n_194) );
INVx2_ASAP7_75t_L g146 ( .A(n_33), .Y(n_146) );
A2O1A1Ixp33_ASAP7_75t_L g497 ( .A1(n_34), .A2(n_489), .B(n_498), .C(n_500), .Y(n_497) );
NAND2xp5_ASAP7_75t_SL g248 ( .A(n_35), .B(n_153), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_36), .B(n_156), .Y(n_178) );
OAI22xp5_ASAP7_75t_L g757 ( .A1(n_37), .A2(n_77), .B1(n_758), .B2(n_759), .Y(n_757) );
CKINVDCx20_ASAP7_75t_R g758 ( .A(n_37), .Y(n_758) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_38), .B(n_173), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_41), .B(n_464), .Y(n_463) );
AOI22xp5_ASAP7_75t_L g753 ( .A1(n_42), .A2(n_754), .B1(n_755), .B2(n_756), .Y(n_753) );
CKINVDCx20_ASAP7_75t_R g754 ( .A(n_42), .Y(n_754) );
CKINVDCx20_ASAP7_75t_R g529 ( .A(n_43), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_44), .B(n_188), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_45), .B(n_465), .Y(n_513) );
A2O1A1Ixp33_ASAP7_75t_L g534 ( .A1(n_46), .A2(n_489), .B(n_498), .C(n_535), .Y(n_534) );
AOI22xp5_ASAP7_75t_L g438 ( .A1(n_47), .A2(n_81), .B1(n_439), .B2(n_440), .Y(n_438) );
CKINVDCx20_ASAP7_75t_R g439 ( .A(n_47), .Y(n_439) );
OAI22xp5_ASAP7_75t_SL g449 ( .A1(n_47), .A2(n_439), .B1(n_450), .B2(n_451), .Y(n_449) );
NAND2xp5_ASAP7_75t_SL g223 ( .A(n_48), .B(n_153), .Y(n_223) );
INVx1_ASAP7_75t_L g563 ( .A(n_49), .Y(n_563) );
AOI22xp33_ASAP7_75t_L g143 ( .A1(n_50), .A2(n_91), .B1(n_144), .B2(n_147), .Y(n_143) );
INVx1_ASAP7_75t_L g536 ( .A(n_51), .Y(n_536) );
NAND2xp5_ASAP7_75t_SL g226 ( .A(n_52), .B(n_153), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_53), .B(n_153), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_54), .B(n_465), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_55), .B(n_215), .Y(n_227) );
AOI22xp33_ASAP7_75t_SL g237 ( .A1(n_57), .A2(n_61), .B1(n_151), .B2(n_153), .Y(n_237) );
CKINVDCx20_ASAP7_75t_R g477 ( .A(n_58), .Y(n_477) );
NAND2xp5_ASAP7_75t_SL g170 ( .A(n_59), .B(n_153), .Y(n_170) );
NAND2xp5_ASAP7_75t_SL g252 ( .A(n_60), .B(n_153), .Y(n_252) );
INVx1_ASAP7_75t_L g163 ( .A(n_62), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_63), .B(n_465), .Y(n_491) );
OAI22xp5_ASAP7_75t_SL g129 ( .A1(n_64), .A2(n_100), .B1(n_130), .B2(n_131), .Y(n_129) );
CKINVDCx20_ASAP7_75t_R g131 ( .A(n_64), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_64), .B(n_550), .Y(n_549) );
A2O1A1Ixp33_ASAP7_75t_L g546 ( .A1(n_65), .A2(n_212), .B(n_215), .C(n_547), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_66), .B(n_153), .Y(n_218) );
INVx1_ASAP7_75t_L g159 ( .A(n_67), .Y(n_159) );
CKINVDCx20_ASAP7_75t_R g119 ( .A(n_68), .Y(n_119) );
NAND2xp5_ASAP7_75t_SL g502 ( .A(n_69), .B(n_188), .Y(n_502) );
AO32x2_ASAP7_75t_L g141 ( .A1(n_70), .A2(n_142), .A3(n_155), .B1(n_161), .B2(n_164), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_71), .B(n_154), .Y(n_526) );
INVx1_ASAP7_75t_L g251 ( .A(n_72), .Y(n_251) );
INVx1_ASAP7_75t_L g186 ( .A(n_73), .Y(n_186) );
CKINVDCx16_ASAP7_75t_R g560 ( .A(n_74), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_75), .B(n_472), .Y(n_471) );
A2O1A1Ixp33_ASAP7_75t_L g484 ( .A1(n_76), .A2(n_468), .B(n_485), .C(n_489), .Y(n_484) );
INVx1_ASAP7_75t_L g759 ( .A(n_77), .Y(n_759) );
NAND2xp5_ASAP7_75t_SL g187 ( .A(n_78), .B(n_151), .Y(n_187) );
CKINVDCx16_ASAP7_75t_R g545 ( .A(n_79), .Y(n_545) );
INVx1_ASAP7_75t_L g114 ( .A(n_80), .Y(n_114) );
CKINVDCx20_ASAP7_75t_R g440 ( .A(n_81), .Y(n_440) );
NAND2xp5_ASAP7_75t_SL g473 ( .A(n_82), .B(n_474), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_84), .B(n_144), .Y(n_176) );
CKINVDCx20_ASAP7_75t_R g505 ( .A(n_85), .Y(n_505) );
NAND2xp5_ASAP7_75t_SL g191 ( .A(n_86), .B(n_151), .Y(n_191) );
INVx2_ASAP7_75t_L g157 ( .A(n_87), .Y(n_157) );
CKINVDCx20_ASAP7_75t_R g493 ( .A(n_88), .Y(n_493) );
NAND2xp5_ASAP7_75t_SL g527 ( .A(n_89), .B(n_148), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_90), .B(n_151), .Y(n_224) );
OR2x2_ASAP7_75t_L g122 ( .A(n_92), .B(n_123), .Y(n_122) );
OR2x2_ASAP7_75t_L g454 ( .A(n_92), .B(n_124), .Y(n_454) );
INVx2_ASAP7_75t_L g751 ( .A(n_92), .Y(n_751) );
AOI22xp33_ASAP7_75t_L g236 ( .A1(n_93), .A2(n_104), .B1(n_151), .B2(n_152), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_94), .B(n_465), .Y(n_496) );
INVx1_ASAP7_75t_L g501 ( .A(n_95), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_96), .B(n_443), .Y(n_442) );
INVxp67_ASAP7_75t_L g548 ( .A(n_97), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_98), .B(n_151), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g113 ( .A(n_99), .B(n_114), .Y(n_113) );
INVx1_ASAP7_75t_L g130 ( .A(n_100), .Y(n_130) );
INVx1_ASAP7_75t_L g486 ( .A(n_101), .Y(n_486) );
INVx1_ASAP7_75t_L g522 ( .A(n_102), .Y(n_522) );
AND2x2_ASAP7_75t_L g538 ( .A(n_103), .B(n_156), .Y(n_538) );
INVx1_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
INVx1_ASAP7_75t_L g771 ( .A(n_108), .Y(n_771) );
AND2x2_ASAP7_75t_L g108 ( .A(n_109), .B(n_110), .Y(n_108) );
AND2x2_ASAP7_75t_L g124 ( .A(n_109), .B(n_125), .Y(n_124) );
INVx1_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
INVx1_ASAP7_75t_SL g112 ( .A(n_113), .Y(n_112) );
OA21x2_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_120), .B(n_445), .Y(n_115) );
BUFx2_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
BUFx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
INVx1_ASAP7_75t_L g770 ( .A(n_118), .Y(n_770) );
INVx2_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
OAI21xp5_ASAP7_75t_L g120 ( .A1(n_121), .A2(n_126), .B(n_442), .Y(n_120) );
INVx2_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
HB1xp67_ASAP7_75t_L g444 ( .A(n_122), .Y(n_444) );
NOR2x2_ASAP7_75t_L g768 ( .A(n_123), .B(n_751), .Y(n_768) );
INVx2_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
OR2x2_ASAP7_75t_L g750 ( .A(n_124), .B(n_751), .Y(n_750) );
AOI22xp5_ASAP7_75t_L g126 ( .A1(n_127), .A2(n_133), .B1(n_134), .B2(n_441), .Y(n_126) );
CKINVDCx20_ASAP7_75t_R g441 ( .A(n_127), .Y(n_441) );
CKINVDCx20_ASAP7_75t_R g128 ( .A(n_129), .Y(n_128) );
INVx1_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
XOR2x2_ASAP7_75t_L g134 ( .A(n_135), .B(n_438), .Y(n_134) );
INVx2_ASAP7_75t_L g450 ( .A(n_135), .Y(n_450) );
AND3x1_ASAP7_75t_L g135 ( .A(n_136), .B(n_358), .C(n_406), .Y(n_135) );
NOR4xp25_ASAP7_75t_L g136 ( .A(n_137), .B(n_286), .C(n_331), .D(n_345), .Y(n_136) );
OAI311xp33_ASAP7_75t_L g137 ( .A1(n_138), .A2(n_202), .A3(n_229), .B1(n_239), .C1(n_254), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g138 ( .A(n_139), .B(n_166), .Y(n_138) );
OAI21xp33_ASAP7_75t_L g239 ( .A1(n_139), .A2(n_240), .B(n_242), .Y(n_239) );
AND2x2_ASAP7_75t_L g347 ( .A(n_139), .B(n_274), .Y(n_347) );
AND2x2_ASAP7_75t_L g404 ( .A(n_139), .B(n_290), .Y(n_404) );
BUFx2_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
AND2x2_ASAP7_75t_L g297 ( .A(n_140), .B(n_195), .Y(n_297) );
AND2x2_ASAP7_75t_L g354 ( .A(n_140), .B(n_302), .Y(n_354) );
INVx1_ASAP7_75t_L g395 ( .A(n_140), .Y(n_395) );
INVx1_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
BUFx6f_ASAP7_75t_L g263 ( .A(n_141), .Y(n_263) );
AND2x2_ASAP7_75t_L g304 ( .A(n_141), .B(n_195), .Y(n_304) );
AND2x2_ASAP7_75t_L g308 ( .A(n_141), .B(n_196), .Y(n_308) );
INVx1_ASAP7_75t_L g320 ( .A(n_141), .Y(n_320) );
OAI22xp5_ASAP7_75t_SL g142 ( .A1(n_143), .A2(n_148), .B1(n_150), .B2(n_154), .Y(n_142) );
INVx1_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
BUFx3_ASAP7_75t_L g147 ( .A(n_145), .Y(n_147) );
BUFx6f_ASAP7_75t_L g153 ( .A(n_145), .Y(n_153) );
AND2x6_ASAP7_75t_L g468 ( .A(n_145), .B(n_469), .Y(n_468) );
INVx2_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx1_ASAP7_75t_L g152 ( .A(n_146), .Y(n_152) );
INVx1_ASAP7_75t_L g216 ( .A(n_146), .Y(n_216) );
HB1xp67_ASAP7_75t_L g503 ( .A(n_147), .Y(n_503) );
INVx2_ASAP7_75t_L g565 ( .A(n_147), .Y(n_565) );
INVx2_ASAP7_75t_L g177 ( .A(n_148), .Y(n_177) );
OAI22xp5_ASAP7_75t_L g197 ( .A1(n_148), .A2(n_198), .B1(n_199), .B2(n_200), .Y(n_197) );
OAI22xp5_ASAP7_75t_L g235 ( .A1(n_148), .A2(n_199), .B1(n_236), .B2(n_237), .Y(n_235) );
INVx4_ASAP7_75t_L g564 ( .A(n_148), .Y(n_564) );
BUFx6f_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx3_ASAP7_75t_L g154 ( .A(n_149), .Y(n_154) );
INVx1_ASAP7_75t_L g173 ( .A(n_149), .Y(n_173) );
BUFx6f_ASAP7_75t_L g193 ( .A(n_149), .Y(n_193) );
AND2x2_ASAP7_75t_L g466 ( .A(n_149), .B(n_216), .Y(n_466) );
INVx1_ASAP7_75t_L g469 ( .A(n_149), .Y(n_469) );
INVx2_ASAP7_75t_L g210 ( .A(n_151), .Y(n_210) );
INVx3_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx3_ASAP7_75t_L g185 ( .A(n_153), .Y(n_185) );
HB1xp67_ASAP7_75t_L g488 ( .A(n_153), .Y(n_488) );
INVx5_ASAP7_75t_L g188 ( .A(n_154), .Y(n_188) );
INVx1_ASAP7_75t_L g475 ( .A(n_155), .Y(n_475) );
INVx2_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
OA21x2_ASAP7_75t_L g167 ( .A1(n_156), .A2(n_168), .B(n_178), .Y(n_167) );
OA21x2_ASAP7_75t_L g182 ( .A1(n_156), .A2(n_183), .B(n_194), .Y(n_182) );
INVx1_ASAP7_75t_L g478 ( .A(n_156), .Y(n_478) );
AOI21xp5_ASAP7_75t_L g495 ( .A1(n_156), .A2(n_496), .B(n_497), .Y(n_495) );
AOI21xp5_ASAP7_75t_L g532 ( .A1(n_156), .A2(n_533), .B(n_534), .Y(n_532) );
AND2x2_ASAP7_75t_SL g156 ( .A(n_157), .B(n_158), .Y(n_156) );
AND2x2_ASAP7_75t_L g165 ( .A(n_157), .B(n_158), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_159), .B(n_160), .Y(n_158) );
NAND3xp33_ASAP7_75t_L g234 ( .A(n_161), .B(n_235), .C(n_238), .Y(n_234) );
OAI21xp5_ASAP7_75t_L g246 ( .A1(n_161), .A2(n_247), .B(n_250), .Y(n_246) );
BUFx3_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
OAI21xp5_ASAP7_75t_L g168 ( .A1(n_162), .A2(n_169), .B(n_174), .Y(n_168) );
OAI21xp5_ASAP7_75t_L g183 ( .A1(n_162), .A2(n_184), .B(n_189), .Y(n_183) );
OAI21xp5_ASAP7_75t_L g207 ( .A1(n_162), .A2(n_208), .B(n_213), .Y(n_207) );
OAI21xp5_ASAP7_75t_L g221 ( .A1(n_162), .A2(n_222), .B(n_225), .Y(n_221) );
AND2x4_ASAP7_75t_L g465 ( .A(n_162), .B(n_466), .Y(n_465) );
INVx4_ASAP7_75t_SL g490 ( .A(n_162), .Y(n_490) );
NAND2x1p5_ASAP7_75t_L g523 ( .A(n_162), .B(n_466), .Y(n_523) );
OA21x2_ASAP7_75t_L g220 ( .A1(n_164), .A2(n_221), .B(n_228), .Y(n_220) );
INVx4_ASAP7_75t_L g238 ( .A(n_164), .Y(n_238) );
AOI21xp5_ASAP7_75t_L g512 ( .A1(n_164), .A2(n_513), .B(n_514), .Y(n_512) );
HB1xp67_ASAP7_75t_L g542 ( .A(n_164), .Y(n_542) );
BUFx6f_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
INVx1_ASAP7_75t_L g201 ( .A(n_165), .Y(n_201) );
AND2x2_ASAP7_75t_L g166 ( .A(n_167), .B(n_179), .Y(n_166) );
AND2x2_ASAP7_75t_L g241 ( .A(n_167), .B(n_195), .Y(n_241) );
INVx2_ASAP7_75t_L g275 ( .A(n_167), .Y(n_275) );
AND2x2_ASAP7_75t_L g290 ( .A(n_167), .B(n_196), .Y(n_290) );
HB1xp67_ASAP7_75t_L g296 ( .A(n_167), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_167), .B(n_302), .Y(n_301) );
OR2x2_ASAP7_75t_L g310 ( .A(n_167), .B(n_273), .Y(n_310) );
INVx1_ASAP7_75t_L g322 ( .A(n_167), .Y(n_322) );
INVx1_ASAP7_75t_L g363 ( .A(n_167), .Y(n_363) );
NOR2xp33_ASAP7_75t_L g416 ( .A(n_167), .B(n_263), .Y(n_416) );
AOI21xp5_ASAP7_75t_L g169 ( .A1(n_170), .A2(n_171), .B(n_172), .Y(n_169) );
INVx1_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
AOI21xp5_ASAP7_75t_L g174 ( .A1(n_175), .A2(n_176), .B(n_177), .Y(n_174) );
O2A1O1Ixp5_ASAP7_75t_L g250 ( .A1(n_177), .A2(n_214), .B(n_251), .C(n_252), .Y(n_250) );
NOR2xp67_ASAP7_75t_L g179 ( .A(n_180), .B(n_195), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
AND2x2_ASAP7_75t_L g240 ( .A(n_181), .B(n_241), .Y(n_240) );
HB1xp67_ASAP7_75t_L g268 ( .A(n_181), .Y(n_268) );
AND2x2_ASAP7_75t_SL g321 ( .A(n_181), .B(n_322), .Y(n_321) );
OR2x2_ASAP7_75t_L g325 ( .A(n_181), .B(n_195), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_181), .B(n_320), .Y(n_383) );
INVx2_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
INVx2_ASAP7_75t_L g273 ( .A(n_182), .Y(n_273) );
HB1xp67_ASAP7_75t_L g289 ( .A(n_182), .Y(n_289) );
OR2x2_ASAP7_75t_L g362 ( .A(n_182), .B(n_363), .Y(n_362) );
O2A1O1Ixp5_ASAP7_75t_SL g184 ( .A1(n_185), .A2(n_186), .B(n_187), .C(n_188), .Y(n_184) );
INVx2_ASAP7_75t_L g199 ( .A(n_188), .Y(n_199) );
AOI21xp5_ASAP7_75t_L g222 ( .A1(n_188), .A2(n_223), .B(n_224), .Y(n_222) );
AOI21xp5_ASAP7_75t_L g247 ( .A1(n_188), .A2(n_248), .B(n_249), .Y(n_247) );
NOR2xp33_ASAP7_75t_L g547 ( .A(n_188), .B(n_548), .Y(n_547) );
AOI21xp5_ASAP7_75t_L g189 ( .A1(n_190), .A2(n_191), .B(n_192), .Y(n_189) );
INVx1_ASAP7_75t_L g212 ( .A(n_192), .Y(n_212) );
INVx4_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
INVx2_ASAP7_75t_L g472 ( .A(n_193), .Y(n_472) );
INVx2_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
BUFx2_ASAP7_75t_L g269 ( .A(n_196), .Y(n_269) );
AND2x2_ASAP7_75t_L g274 ( .A(n_196), .B(n_275), .Y(n_274) );
O2A1O1Ixp33_ASAP7_75t_L g213 ( .A1(n_199), .A2(n_214), .B(n_217), .C(n_218), .Y(n_213) );
AOI21xp5_ASAP7_75t_L g225 ( .A1(n_199), .A2(n_226), .B(n_227), .Y(n_225) );
INVx2_ASAP7_75t_L g206 ( .A(n_201), .Y(n_206) );
NOR2xp33_ASAP7_75t_L g528 ( .A(n_201), .B(n_529), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_202), .B(n_257), .Y(n_420) );
INVx1_ASAP7_75t_SL g202 ( .A(n_203), .Y(n_202) );
OR2x2_ASAP7_75t_L g390 ( .A(n_203), .B(n_231), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_204), .B(n_220), .Y(n_203) );
AND2x2_ASAP7_75t_L g266 ( .A(n_204), .B(n_257), .Y(n_266) );
INVx2_ASAP7_75t_L g278 ( .A(n_204), .Y(n_278) );
AND2x2_ASAP7_75t_L g312 ( .A(n_204), .B(n_260), .Y(n_312) );
AND2x2_ASAP7_75t_L g379 ( .A(n_204), .B(n_380), .Y(n_379) );
INVx2_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_205), .B(n_245), .Y(n_244) );
AND2x2_ASAP7_75t_L g259 ( .A(n_205), .B(n_260), .Y(n_259) );
AND2x2_ASAP7_75t_L g299 ( .A(n_205), .B(n_220), .Y(n_299) );
AND2x2_ASAP7_75t_L g316 ( .A(n_205), .B(n_317), .Y(n_316) );
OA21x2_ASAP7_75t_L g205 ( .A1(n_206), .A2(n_207), .B(n_219), .Y(n_205) );
OA21x2_ASAP7_75t_L g245 ( .A1(n_206), .A2(n_246), .B(n_253), .Y(n_245) );
O2A1O1Ixp33_ASAP7_75t_L g208 ( .A1(n_209), .A2(n_210), .B(n_211), .C(n_212), .Y(n_208) );
AOI21xp5_ASAP7_75t_L g515 ( .A1(n_210), .A2(n_516), .B(n_517), .Y(n_515) );
AOI21xp5_ASAP7_75t_L g525 ( .A1(n_210), .A2(n_526), .B(n_527), .Y(n_525) );
O2A1O1Ixp33_ASAP7_75t_L g485 ( .A1(n_212), .A2(n_486), .B(n_487), .C(n_488), .Y(n_485) );
AOI21xp5_ASAP7_75t_L g470 ( .A1(n_214), .A2(n_471), .B(n_473), .Y(n_470) );
INVx2_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
AND2x2_ASAP7_75t_L g242 ( .A(n_220), .B(n_243), .Y(n_242) );
INVx3_ASAP7_75t_L g260 ( .A(n_220), .Y(n_260) );
AND2x2_ASAP7_75t_L g265 ( .A(n_220), .B(n_245), .Y(n_265) );
AND2x2_ASAP7_75t_L g338 ( .A(n_220), .B(n_317), .Y(n_338) );
AND2x2_ASAP7_75t_L g403 ( .A(n_220), .B(n_393), .Y(n_403) );
OAI311xp33_ASAP7_75t_L g286 ( .A1(n_229), .A2(n_287), .A3(n_291), .B1(n_293), .C1(n_313), .Y(n_286) );
INVx1_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
AND2x2_ASAP7_75t_L g298 ( .A(n_230), .B(n_299), .Y(n_298) );
AND2x2_ASAP7_75t_L g357 ( .A(n_230), .B(n_265), .Y(n_357) );
AND2x2_ASAP7_75t_L g431 ( .A(n_230), .B(n_312), .Y(n_431) );
INVx2_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
NOR2xp33_ASAP7_75t_L g243 ( .A(n_231), .B(n_244), .Y(n_243) );
INVx1_ASAP7_75t_L g366 ( .A(n_231), .Y(n_366) );
INVx2_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
INVx3_ASAP7_75t_L g257 ( .A(n_232), .Y(n_257) );
NOR2x1_ASAP7_75t_L g329 ( .A(n_232), .B(n_330), .Y(n_329) );
AND2x2_ASAP7_75t_L g386 ( .A(n_232), .B(n_260), .Y(n_386) );
AND2x4_ASAP7_75t_L g232 ( .A(n_233), .B(n_234), .Y(n_232) );
INVx1_ASAP7_75t_L g283 ( .A(n_233), .Y(n_283) );
AO21x1_ASAP7_75t_L g282 ( .A1(n_235), .A2(n_238), .B(n_283), .Y(n_282) );
AO21x2_ASAP7_75t_L g482 ( .A1(n_238), .A2(n_483), .B(n_492), .Y(n_482) );
NOR2xp33_ASAP7_75t_L g492 ( .A(n_238), .B(n_493), .Y(n_492) );
NOR2xp33_ASAP7_75t_L g504 ( .A(n_238), .B(n_505), .Y(n_504) );
AO21x2_ASAP7_75t_L g520 ( .A1(n_238), .A2(n_521), .B(n_528), .Y(n_520) );
INVx3_ASAP7_75t_L g550 ( .A(n_238), .Y(n_550) );
AND2x2_ASAP7_75t_L g261 ( .A(n_241), .B(n_262), .Y(n_261) );
AND2x2_ASAP7_75t_L g314 ( .A(n_241), .B(n_315), .Y(n_314) );
AND2x2_ASAP7_75t_L g394 ( .A(n_241), .B(n_395), .Y(n_394) );
AOI221xp5_ASAP7_75t_L g293 ( .A1(n_242), .A2(n_274), .B1(n_294), .B2(n_298), .C(n_300), .Y(n_293) );
INVx1_ASAP7_75t_L g418 ( .A(n_243), .Y(n_418) );
OR2x2_ASAP7_75t_L g384 ( .A(n_244), .B(n_385), .Y(n_384) );
AND2x2_ASAP7_75t_L g279 ( .A(n_245), .B(n_260), .Y(n_279) );
OR2x2_ASAP7_75t_L g281 ( .A(n_245), .B(n_282), .Y(n_281) );
INVx1_ASAP7_75t_L g306 ( .A(n_245), .Y(n_306) );
INVx2_ASAP7_75t_L g317 ( .A(n_245), .Y(n_317) );
AND2x2_ASAP7_75t_L g344 ( .A(n_245), .B(n_282), .Y(n_344) );
HB1xp67_ASAP7_75t_L g373 ( .A(n_245), .Y(n_373) );
AOI221xp5_ASAP7_75t_L g254 ( .A1(n_255), .A2(n_261), .B1(n_264), .B2(n_267), .C(n_270), .Y(n_254) );
INVx1_ASAP7_75t_SL g255 ( .A(n_256), .Y(n_255) );
OR2x2_ASAP7_75t_L g256 ( .A(n_257), .B(n_258), .Y(n_256) );
AND2x2_ASAP7_75t_L g355 ( .A(n_257), .B(n_265), .Y(n_355) );
AND2x2_ASAP7_75t_L g405 ( .A(n_257), .B(n_259), .Y(n_405) );
INVx2_ASAP7_75t_SL g258 ( .A(n_259), .Y(n_258) );
AND2x2_ASAP7_75t_L g292 ( .A(n_259), .B(n_263), .Y(n_292) );
AND2x2_ASAP7_75t_L g371 ( .A(n_259), .B(n_344), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_260), .B(n_306), .Y(n_305) );
INVx2_ASAP7_75t_L g330 ( .A(n_260), .Y(n_330) );
OAI21xp33_ASAP7_75t_L g340 ( .A1(n_261), .A2(n_341), .B(n_343), .Y(n_340) );
OR2x2_ASAP7_75t_L g284 ( .A(n_262), .B(n_285), .Y(n_284) );
OR2x2_ASAP7_75t_L g350 ( .A(n_262), .B(n_310), .Y(n_350) );
NOR2xp33_ASAP7_75t_L g361 ( .A(n_262), .B(n_362), .Y(n_361) );
INVx2_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
AND2x2_ASAP7_75t_L g327 ( .A(n_263), .B(n_296), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_263), .B(n_410), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_264), .B(n_290), .Y(n_400) );
AND2x2_ASAP7_75t_L g264 ( .A(n_265), .B(n_266), .Y(n_264) );
AND2x2_ASAP7_75t_L g323 ( .A(n_265), .B(n_278), .Y(n_323) );
INVx1_ASAP7_75t_L g339 ( .A(n_266), .Y(n_339) );
NOR2xp33_ASAP7_75t_L g267 ( .A(n_268), .B(n_269), .Y(n_267) );
OAI22xp5_ASAP7_75t_L g270 ( .A1(n_271), .A2(n_276), .B1(n_280), .B2(n_284), .Y(n_270) );
INVx2_ASAP7_75t_SL g271 ( .A(n_272), .Y(n_271) );
AND2x2_ASAP7_75t_L g272 ( .A(n_273), .B(n_274), .Y(n_272) );
INVx2_ASAP7_75t_L g302 ( .A(n_273), .Y(n_302) );
INVx1_ASAP7_75t_L g315 ( .A(n_273), .Y(n_315) );
INVx1_ASAP7_75t_L g285 ( .A(n_274), .Y(n_285) );
AND2x2_ASAP7_75t_L g356 ( .A(n_274), .B(n_302), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_274), .B(n_382), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_277), .B(n_279), .Y(n_276) );
OR2x2_ASAP7_75t_L g280 ( .A(n_277), .B(n_281), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_277), .B(n_393), .Y(n_392) );
NOR2xp67_ASAP7_75t_L g424 ( .A(n_277), .B(n_425), .Y(n_424) );
INVx3_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
AND2x2_ASAP7_75t_L g427 ( .A(n_279), .B(n_379), .Y(n_427) );
INVx1_ASAP7_75t_SL g393 ( .A(n_281), .Y(n_393) );
AND2x2_ASAP7_75t_L g333 ( .A(n_282), .B(n_317), .Y(n_333) );
INVx1_ASAP7_75t_L g380 ( .A(n_282), .Y(n_380) );
OAI222xp33_ASAP7_75t_L g421 ( .A1(n_287), .A2(n_377), .B1(n_422), .B2(n_423), .C1(n_426), .C2(n_428), .Y(n_421) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
AND2x2_ASAP7_75t_L g288 ( .A(n_289), .B(n_290), .Y(n_288) );
INVx1_ASAP7_75t_L g342 ( .A(n_289), .Y(n_342) );
AND2x2_ASAP7_75t_L g353 ( .A(n_290), .B(n_354), .Y(n_353) );
NAND2xp5_ASAP7_75t_SL g422 ( .A(n_290), .B(n_395), .Y(n_422) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_292), .B(n_375), .Y(n_374) );
INVx1_ASAP7_75t_L g397 ( .A(n_294), .Y(n_397) );
AND2x2_ASAP7_75t_L g294 ( .A(n_295), .B(n_297), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
INVx1_ASAP7_75t_SL g335 ( .A(n_297), .Y(n_335) );
AND2x2_ASAP7_75t_L g414 ( .A(n_297), .B(n_375), .Y(n_414) );
AND2x2_ASAP7_75t_L g437 ( .A(n_297), .B(n_321), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_299), .B(n_333), .Y(n_332) );
OAI32xp33_ASAP7_75t_L g300 ( .A1(n_301), .A2(n_303), .A3(n_305), .B1(n_307), .B2(n_311), .Y(n_300) );
BUFx2_ASAP7_75t_L g375 ( .A(n_302), .Y(n_375) );
NOR2xp33_ASAP7_75t_L g402 ( .A(n_303), .B(n_321), .Y(n_402) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
AND2x2_ASAP7_75t_L g341 ( .A(n_304), .B(n_342), .Y(n_341) );
AND2x4_ASAP7_75t_L g409 ( .A(n_304), .B(n_410), .Y(n_409) );
OR2x2_ASAP7_75t_L g398 ( .A(n_305), .B(n_399), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_308), .B(n_309), .Y(n_307) );
AND2x2_ASAP7_75t_L g369 ( .A(n_308), .B(n_342), .Y(n_369) );
INVx2_ASAP7_75t_SL g309 ( .A(n_310), .Y(n_309) );
OAI221xp5_ASAP7_75t_SL g331 ( .A1(n_310), .A2(n_332), .B1(n_334), .B2(n_336), .C(n_340), .Y(n_331) );
INVx2_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
AND2x2_ASAP7_75t_L g343 ( .A(n_312), .B(n_344), .Y(n_343) );
AND2x2_ASAP7_75t_L g349 ( .A(n_312), .B(n_333), .Y(n_349) );
AOI221xp5_ASAP7_75t_L g313 ( .A1(n_314), .A2(n_316), .B1(n_318), .B2(n_323), .C(n_324), .Y(n_313) );
INVx1_ASAP7_75t_L g432 ( .A(n_314), .Y(n_432) );
NAND2xp5_ASAP7_75t_SL g408 ( .A(n_315), .B(n_409), .Y(n_408) );
NAND2x1p5_ASAP7_75t_L g328 ( .A(n_316), .B(n_329), .Y(n_328) );
AND2x2_ASAP7_75t_L g318 ( .A(n_319), .B(n_321), .Y(n_318) );
HB1xp67_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_321), .B(n_335), .Y(n_334) );
INVx2_ASAP7_75t_L g387 ( .A(n_321), .Y(n_387) );
BUFx3_ASAP7_75t_L g410 ( .A(n_322), .Y(n_410) );
INVx1_ASAP7_75t_SL g351 ( .A(n_323), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_323), .B(n_365), .Y(n_364) );
AOI21xp33_ASAP7_75t_SL g324 ( .A1(n_325), .A2(n_326), .B(n_328), .Y(n_324) );
OAI221xp5_ASAP7_75t_L g429 ( .A1(n_325), .A2(n_426), .B1(n_430), .B2(n_432), .C(n_433), .Y(n_429) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
AND2x2_ASAP7_75t_L g372 ( .A(n_330), .B(n_333), .Y(n_372) );
INVx1_ASAP7_75t_L g436 ( .A(n_330), .Y(n_436) );
INVx2_ASAP7_75t_L g425 ( .A(n_333), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_333), .B(n_436), .Y(n_435) );
OR2x2_ASAP7_75t_L g336 ( .A(n_337), .B(n_339), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
AND2x2_ASAP7_75t_L g378 ( .A(n_338), .B(n_379), .Y(n_378) );
OAI221xp5_ASAP7_75t_SL g345 ( .A1(n_346), .A2(n_348), .B1(n_350), .B2(n_351), .C(n_352), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
INVx1_ASAP7_75t_SL g348 ( .A(n_349), .Y(n_348) );
AOI22xp33_ASAP7_75t_L g352 ( .A1(n_353), .A2(n_355), .B1(n_356), .B2(n_357), .Y(n_352) );
AOI22xp5_ASAP7_75t_L g415 ( .A1(n_354), .A2(n_416), .B1(n_417), .B2(n_419), .Y(n_415) );
OAI21xp5_ASAP7_75t_L g433 ( .A1(n_357), .A2(n_434), .B(n_437), .Y(n_433) );
NOR4xp25_ASAP7_75t_SL g358 ( .A(n_359), .B(n_367), .C(n_376), .D(n_396), .Y(n_358) );
NOR2xp33_ASAP7_75t_L g359 ( .A(n_360), .B(n_364), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
OAI22xp5_ASAP7_75t_L g367 ( .A1(n_368), .A2(n_370), .B1(n_373), .B2(n_374), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
NOR2xp33_ASAP7_75t_L g370 ( .A(n_371), .B(n_372), .Y(n_370) );
INVx1_ASAP7_75t_L g412 ( .A(n_372), .Y(n_412) );
OAI221xp5_ASAP7_75t_L g376 ( .A1(n_377), .A2(n_381), .B1(n_384), .B2(n_387), .C(n_388), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g399 ( .A(n_379), .Y(n_399) );
INVx1_ASAP7_75t_SL g382 ( .A(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
OAI21xp5_ASAP7_75t_SL g388 ( .A1(n_389), .A2(n_391), .B(n_394), .Y(n_388) );
INVx1_ASAP7_75t_SL g389 ( .A(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
OAI211xp5_ASAP7_75t_L g396 ( .A1(n_397), .A2(n_398), .B(n_400), .C(n_401), .Y(n_396) );
AOI22xp5_ASAP7_75t_L g401 ( .A1(n_402), .A2(n_403), .B1(n_404), .B2(n_405), .Y(n_401) );
CKINVDCx14_ASAP7_75t_R g411 ( .A(n_405), .Y(n_411) );
NOR3xp33_ASAP7_75t_L g406 ( .A(n_407), .B(n_421), .C(n_429), .Y(n_406) );
OAI221xp5_ASAP7_75t_L g407 ( .A1(n_408), .A2(n_411), .B1(n_412), .B2(n_413), .C(n_415), .Y(n_407) );
INVxp67_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_SL g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
CKINVDCx16_ASAP7_75t_R g430 ( .A(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
NAND3xp33_ASAP7_75t_L g445 ( .A(n_442), .B(n_446), .C(n_769), .Y(n_445) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
OAI22xp5_ASAP7_75t_SL g447 ( .A1(n_448), .A2(n_452), .B1(n_455), .B2(n_748), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
OAI22xp5_ASAP7_75t_SL g762 ( .A1(n_449), .A2(n_763), .B1(n_764), .B2(n_765), .Y(n_762) );
INVx2_ASAP7_75t_L g451 ( .A(n_450), .Y(n_451) );
INVx2_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx2_ASAP7_75t_L g763 ( .A(n_453), .Y(n_763) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
BUFx2_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVx1_ASAP7_75t_L g764 ( .A(n_456), .Y(n_764) );
AND3x1_ASAP7_75t_L g456 ( .A(n_457), .B(n_652), .C(n_709), .Y(n_456) );
NOR3xp33_ASAP7_75t_L g457 ( .A(n_458), .B(n_597), .C(n_633), .Y(n_457) );
OAI211xp5_ASAP7_75t_L g458 ( .A1(n_459), .A2(n_506), .B(n_552), .C(n_584), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_460), .B(n_479), .Y(n_459) );
HB1xp67_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
AND2x4_ASAP7_75t_L g555 ( .A(n_461), .B(n_556), .Y(n_555) );
INVx5_ASAP7_75t_L g583 ( .A(n_461), .Y(n_583) );
AND2x2_ASAP7_75t_L g656 ( .A(n_461), .B(n_572), .Y(n_656) );
AND2x2_ASAP7_75t_L g694 ( .A(n_461), .B(n_600), .Y(n_694) );
AND2x2_ASAP7_75t_L g714 ( .A(n_461), .B(n_557), .Y(n_714) );
OR2x6_ASAP7_75t_L g461 ( .A(n_462), .B(n_476), .Y(n_461) );
AOI21xp5_ASAP7_75t_SL g462 ( .A1(n_463), .A2(n_467), .B(n_475), .Y(n_462) );
BUFx2_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
INVx5_ASAP7_75t_L g499 ( .A(n_468), .Y(n_499) );
INVx2_ASAP7_75t_L g474 ( .A(n_472), .Y(n_474) );
O2A1O1Ixp33_ASAP7_75t_L g500 ( .A1(n_474), .A2(n_501), .B(n_502), .C(n_503), .Y(n_500) );
O2A1O1Ixp33_ASAP7_75t_L g535 ( .A1(n_474), .A2(n_503), .B(n_536), .C(n_537), .Y(n_535) );
NOR2xp33_ASAP7_75t_L g476 ( .A(n_477), .B(n_478), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_479), .B(n_587), .Y(n_586) );
AND2x2_ASAP7_75t_L g479 ( .A(n_480), .B(n_494), .Y(n_479) );
HB1xp67_ASAP7_75t_L g595 ( .A(n_480), .Y(n_595) );
AND2x2_ASAP7_75t_L g609 ( .A(n_480), .B(n_556), .Y(n_609) );
INVx1_ASAP7_75t_L g632 ( .A(n_480), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_480), .B(n_583), .Y(n_671) );
OR2x2_ASAP7_75t_L g708 ( .A(n_480), .B(n_554), .Y(n_708) );
INVx2_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
HB1xp67_ASAP7_75t_L g644 ( .A(n_481), .Y(n_644) );
AND2x2_ASAP7_75t_L g651 ( .A(n_481), .B(n_557), .Y(n_651) );
INVx2_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
AND2x2_ASAP7_75t_L g572 ( .A(n_482), .B(n_557), .Y(n_572) );
BUFx2_ASAP7_75t_L g600 ( .A(n_482), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_484), .B(n_491), .Y(n_483) );
INVx1_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
O2A1O1Ixp33_ASAP7_75t_L g544 ( .A1(n_490), .A2(n_499), .B(n_545), .C(n_546), .Y(n_544) );
O2A1O1Ixp33_ASAP7_75t_SL g559 ( .A1(n_490), .A2(n_499), .B(n_560), .C(n_561), .Y(n_559) );
INVx5_ASAP7_75t_L g554 ( .A(n_494), .Y(n_554) );
BUFx2_ASAP7_75t_L g576 ( .A(n_494), .Y(n_576) );
AND2x2_ASAP7_75t_L g733 ( .A(n_494), .B(n_587), .Y(n_733) );
OR2x6_ASAP7_75t_L g494 ( .A(n_495), .B(n_504), .Y(n_494) );
INVx2_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
INVx1_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
NAND2xp33_ASAP7_75t_L g507 ( .A(n_508), .B(n_539), .Y(n_507) );
OAI221xp5_ASAP7_75t_L g633 ( .A1(n_508), .A2(n_634), .B1(n_641), .B2(n_642), .C(n_645), .Y(n_633) );
OR2x2_ASAP7_75t_L g508 ( .A(n_509), .B(n_518), .Y(n_508) );
AND2x2_ASAP7_75t_L g540 ( .A(n_509), .B(n_541), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_509), .B(n_628), .Y(n_627) );
INVx1_ASAP7_75t_SL g509 ( .A(n_510), .Y(n_509) );
AND2x2_ASAP7_75t_L g568 ( .A(n_510), .B(n_519), .Y(n_568) );
NAND2xp5_ASAP7_75t_SL g578 ( .A(n_510), .B(n_520), .Y(n_578) );
OR2x2_ASAP7_75t_L g589 ( .A(n_510), .B(n_541), .Y(n_589) );
AND2x2_ASAP7_75t_L g592 ( .A(n_510), .B(n_580), .Y(n_592) );
AND2x2_ASAP7_75t_L g608 ( .A(n_510), .B(n_530), .Y(n_608) );
OR2x2_ASAP7_75t_L g624 ( .A(n_510), .B(n_520), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_510), .B(n_541), .Y(n_686) );
INVx2_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_511), .B(n_530), .Y(n_678) );
AND2x2_ASAP7_75t_L g681 ( .A(n_511), .B(n_520), .Y(n_681) );
OR2x2_ASAP7_75t_L g602 ( .A(n_518), .B(n_589), .Y(n_602) );
INVx2_ASAP7_75t_L g628 ( .A(n_518), .Y(n_628) );
OR2x2_ASAP7_75t_L g518 ( .A(n_519), .B(n_530), .Y(n_518) );
AND2x2_ASAP7_75t_L g551 ( .A(n_519), .B(n_531), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_519), .B(n_541), .Y(n_607) );
OR2x2_ASAP7_75t_L g618 ( .A(n_519), .B(n_531), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_519), .B(n_580), .Y(n_677) );
OAI221xp5_ASAP7_75t_L g710 ( .A1(n_519), .A2(n_711), .B1(n_713), .B2(n_715), .C(n_718), .Y(n_710) );
INVx5_ASAP7_75t_SL g519 ( .A(n_520), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_520), .B(n_541), .Y(n_649) );
OAI21xp5_ASAP7_75t_L g521 ( .A1(n_522), .A2(n_523), .B(n_524), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_530), .B(n_580), .Y(n_579) );
NOR2xp33_ASAP7_75t_L g590 ( .A(n_530), .B(n_591), .Y(n_590) );
AND2x2_ASAP7_75t_L g596 ( .A(n_530), .B(n_568), .Y(n_596) );
OR2x2_ASAP7_75t_L g640 ( .A(n_530), .B(n_541), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_530), .B(n_592), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_530), .B(n_685), .Y(n_684) );
AND2x2_ASAP7_75t_L g705 ( .A(n_530), .B(n_706), .Y(n_705) );
INVx5_ASAP7_75t_SL g530 ( .A(n_531), .Y(n_530) );
AND2x2_ASAP7_75t_SL g569 ( .A(n_531), .B(n_540), .Y(n_569) );
O2A1O1Ixp33_ASAP7_75t_SL g573 ( .A1(n_531), .A2(n_574), .B(n_577), .C(n_581), .Y(n_573) );
OR2x2_ASAP7_75t_L g611 ( .A(n_531), .B(n_607), .Y(n_611) );
OR2x2_ASAP7_75t_L g647 ( .A(n_531), .B(n_589), .Y(n_647) );
OAI311xp33_ASAP7_75t_L g653 ( .A1(n_531), .A2(n_592), .A3(n_654), .B1(n_657), .C1(n_664), .Y(n_653) );
AND2x2_ASAP7_75t_L g704 ( .A(n_531), .B(n_541), .Y(n_704) );
AND2x2_ASAP7_75t_L g712 ( .A(n_531), .B(n_567), .Y(n_712) );
HB1xp67_ASAP7_75t_L g730 ( .A(n_531), .Y(n_730) );
AND2x2_ASAP7_75t_L g747 ( .A(n_531), .B(n_568), .Y(n_747) );
OR2x6_ASAP7_75t_L g531 ( .A(n_532), .B(n_538), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_540), .B(n_551), .Y(n_539) );
AND2x2_ASAP7_75t_L g575 ( .A(n_540), .B(n_576), .Y(n_575) );
INVx2_ASAP7_75t_L g731 ( .A(n_540), .Y(n_731) );
AND2x2_ASAP7_75t_L g567 ( .A(n_541), .B(n_568), .Y(n_567) );
INVx3_ASAP7_75t_L g580 ( .A(n_541), .Y(n_580) );
HB1xp67_ASAP7_75t_L g623 ( .A(n_541), .Y(n_623) );
INVxp67_ASAP7_75t_L g662 ( .A(n_541), .Y(n_662) );
OA21x2_ASAP7_75t_L g541 ( .A1(n_542), .A2(n_543), .B(n_549), .Y(n_541) );
OA21x2_ASAP7_75t_L g557 ( .A1(n_550), .A2(n_558), .B(n_566), .Y(n_557) );
AND2x2_ASAP7_75t_L g740 ( .A(n_551), .B(n_588), .Y(n_740) );
AOI221xp5_ASAP7_75t_L g552 ( .A1(n_553), .A2(n_567), .B1(n_569), .B2(n_570), .C(n_573), .Y(n_552) );
AND2x2_ASAP7_75t_L g553 ( .A(n_554), .B(n_555), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_554), .B(n_572), .Y(n_571) );
AND2x2_ASAP7_75t_L g593 ( .A(n_554), .B(n_583), .Y(n_593) );
AND2x2_ASAP7_75t_L g601 ( .A(n_554), .B(n_556), .Y(n_601) );
OR2x2_ASAP7_75t_L g613 ( .A(n_554), .B(n_614), .Y(n_613) );
AND2x2_ASAP7_75t_L g631 ( .A(n_554), .B(n_632), .Y(n_631) );
AND2x2_ASAP7_75t_L g655 ( .A(n_554), .B(n_656), .Y(n_655) );
HB1xp67_ASAP7_75t_L g675 ( .A(n_554), .Y(n_675) );
AND2x2_ASAP7_75t_L g727 ( .A(n_554), .B(n_651), .Y(n_727) );
OAI31xp33_ASAP7_75t_L g735 ( .A1(n_554), .A2(n_604), .A3(n_703), .B(n_736), .Y(n_735) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_555), .B(n_631), .Y(n_630) );
INVx1_ASAP7_75t_SL g699 ( .A(n_555), .Y(n_699) );
NOR2xp33_ASAP7_75t_L g707 ( .A(n_555), .B(n_708), .Y(n_707) );
AND2x4_ASAP7_75t_L g587 ( .A(n_556), .B(n_583), .Y(n_587) );
INVx1_ASAP7_75t_L g674 ( .A(n_556), .Y(n_674) );
INVx2_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
AND2x2_ASAP7_75t_L g724 ( .A(n_557), .B(n_583), .Y(n_724) );
NOR2xp33_ASAP7_75t_L g562 ( .A(n_563), .B(n_564), .Y(n_562) );
INVx1_ASAP7_75t_SL g734 ( .A(n_567), .Y(n_734) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_568), .B(n_639), .Y(n_638) );
AOI22xp5_ASAP7_75t_L g718 ( .A1(n_569), .A2(n_681), .B1(n_719), .B2(n_722), .Y(n_718) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
AND2x2_ASAP7_75t_L g582 ( .A(n_572), .B(n_583), .Y(n_582) );
INVx1_ASAP7_75t_L g641 ( .A(n_572), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g746 ( .A(n_572), .B(n_593), .Y(n_746) );
INVx1_ASAP7_75t_SL g574 ( .A(n_575), .Y(n_574) );
AND2x2_ASAP7_75t_L g716 ( .A(n_575), .B(n_717), .Y(n_716) );
AOI21xp5_ASAP7_75t_L g634 ( .A1(n_576), .A2(n_635), .B(n_637), .Y(n_634) );
OR2x2_ASAP7_75t_L g642 ( .A(n_576), .B(n_643), .Y(n_642) );
AND2x2_ASAP7_75t_L g663 ( .A(n_576), .B(n_651), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_576), .B(n_674), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_576), .B(n_714), .Y(n_713) );
OAI221xp5_ASAP7_75t_SL g690 ( .A1(n_577), .A2(n_691), .B1(n_696), .B2(n_699), .C(n_700), .Y(n_690) );
OR2x2_ASAP7_75t_L g577 ( .A(n_578), .B(n_579), .Y(n_577) );
OR2x2_ASAP7_75t_L g667 ( .A(n_578), .B(n_640), .Y(n_667) );
INVx1_ASAP7_75t_L g706 ( .A(n_578), .Y(n_706) );
INVx2_ASAP7_75t_L g682 ( .A(n_579), .Y(n_682) );
INVx1_ASAP7_75t_L g616 ( .A(n_580), .Y(n_616) );
INVx1_ASAP7_75t_SL g581 ( .A(n_582), .Y(n_581) );
INVx2_ASAP7_75t_L g621 ( .A(n_583), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_583), .B(n_644), .Y(n_643) );
AND2x2_ASAP7_75t_L g650 ( .A(n_583), .B(n_651), .Y(n_650) );
OR2x2_ASAP7_75t_L g738 ( .A(n_583), .B(n_708), .Y(n_738) );
AOI222xp33_ASAP7_75t_L g584 ( .A1(n_585), .A2(n_588), .B1(n_590), .B2(n_593), .C1(n_594), .C2(n_596), .Y(n_584) );
INVxp67_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
AND2x2_ASAP7_75t_L g594 ( .A(n_587), .B(n_595), .Y(n_594) );
AOI22xp33_ASAP7_75t_L g664 ( .A1(n_587), .A2(n_637), .B1(n_665), .B2(n_666), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_587), .B(n_721), .Y(n_720) );
INVx1_ASAP7_75t_SL g588 ( .A(n_589), .Y(n_588) );
INVx1_ASAP7_75t_SL g591 ( .A(n_592), .Y(n_591) );
OAI21xp33_ASAP7_75t_SL g625 ( .A1(n_596), .A2(n_626), .B(n_629), .Y(n_625) );
OAI211xp5_ASAP7_75t_SL g597 ( .A1(n_598), .A2(n_602), .B(n_603), .C(n_625), .Y(n_597) );
INVxp67_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
AND2x2_ASAP7_75t_L g599 ( .A(n_600), .B(n_601), .Y(n_599) );
AOI221xp5_ASAP7_75t_L g603 ( .A1(n_601), .A2(n_604), .B1(n_609), .B2(n_610), .C(n_612), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_601), .B(n_689), .Y(n_688) );
INVxp67_ASAP7_75t_L g695 ( .A(n_601), .Y(n_695) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_606), .B(n_608), .Y(n_605) );
AND2x2_ASAP7_75t_L g697 ( .A(n_606), .B(n_698), .Y(n_697) );
INVx1_ASAP7_75t_SL g606 ( .A(n_607), .Y(n_606) );
INVx1_ASAP7_75t_L g614 ( .A(n_609), .Y(n_614) );
AND2x2_ASAP7_75t_L g620 ( .A(n_609), .B(n_621), .Y(n_620) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
OAI22xp5_ASAP7_75t_L g612 ( .A1(n_613), .A2(n_615), .B1(n_619), .B2(n_622), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_616), .B(n_617), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_616), .B(n_628), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_617), .B(n_662), .Y(n_661) );
INVx1_ASAP7_75t_SL g617 ( .A(n_618), .Y(n_617) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
INVx1_ASAP7_75t_L g717 ( .A(n_621), .Y(n_717) );
AND2x2_ASAP7_75t_L g736 ( .A(n_621), .B(n_651), .Y(n_736) );
OR2x2_ASAP7_75t_L g622 ( .A(n_623), .B(n_624), .Y(n_622) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g744 ( .A(n_628), .B(n_685), .Y(n_744) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
NOR2xp33_ASAP7_75t_L g742 ( .A(n_631), .B(n_699), .Y(n_742) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
INVx1_ASAP7_75t_L g665 ( .A(n_643), .Y(n_665) );
BUFx2_ASAP7_75t_L g689 ( .A(n_644), .Y(n_689) );
OAI21xp5_ASAP7_75t_SL g645 ( .A1(n_646), .A2(n_648), .B(n_650), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
NOR3xp33_ASAP7_75t_L g652 ( .A(n_653), .B(n_668), .C(n_690), .Y(n_652) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
OAI21xp5_ASAP7_75t_L g657 ( .A1(n_658), .A2(n_660), .B(n_663), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
INVx1_ASAP7_75t_SL g666 ( .A(n_667), .Y(n_666) );
A2O1A1Ixp33_ASAP7_75t_SL g668 ( .A1(n_669), .A2(n_672), .B(n_676), .C(n_679), .Y(n_668) );
NAND2xp5_ASAP7_75t_SL g701 ( .A(n_669), .B(n_702), .Y(n_701) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
NOR2xp67_ASAP7_75t_SL g673 ( .A(n_674), .B(n_675), .Y(n_673) );
OR2x2_ASAP7_75t_L g676 ( .A(n_677), .B(n_678), .Y(n_676) );
INVx1_ASAP7_75t_SL g698 ( .A(n_678), .Y(n_698) );
OAI21xp5_ASAP7_75t_L g679 ( .A1(n_680), .A2(n_683), .B(n_687), .Y(n_679) );
AND2x4_ASAP7_75t_L g680 ( .A(n_681), .B(n_682), .Y(n_680) );
AND2x2_ASAP7_75t_L g703 ( .A(n_681), .B(n_704), .Y(n_703) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
INVx1_ASAP7_75t_SL g685 ( .A(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
NOR2xp33_ASAP7_75t_L g692 ( .A(n_693), .B(n_695), .Y(n_692) );
INVx2_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
AOI22xp33_ASAP7_75t_L g700 ( .A1(n_701), .A2(n_703), .B1(n_705), .B2(n_707), .Y(n_700) );
INVx2_ASAP7_75t_SL g721 ( .A(n_708), .Y(n_721) );
NOR3xp33_ASAP7_75t_L g709 ( .A(n_710), .B(n_725), .C(n_737), .Y(n_709) );
INVx1_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
INVxp67_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
INVxp67_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_721), .B(n_724), .Y(n_723) );
INVx1_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
OAI221xp5_ASAP7_75t_L g725 ( .A1(n_726), .A2(n_728), .B1(n_732), .B2(n_734), .C(n_735), .Y(n_725) );
A2O1A1Ixp33_ASAP7_75t_L g737 ( .A1(n_726), .A2(n_738), .B(n_739), .C(n_741), .Y(n_737) );
INVx1_ASAP7_75t_SL g726 ( .A(n_727), .Y(n_726) );
INVxp67_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
NOR2xp33_ASAP7_75t_L g729 ( .A(n_730), .B(n_731), .Y(n_729) );
INVx1_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
INVx1_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
AOI22xp5_ASAP7_75t_L g741 ( .A1(n_742), .A2(n_743), .B1(n_745), .B2(n_747), .Y(n_741) );
INVx1_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
INVx1_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
INVx2_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
INVx2_ASAP7_75t_L g765 ( .A(n_749), .Y(n_765) );
INVx1_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
INVx1_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
INVx1_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
INVx1_ASAP7_75t_L g760 ( .A(n_757), .Y(n_760) );
INVx1_ASAP7_75t_SL g766 ( .A(n_767), .Y(n_766) );
INVx3_ASAP7_75t_SL g767 ( .A(n_768), .Y(n_767) );
CKINVDCx20_ASAP7_75t_R g769 ( .A(n_770), .Y(n_769) );
endmodule