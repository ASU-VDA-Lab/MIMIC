module real_jpeg_18296_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_247;
wire n_146;
wire n_78;
wire n_83;
wire n_249;
wire n_215;
wire n_176;
wire n_166;
wire n_292;
wire n_221;
wire n_286;
wire n_288;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_281;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_237;
wire n_174;
wire n_87;
wire n_197;
wire n_105;
wire n_40;
wire n_299;
wire n_173;
wire n_243;
wire n_115;
wire n_255;
wire n_98;
wire n_27;
wire n_200;
wire n_56;
wire n_48;
wire n_164;
wire n_184;
wire n_275;
wire n_293;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_139;
wire n_188;
wire n_33;
wire n_65;
wire n_142;
wire n_175;
wire n_76;
wire n_238;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_290;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_211;
wire n_160;
wire n_45;
wire n_285;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_294;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_298;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_296;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_195;
wire n_61;
wire n_110;
wire n_205;
wire n_258;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_150;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_70;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_259;
wire n_225;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_297;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_187;
wire n_75;
wire n_97;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_128;
wire n_202;
wire n_213;
wire n_167;
wire n_179;
wire n_216;
wire n_133;
wire n_244;
wire n_295;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_210;
wire n_127;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_283;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_253;
wire n_96;
wire n_269;
wire n_273;
wire n_89;
wire n_16;

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_0),
.A2(n_15),
.B(n_298),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_0),
.B(n_299),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_1),
.Y(n_299)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_2),
.B(n_38),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_2),
.B(n_55),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_2),
.B(n_46),
.Y(n_62)
);

AND2x4_ASAP7_75t_L g84 ( 
.A(n_2),
.B(n_85),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_2),
.B(n_98),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_2),
.B(n_113),
.Y(n_112)
);

NAND2x1_ASAP7_75t_SL g133 ( 
.A(n_2),
.B(n_134),
.Y(n_133)
);

NAND2x1_ASAP7_75t_L g171 ( 
.A(n_2),
.B(n_172),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_4),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_5),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_5),
.Y(n_55)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_5),
.Y(n_66)
);

INVx2_ASAP7_75t_SL g35 ( 
.A(n_6),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_6),
.B(n_80),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_6),
.B(n_46),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_6),
.B(n_89),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g201 ( 
.A(n_6),
.B(n_202),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_6),
.B(n_251),
.Y(n_250)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_7),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_7),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g294 ( 
.A(n_7),
.Y(n_294)
);

AND2x2_ASAP7_75t_SL g25 ( 
.A(n_8),
.B(n_26),
.Y(n_25)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_8),
.B(n_44),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_8),
.B(n_64),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_8),
.B(n_69),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_8),
.B(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_8),
.Y(n_129)
);

AND2x2_ASAP7_75t_SL g162 ( 
.A(n_8),
.B(n_163),
.Y(n_162)
);

AND2x2_ASAP7_75t_SL g210 ( 
.A(n_8),
.B(n_211),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_9),
.B(n_176),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_9),
.B(n_215),
.Y(n_214)
);

AND2x2_ASAP7_75t_L g236 ( 
.A(n_9),
.B(n_237),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_9),
.B(n_292),
.Y(n_291)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_10),
.Y(n_134)
);

INVx6_ASAP7_75t_L g164 ( 
.A(n_10),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_11),
.Y(n_86)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_12),
.Y(n_46)
);

BUFx4f_ASAP7_75t_L g217 ( 
.A(n_12),
.Y(n_217)
);

BUFx8_ASAP7_75t_L g172 ( 
.A(n_13),
.Y(n_172)
);

BUFx5_ASAP7_75t_L g211 ( 
.A(n_13),
.Y(n_211)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_13),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_265),
.Y(n_15)
);

AOI21xp5_ASAP7_75t_L g16 ( 
.A1(n_17),
.A2(n_223),
.B(n_259),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_188),
.Y(n_18)
);

OAI21xp5_ASAP7_75t_SL g19 ( 
.A1(n_20),
.A2(n_150),
.B(n_187),
.Y(n_19)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_122),
.B(n_149),
.Y(n_20)
);

OAI21xp5_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_94),
.B(n_121),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_57),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_23),
.B(n_57),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_42),
.C(n_51),
.Y(n_23)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_24),
.B(n_105),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_30),
.B1(n_40),
.B2(n_41),
.Y(n_24)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_25),
.A2(n_40),
.B1(n_139),
.B2(n_142),
.Y(n_138)
);

O2A1O1Ixp5_ASAP7_75t_L g157 ( 
.A1(n_25),
.A2(n_103),
.B(n_112),
.C(n_140),
.Y(n_157)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_31),
.A2(n_32),
.B1(n_36),
.B2(n_37),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_31),
.A2(n_32),
.B1(n_128),
.B2(n_135),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_31),
.B(n_135),
.C(n_195),
.Y(n_231)
);

CKINVDCx14_ASAP7_75t_R g31 ( 
.A(n_32),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_32),
.B(n_36),
.C(n_40),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_32),
.B(n_289),
.Y(n_288)
);

OR2x4_ASAP7_75t_SL g32 ( 
.A(n_33),
.B(n_35),
.Y(n_32)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_33),
.Y(n_113)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_33),
.Y(n_237)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_34),
.Y(n_71)
);

OR2x2_ASAP7_75t_L g48 ( 
.A(n_35),
.B(n_49),
.Y(n_48)
);

OR2x2_ASAP7_75t_L g180 ( 
.A(n_35),
.B(n_181),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_36),
.A2(n_37),
.B1(n_162),
.B2(n_165),
.Y(n_257)
);

INVx2_ASAP7_75t_SL g36 ( 
.A(n_37),
.Y(n_36)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_37),
.B(n_200),
.Y(n_199)
);

AO21x1_ASAP7_75t_L g245 ( 
.A1(n_37),
.A2(n_246),
.B(n_247),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_37),
.B(n_79),
.C(n_162),
.Y(n_278)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_42),
.A2(n_51),
.B1(n_52),
.B2(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_42),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_42),
.A2(n_43),
.B(n_47),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_47),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_43),
.A2(n_53),
.B1(n_54),
.B2(n_56),
.Y(n_52)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_47),
.A2(n_48),
.B1(n_61),
.B2(n_62),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_47),
.A2(n_48),
.B1(n_213),
.B2(n_214),
.Y(n_212)
);

INVx1_ASAP7_75t_SL g47 ( 
.A(n_48),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_48),
.B(n_210),
.C(n_214),
.Y(n_233)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_53),
.A2(n_54),
.B1(n_100),
.B2(n_101),
.Y(n_254)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_L g72 ( 
.A1(n_54),
.A2(n_62),
.B(n_73),
.Y(n_72)
);

NAND2x1_ASAP7_75t_L g73 ( 
.A(n_54),
.B(n_62),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_54),
.B(n_100),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g287 ( 
.A1(n_54),
.A2(n_100),
.B(n_250),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_76),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_58),
.B(n_77),
.C(n_93),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_67),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_60),
.A2(n_109),
.B(n_114),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_60),
.A2(n_68),
.B(n_75),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_63),
.Y(n_60)
);

INVx2_ASAP7_75t_SL g61 ( 
.A(n_62),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_63),
.A2(n_100),
.B1(n_101),
.B2(n_102),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_63),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_66),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_68),
.A2(n_72),
.B1(n_74),
.B2(n_75),
.Y(n_67)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_68),
.Y(n_74)
);

O2A1O1Ixp33_ASAP7_75t_SL g96 ( 
.A1(n_68),
.A2(n_97),
.B(n_99),
.C(n_103),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_68),
.B(n_97),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_68),
.A2(n_74),
.B1(n_97),
.B2(n_118),
.Y(n_117)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_72),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_72),
.A2(n_75),
.B1(n_132),
.B2(n_133),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_73),
.B(n_127),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_73),
.B(n_128),
.C(n_133),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_77),
.A2(n_78),
.B1(n_92),
.B2(n_93),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_82),
.B1(n_83),
.B2(n_91),
.Y(n_78)
);

INVx1_ASAP7_75t_SL g91 ( 
.A(n_79),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_79),
.B(n_84),
.C(n_146),
.Y(n_145)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_87),
.Y(n_83)
);

AOI22x1_ASAP7_75t_SL g234 ( 
.A1(n_84),
.A2(n_235),
.B1(n_236),
.B2(n_238),
.Y(n_234)
);

INVx2_ASAP7_75t_SL g235 ( 
.A(n_84),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_84),
.B(n_233),
.C(n_236),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_84),
.B(n_209),
.Y(n_280)
);

BUFx5_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_86),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_86),
.Y(n_184)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_87),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_SL g160 ( 
.A(n_87),
.B(n_161),
.Y(n_160)
);

BUFx2_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_91),
.B(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_95),
.A2(n_107),
.B(n_120),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_104),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_96),
.B(n_104),
.Y(n_120)
);

INVx1_ASAP7_75t_SL g118 ( 
.A(n_97),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_97),
.B(n_111),
.Y(n_169)
);

MAJx2_ASAP7_75t_L g195 ( 
.A(n_97),
.B(n_112),
.C(n_171),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_97),
.A2(n_118),
.B1(n_199),
.B2(n_203),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g247 ( 
.A(n_97),
.B(n_201),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_99),
.B(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_SL g101 ( 
.A(n_100),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_100),
.A2(n_101),
.B1(n_162),
.B2(n_165),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_100),
.B(n_146),
.C(n_162),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_106),
.B(n_116),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_106),
.B(n_116),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_115),
.B(n_119),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_110),
.B(n_111),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_110),
.B(n_111),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_111),
.A2(n_112),
.B1(n_140),
.B2(n_141),
.Y(n_139)
);

INVx2_ASAP7_75t_SL g111 ( 
.A(n_112),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_118),
.B(n_200),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_124),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_123),
.B(n_124),
.Y(n_149)
);

XOR2x2_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_137),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_136),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_126),
.B(n_136),
.C(n_137),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_128),
.A2(n_132),
.B1(n_133),
.B2(n_135),
.Y(n_127)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_128),
.Y(n_135)
);

OR2x2_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_130),
.Y(n_128)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_SL g132 ( 
.A(n_133),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_SL g137 ( 
.A(n_138),
.B(n_143),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_138),
.B(n_144),
.C(n_148),
.Y(n_154)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_139),
.Y(n_142)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_140),
.Y(n_141)
);

AO22x1_ASAP7_75t_L g289 ( 
.A1(n_140),
.A2(n_141),
.B1(n_290),
.B2(n_291),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_144),
.A2(n_145),
.B1(n_147),
.B2(n_148),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

NOR2xp67_ASAP7_75t_SL g150 ( 
.A(n_151),
.B(n_152),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_151),
.B(n_152),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_166),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_155),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_154),
.B(n_155),
.C(n_166),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_160),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_158),
.Y(n_156)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_157),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_158),
.B(n_160),
.C(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_159),
.B(n_287),
.Y(n_286)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_162),
.Y(n_165)
);

INVx3_ASAP7_75t_SL g163 ( 
.A(n_164),
.Y(n_163)
);

INVx4_ASAP7_75t_L g202 ( 
.A(n_164),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_SL g166 ( 
.A(n_167),
.B(n_186),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_174),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_168),
.B(n_174),
.C(n_186),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_169),
.A2(n_170),
.B1(n_171),
.B2(n_173),
.Y(n_168)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_169),
.Y(n_173)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_175),
.A2(n_180),
.B(n_185),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_175),
.B(n_180),
.Y(n_185)
);

BUFx2_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_185),
.A2(n_219),
.B1(n_220),
.B2(n_221),
.Y(n_218)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_185),
.Y(n_221)
);

OR2x2_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_190),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_189),
.B(n_190),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_206),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_191),
.B(n_207),
.C(n_222),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_204),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_193),
.A2(n_194),
.B1(n_197),
.B2(n_198),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_194),
.B(n_197),
.C(n_204),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_196),
.Y(n_194)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_199),
.Y(n_203)
);

INVx1_ASAP7_75t_SL g200 ( 
.A(n_201),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_222),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_218),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_208),
.B(n_220),
.C(n_221),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_212),
.Y(n_208)
);

INVx1_ASAP7_75t_SL g209 ( 
.A(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_223),
.Y(n_260)
);

OR2x2_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_258),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_224),
.B(n_258),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_226),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_225),
.B(n_227),
.C(n_242),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_227),
.A2(n_228),
.B1(n_241),
.B2(n_242),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_230),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_229),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_231),
.A2(n_232),
.B1(n_239),
.B2(n_240),
.Y(n_230)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_231),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_231),
.B(n_270),
.C(n_271),
.Y(n_269)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_232),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_234),
.Y(n_232)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_236),
.Y(n_238)
);

HB1xp67_ASAP7_75t_L g271 ( 
.A(n_239),
.Y(n_271)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

XNOR2x1_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_255),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_244),
.A2(n_245),
.B1(n_248),
.B2(n_249),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_245),
.B(n_248),
.C(n_256),
.Y(n_283)
);

INVx1_ASAP7_75t_SL g248 ( 
.A(n_249),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_254),
.Y(n_249)
);

INVx5_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_261),
.Y(n_259)
);

INVxp33_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_263),
.B(n_264),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_296),
.Y(n_265)
);

NOR2x1_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_268),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_267),
.B(n_268),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_272),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_284),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_283),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_275),
.A2(n_276),
.B1(n_281),
.B2(n_282),
.Y(n_274)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_275),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_276),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_277),
.A2(n_278),
.B1(n_279),
.B2(n_280),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

XOR2x1_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_295),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_288),
.Y(n_285)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx6_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVxp33_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);


endmodule