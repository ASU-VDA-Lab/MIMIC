module fake_jpeg_2837_n_577 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_577);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_577;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx13_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

BUFx16f_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_12),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

BUFx10_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

INVxp67_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

BUFx12_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_9),
.Y(n_45)
);

BUFx4f_ASAP7_75t_L g46 ( 
.A(n_6),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_10),
.B(n_6),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_18),
.Y(n_48)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_8),
.Y(n_49)
);

BUFx16f_ASAP7_75t_L g50 ( 
.A(n_8),
.Y(n_50)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_13),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_16),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_16),
.B(n_9),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_50),
.Y(n_54)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_54),
.Y(n_111)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_29),
.Y(n_55)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_55),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_33),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_56),
.B(n_62),
.Y(n_116)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_25),
.Y(n_57)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_57),
.Y(n_141)
);

INVx13_ASAP7_75t_L g58 ( 
.A(n_50),
.Y(n_58)
);

INVx13_ASAP7_75t_L g110 ( 
.A(n_58),
.Y(n_110)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_25),
.Y(n_59)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_59),
.Y(n_142)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_50),
.Y(n_60)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_60),
.Y(n_113)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_33),
.Y(n_61)
);

BUFx4f_ASAP7_75t_SL g137 ( 
.A(n_61),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_53),
.B(n_47),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_50),
.Y(n_63)
);

INVx5_ASAP7_75t_L g121 ( 
.A(n_63),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_22),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_64),
.Y(n_112)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_65),
.Y(n_118)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_66),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_22),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_67),
.Y(n_130)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_19),
.Y(n_68)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_68),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_53),
.B(n_18),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_69),
.B(n_70),
.Y(n_124)
);

INVx1_ASAP7_75t_SL g70 ( 
.A(n_20),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_21),
.Y(n_71)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_71),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_22),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_72),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_47),
.B(n_29),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_73),
.B(n_92),
.Y(n_134)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_40),
.Y(n_74)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_74),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_33),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_75),
.B(n_94),
.Y(n_128)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_76),
.Y(n_149)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_19),
.Y(n_77)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_77),
.Y(n_138)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_49),
.Y(n_78)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_78),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_28),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_79),
.Y(n_145)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_40),
.Y(n_80)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_80),
.Y(n_127)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_21),
.Y(n_81)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_81),
.Y(n_117)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_46),
.Y(n_82)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_82),
.Y(n_132)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_39),
.Y(n_83)
);

INVx5_ASAP7_75t_L g159 ( 
.A(n_83),
.Y(n_159)
);

BUFx5_ASAP7_75t_L g84 ( 
.A(n_33),
.Y(n_84)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_84),
.Y(n_126)
);

BUFx16f_ASAP7_75t_L g85 ( 
.A(n_20),
.Y(n_85)
);

BUFx24_ASAP7_75t_L g109 ( 
.A(n_85),
.Y(n_109)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_39),
.Y(n_86)
);

INVx5_ASAP7_75t_L g172 ( 
.A(n_86),
.Y(n_172)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_26),
.Y(n_87)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_87),
.Y(n_140)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_51),
.Y(n_88)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_88),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_28),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_89),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_28),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_90),
.Y(n_154)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_46),
.Y(n_91)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_91),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_30),
.B(n_18),
.Y(n_92)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_35),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_93),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_30),
.B(n_15),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_21),
.Y(n_95)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_95),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_52),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_96),
.B(n_97),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_52),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_35),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_98),
.Y(n_168)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_26),
.Y(n_99)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_99),
.Y(n_158)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_51),
.Y(n_100)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_100),
.Y(n_165)
);

BUFx5_ASAP7_75t_L g101 ( 
.A(n_31),
.Y(n_101)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_101),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_35),
.Y(n_102)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_102),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_52),
.Y(n_103)
);

INVx6_ASAP7_75t_L g146 ( 
.A(n_103),
.Y(n_146)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_46),
.Y(n_104)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_104),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_39),
.Y(n_105)
);

INVx6_ASAP7_75t_L g160 ( 
.A(n_105),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_43),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_106),
.B(n_48),
.Y(n_155)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_24),
.Y(n_107)
);

INVx8_ASAP7_75t_L g150 ( 
.A(n_107),
.Y(n_150)
);

BUFx5_ASAP7_75t_L g108 ( 
.A(n_31),
.Y(n_108)
);

INVx11_ASAP7_75t_L g163 ( 
.A(n_108),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_85),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_114),
.B(n_148),
.Y(n_174)
);

BUFx12_ASAP7_75t_L g115 ( 
.A(n_58),
.Y(n_115)
);

BUFx12f_ASAP7_75t_L g220 ( 
.A(n_115),
.Y(n_220)
);

AOI21xp33_ASAP7_75t_SL g122 ( 
.A1(n_54),
.A2(n_60),
.B(n_63),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_122),
.B(n_32),
.C(n_20),
.Y(n_203)
);

HB1xp67_ASAP7_75t_L g129 ( 
.A(n_70),
.Y(n_129)
);

BUFx2_ASAP7_75t_L g234 ( 
.A(n_129),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_103),
.A2(n_93),
.B1(n_64),
.B2(n_72),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_139),
.A2(n_151),
.B1(n_41),
.B2(n_34),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_107),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_67),
.A2(n_23),
.B1(n_48),
.B2(n_46),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_155),
.B(n_61),
.Y(n_176)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_57),
.Y(n_156)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_156),
.Y(n_177)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_59),
.Y(n_161)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_161),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_76),
.A2(n_23),
.B1(n_88),
.B2(n_100),
.Y(n_162)
);

OA22x2_ASAP7_75t_L g178 ( 
.A1(n_162),
.A2(n_81),
.B1(n_71),
.B2(n_95),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_105),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_164),
.B(n_84),
.Y(n_185)
);

INVx11_ASAP7_75t_L g169 ( 
.A(n_61),
.Y(n_169)
);

INVx4_ASAP7_75t_L g221 ( 
.A(n_169),
.Y(n_221)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_78),
.Y(n_170)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_170),
.Y(n_208)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_79),
.Y(n_171)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_171),
.Y(n_213)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_118),
.Y(n_173)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_173),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_134),
.B(n_124),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_175),
.B(n_176),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_178),
.A2(n_229),
.B1(n_44),
.B2(n_2),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_162),
.A2(n_90),
.B1(n_102),
.B2(n_89),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_179),
.A2(n_184),
.B1(n_206),
.B2(n_209),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_112),
.Y(n_180)
);

BUFx2_ASAP7_75t_L g245 ( 
.A(n_180),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_116),
.B(n_86),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_181),
.B(n_182),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_116),
.B(n_83),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_124),
.B(n_39),
.Y(n_183)
);

OR2x2_ASAP7_75t_L g254 ( 
.A(n_183),
.B(n_211),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_120),
.A2(n_98),
.B1(n_24),
.B2(n_27),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_185),
.B(n_186),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_128),
.B(n_42),
.Y(n_186)
);

INVx6_ASAP7_75t_L g187 ( 
.A(n_112),
.Y(n_187)
);

BUFx2_ASAP7_75t_L g255 ( 
.A(n_187),
.Y(n_255)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_159),
.Y(n_188)
);

INVx4_ASAP7_75t_L g239 ( 
.A(n_188),
.Y(n_239)
);

INVx6_ASAP7_75t_L g189 ( 
.A(n_130),
.Y(n_189)
);

INVx4_ASAP7_75t_L g241 ( 
.A(n_189),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_128),
.B(n_42),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_190),
.B(n_193),
.Y(n_256)
);

BUFx16f_ASAP7_75t_L g191 ( 
.A(n_109),
.Y(n_191)
);

BUFx12f_ASAP7_75t_L g269 ( 
.A(n_191),
.Y(n_269)
);

BUFx10_ASAP7_75t_L g192 ( 
.A(n_115),
.Y(n_192)
);

INVx4_ASAP7_75t_L g277 ( 
.A(n_192),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_125),
.B(n_37),
.Y(n_193)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_157),
.Y(n_195)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_195),
.Y(n_268)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_130),
.Y(n_196)
);

INVx3_ASAP7_75t_L g252 ( 
.A(n_196),
.Y(n_252)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_129),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_197),
.B(n_199),
.Y(n_287)
);

INVx6_ASAP7_75t_L g198 ( 
.A(n_136),
.Y(n_198)
);

INVx3_ASAP7_75t_L g275 ( 
.A(n_198),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_133),
.B(n_37),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_157),
.Y(n_200)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_200),
.Y(n_237)
);

CKINVDCx14_ASAP7_75t_SL g201 ( 
.A(n_110),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_201),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_138),
.B(n_32),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_202),
.B(n_205),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g284 ( 
.A(n_203),
.B(n_228),
.Y(n_284)
);

BUFx3_ASAP7_75t_L g204 ( 
.A(n_111),
.Y(n_204)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_204),
.Y(n_274)
);

OR2x2_ASAP7_75t_L g205 ( 
.A(n_140),
.B(n_36),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_123),
.A2(n_24),
.B1(n_45),
.B2(n_36),
.Y(n_206)
);

INVx8_ASAP7_75t_L g207 ( 
.A(n_160),
.Y(n_207)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_207),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_127),
.A2(n_45),
.B1(n_27),
.B2(n_41),
.Y(n_209)
);

INVx8_ASAP7_75t_L g210 ( 
.A(n_160),
.Y(n_210)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_210),
.Y(n_282)
);

CKINVDCx9p33_ASAP7_75t_R g211 ( 
.A(n_109),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_158),
.Y(n_212)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_212),
.Y(n_238)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_172),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g265 ( 
.A(n_214),
.Y(n_265)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_136),
.Y(n_215)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_215),
.Y(n_242)
);

INVx6_ASAP7_75t_L g216 ( 
.A(n_168),
.Y(n_216)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_216),
.Y(n_246)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_132),
.Y(n_217)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_217),
.Y(n_264)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_144),
.Y(n_218)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_218),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_L g249 ( 
.A1(n_219),
.A2(n_163),
.B1(n_166),
.B2(n_145),
.Y(n_249)
);

BUFx5_ASAP7_75t_L g222 ( 
.A(n_110),
.Y(n_222)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_222),
.Y(n_280)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_152),
.Y(n_223)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_223),
.Y(n_286)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_141),
.Y(n_224)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_224),
.Y(n_288)
);

A2O1A1Ixp33_ASAP7_75t_L g225 ( 
.A1(n_137),
.A2(n_108),
.B(n_101),
.C(n_41),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_225),
.B(n_41),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_142),
.B(n_17),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_226),
.B(n_227),
.Y(n_279)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_149),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_153),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_135),
.B(n_17),
.Y(n_229)
);

INVx2_ASAP7_75t_SL g230 ( 
.A(n_143),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_230),
.Y(n_240)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_165),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_231),
.Y(n_258)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_113),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_232),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_137),
.B(n_0),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_233),
.B(n_235),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_145),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_203),
.A2(n_183),
.B1(n_205),
.B2(n_179),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g329 ( 
.A1(n_243),
.A2(n_249),
.B1(n_259),
.B2(n_273),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_178),
.A2(n_167),
.B1(n_150),
.B2(n_119),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_244),
.B(n_250),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_178),
.A2(n_167),
.B1(n_150),
.B2(n_119),
.Y(n_250)
);

AND2x2_ASAP7_75t_L g296 ( 
.A(n_251),
.B(n_263),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_184),
.A2(n_146),
.B1(n_154),
.B2(n_147),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_257),
.B(n_261),
.Y(n_319)
);

AOI22xp33_ASAP7_75t_L g259 ( 
.A1(n_206),
.A2(n_209),
.B1(n_154),
.B2(n_168),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_187),
.A2(n_146),
.B1(n_147),
.B2(n_117),
.Y(n_261)
);

AO22x1_ASAP7_75t_SL g263 ( 
.A1(n_225),
.A2(n_126),
.B1(n_131),
.B2(n_41),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_174),
.B(n_213),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_272),
.B(n_283),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_189),
.A2(n_121),
.B1(n_44),
.B2(n_34),
.Y(n_273)
);

AND2x2_ASAP7_75t_L g308 ( 
.A(n_276),
.B(n_285),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_177),
.B(n_44),
.C(n_2),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_281),
.B(n_211),
.C(n_191),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_194),
.B(n_1),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_198),
.A2(n_44),
.B1(n_3),
.B2(n_4),
.Y(n_285)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_246),
.Y(n_289)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_289),
.Y(n_361)
);

INVx13_ASAP7_75t_L g290 ( 
.A(n_269),
.Y(n_290)
);

INVx1_ASAP7_75t_SL g377 ( 
.A(n_290),
.Y(n_377)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_246),
.Y(n_291)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_291),
.Y(n_337)
);

AND2x2_ASAP7_75t_SL g292 ( 
.A(n_284),
.B(n_201),
.Y(n_292)
);

AND2x2_ASAP7_75t_L g368 ( 
.A(n_292),
.B(n_314),
.Y(n_368)
);

OAI21xp5_ASAP7_75t_L g293 ( 
.A1(n_248),
.A2(n_272),
.B(n_284),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_L g356 ( 
.A1(n_293),
.A2(n_303),
.B(n_311),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_268),
.B(n_234),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_294),
.B(n_299),
.Y(n_352)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_275),
.Y(n_295)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_295),
.Y(n_338)
);

BUFx12f_ASAP7_75t_L g297 ( 
.A(n_252),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_297),
.B(n_316),
.Y(n_348)
);

INVx13_ASAP7_75t_L g298 ( 
.A(n_269),
.Y(n_298)
);

CKINVDCx16_ASAP7_75t_R g367 ( 
.A(n_298),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_237),
.B(n_234),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g366 ( 
.A(n_300),
.B(n_274),
.Y(n_366)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_238),
.Y(n_301)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_301),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_247),
.B(n_208),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_302),
.B(n_321),
.Y(n_340)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_251),
.A2(n_191),
.B(n_230),
.Y(n_303)
);

INVx5_ASAP7_75t_L g304 ( 
.A(n_252),
.Y(n_304)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_304),
.Y(n_357)
);

INVx13_ASAP7_75t_L g305 ( 
.A(n_269),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_305),
.Y(n_379)
);

INVx3_ASAP7_75t_L g306 ( 
.A(n_278),
.Y(n_306)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_306),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_284),
.B(n_214),
.C(n_188),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_307),
.B(n_265),
.C(n_264),
.Y(n_349)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_238),
.Y(n_309)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_309),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_237),
.B(n_232),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g359 ( 
.A(n_310),
.B(n_315),
.Y(n_359)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_254),
.A2(n_276),
.B(n_253),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g313 ( 
.A1(n_254),
.A2(n_221),
.B(n_222),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_L g362 ( 
.A1(n_313),
.A2(n_326),
.B(n_265),
.Y(n_362)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_288),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_SL g315 ( 
.A(n_267),
.B(n_204),
.Y(n_315)
);

AOI32xp33_ASAP7_75t_L g316 ( 
.A1(n_271),
.A2(n_221),
.A3(n_210),
.B1(n_207),
.B2(n_192),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_256),
.B(n_220),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_317),
.B(n_318),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_236),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_279),
.B(n_220),
.Y(n_320)
);

OAI21xp33_ASAP7_75t_SL g346 ( 
.A1(n_320),
.A2(n_334),
.B(n_336),
.Y(n_346)
);

INVx3_ASAP7_75t_L g321 ( 
.A(n_278),
.Y(n_321)
);

BUFx3_ASAP7_75t_L g323 ( 
.A(n_277),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_323),
.B(n_325),
.Y(n_347)
);

INVx13_ASAP7_75t_L g324 ( 
.A(n_269),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_324),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_271),
.B(n_216),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_SL g326 ( 
.A1(n_262),
.A2(n_192),
.B(n_220),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_283),
.B(n_235),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_327),
.B(n_328),
.Y(n_351)
);

NOR2x1_ASAP7_75t_L g328 ( 
.A(n_262),
.B(n_288),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_287),
.B(n_215),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_SL g341 ( 
.A(n_330),
.B(n_250),
.Y(n_341)
);

INVx13_ASAP7_75t_L g331 ( 
.A(n_280),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_331),
.Y(n_350)
);

INVx13_ASAP7_75t_L g332 ( 
.A(n_280),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_332),
.Y(n_354)
);

INVx4_ASAP7_75t_L g333 ( 
.A(n_239),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_333),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_266),
.B(n_196),
.Y(n_334)
);

INVx13_ASAP7_75t_L g335 ( 
.A(n_277),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_335),
.Y(n_371)
);

AND2x2_ASAP7_75t_L g336 ( 
.A(n_263),
.B(n_180),
.Y(n_336)
);

HB1xp67_ASAP7_75t_L g386 ( 
.A(n_341),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_296),
.A2(n_263),
.B1(n_244),
.B2(n_257),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g392 ( 
.A1(n_342),
.A2(n_343),
.B1(n_344),
.B2(n_369),
.Y(n_392)
);

OAI22xp33_ASAP7_75t_SL g343 ( 
.A1(n_328),
.A2(n_260),
.B1(n_240),
.B2(n_282),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_296),
.A2(n_275),
.B1(n_242),
.B2(n_282),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_293),
.B(n_286),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g404 ( 
.A(n_345),
.B(n_349),
.Y(n_404)
);

MAJx2_ASAP7_75t_L g353 ( 
.A(n_302),
.B(n_281),
.C(n_286),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_353),
.B(n_375),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_307),
.B(n_270),
.C(n_264),
.Y(n_358)
);

XOR2x2_ASAP7_75t_L g412 ( 
.A(n_358),
.B(n_365),
.Y(n_412)
);

AND2x2_ASAP7_75t_L g398 ( 
.A(n_362),
.B(n_346),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_336),
.A2(n_274),
.B1(n_261),
.B2(n_239),
.Y(n_363)
);

OAI21xp5_ASAP7_75t_SL g410 ( 
.A1(n_363),
.A2(n_313),
.B(n_354),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_322),
.B(n_270),
.Y(n_365)
);

INVxp67_ASAP7_75t_L g393 ( 
.A(n_366),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_296),
.A2(n_242),
.B1(n_241),
.B2(n_255),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_312),
.A2(n_255),
.B1(n_241),
.B2(n_245),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_L g411 ( 
.A1(n_370),
.A2(n_301),
.B1(n_314),
.B2(n_289),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_322),
.B(n_258),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_SL g382 ( 
.A(n_372),
.B(n_374),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_304),
.Y(n_374)
);

BUFx24_ASAP7_75t_SL g375 ( 
.A(n_315),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_312),
.A2(n_245),
.B1(n_236),
.B2(n_5),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_376),
.B(n_318),
.Y(n_383)
);

AOI22xp33_ASAP7_75t_SL g380 ( 
.A1(n_379),
.A2(n_329),
.B1(n_336),
.B2(n_308),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_L g417 ( 
.A1(n_380),
.A2(n_383),
.B1(n_394),
.B2(n_409),
.Y(n_417)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_355),
.Y(n_381)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_381),
.Y(n_419)
);

INVx2_ASAP7_75t_SL g385 ( 
.A(n_355),
.Y(n_385)
);

INVx1_ASAP7_75t_SL g444 ( 
.A(n_385),
.Y(n_444)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_378),
.Y(n_387)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_387),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_SL g388 ( 
.A(n_359),
.B(n_364),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_SL g422 ( 
.A(n_388),
.B(n_390),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_347),
.B(n_325),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_389),
.B(n_395),
.Y(n_425)
);

OAI21xp33_ASAP7_75t_SL g390 ( 
.A1(n_348),
.A2(n_351),
.B(n_326),
.Y(n_390)
);

BUFx3_ASAP7_75t_L g391 ( 
.A(n_377),
.Y(n_391)
);

INVx5_ASAP7_75t_L g432 ( 
.A(n_391),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_L g394 ( 
.A1(n_351),
.A2(n_319),
.B1(n_308),
.B2(n_329),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_347),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_352),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_396),
.B(n_400),
.Y(n_428)
);

OAI21xp5_ASAP7_75t_L g397 ( 
.A1(n_362),
.A2(n_303),
.B(n_311),
.Y(n_397)
);

AOI21xp5_ASAP7_75t_SL g443 ( 
.A1(n_397),
.A2(n_403),
.B(n_361),
.Y(n_443)
);

INVxp67_ASAP7_75t_L g441 ( 
.A(n_398),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_SL g399 ( 
.A(n_345),
.B(n_330),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_SL g433 ( 
.A(n_399),
.B(n_401),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_340),
.B(n_327),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_365),
.B(n_323),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_372),
.B(n_309),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_402),
.B(n_413),
.Y(n_418)
);

OAI21xp5_ASAP7_75t_L g403 ( 
.A1(n_356),
.A2(n_368),
.B(n_340),
.Y(n_403)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_361),
.Y(n_405)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_405),
.Y(n_424)
);

AND2x6_ASAP7_75t_L g406 ( 
.A(n_356),
.B(n_316),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_406),
.B(n_407),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_350),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_378),
.Y(n_408)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_408),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_L g409 ( 
.A1(n_363),
.A2(n_366),
.B1(n_319),
.B2(n_370),
.Y(n_409)
);

AOI21xp5_ASAP7_75t_L g429 ( 
.A1(n_410),
.A2(n_344),
.B(n_369),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_411),
.B(n_415),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_339),
.B(n_333),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_337),
.Y(n_414)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_414),
.Y(n_430)
);

AND2x6_ASAP7_75t_L g415 ( 
.A(n_353),
.B(n_292),
.Y(n_415)
);

INVx5_ASAP7_75t_SL g416 ( 
.A(n_379),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_416),
.B(n_367),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_SL g421 ( 
.A(n_404),
.B(n_349),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_SL g476 ( 
.A(n_421),
.B(n_439),
.Y(n_476)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_423),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_393),
.B(n_358),
.C(n_292),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_426),
.B(n_450),
.C(n_414),
.Y(n_469)
);

AND2x2_ASAP7_75t_L g451 ( 
.A(n_429),
.B(n_443),
.Y(n_451)
);

NOR2x1_ASAP7_75t_R g434 ( 
.A(n_397),
.B(n_342),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_434),
.B(n_442),
.Y(n_464)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_385),
.Y(n_435)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_435),
.Y(n_459)
);

XOR2xp5_ASAP7_75t_L g436 ( 
.A(n_404),
.B(n_368),
.Y(n_436)
);

XOR2xp5_ASAP7_75t_L g452 ( 
.A(n_436),
.B(n_445),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_392),
.A2(n_308),
.B1(n_341),
.B2(n_368),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_L g457 ( 
.A1(n_438),
.A2(n_409),
.B1(n_398),
.B2(n_392),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_SL g439 ( 
.A(n_384),
.B(n_300),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_394),
.A2(n_376),
.B1(n_360),
.B2(n_337),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_SL g460 ( 
.A1(n_440),
.A2(n_395),
.B1(n_383),
.B2(n_382),
.Y(n_460)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_385),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_L g445 ( 
.A(n_412),
.B(n_373),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_381),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_446),
.B(n_449),
.Y(n_471)
);

XOR2xp5_ASAP7_75t_L g447 ( 
.A(n_412),
.B(n_373),
.Y(n_447)
);

XOR2xp5_ASAP7_75t_L g453 ( 
.A(n_447),
.B(n_448),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_393),
.B(n_338),
.Y(n_448)
);

CKINVDCx16_ASAP7_75t_R g449 ( 
.A(n_403),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_386),
.B(n_338),
.C(n_357),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_L g454 ( 
.A(n_447),
.B(n_398),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_L g482 ( 
.A(n_454),
.B(n_461),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_433),
.B(n_396),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_SL g489 ( 
.A(n_455),
.B(n_472),
.Y(n_489)
);

OAI22xp5_ASAP7_75t_L g481 ( 
.A1(n_457),
.A2(n_463),
.B1(n_429),
.B2(n_437),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_SL g458 ( 
.A(n_422),
.B(n_388),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g499 ( 
.A(n_458),
.B(n_462),
.Y(n_499)
);

AOI22xp5_ASAP7_75t_L g480 ( 
.A1(n_460),
.A2(n_440),
.B1(n_441),
.B2(n_437),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_421),
.B(n_415),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_425),
.Y(n_462)
);

AOI22xp5_ASAP7_75t_L g463 ( 
.A1(n_417),
.A2(n_389),
.B1(n_400),
.B2(n_406),
.Y(n_463)
);

XOR2xp5_ASAP7_75t_L g465 ( 
.A(n_445),
.B(n_436),
.Y(n_465)
);

XOR2xp5_ASAP7_75t_L g483 ( 
.A(n_465),
.B(n_466),
.Y(n_483)
);

XOR2xp5_ASAP7_75t_L g466 ( 
.A(n_439),
.B(n_410),
.Y(n_466)
);

XNOR2xp5_ASAP7_75t_L g467 ( 
.A(n_426),
.B(n_450),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_L g487 ( 
.A(n_467),
.B(n_468),
.Y(n_487)
);

XNOR2xp5_ASAP7_75t_L g468 ( 
.A(n_448),
.B(n_387),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_L g493 ( 
.A(n_469),
.B(n_473),
.Y(n_493)
);

OAI21xp5_ASAP7_75t_SL g470 ( 
.A1(n_431),
.A2(n_407),
.B(n_377),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_470),
.B(n_419),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_418),
.B(n_371),
.Y(n_472)
);

XNOR2xp5_ASAP7_75t_L g473 ( 
.A(n_428),
.B(n_408),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_SL g474 ( 
.A(n_431),
.B(n_357),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_SL g495 ( 
.A(n_474),
.B(n_477),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_441),
.B(n_295),
.C(n_306),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_475),
.B(n_391),
.C(n_405),
.Y(n_494)
);

CKINVDCx20_ASAP7_75t_R g477 ( 
.A(n_425),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_428),
.B(n_432),
.Y(n_478)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_478),
.Y(n_496)
);

XNOR2xp5_ASAP7_75t_L g479 ( 
.A(n_438),
.B(n_291),
.Y(n_479)
);

XOR2xp5_ASAP7_75t_L g485 ( 
.A(n_479),
.B(n_443),
.Y(n_485)
);

OAI22xp5_ASAP7_75t_SL g520 ( 
.A1(n_480),
.A2(n_488),
.B1(n_297),
.B2(n_298),
.Y(n_520)
);

AOI22xp5_ASAP7_75t_L g522 ( 
.A1(n_481),
.A2(n_297),
.B1(n_4),
.B2(n_5),
.Y(n_522)
);

AOI22xp5_ASAP7_75t_L g484 ( 
.A1(n_456),
.A2(n_430),
.B1(n_420),
.B2(n_427),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_SL g506 ( 
.A(n_484),
.B(n_486),
.Y(n_506)
);

XOR2xp5_ASAP7_75t_L g508 ( 
.A(n_485),
.B(n_500),
.Y(n_508)
);

BUFx2_ASAP7_75t_L g486 ( 
.A(n_459),
.Y(n_486)
);

CKINVDCx20_ASAP7_75t_R g521 ( 
.A(n_486),
.Y(n_521)
);

AOI22xp5_ASAP7_75t_L g488 ( 
.A1(n_463),
.A2(n_434),
.B1(n_444),
.B2(n_416),
.Y(n_488)
);

OAI21xp5_ASAP7_75t_SL g516 ( 
.A1(n_490),
.A2(n_498),
.B(n_324),
.Y(n_516)
);

OAI22xp5_ASAP7_75t_L g491 ( 
.A1(n_457),
.A2(n_444),
.B1(n_424),
.B2(n_432),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_491),
.B(n_451),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_469),
.B(n_467),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_492),
.B(n_503),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g509 ( 
.A(n_494),
.B(n_497),
.C(n_502),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_452),
.B(n_465),
.C(n_453),
.Y(n_497)
);

OAI21xp5_ASAP7_75t_L g498 ( 
.A1(n_464),
.A2(n_321),
.B(n_290),
.Y(n_498)
);

XOR2xp5_ASAP7_75t_L g500 ( 
.A(n_452),
.B(n_332),
.Y(n_500)
);

INVxp67_ASAP7_75t_L g501 ( 
.A(n_475),
.Y(n_501)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_501),
.Y(n_507)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_453),
.B(n_335),
.C(n_331),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_471),
.B(n_297),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_473),
.Y(n_504)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_504),
.Y(n_511)
);

INVxp67_ASAP7_75t_L g524 ( 
.A(n_505),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_506),
.B(n_512),
.Y(n_529)
);

AOI22xp5_ASAP7_75t_SL g510 ( 
.A1(n_495),
.A2(n_451),
.B1(n_466),
.B2(n_461),
.Y(n_510)
);

OAI22xp5_ASAP7_75t_SL g533 ( 
.A1(n_510),
.A2(n_522),
.B1(n_523),
.B2(n_483),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_499),
.B(n_468),
.Y(n_512)
);

NOR2x1_ASAP7_75t_L g513 ( 
.A(n_488),
.B(n_485),
.Y(n_513)
);

AOI21xp5_ASAP7_75t_L g525 ( 
.A1(n_513),
.A2(n_514),
.B(n_517),
.Y(n_525)
);

AOI21xp5_ASAP7_75t_L g514 ( 
.A1(n_498),
.A2(n_479),
.B(n_454),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_496),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_515),
.B(n_516),
.Y(n_527)
);

AOI21xp5_ASAP7_75t_L g517 ( 
.A1(n_501),
.A2(n_476),
.B(n_305),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_493),
.B(n_476),
.Y(n_519)
);

XNOR2xp5_ASAP7_75t_L g532 ( 
.A(n_519),
.B(n_483),
.Y(n_532)
);

AOI22xp5_ASAP7_75t_L g530 ( 
.A1(n_520),
.A2(n_502),
.B1(n_500),
.B2(n_482),
.Y(n_530)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_494),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_523),
.B(n_493),
.C(n_487),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_526),
.B(n_533),
.Y(n_544)
);

XOR2xp5_ASAP7_75t_L g528 ( 
.A(n_509),
.B(n_482),
.Y(n_528)
);

XOR2xp5_ASAP7_75t_L g547 ( 
.A(n_528),
.B(n_532),
.Y(n_547)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_530),
.Y(n_542)
);

OAI21xp5_ASAP7_75t_SL g531 ( 
.A1(n_518),
.A2(n_487),
.B(n_497),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_SL g546 ( 
.A(n_531),
.B(n_534),
.Y(n_546)
);

OAI22xp5_ASAP7_75t_SL g534 ( 
.A1(n_515),
.A2(n_489),
.B1(n_4),
.B2(n_5),
.Y(n_534)
);

OAI22x1_ASAP7_75t_L g535 ( 
.A1(n_505),
.A2(n_1),
.B1(n_5),
.B2(n_6),
.Y(n_535)
);

AOI21xp5_ASAP7_75t_L g543 ( 
.A1(n_535),
.A2(n_539),
.B(n_521),
.Y(n_543)
);

XNOR2xp5_ASAP7_75t_L g536 ( 
.A(n_509),
.B(n_7),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_SL g548 ( 
.A(n_536),
.B(n_537),
.Y(n_548)
);

MAJIxp5_ASAP7_75t_L g537 ( 
.A(n_507),
.B(n_7),
.C(n_8),
.Y(n_537)
);

XOR2xp5_ASAP7_75t_L g538 ( 
.A(n_517),
.B(n_10),
.Y(n_538)
);

OAI21x1_ASAP7_75t_L g552 ( 
.A1(n_538),
.A2(n_514),
.B(n_513),
.Y(n_552)
);

OAI21xp5_ASAP7_75t_SL g539 ( 
.A1(n_518),
.A2(n_10),
.B(n_11),
.Y(n_539)
);

XNOR2xp5_ASAP7_75t_L g540 ( 
.A(n_507),
.B(n_512),
.Y(n_540)
);

MAJIxp5_ASAP7_75t_L g541 ( 
.A(n_540),
.B(n_516),
.C(n_511),
.Y(n_541)
);

XNOR2xp5_ASAP7_75t_L g555 ( 
.A(n_541),
.B(n_553),
.Y(n_555)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_543),
.Y(n_562)
);

O2A1O1Ixp33_ASAP7_75t_SL g545 ( 
.A1(n_527),
.A2(n_511),
.B(n_513),
.C(n_510),
.Y(n_545)
);

INVxp33_ASAP7_75t_L g558 ( 
.A(n_545),
.Y(n_558)
);

OAI22xp5_ASAP7_75t_L g549 ( 
.A1(n_524),
.A2(n_522),
.B1(n_521),
.B2(n_506),
.Y(n_549)
);

AOI22xp5_ASAP7_75t_L g556 ( 
.A1(n_549),
.A2(n_551),
.B1(n_535),
.B2(n_525),
.Y(n_556)
);

CKINVDCx16_ASAP7_75t_R g550 ( 
.A(n_529),
.Y(n_550)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_550),
.Y(n_557)
);

INVx3_ASAP7_75t_L g551 ( 
.A(n_524),
.Y(n_551)
);

OAI21x1_ASAP7_75t_L g559 ( 
.A1(n_552),
.A2(n_530),
.B(n_508),
.Y(n_559)
);

MAJIxp5_ASAP7_75t_L g553 ( 
.A(n_526),
.B(n_508),
.C(n_520),
.Y(n_553)
);

MAJIxp5_ASAP7_75t_L g554 ( 
.A(n_547),
.B(n_528),
.C(n_540),
.Y(n_554)
);

MAJIxp5_ASAP7_75t_L g565 ( 
.A(n_554),
.B(n_553),
.C(n_541),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_556),
.Y(n_566)
);

AOI21xp5_ASAP7_75t_L g567 ( 
.A1(n_559),
.A2(n_560),
.B(n_561),
.Y(n_567)
);

OAI21xp5_ASAP7_75t_SL g560 ( 
.A1(n_544),
.A2(n_519),
.B(n_532),
.Y(n_560)
);

MAJIxp5_ASAP7_75t_L g561 ( 
.A(n_547),
.B(n_536),
.C(n_537),
.Y(n_561)
);

NOR2xp33_ASAP7_75t_L g563 ( 
.A(n_555),
.B(n_546),
.Y(n_563)
);

AOI21xp5_ASAP7_75t_L g570 ( 
.A1(n_563),
.A2(n_558),
.B(n_548),
.Y(n_570)
);

OAI22xp5_ASAP7_75t_L g564 ( 
.A1(n_562),
.A2(n_542),
.B1(n_551),
.B2(n_543),
.Y(n_564)
);

AOI21xp33_ASAP7_75t_L g569 ( 
.A1(n_564),
.A2(n_557),
.B(n_558),
.Y(n_569)
);

XNOR2xp5_ASAP7_75t_L g568 ( 
.A(n_565),
.B(n_554),
.Y(n_568)
);

MAJIxp5_ASAP7_75t_L g571 ( 
.A(n_568),
.B(n_570),
.C(n_565),
.Y(n_571)
);

AOI322xp5_ASAP7_75t_L g572 ( 
.A1(n_569),
.A2(n_566),
.A3(n_567),
.B1(n_545),
.B2(n_538),
.C1(n_14),
.C2(n_12),
.Y(n_572)
);

OAI21xp5_ASAP7_75t_L g573 ( 
.A1(n_571),
.A2(n_572),
.B(n_10),
.Y(n_573)
);

MAJIxp5_ASAP7_75t_L g574 ( 
.A(n_573),
.B(n_14),
.C(n_11),
.Y(n_574)
);

OAI21xp5_ASAP7_75t_SL g575 ( 
.A1(n_574),
.A2(n_11),
.B(n_12),
.Y(n_575)
);

XNOR2xp5_ASAP7_75t_L g576 ( 
.A(n_575),
.B(n_11),
.Y(n_576)
);

FAx1_ASAP7_75t_SL g577 ( 
.A(n_576),
.B(n_14),
.CI(n_211),
.CON(n_577),
.SN(n_577)
);


endmodule