module real_aes_6812_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_704, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_704;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_357;
wire n_287;
wire n_635;
wire n_503;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_417;
wire n_182;
wire n_363;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_527;
wire n_502;
wire n_600;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_404;
wire n_147;
wire n_288;
wire n_598;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_481;
wire n_148;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_637;
wire n_526;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_105;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g155 ( .A1(n_0), .A2(n_156), .B(n_157), .C(n_161), .Y(n_155) );
CKINVDCx20_ASAP7_75t_R g687 ( .A(n_1), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_2), .B(n_150), .Y(n_163) );
INVx1_ASAP7_75t_L g406 ( .A(n_3), .Y(n_406) );
NAND2xp5_ASAP7_75t_SL g134 ( .A(n_4), .B(n_135), .Y(n_134) );
A2O1A1Ixp33_ASAP7_75t_L g448 ( .A1(n_5), .A2(n_124), .B(n_141), .C(n_449), .Y(n_448) );
AOI21xp5_ASAP7_75t_L g469 ( .A1(n_6), .A2(n_144), .B(n_470), .Y(n_469) );
AOI21xp5_ASAP7_75t_L g245 ( .A1(n_7), .A2(n_144), .B(n_246), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_8), .B(n_150), .Y(n_476) );
AO21x2_ASAP7_75t_L g202 ( .A1(n_9), .A2(n_116), .B(n_203), .Y(n_202) );
AND2x6_ASAP7_75t_L g141 ( .A(n_10), .B(n_142), .Y(n_141) );
A2O1A1Ixp33_ASAP7_75t_L g220 ( .A1(n_11), .A2(n_124), .B(n_141), .C(n_221), .Y(n_220) );
INVx1_ASAP7_75t_L g441 ( .A(n_12), .Y(n_441) );
NOR2xp33_ASAP7_75t_L g407 ( .A(n_13), .B(n_40), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_13), .B(n_40), .Y(n_695) );
NAND2xp5_ASAP7_75t_SL g451 ( .A(n_14), .B(n_160), .Y(n_451) );
INVx1_ASAP7_75t_L g121 ( .A(n_15), .Y(n_121) );
NAND2xp5_ASAP7_75t_SL g209 ( .A(n_16), .B(n_135), .Y(n_209) );
A2O1A1Ixp33_ASAP7_75t_L g459 ( .A1(n_17), .A2(n_136), .B(n_460), .C(n_462), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_18), .B(n_150), .Y(n_463) );
OAI22xp5_ASAP7_75t_SL g106 ( .A1(n_19), .A2(n_107), .B1(n_108), .B2(n_400), .Y(n_106) );
CKINVDCx20_ASAP7_75t_R g400 ( .A(n_19), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_20), .B(n_193), .Y(n_510) );
A2O1A1Ixp33_ASAP7_75t_L g186 ( .A1(n_21), .A2(n_124), .B(n_187), .C(n_192), .Y(n_186) );
A2O1A1Ixp33_ASAP7_75t_L g430 ( .A1(n_22), .A2(n_159), .B(n_211), .C(n_431), .Y(n_430) );
NAND2xp5_ASAP7_75t_SL g483 ( .A(n_23), .B(n_160), .Y(n_483) );
NAND2xp5_ASAP7_75t_SL g492 ( .A(n_24), .B(n_160), .Y(n_492) );
CKINVDCx16_ASAP7_75t_R g479 ( .A(n_25), .Y(n_479) );
INVx1_ASAP7_75t_L g491 ( .A(n_26), .Y(n_491) );
A2O1A1Ixp33_ASAP7_75t_L g205 ( .A1(n_27), .A2(n_124), .B(n_192), .C(n_206), .Y(n_205) );
BUFx6f_ASAP7_75t_L g128 ( .A(n_28), .Y(n_128) );
CKINVDCx20_ASAP7_75t_R g447 ( .A(n_29), .Y(n_447) );
INVx1_ASAP7_75t_L g508 ( .A(n_30), .Y(n_508) );
AOI21xp5_ASAP7_75t_L g151 ( .A1(n_31), .A2(n_144), .B(n_152), .Y(n_151) );
INVx2_ASAP7_75t_L g126 ( .A(n_32), .Y(n_126) );
A2O1A1Ixp33_ASAP7_75t_L g170 ( .A1(n_33), .A2(n_139), .B(n_171), .C(n_172), .Y(n_170) );
CKINVDCx20_ASAP7_75t_R g454 ( .A(n_34), .Y(n_454) );
A2O1A1Ixp33_ASAP7_75t_L g472 ( .A1(n_35), .A2(n_159), .B(n_473), .C(n_475), .Y(n_472) );
INVxp67_ASAP7_75t_L g509 ( .A(n_36), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_37), .B(n_208), .Y(n_207) );
CKINVDCx14_ASAP7_75t_R g471 ( .A(n_38), .Y(n_471) );
A2O1A1Ixp33_ASAP7_75t_L g489 ( .A1(n_39), .A2(n_124), .B(n_192), .C(n_490), .Y(n_489) );
A2O1A1Ixp33_ASAP7_75t_L g438 ( .A1(n_41), .A2(n_161), .B(n_439), .C(n_440), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_42), .B(n_185), .Y(n_184) );
CKINVDCx20_ASAP7_75t_R g225 ( .A(n_43), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_44), .B(n_135), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_45), .B(n_144), .Y(n_204) );
CKINVDCx20_ASAP7_75t_R g494 ( .A(n_46), .Y(n_494) );
CKINVDCx20_ASAP7_75t_R g505 ( .A(n_47), .Y(n_505) );
A2O1A1Ixp33_ASAP7_75t_L g231 ( .A1(n_48), .A2(n_139), .B(n_171), .C(n_232), .Y(n_231) );
CKINVDCx20_ASAP7_75t_R g409 ( .A(n_49), .Y(n_409) );
INVx1_ASAP7_75t_L g158 ( .A(n_50), .Y(n_158) );
OAI222xp33_ASAP7_75t_L g413 ( .A1(n_51), .A2(n_414), .B1(n_681), .B2(n_684), .C1(n_685), .C2(n_687), .Y(n_413) );
CKINVDCx20_ASAP7_75t_R g684 ( .A(n_51), .Y(n_684) );
INVx1_ASAP7_75t_L g233 ( .A(n_52), .Y(n_233) );
INVx1_ASAP7_75t_L g429 ( .A(n_53), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_54), .B(n_144), .Y(n_230) );
CKINVDCx20_ASAP7_75t_R g196 ( .A(n_55), .Y(n_196) );
CKINVDCx14_ASAP7_75t_R g437 ( .A(n_56), .Y(n_437) );
INVx1_ASAP7_75t_L g142 ( .A(n_57), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_58), .B(n_144), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_59), .B(n_150), .Y(n_251) );
A2O1A1Ixp33_ASAP7_75t_L g248 ( .A1(n_60), .A2(n_131), .B(n_191), .C(n_249), .Y(n_248) );
INVx1_ASAP7_75t_L g120 ( .A(n_61), .Y(n_120) );
INVx1_ASAP7_75t_SL g474 ( .A(n_62), .Y(n_474) );
CKINVDCx20_ASAP7_75t_R g104 ( .A(n_63), .Y(n_104) );
NAND2xp5_ASAP7_75t_SL g176 ( .A(n_64), .B(n_135), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_65), .B(n_150), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_66), .B(n_136), .Y(n_222) );
INVx1_ASAP7_75t_L g482 ( .A(n_67), .Y(n_482) );
CKINVDCx16_ASAP7_75t_R g153 ( .A(n_68), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_69), .B(n_175), .Y(n_188) );
A2O1A1Ixp33_ASAP7_75t_L g123 ( .A1(n_70), .A2(n_124), .B(n_129), .C(n_139), .Y(n_123) );
CKINVDCx16_ASAP7_75t_R g247 ( .A(n_71), .Y(n_247) );
INVx1_ASAP7_75t_L g700 ( .A(n_72), .Y(n_700) );
AOI21xp5_ASAP7_75t_L g435 ( .A1(n_73), .A2(n_144), .B(n_436), .Y(n_435) );
CKINVDCx20_ASAP7_75t_R g485 ( .A(n_74), .Y(n_485) );
AOI21xp5_ASAP7_75t_L g456 ( .A1(n_75), .A2(n_144), .B(n_457), .Y(n_456) );
AOI21xp5_ASAP7_75t_L g503 ( .A1(n_76), .A2(n_185), .B(n_504), .Y(n_503) );
INVx1_ASAP7_75t_L g458 ( .A(n_77), .Y(n_458) );
CKINVDCx16_ASAP7_75t_R g488 ( .A(n_78), .Y(n_488) );
NAND2xp5_ASAP7_75t_SL g189 ( .A(n_79), .B(n_174), .Y(n_189) );
CKINVDCx20_ASAP7_75t_R g180 ( .A(n_80), .Y(n_180) );
AOI21xp5_ASAP7_75t_L g427 ( .A1(n_81), .A2(n_144), .B(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g461 ( .A(n_82), .Y(n_461) );
INVx2_ASAP7_75t_L g118 ( .A(n_83), .Y(n_118) );
INVx1_ASAP7_75t_L g450 ( .A(n_84), .Y(n_450) );
CKINVDCx20_ASAP7_75t_R g148 ( .A(n_85), .Y(n_148) );
NAND2xp5_ASAP7_75t_SL g223 ( .A(n_86), .B(n_160), .Y(n_223) );
OR2x2_ASAP7_75t_L g403 ( .A(n_87), .B(n_404), .Y(n_403) );
OR2x2_ASAP7_75t_L g416 ( .A(n_87), .B(n_405), .Y(n_416) );
INVx2_ASAP7_75t_L g419 ( .A(n_87), .Y(n_419) );
A2O1A1Ixp33_ASAP7_75t_L g480 ( .A1(n_88), .A2(n_124), .B(n_139), .C(n_481), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_89), .B(n_144), .Y(n_169) );
INVx1_ASAP7_75t_L g173 ( .A(n_90), .Y(n_173) );
AOI22xp33_ASAP7_75t_SL g99 ( .A1(n_91), .A2(n_100), .B1(n_690), .B2(n_701), .Y(n_99) );
INVxp67_ASAP7_75t_L g250 ( .A(n_92), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_93), .B(n_116), .Y(n_442) );
INVx1_ASAP7_75t_L g130 ( .A(n_94), .Y(n_130) );
INVx1_ASAP7_75t_L g218 ( .A(n_95), .Y(n_218) );
INVx2_ASAP7_75t_L g432 ( .A(n_96), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_97), .B(n_700), .Y(n_699) );
AND2x2_ASAP7_75t_L g235 ( .A(n_98), .B(n_178), .Y(n_235) );
OAI21xp5_ASAP7_75t_L g100 ( .A1(n_101), .A2(n_105), .B(n_412), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
INVx1_ASAP7_75t_SL g102 ( .A(n_103), .Y(n_102) );
BUFx2_ASAP7_75t_L g689 ( .A(n_103), .Y(n_689) );
INVx2_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
AOI21xp5_ASAP7_75t_L g105 ( .A1(n_106), .A2(n_401), .B(n_408), .Y(n_105) );
INVx1_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
AOI22xp5_ASAP7_75t_L g681 ( .A1(n_108), .A2(n_415), .B1(n_682), .B2(n_683), .Y(n_681) );
INVx2_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
AOI22xp5_ASAP7_75t_L g414 ( .A1(n_109), .A2(n_415), .B1(n_417), .B2(n_420), .Y(n_414) );
NAND2x1p5_ASAP7_75t_L g109 ( .A(n_110), .B(n_343), .Y(n_109) );
AND4x1_ASAP7_75t_L g110 ( .A(n_111), .B(n_283), .C(n_298), .D(n_323), .Y(n_110) );
NOR2xp33_ASAP7_75t_SL g111 ( .A(n_112), .B(n_256), .Y(n_111) );
OAI21xp33_ASAP7_75t_L g112 ( .A1(n_113), .A2(n_164), .B(n_236), .Y(n_112) );
AND2x2_ASAP7_75t_L g286 ( .A(n_113), .B(n_182), .Y(n_286) );
AND2x2_ASAP7_75t_L g299 ( .A(n_113), .B(n_181), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_113), .B(n_165), .Y(n_349) );
INVx1_ASAP7_75t_L g353 ( .A(n_113), .Y(n_353) );
AND2x2_ASAP7_75t_L g113 ( .A(n_114), .B(n_149), .Y(n_113) );
INVx2_ASAP7_75t_L g270 ( .A(n_114), .Y(n_270) );
BUFx2_ASAP7_75t_L g297 ( .A(n_114), .Y(n_297) );
AO21x2_ASAP7_75t_L g114 ( .A1(n_115), .A2(n_122), .B(n_147), .Y(n_114) );
NOR2xp33_ASAP7_75t_L g147 ( .A(n_115), .B(n_148), .Y(n_147) );
INVx3_ASAP7_75t_L g150 ( .A(n_115), .Y(n_150) );
NOR2xp33_ASAP7_75t_L g179 ( .A(n_115), .B(n_180), .Y(n_179) );
AO21x2_ASAP7_75t_L g216 ( .A1(n_115), .A2(n_217), .B(n_224), .Y(n_216) );
NOR2xp33_ASAP7_75t_L g453 ( .A(n_115), .B(n_454), .Y(n_453) );
AO21x2_ASAP7_75t_L g477 ( .A1(n_115), .A2(n_478), .B(n_484), .Y(n_477) );
NOR2xp33_ASAP7_75t_L g493 ( .A(n_115), .B(n_494), .Y(n_493) );
INVx4_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
AOI21xp5_ASAP7_75t_L g203 ( .A1(n_116), .A2(n_204), .B(n_205), .Y(n_203) );
HB1xp67_ASAP7_75t_L g244 ( .A(n_116), .Y(n_244) );
BUFx6f_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
INVx1_ASAP7_75t_L g226 ( .A(n_117), .Y(n_226) );
AND2x2_ASAP7_75t_L g117 ( .A(n_118), .B(n_119), .Y(n_117) );
AND2x2_ASAP7_75t_SL g178 ( .A(n_118), .B(n_119), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g119 ( .A(n_120), .B(n_121), .Y(n_119) );
NAND2xp5_ASAP7_75t_L g122 ( .A(n_123), .B(n_143), .Y(n_122) );
INVx5_ASAP7_75t_L g154 ( .A(n_124), .Y(n_154) );
AND2x6_ASAP7_75t_L g124 ( .A(n_125), .B(n_127), .Y(n_124) );
BUFx6f_ASAP7_75t_L g138 ( .A(n_125), .Y(n_138) );
BUFx3_ASAP7_75t_L g162 ( .A(n_125), .Y(n_162) );
INVx2_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
INVx1_ASAP7_75t_L g146 ( .A(n_126), .Y(n_146) );
INVx1_ASAP7_75t_L g212 ( .A(n_126), .Y(n_212) );
INVx1_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
BUFx6f_ASAP7_75t_L g133 ( .A(n_128), .Y(n_133) );
INVx3_ASAP7_75t_L g136 ( .A(n_128), .Y(n_136) );
AND2x2_ASAP7_75t_L g145 ( .A(n_128), .B(n_146), .Y(n_145) );
BUFx6f_ASAP7_75t_L g160 ( .A(n_128), .Y(n_160) );
INVx1_ASAP7_75t_L g208 ( .A(n_128), .Y(n_208) );
O2A1O1Ixp33_ASAP7_75t_L g129 ( .A1(n_130), .A2(n_131), .B(n_134), .C(n_137), .Y(n_129) );
INVx1_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
NOR2xp33_ASAP7_75t_L g431 ( .A(n_132), .B(n_432), .Y(n_431) );
NOR2xp33_ASAP7_75t_L g460 ( .A(n_132), .B(n_461), .Y(n_460) );
OAI22xp33_ASAP7_75t_L g507 ( .A1(n_132), .A2(n_135), .B1(n_508), .B2(n_509), .Y(n_507) );
INVx4_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
INVx2_ASAP7_75t_L g175 ( .A(n_133), .Y(n_175) );
INVx2_ASAP7_75t_L g156 ( .A(n_135), .Y(n_156) );
NOR2xp33_ASAP7_75t_L g249 ( .A(n_135), .B(n_250), .Y(n_249) );
O2A1O1Ixp33_ASAP7_75t_L g490 ( .A1(n_135), .A2(n_190), .B(n_491), .C(n_492), .Y(n_490) );
INVx5_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
NOR2xp33_ASAP7_75t_L g440 ( .A(n_136), .B(n_441), .Y(n_440) );
HB1xp67_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
INVx3_ASAP7_75t_L g475 ( .A(n_138), .Y(n_475) );
INVx1_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
O2A1O1Ixp33_ASAP7_75t_SL g152 ( .A1(n_140), .A2(n_153), .B(n_154), .C(n_155), .Y(n_152) );
O2A1O1Ixp33_ASAP7_75t_L g246 ( .A1(n_140), .A2(n_154), .B(n_247), .C(n_248), .Y(n_246) );
O2A1O1Ixp33_ASAP7_75t_SL g428 ( .A1(n_140), .A2(n_154), .B(n_429), .C(n_430), .Y(n_428) );
O2A1O1Ixp33_ASAP7_75t_SL g436 ( .A1(n_140), .A2(n_154), .B(n_437), .C(n_438), .Y(n_436) );
O2A1O1Ixp33_ASAP7_75t_SL g457 ( .A1(n_140), .A2(n_154), .B(n_458), .C(n_459), .Y(n_457) );
O2A1O1Ixp33_ASAP7_75t_L g470 ( .A1(n_140), .A2(n_154), .B(n_471), .C(n_472), .Y(n_470) );
O2A1O1Ixp33_ASAP7_75t_SL g504 ( .A1(n_140), .A2(n_154), .B(n_505), .C(n_506), .Y(n_504) );
INVx4_ASAP7_75t_SL g140 ( .A(n_141), .Y(n_140) );
AND2x4_ASAP7_75t_L g144 ( .A(n_141), .B(n_145), .Y(n_144) );
BUFx3_ASAP7_75t_L g192 ( .A(n_141), .Y(n_192) );
NAND2x1p5_ASAP7_75t_L g219 ( .A(n_141), .B(n_145), .Y(n_219) );
BUFx2_ASAP7_75t_L g185 ( .A(n_144), .Y(n_185) );
INVx1_ASAP7_75t_L g191 ( .A(n_146), .Y(n_191) );
AND2x2_ASAP7_75t_L g237 ( .A(n_149), .B(n_182), .Y(n_237) );
INVx2_ASAP7_75t_L g253 ( .A(n_149), .Y(n_253) );
AND2x2_ASAP7_75t_L g262 ( .A(n_149), .B(n_181), .Y(n_262) );
AND2x2_ASAP7_75t_L g341 ( .A(n_149), .B(n_270), .Y(n_341) );
OA21x2_ASAP7_75t_L g149 ( .A1(n_150), .A2(n_151), .B(n_163), .Y(n_149) );
INVx2_ASAP7_75t_L g171 ( .A(n_154), .Y(n_171) );
NOR2xp33_ASAP7_75t_L g157 ( .A(n_158), .B(n_159), .Y(n_157) );
NOR2xp33_ASAP7_75t_L g473 ( .A(n_159), .B(n_474), .Y(n_473) );
INVx4_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
INVx2_ASAP7_75t_L g439 ( .A(n_160), .Y(n_439) );
INVx2_ASAP7_75t_L g452 ( .A(n_161), .Y(n_452) );
INVx2_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
HB1xp67_ASAP7_75t_L g177 ( .A(n_162), .Y(n_177) );
INVx1_ASAP7_75t_L g462 ( .A(n_162), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_165), .B(n_198), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_165), .B(n_268), .Y(n_306) );
INVx1_ASAP7_75t_L g394 ( .A(n_165), .Y(n_394) );
AND2x2_ASAP7_75t_L g165 ( .A(n_166), .B(n_181), .Y(n_165) );
AND2x2_ASAP7_75t_L g252 ( .A(n_166), .B(n_253), .Y(n_252) );
OR2x2_ASAP7_75t_L g266 ( .A(n_166), .B(n_267), .Y(n_266) );
HB1xp67_ASAP7_75t_L g295 ( .A(n_166), .Y(n_295) );
OR2x2_ASAP7_75t_L g327 ( .A(n_166), .B(n_269), .Y(n_327) );
AND2x2_ASAP7_75t_L g335 ( .A(n_166), .B(n_336), .Y(n_335) );
AND2x2_ASAP7_75t_L g368 ( .A(n_166), .B(n_337), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_166), .B(n_237), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_166), .B(n_297), .Y(n_393) );
AND2x2_ASAP7_75t_L g399 ( .A(n_166), .B(n_286), .Y(n_399) );
INVx5_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
BUFx2_ASAP7_75t_L g259 ( .A(n_167), .Y(n_259) );
AND2x2_ASAP7_75t_L g289 ( .A(n_167), .B(n_269), .Y(n_289) );
AND2x2_ASAP7_75t_L g322 ( .A(n_167), .B(n_282), .Y(n_322) );
AND2x2_ASAP7_75t_L g342 ( .A(n_167), .B(n_182), .Y(n_342) );
AND2x2_ASAP7_75t_L g376 ( .A(n_167), .B(n_242), .Y(n_376) );
OR2x6_ASAP7_75t_L g167 ( .A(n_168), .B(n_179), .Y(n_167) );
AOI21xp5_ASAP7_75t_L g168 ( .A1(n_169), .A2(n_170), .B(n_178), .Y(n_168) );
O2A1O1Ixp33_ASAP7_75t_L g172 ( .A1(n_173), .A2(n_174), .B(n_176), .C(n_177), .Y(n_172) );
O2A1O1Ixp33_ASAP7_75t_L g232 ( .A1(n_174), .A2(n_177), .B(n_233), .C(n_234), .Y(n_232) );
O2A1O1Ixp5_ASAP7_75t_L g449 ( .A1(n_174), .A2(n_450), .B(n_451), .C(n_452), .Y(n_449) );
O2A1O1Ixp33_ASAP7_75t_L g481 ( .A1(n_174), .A2(n_452), .B(n_482), .C(n_483), .Y(n_481) );
INVx2_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
INVx2_ASAP7_75t_L g194 ( .A(n_178), .Y(n_194) );
INVx1_ASAP7_75t_L g197 ( .A(n_178), .Y(n_197) );
AOI21xp5_ASAP7_75t_L g229 ( .A1(n_178), .A2(n_230), .B(n_231), .Y(n_229) );
OA21x2_ASAP7_75t_L g434 ( .A1(n_178), .A2(n_435), .B(n_442), .Y(n_434) );
O2A1O1Ixp33_ASAP7_75t_L g487 ( .A1(n_178), .A2(n_219), .B(n_488), .C(n_489), .Y(n_487) );
AND2x4_ASAP7_75t_L g282 ( .A(n_181), .B(n_253), .Y(n_282) );
AND2x2_ASAP7_75t_L g293 ( .A(n_181), .B(n_289), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_181), .B(n_269), .Y(n_332) );
INVx2_ASAP7_75t_L g347 ( .A(n_181), .Y(n_347) );
NOR2xp33_ASAP7_75t_L g370 ( .A(n_181), .B(n_281), .Y(n_370) );
AND2x2_ASAP7_75t_L g389 ( .A(n_181), .B(n_341), .Y(n_389) );
INVx5_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
HB1xp67_ASAP7_75t_L g288 ( .A(n_182), .Y(n_288) );
AND2x2_ASAP7_75t_L g296 ( .A(n_182), .B(n_297), .Y(n_296) );
AND2x4_ASAP7_75t_L g337 ( .A(n_182), .B(n_253), .Y(n_337) );
OR2x6_ASAP7_75t_L g182 ( .A(n_183), .B(n_195), .Y(n_182) );
AOI21xp5_ASAP7_75t_SL g183 ( .A1(n_184), .A2(n_186), .B(n_193), .Y(n_183) );
AOI21xp5_ASAP7_75t_L g187 ( .A1(n_188), .A2(n_189), .B(n_190), .Y(n_187) );
INVx2_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
NAND2xp5_ASAP7_75t_SL g506 ( .A(n_191), .B(n_507), .Y(n_506) );
INVx1_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
NOR2xp33_ASAP7_75t_L g484 ( .A(n_194), .B(n_485), .Y(n_484) );
NOR2xp33_ASAP7_75t_L g195 ( .A(n_196), .B(n_197), .Y(n_195) );
AO21x2_ASAP7_75t_L g445 ( .A1(n_197), .A2(n_446), .B(n_453), .Y(n_445) );
INVx1_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_200), .B(n_213), .Y(n_199) );
AND2x2_ASAP7_75t_L g260 ( .A(n_200), .B(n_243), .Y(n_260) );
INVx1_ASAP7_75t_SL g200 ( .A(n_201), .Y(n_200) );
NAND2xp5_ASAP7_75t_SL g240 ( .A(n_201), .B(n_216), .Y(n_240) );
OR2x2_ASAP7_75t_L g273 ( .A(n_201), .B(n_243), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_201), .B(n_243), .Y(n_278) );
AND2x2_ASAP7_75t_L g305 ( .A(n_201), .B(n_242), .Y(n_305) );
AND2x2_ASAP7_75t_L g357 ( .A(n_201), .B(n_215), .Y(n_357) );
INVx2_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_202), .B(n_227), .Y(n_265) );
AND2x2_ASAP7_75t_L g301 ( .A(n_202), .B(n_216), .Y(n_301) );
AOI21xp5_ASAP7_75t_L g206 ( .A1(n_207), .A2(n_209), .B(n_210), .Y(n_206) );
AOI21xp5_ASAP7_75t_L g221 ( .A1(n_210), .A2(n_222), .B(n_223), .Y(n_221) );
INVx2_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
INVx3_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_213), .B(n_365), .Y(n_364) );
INVx2_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
OR2x2_ASAP7_75t_L g291 ( .A(n_214), .B(n_273), .Y(n_291) );
OR2x2_ASAP7_75t_L g214 ( .A(n_215), .B(n_227), .Y(n_214) );
OAI322xp33_ASAP7_75t_L g256 ( .A1(n_215), .A2(n_257), .A3(n_261), .B1(n_263), .B2(n_266), .C1(n_271), .C2(n_279), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_215), .B(n_242), .Y(n_264) );
OR2x2_ASAP7_75t_L g274 ( .A(n_215), .B(n_228), .Y(n_274) );
AND2x2_ASAP7_75t_L g276 ( .A(n_215), .B(n_228), .Y(n_276) );
NOR2xp33_ASAP7_75t_L g277 ( .A(n_215), .B(n_278), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_215), .B(n_243), .Y(n_338) );
NOR2xp33_ASAP7_75t_L g371 ( .A(n_215), .B(n_372), .Y(n_371) );
INVx5_ASAP7_75t_SL g215 ( .A(n_216), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_216), .B(n_260), .Y(n_386) );
OAI21xp5_ASAP7_75t_L g217 ( .A1(n_218), .A2(n_219), .B(n_220), .Y(n_217) );
OAI21xp5_ASAP7_75t_L g446 ( .A1(n_219), .A2(n_447), .B(n_448), .Y(n_446) );
OAI21xp5_ASAP7_75t_L g478 ( .A1(n_219), .A2(n_479), .B(n_480), .Y(n_478) );
NOR2xp33_ASAP7_75t_L g224 ( .A(n_225), .B(n_226), .Y(n_224) );
INVx2_ASAP7_75t_L g502 ( .A(n_226), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_227), .B(n_242), .Y(n_241) );
AND2x2_ASAP7_75t_L g254 ( .A(n_227), .B(n_255), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_227), .B(n_305), .Y(n_304) );
OR2x2_ASAP7_75t_L g316 ( .A(n_227), .B(n_243), .Y(n_316) );
AOI211xp5_ASAP7_75t_SL g344 ( .A1(n_227), .A2(n_345), .B(n_348), .C(n_360), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_227), .B(n_351), .Y(n_350) );
AND2x2_ASAP7_75t_L g382 ( .A(n_227), .B(n_357), .Y(n_382) );
INVx5_ASAP7_75t_SL g227 ( .A(n_228), .Y(n_227) );
AND2x2_ASAP7_75t_L g310 ( .A(n_228), .B(n_243), .Y(n_310) );
HB1xp67_ASAP7_75t_L g319 ( .A(n_228), .Y(n_319) );
AND2x2_ASAP7_75t_L g359 ( .A(n_228), .B(n_357), .Y(n_359) );
AND2x2_ASAP7_75t_SL g390 ( .A(n_228), .B(n_260), .Y(n_390) );
AND2x2_ASAP7_75t_L g397 ( .A(n_228), .B(n_356), .Y(n_397) );
OR2x6_ASAP7_75t_L g228 ( .A(n_229), .B(n_235), .Y(n_228) );
AOI22xp33_ASAP7_75t_L g236 ( .A1(n_237), .A2(n_238), .B1(n_252), .B2(n_254), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_237), .B(n_259), .Y(n_307) );
INVx2_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
OR2x2_ASAP7_75t_L g239 ( .A(n_240), .B(n_241), .Y(n_239) );
INVx1_ASAP7_75t_L g255 ( .A(n_240), .Y(n_255) );
OR2x2_ASAP7_75t_L g315 ( .A(n_240), .B(n_316), .Y(n_315) );
OAI221xp5_ASAP7_75t_SL g363 ( .A1(n_240), .A2(n_364), .B1(n_366), .B2(n_367), .C(n_369), .Y(n_363) );
INVx2_ASAP7_75t_L g302 ( .A(n_241), .Y(n_302) );
AND2x2_ASAP7_75t_L g275 ( .A(n_242), .B(n_276), .Y(n_275) );
INVx1_ASAP7_75t_L g365 ( .A(n_242), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_242), .B(n_357), .Y(n_378) );
INVx3_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
INVxp67_ASAP7_75t_L g320 ( .A(n_243), .Y(n_320) );
AND2x2_ASAP7_75t_L g356 ( .A(n_243), .B(n_357), .Y(n_356) );
OA21x2_ASAP7_75t_L g243 ( .A1(n_244), .A2(n_245), .B(n_251), .Y(n_243) );
OA21x2_ASAP7_75t_L g426 ( .A1(n_244), .A2(n_427), .B(n_433), .Y(n_426) );
OA21x2_ASAP7_75t_L g455 ( .A1(n_244), .A2(n_456), .B(n_463), .Y(n_455) );
OA21x2_ASAP7_75t_L g468 ( .A1(n_244), .A2(n_469), .B(n_476), .Y(n_468) );
AND2x2_ASAP7_75t_L g358 ( .A(n_252), .B(n_297), .Y(n_358) );
AND2x2_ASAP7_75t_L g268 ( .A(n_253), .B(n_269), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_253), .B(n_326), .Y(n_325) );
NOR2xp33_ASAP7_75t_SL g339 ( .A(n_255), .B(n_302), .Y(n_339) );
INVx1_ASAP7_75t_SL g257 ( .A(n_258), .Y(n_257) );
AND2x2_ASAP7_75t_L g345 ( .A(n_258), .B(n_346), .Y(n_345) );
AND2x2_ASAP7_75t_L g258 ( .A(n_259), .B(n_260), .Y(n_258) );
OR2x2_ASAP7_75t_L g331 ( .A(n_259), .B(n_332), .Y(n_331) );
AND2x2_ASAP7_75t_L g396 ( .A(n_259), .B(n_341), .Y(n_396) );
INVx2_ASAP7_75t_L g329 ( .A(n_260), .Y(n_329) );
NAND4xp25_ASAP7_75t_SL g392 ( .A(n_261), .B(n_393), .C(n_394), .D(n_395), .Y(n_392) );
INVx1_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_262), .B(n_326), .Y(n_361) );
OR2x2_ASAP7_75t_L g263 ( .A(n_264), .B(n_265), .Y(n_263) );
INVx1_ASAP7_75t_SL g398 ( .A(n_265), .Y(n_398) );
O2A1O1Ixp33_ASAP7_75t_SL g360 ( .A1(n_266), .A2(n_329), .B(n_333), .C(n_361), .Y(n_360) );
INVx1_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
AND2x2_ASAP7_75t_L g355 ( .A(n_268), .B(n_347), .Y(n_355) );
HB1xp67_ASAP7_75t_L g281 ( .A(n_269), .Y(n_281) );
INVx1_ASAP7_75t_L g336 ( .A(n_269), .Y(n_336) );
INVx2_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
HB1xp67_ASAP7_75t_L g313 ( .A(n_270), .Y(n_313) );
AOI211xp5_ASAP7_75t_L g271 ( .A1(n_272), .A2(n_274), .B(n_275), .C(n_277), .Y(n_271) );
AND2x2_ASAP7_75t_L g292 ( .A(n_272), .B(n_276), .Y(n_292) );
OAI322xp33_ASAP7_75t_SL g330 ( .A1(n_272), .A2(n_331), .A3(n_333), .B1(n_334), .B2(n_338), .C1(n_339), .C2(n_340), .Y(n_330) );
INVx1_ASAP7_75t_SL g272 ( .A(n_273), .Y(n_272) );
OR2x2_ASAP7_75t_L g352 ( .A(n_274), .B(n_278), .Y(n_352) );
INVx1_ASAP7_75t_L g333 ( .A(n_276), .Y(n_333) );
INVx1_ASAP7_75t_SL g351 ( .A(n_278), .Y(n_351) );
INVx2_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
AND2x2_ASAP7_75t_L g280 ( .A(n_281), .B(n_282), .Y(n_280) );
AOI222xp33_ASAP7_75t_L g283 ( .A1(n_284), .A2(n_290), .B1(n_292), .B2(n_293), .C1(n_294), .C2(n_704), .Y(n_283) );
NAND2xp5_ASAP7_75t_SL g284 ( .A(n_285), .B(n_287), .Y(n_284) );
OAI322xp33_ASAP7_75t_L g373 ( .A1(n_285), .A2(n_347), .A3(n_352), .B1(n_374), .B2(n_375), .C1(n_377), .C2(n_378), .Y(n_373) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
AOI221xp5_ASAP7_75t_L g323 ( .A1(n_286), .A2(n_300), .B1(n_324), .B2(n_328), .C(n_330), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_288), .B(n_289), .Y(n_287) );
INVx1_ASAP7_75t_SL g290 ( .A(n_291), .Y(n_290) );
OAI222xp33_ASAP7_75t_L g303 ( .A1(n_291), .A2(n_304), .B1(n_306), .B2(n_307), .C1(n_308), .C2(n_311), .Y(n_303) );
AOI22xp5_ASAP7_75t_L g369 ( .A1(n_293), .A2(n_300), .B1(n_370), .B2(n_371), .Y(n_369) );
AND2x2_ASAP7_75t_L g294 ( .A(n_295), .B(n_296), .Y(n_294) );
AOI211xp5_ASAP7_75t_L g298 ( .A1(n_299), .A2(n_300), .B(n_303), .C(n_314), .Y(n_298) );
O2A1O1Ixp33_ASAP7_75t_L g379 ( .A1(n_300), .A2(n_337), .B(n_380), .C(n_383), .Y(n_379) );
AND2x4_ASAP7_75t_L g300 ( .A(n_301), .B(n_302), .Y(n_300) );
AND2x2_ASAP7_75t_L g309 ( .A(n_301), .B(n_310), .Y(n_309) );
INVx1_ASAP7_75t_SL g372 ( .A(n_305), .Y(n_372) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_312), .B(n_337), .Y(n_366) );
BUFx2_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
AOI21xp33_ASAP7_75t_L g314 ( .A1(n_315), .A2(n_317), .B(n_321), .Y(n_314) );
OAI221xp5_ASAP7_75t_SL g383 ( .A1(n_315), .A2(n_384), .B1(n_385), .B2(n_386), .C(n_387), .Y(n_383) );
INVxp33_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
NOR2xp33_ASAP7_75t_L g318 ( .A(n_319), .B(n_320), .Y(n_318) );
NOR2xp33_ASAP7_75t_L g328 ( .A(n_319), .B(n_329), .Y(n_328) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_326), .B(n_337), .Y(n_377) );
INVx2_ASAP7_75t_SL g326 ( .A(n_327), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_335), .B(n_337), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_341), .B(n_342), .Y(n_340) );
AND2x2_ASAP7_75t_L g388 ( .A(n_341), .B(n_347), .Y(n_388) );
AND4x1_ASAP7_75t_L g343 ( .A(n_344), .B(n_362), .C(n_379), .D(n_391), .Y(n_343) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
OAI221xp5_ASAP7_75t_SL g348 ( .A1(n_349), .A2(n_350), .B1(n_352), .B2(n_353), .C(n_354), .Y(n_348) );
AOI22xp5_ASAP7_75t_L g354 ( .A1(n_355), .A2(n_356), .B1(n_358), .B2(n_359), .Y(n_354) );
INVx1_ASAP7_75t_L g384 ( .A(n_355), .Y(n_384) );
INVx1_ASAP7_75t_SL g374 ( .A(n_359), .Y(n_374) );
NOR2xp33_ASAP7_75t_SL g362 ( .A(n_363), .B(n_373), .Y(n_362) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
NOR2xp33_ASAP7_75t_L g380 ( .A(n_375), .B(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
AOI22xp33_ASAP7_75t_L g387 ( .A1(n_382), .A2(n_388), .B1(n_389), .B2(n_390), .Y(n_387) );
AOI22xp5_ASAP7_75t_L g391 ( .A1(n_392), .A2(n_397), .B1(n_398), .B2(n_399), .Y(n_391) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx1_ASAP7_75t_SL g401 ( .A(n_402), .Y(n_401) );
INVx1_ASAP7_75t_SL g402 ( .A(n_403), .Y(n_402) );
INVx2_ASAP7_75t_L g411 ( .A(n_403), .Y(n_411) );
NOR2x2_ASAP7_75t_L g686 ( .A(n_404), .B(n_419), .Y(n_686) );
INVx2_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
OR2x2_ASAP7_75t_L g418 ( .A(n_405), .B(n_419), .Y(n_418) );
AND2x2_ASAP7_75t_L g405 ( .A(n_406), .B(n_407), .Y(n_405) );
NAND3xp33_ASAP7_75t_SL g697 ( .A(n_406), .B(n_419), .C(n_698), .Y(n_697) );
OAI21xp5_ASAP7_75t_SL g412 ( .A1(n_408), .A2(n_413), .B(n_688), .Y(n_412) );
NOR2xp33_ASAP7_75t_L g408 ( .A(n_409), .B(n_410), .Y(n_408) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx6_ASAP7_75t_L g682 ( .A(n_418), .Y(n_682) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
BUFx2_ASAP7_75t_L g683 ( .A(n_421), .Y(n_683) );
AND2x2_ASAP7_75t_L g421 ( .A(n_422), .B(n_607), .Y(n_421) );
NOR4xp25_ASAP7_75t_L g422 ( .A(n_423), .B(n_549), .C(n_579), .D(n_589), .Y(n_422) );
OAI211xp5_ASAP7_75t_L g423 ( .A1(n_424), .A2(n_464), .B(n_512), .C(n_539), .Y(n_423) );
OAI222xp33_ASAP7_75t_L g634 ( .A1(n_424), .A2(n_554), .B1(n_635), .B2(n_636), .C1(n_637), .C2(n_638), .Y(n_634) );
OR2x2_ASAP7_75t_L g424 ( .A(n_425), .B(n_443), .Y(n_424) );
AOI33xp33_ASAP7_75t_L g560 ( .A1(n_425), .A2(n_547), .A3(n_548), .B1(n_561), .B2(n_566), .B3(n_568), .Y(n_560) );
OAI211xp5_ASAP7_75t_SL g617 ( .A1(n_425), .A2(n_618), .B(n_620), .C(n_622), .Y(n_617) );
OR2x2_ASAP7_75t_L g633 ( .A(n_425), .B(n_619), .Y(n_633) );
INVx1_ASAP7_75t_L g666 ( .A(n_425), .Y(n_666) );
OR2x2_ASAP7_75t_L g425 ( .A(n_426), .B(n_434), .Y(n_425) );
INVx2_ASAP7_75t_L g543 ( .A(n_426), .Y(n_543) );
AND2x2_ASAP7_75t_L g559 ( .A(n_426), .B(n_455), .Y(n_559) );
HB1xp67_ASAP7_75t_L g594 ( .A(n_426), .Y(n_594) );
AND2x2_ASAP7_75t_L g623 ( .A(n_426), .B(n_434), .Y(n_623) );
INVx2_ASAP7_75t_L g523 ( .A(n_434), .Y(n_523) );
BUFx3_ASAP7_75t_L g531 ( .A(n_434), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_434), .B(n_534), .Y(n_533) );
AND2x2_ASAP7_75t_L g542 ( .A(n_434), .B(n_543), .Y(n_542) );
NOR2xp33_ASAP7_75t_L g571 ( .A(n_434), .B(n_444), .Y(n_571) );
AND2x2_ASAP7_75t_L g640 ( .A(n_434), .B(n_574), .Y(n_640) );
INVx2_ASAP7_75t_SL g534 ( .A(n_443), .Y(n_534) );
OR2x2_ASAP7_75t_L g443 ( .A(n_444), .B(n_455), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_444), .B(n_523), .Y(n_522) );
INVx1_ASAP7_75t_L g576 ( .A(n_444), .Y(n_576) );
AND2x2_ASAP7_75t_L g587 ( .A(n_444), .B(n_543), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_444), .B(n_572), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_444), .B(n_574), .Y(n_619) );
AND2x2_ASAP7_75t_L g678 ( .A(n_444), .B(n_623), .Y(n_678) );
INVx4_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
AND2x2_ASAP7_75t_L g548 ( .A(n_445), .B(n_455), .Y(n_548) );
AND2x2_ASAP7_75t_L g558 ( .A(n_445), .B(n_559), .Y(n_558) );
BUFx3_ASAP7_75t_L g580 ( .A(n_445), .Y(n_580) );
AND3x2_ASAP7_75t_L g639 ( .A(n_445), .B(n_640), .C(n_641), .Y(n_639) );
HB1xp67_ASAP7_75t_L g530 ( .A(n_455), .Y(n_530) );
INVx1_ASAP7_75t_SL g574 ( .A(n_455), .Y(n_574) );
NAND3xp33_ASAP7_75t_L g586 ( .A(n_455), .B(n_523), .C(n_587), .Y(n_586) );
NOR2xp33_ASAP7_75t_L g464 ( .A(n_465), .B(n_495), .Y(n_464) );
A2O1A1Ixp33_ASAP7_75t_L g609 ( .A1(n_465), .A2(n_558), .B(n_610), .C(n_612), .Y(n_609) );
INVx1_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
NAND2xp5_ASAP7_75t_SL g466 ( .A(n_467), .B(n_486), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_467), .B(n_616), .Y(n_615) );
INVx2_ASAP7_75t_SL g626 ( .A(n_467), .Y(n_626) );
AND2x2_ASAP7_75t_L g647 ( .A(n_467), .B(n_497), .Y(n_647) );
NOR2xp33_ASAP7_75t_L g675 ( .A(n_467), .B(n_556), .Y(n_675) );
AND2x2_ASAP7_75t_L g467 ( .A(n_468), .B(n_477), .Y(n_467) );
AND2x2_ASAP7_75t_L g520 ( .A(n_468), .B(n_511), .Y(n_520) );
INVx2_ASAP7_75t_L g527 ( .A(n_468), .Y(n_527) );
AND2x2_ASAP7_75t_L g547 ( .A(n_468), .B(n_497), .Y(n_547) );
AND2x2_ASAP7_75t_L g597 ( .A(n_468), .B(n_486), .Y(n_597) );
INVx1_ASAP7_75t_L g601 ( .A(n_468), .Y(n_601) );
INVx2_ASAP7_75t_SL g511 ( .A(n_477), .Y(n_511) );
BUFx2_ASAP7_75t_L g537 ( .A(n_477), .Y(n_537) );
AND2x2_ASAP7_75t_L g664 ( .A(n_477), .B(n_486), .Y(n_664) );
INVx3_ASAP7_75t_SL g497 ( .A(n_486), .Y(n_497) );
AND2x2_ASAP7_75t_L g519 ( .A(n_486), .B(n_520), .Y(n_519) );
AND2x4_ASAP7_75t_L g526 ( .A(n_486), .B(n_527), .Y(n_526) );
OR2x2_ASAP7_75t_L g556 ( .A(n_486), .B(n_516), .Y(n_556) );
OR2x2_ASAP7_75t_L g565 ( .A(n_486), .B(n_511), .Y(n_565) );
HB1xp67_ASAP7_75t_L g583 ( .A(n_486), .Y(n_583) );
AND2x2_ASAP7_75t_L g588 ( .A(n_486), .B(n_541), .Y(n_588) );
AND2x2_ASAP7_75t_L g616 ( .A(n_486), .B(n_499), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_486), .B(n_652), .Y(n_651) );
OR2x2_ASAP7_75t_L g654 ( .A(n_486), .B(n_498), .Y(n_654) );
OR2x6_ASAP7_75t_L g486 ( .A(n_487), .B(n_493), .Y(n_486) );
INVx1_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
OR2x2_ASAP7_75t_L g496 ( .A(n_497), .B(n_498), .Y(n_496) );
AND2x2_ASAP7_75t_L g578 ( .A(n_497), .B(n_527), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_497), .B(n_520), .Y(n_606) );
AND2x2_ASAP7_75t_L g624 ( .A(n_497), .B(n_541), .Y(n_624) );
OR2x2_ASAP7_75t_L g498 ( .A(n_499), .B(n_511), .Y(n_498) );
AND2x2_ASAP7_75t_L g525 ( .A(n_499), .B(n_511), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_499), .B(n_554), .Y(n_553) );
BUFx3_ASAP7_75t_L g563 ( .A(n_499), .Y(n_563) );
OR2x2_ASAP7_75t_L g611 ( .A(n_499), .B(n_531), .Y(n_611) );
OA21x2_ASAP7_75t_L g499 ( .A1(n_500), .A2(n_503), .B(n_510), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
AO21x2_ASAP7_75t_L g516 ( .A1(n_501), .A2(n_517), .B(n_518), .Y(n_516) );
INVx1_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
INVx1_ASAP7_75t_L g517 ( .A(n_503), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_510), .Y(n_518) );
AND2x2_ASAP7_75t_L g546 ( .A(n_511), .B(n_516), .Y(n_546) );
INVx1_ASAP7_75t_L g554 ( .A(n_511), .Y(n_554) );
AND2x2_ASAP7_75t_L g649 ( .A(n_511), .B(n_527), .Y(n_649) );
AOI222xp33_ASAP7_75t_L g512 ( .A1(n_513), .A2(n_521), .B1(n_524), .B2(n_528), .C1(n_532), .C2(n_535), .Y(n_512) );
INVx1_ASAP7_75t_L g644 ( .A(n_513), .Y(n_644) );
AND2x2_ASAP7_75t_L g513 ( .A(n_514), .B(n_519), .Y(n_513) );
AND2x2_ASAP7_75t_L g540 ( .A(n_514), .B(n_541), .Y(n_540) );
AND2x2_ASAP7_75t_L g551 ( .A(n_514), .B(n_520), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_514), .B(n_542), .Y(n_567) );
OAI222xp33_ASAP7_75t_L g589 ( .A1(n_514), .A2(n_590), .B1(n_595), .B2(n_596), .C1(n_604), .C2(n_606), .Y(n_589) );
INVx2_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
INVx1_ASAP7_75t_SL g515 ( .A(n_516), .Y(n_515) );
AND2x2_ASAP7_75t_L g577 ( .A(n_516), .B(n_578), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_516), .B(n_597), .Y(n_637) );
AND2x2_ASAP7_75t_L g648 ( .A(n_516), .B(n_649), .Y(n_648) );
INVx1_ASAP7_75t_L g656 ( .A(n_519), .Y(n_656) );
NAND2xp5_ASAP7_75t_SL g635 ( .A(n_521), .B(n_572), .Y(n_635) );
INVx1_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
NOR2xp33_ASAP7_75t_L g575 ( .A(n_523), .B(n_576), .Y(n_575) );
AND2x2_ASAP7_75t_L g593 ( .A(n_523), .B(n_594), .Y(n_593) );
AND2x2_ASAP7_75t_L g524 ( .A(n_525), .B(n_526), .Y(n_524) );
INVx3_ASAP7_75t_L g538 ( .A(n_526), .Y(n_538) );
O2A1O1Ixp33_ASAP7_75t_L g628 ( .A1(n_526), .A2(n_629), .B(n_632), .C(n_634), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_526), .B(n_563), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_526), .B(n_546), .Y(n_668) );
AND2x2_ASAP7_75t_L g541 ( .A(n_527), .B(n_537), .Y(n_541) );
INVx1_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_530), .B(n_531), .Y(n_529) );
INVx1_ASAP7_75t_L g568 ( .A(n_530), .Y(n_568) );
NAND2xp5_ASAP7_75t_SL g557 ( .A(n_531), .B(n_558), .Y(n_557) );
OR2x2_ASAP7_75t_L g620 ( .A(n_531), .B(n_621), .Y(n_620) );
AND2x2_ASAP7_75t_L g659 ( .A(n_531), .B(n_559), .Y(n_659) );
INVx1_ASAP7_75t_L g671 ( .A(n_531), .Y(n_671) );
INVx1_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_534), .B(n_673), .Y(n_672) );
INVx1_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
OR2x2_ASAP7_75t_L g536 ( .A(n_537), .B(n_538), .Y(n_536) );
INVx1_ASAP7_75t_L g652 ( .A(n_537), .Y(n_652) );
A2O1A1Ixp33_ASAP7_75t_SL g539 ( .A1(n_540), .A2(n_542), .B(n_544), .C(n_548), .Y(n_539) );
AOI22xp33_ASAP7_75t_L g584 ( .A1(n_540), .A2(n_570), .B1(n_585), .B2(n_588), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_541), .B(n_555), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_541), .B(n_563), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_542), .B(n_600), .Y(n_599) );
INVx1_ASAP7_75t_SL g605 ( .A(n_542), .Y(n_605) );
AND2x2_ASAP7_75t_L g612 ( .A(n_542), .B(n_592), .Y(n_612) );
INVx2_ASAP7_75t_L g573 ( .A(n_543), .Y(n_573) );
INVxp67_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_546), .B(n_547), .Y(n_545) );
NOR4xp25_ASAP7_75t_L g550 ( .A(n_547), .B(n_551), .C(n_552), .D(n_555), .Y(n_550) );
INVx1_ASAP7_75t_SL g621 ( .A(n_548), .Y(n_621) );
AND2x2_ASAP7_75t_L g665 ( .A(n_548), .B(n_666), .Y(n_665) );
OAI211xp5_ASAP7_75t_SL g549 ( .A1(n_550), .A2(n_557), .B(n_560), .C(n_569), .Y(n_549) );
INVx1_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
INVx1_ASAP7_75t_SL g555 ( .A(n_556), .Y(n_555) );
NOR2xp33_ASAP7_75t_L g677 ( .A(n_556), .B(n_626), .Y(n_677) );
AOI22xp5_ASAP7_75t_L g676 ( .A1(n_558), .A2(n_677), .B1(n_678), .B2(n_679), .Y(n_676) );
INVx1_ASAP7_75t_SL g631 ( .A(n_559), .Y(n_631) );
AND2x2_ASAP7_75t_L g670 ( .A(n_559), .B(n_671), .Y(n_670) );
INVx1_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_563), .B(n_564), .Y(n_562) );
NAND2xp5_ASAP7_75t_SL g663 ( .A(n_563), .B(n_664), .Y(n_663) );
INVx1_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
INVx1_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
NOR2xp33_ASAP7_75t_L g582 ( .A(n_567), .B(n_583), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_568), .B(n_593), .Y(n_653) );
OAI21xp5_ASAP7_75t_SL g569 ( .A1(n_570), .A2(n_575), .B(n_577), .Y(n_569) );
AND2x2_ASAP7_75t_L g570 ( .A(n_571), .B(n_572), .Y(n_570) );
INVx1_ASAP7_75t_L g645 ( .A(n_572), .Y(n_645) );
AND2x2_ASAP7_75t_L g572 ( .A(n_573), .B(n_574), .Y(n_572) );
INVx2_ASAP7_75t_L g673 ( .A(n_573), .Y(n_673) );
HB1xp67_ASAP7_75t_L g600 ( .A(n_574), .Y(n_600) );
OAI21xp33_ASAP7_75t_L g579 ( .A1(n_580), .A2(n_581), .B(n_584), .Y(n_579) );
CKINVDCx16_ASAP7_75t_R g592 ( .A(n_580), .Y(n_592) );
OR2x2_ASAP7_75t_L g630 ( .A(n_580), .B(n_631), .Y(n_630) );
INVx1_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
AOI21xp33_ASAP7_75t_SL g625 ( .A1(n_583), .A2(n_626), .B(n_627), .Y(n_625) );
INVx1_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
AOI221xp5_ASAP7_75t_L g613 ( .A1(n_587), .A2(n_614), .B1(n_617), .B2(n_624), .C(n_625), .Y(n_613) );
INVx1_ASAP7_75t_SL g657 ( .A(n_588), .Y(n_657) );
INVx1_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
AND2x2_ASAP7_75t_L g591 ( .A(n_592), .B(n_593), .Y(n_591) );
OR2x2_ASAP7_75t_L g604 ( .A(n_592), .B(n_605), .Y(n_604) );
INVxp67_ASAP7_75t_L g641 ( .A(n_594), .Y(n_641) );
AOI22xp5_ASAP7_75t_L g596 ( .A1(n_597), .A2(n_598), .B1(n_601), .B2(n_602), .Y(n_596) );
INVx1_ASAP7_75t_L g636 ( .A(n_597), .Y(n_636) );
INVxp67_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_600), .B(n_623), .Y(n_622) );
INVx1_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
NOR4xp25_ASAP7_75t_L g607 ( .A(n_608), .B(n_642), .C(n_655), .D(n_667), .Y(n_607) );
NAND3xp33_ASAP7_75t_SL g608 ( .A(n_609), .B(n_613), .C(n_628), .Y(n_608) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
NOR2xp33_ASAP7_75t_L g629 ( .A(n_611), .B(n_630), .Y(n_629) );
INVx1_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_618), .B(n_623), .Y(n_627) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
OAI221xp5_ASAP7_75t_SL g655 ( .A1(n_630), .A2(n_656), .B1(n_657), .B2(n_658), .C(n_660), .Y(n_655) );
O2A1O1Ixp33_ASAP7_75t_L g646 ( .A1(n_632), .A2(n_647), .B(n_648), .C(n_650), .Y(n_646) );
INVx2_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
OAI22xp5_ASAP7_75t_L g650 ( .A1(n_633), .A2(n_651), .B1(n_653), .B2(n_654), .Y(n_650) );
INVx2_ASAP7_75t_SL g638 ( .A(n_639), .Y(n_638) );
A2O1A1Ixp33_ASAP7_75t_L g642 ( .A1(n_643), .A2(n_644), .B(n_645), .C(n_646), .Y(n_642) );
INVx1_ASAP7_75t_L g661 ( .A(n_654), .Y(n_661) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
OAI21xp5_ASAP7_75t_SL g660 ( .A1(n_661), .A2(n_662), .B(n_665), .Y(n_660) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
OAI221xp5_ASAP7_75t_SL g667 ( .A1(n_668), .A2(n_669), .B1(n_672), .B2(n_674), .C(n_676), .Y(n_667) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
INVxp67_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
INVx3_ASAP7_75t_SL g685 ( .A(n_686), .Y(n_685) );
BUFx2_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
CKINVDCx9p33_ASAP7_75t_R g692 ( .A(n_693), .Y(n_692) );
INVx1_ASAP7_75t_L g702 ( .A(n_693), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_694), .B(n_696), .Y(n_693) );
CKINVDCx20_ASAP7_75t_R g694 ( .A(n_695), .Y(n_694) );
CKINVDCx14_ASAP7_75t_R g696 ( .A(n_697), .Y(n_696) );
INVx1_ASAP7_75t_SL g698 ( .A(n_699), .Y(n_698) );
INVx1_ASAP7_75t_SL g701 ( .A(n_702), .Y(n_701) );
endmodule