module real_jpeg_4920_n_29 (n_17, n_8, n_0, n_21, n_168, n_2, n_10, n_9, n_12, n_24, n_165, n_166, n_170, n_6, n_28, n_171, n_169, n_167, n_23, n_11, n_14, n_172, n_25, n_163, n_7, n_22, n_18, n_3, n_5, n_4, n_1, n_26, n_27, n_20, n_19, n_164, n_16, n_15, n_13, n_29);

input n_17;
input n_8;
input n_0;
input n_21;
input n_168;
input n_2;
input n_10;
input n_9;
input n_12;
input n_24;
input n_165;
input n_166;
input n_170;
input n_6;
input n_28;
input n_171;
input n_169;
input n_167;
input n_23;
input n_11;
input n_14;
input n_172;
input n_25;
input n_163;
input n_7;
input n_22;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_26;
input n_27;
input n_20;
input n_19;
input n_164;
input n_16;
input n_15;
input n_13;

output n_29;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_47;
wire n_131;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_56;
wire n_48;
wire n_140;
wire n_126;
wire n_113;
wire n_120;
wire n_155;
wire n_93;
wire n_141;
wire n_95;
wire n_139;
wire n_33;
wire n_65;
wire n_142;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_66;
wire n_136;
wire n_44;
wire n_62;
wire n_121;
wire n_106;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_148;
wire n_118;
wire n_123;
wire n_116;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_134;
wire n_72;
wire n_159;
wire n_151;
wire n_100;
wire n_51;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_150;
wire n_80;
wire n_41;
wire n_32;
wire n_74;
wire n_30;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_92;
wire n_97;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_138;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g75 ( 
.A(n_0),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_0),
.B(n_89),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_1),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_2),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_3),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_4),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_5),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_6),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_7),
.B(n_42),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_7),
.B(n_42),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_8),
.B(n_64),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_8),
.B(n_64),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_9),
.B(n_101),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_9),
.B(n_101),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_10),
.B(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_10),
.B(n_54),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_11),
.B(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_12),
.Y(n_85)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_13),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_14),
.B(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_14),
.B(n_57),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_15),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_16),
.B(n_127),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_16),
.B(n_127),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_17),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_18),
.B(n_145),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_18),
.B(n_145),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_19),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_20),
.B(n_88),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_20),
.B(n_88),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_21),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_22),
.B(n_48),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_22),
.B(n_48),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_23),
.Y(n_122)
);

OR2x2_ASAP7_75t_L g115 ( 
.A(n_24),
.B(n_116),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_24),
.B(n_116),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_25),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_26),
.B(n_32),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_26),
.B(n_141),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_26),
.B(n_141),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_26),
.B(n_32),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_26),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_27),
.B(n_69),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_27),
.B(n_69),
.Y(n_94)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_28),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_151),
.Y(n_29)
);

OAI21xp5_ASAP7_75t_L g30 ( 
.A1(n_31),
.A2(n_37),
.B(n_150),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_34),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_34),
.B(n_58),
.Y(n_57)
);

BUFx8_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_35),
.B(n_70),
.Y(n_69)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_35),
.Y(n_124)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

AOI21xp5_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_139),
.B(n_147),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_SL g38 ( 
.A1(n_39),
.A2(n_118),
.B(n_133),
.Y(n_38)
);

A2O1A1Ixp33_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_59),
.B(n_106),
.C(n_115),
.Y(n_39)
);

NOR4xp25_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_47),
.C(n_53),
.D(n_56),
.Y(n_40)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_41),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_44),
.Y(n_42)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_46),
.Y(n_143)
);

INVx11_ASAP7_75t_L g159 ( 
.A(n_46),
.Y(n_159)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_47),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_50),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_50),
.B(n_55),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_50),
.B(n_117),
.Y(n_116)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_52),
.B(n_81),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_53),
.A2(n_110),
.B(n_111),
.Y(n_109)
);

OAI21x1_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_100),
.B(n_105),
.Y(n_59)
);

AOI21xp5_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_95),
.B(n_99),
.Y(n_60)
);

AO221x1_ASAP7_75t_L g61 ( 
.A1(n_62),
.A2(n_71),
.B1(n_92),
.B2(n_93),
.C(n_94),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_68),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_66),
.Y(n_64)
);

OR2x2_ASAP7_75t_L g96 ( 
.A(n_66),
.B(n_97),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_66),
.B(n_128),
.Y(n_127)
);

BUFx12_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_68),
.Y(n_92)
);

AO21x1_ASAP7_75t_L g71 ( 
.A1(n_72),
.A2(n_77),
.B(n_91),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_73),
.B(n_76),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_73),
.B(n_76),
.Y(n_91)
);

OR2x2_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_75),
.Y(n_73)
);

OR2x2_ASAP7_75t_L g83 ( 
.A(n_75),
.B(n_84),
.Y(n_83)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_75),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_87),
.B(n_90),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_82),
.B(n_86),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_83),
.B(n_85),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_83),
.B(n_85),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_96),
.B(n_98),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_96),
.B(n_98),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_103),
.Y(n_101)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

A2O1A1O1Ixp25_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_109),
.B(n_112),
.C(n_113),
.D(n_114),
.Y(n_107)
);

NAND3xp33_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_125),
.C(n_129),
.Y(n_118)
);

A2O1A1O1Ixp25_ASAP7_75t_L g133 ( 
.A1(n_119),
.A2(n_129),
.B(n_134),
.C(n_137),
.D(n_138),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_121),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_120),
.B(n_121),
.Y(n_138)
);

OR2x2_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_123),
.Y(n_121)
);

OR2x2_ASAP7_75t_L g130 ( 
.A(n_123),
.B(n_131),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_123),
.B(n_146),
.Y(n_145)
);

INVx8_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_126),
.A2(n_135),
.B(n_136),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_130),
.B(n_132),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_130),
.B(n_132),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_144),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_143),
.Y(n_141)
);

OAI21xp33_ASAP7_75t_L g147 ( 
.A1(n_144),
.A2(n_148),
.B(n_149),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_161),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_153),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_154),
.B(n_160),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_154),
.B(n_160),
.Y(n_161)
);

OR2x2_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_156),
.Y(n_154)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_158),
.Y(n_157)
);

BUFx3_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_163),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_164),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_165),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_166),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_167),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_168),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_169),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_170),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_171),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_172),
.Y(n_102)
);


endmodule