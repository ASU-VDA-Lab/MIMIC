module fake_jpeg_2154_n_327 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_327);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_327;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_15),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_10),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

CKINVDCx14_ASAP7_75t_R g23 ( 
.A(n_16),
.Y(n_23)
);

BUFx4f_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_13),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_5),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

BUFx12_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_0),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_9),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_5),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_13),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_14),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_9),
.Y(n_44)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_2),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_8),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_48),
.Y(n_97)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_49),
.Y(n_119)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_47),
.Y(n_50)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_50),
.Y(n_116)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_51),
.Y(n_103)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

INVx11_ASAP7_75t_L g145 ( 
.A(n_52),
.Y(n_145)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_22),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_53),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_28),
.B(n_12),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_54),
.B(n_69),
.Y(n_137)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_28),
.Y(n_55)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_55),
.Y(n_105)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_56),
.Y(n_123)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_32),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g96 ( 
.A(n_57),
.Y(n_96)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g142 ( 
.A(n_58),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_22),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_59),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_23),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_60),
.B(n_67),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g132 ( 
.A(n_61),
.Y(n_132)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_62),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_63),
.Y(n_141)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_34),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_64),
.Y(n_147)
);

OR2x2_ASAP7_75t_SL g65 ( 
.A(n_41),
.B(n_0),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_65),
.B(n_35),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_66),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_17),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_68),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_18),
.B(n_0),
.Y(n_69)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_29),
.Y(n_70)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_70),
.Y(n_148)
);

INVx11_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_71),
.Y(n_129)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_21),
.Y(n_72)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_72),
.Y(n_109)
);

BUFx5_ASAP7_75t_L g73 ( 
.A(n_21),
.Y(n_73)
);

INVx13_ASAP7_75t_L g100 ( 
.A(n_73),
.Y(n_100)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_34),
.Y(n_74)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_74),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_17),
.B(n_1),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_75),
.B(n_85),
.Y(n_138)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_29),
.Y(n_76)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_76),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_19),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_77),
.B(n_78),
.Y(n_113)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_21),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_26),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_79),
.B(n_83),
.Y(n_101)
);

BUFx16f_ASAP7_75t_L g80 ( 
.A(n_21),
.Y(n_80)
);

CKINVDCx12_ASAP7_75t_R g124 ( 
.A(n_80),
.Y(n_124)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_19),
.Y(n_81)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_81),
.Y(n_115)
);

AOI21xp33_ASAP7_75t_SL g82 ( 
.A1(n_24),
.A2(n_2),
.B(n_4),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_82),
.B(n_84),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_26),
.Y(n_83)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_24),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_46),
.B(n_6),
.Y(n_85)
);

BUFx5_ASAP7_75t_L g86 ( 
.A(n_24),
.Y(n_86)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_86),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_42),
.B(n_6),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_87),
.B(n_51),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_20),
.Y(n_88)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_88),
.Y(n_126)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_20),
.Y(n_89)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_89),
.Y(n_140)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_18),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_90),
.B(n_92),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_42),
.B(n_7),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_91),
.B(n_93),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_25),
.Y(n_92)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_27),
.Y(n_93)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_27),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_94),
.B(n_44),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_98),
.B(n_128),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_89),
.B(n_41),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_102),
.B(n_110),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_59),
.A2(n_33),
.B1(n_36),
.B2(n_40),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_106),
.A2(n_108),
.B1(n_139),
.B2(n_129),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_52),
.A2(n_46),
.B1(n_44),
.B2(n_38),
.Y(n_107)
);

OA22x2_ASAP7_75t_L g150 ( 
.A1(n_107),
.A2(n_133),
.B1(n_135),
.B2(n_56),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_88),
.A2(n_33),
.B1(n_40),
.B2(n_36),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_77),
.B(n_38),
.Y(n_110)
);

CKINVDCx14_ASAP7_75t_R g182 ( 
.A(n_117),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_80),
.B(n_37),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_121),
.B(n_127),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_61),
.A2(n_25),
.B1(n_30),
.B2(n_37),
.Y(n_122)
);

OR2x2_ASAP7_75t_L g153 ( 
.A(n_122),
.B(n_146),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_93),
.B(n_31),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_92),
.B(n_31),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_72),
.A2(n_35),
.B1(n_30),
.B2(n_11),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_51),
.B(n_7),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_134),
.B(n_74),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_63),
.A2(n_7),
.B1(n_8),
.B2(n_11),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_70),
.B(n_12),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_136),
.B(n_144),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_62),
.A2(n_12),
.B1(n_66),
.B2(n_78),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_53),
.B(n_76),
.Y(n_146)
);

INVx5_ASAP7_75t_L g149 ( 
.A(n_132),
.Y(n_149)
);

INVx1_ASAP7_75t_SL g208 ( 
.A(n_149),
.Y(n_208)
);

A2O1A1Ixp33_ASAP7_75t_SL g222 ( 
.A1(n_150),
.A2(n_190),
.B(n_181),
.C(n_184),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_101),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_152),
.B(n_173),
.Y(n_195)
);

INVx8_ASAP7_75t_L g154 ( 
.A(n_142),
.Y(n_154)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_154),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_130),
.A2(n_58),
.B1(n_64),
.B2(n_74),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_155),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_131),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_156),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_157),
.B(n_159),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_137),
.B(n_120),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_158),
.B(n_164),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_95),
.B(n_111),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_105),
.B(n_58),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_160),
.B(n_171),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_130),
.A2(n_64),
.B1(n_120),
.B2(n_113),
.Y(n_161)
);

INVxp33_ASAP7_75t_L g201 ( 
.A(n_161),
.Y(n_201)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_114),
.Y(n_162)
);

HB1xp67_ASAP7_75t_L g200 ( 
.A(n_162),
.Y(n_200)
);

OAI32xp33_ASAP7_75t_L g163 ( 
.A1(n_138),
.A2(n_97),
.A3(n_143),
.B1(n_115),
.B2(n_140),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_163),
.B(n_166),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_148),
.B(n_126),
.Y(n_164)
);

OR2x2_ASAP7_75t_SL g165 ( 
.A(n_116),
.B(n_119),
.Y(n_165)
);

CKINVDCx14_ASAP7_75t_R g221 ( 
.A(n_165),
.Y(n_221)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_113),
.B(n_118),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_125),
.Y(n_167)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_167),
.Y(n_203)
);

INVx8_ASAP7_75t_L g168 ( 
.A(n_142),
.Y(n_168)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_168),
.Y(n_211)
);

INVxp33_ASAP7_75t_L g220 ( 
.A(n_170),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_123),
.B(n_132),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_135),
.B(n_107),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_L g174 ( 
.A1(n_131),
.A2(n_104),
.B1(n_141),
.B2(n_145),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_174),
.A2(n_184),
.B1(n_188),
.B2(n_191),
.Y(n_193)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_123),
.Y(n_175)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_175),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_104),
.B(n_99),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_176),
.B(n_180),
.Y(n_202)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_99),
.Y(n_177)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_177),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_112),
.B(n_103),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_178),
.B(n_179),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_112),
.B(n_103),
.Y(n_179)
);

OR2x2_ASAP7_75t_SL g180 ( 
.A(n_119),
.B(n_124),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_147),
.B(n_141),
.C(n_129),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_181),
.B(n_165),
.C(n_166),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_133),
.A2(n_147),
.B1(n_109),
.B2(n_100),
.Y(n_184)
);

INVx8_ASAP7_75t_L g185 ( 
.A(n_142),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_185),
.B(n_186),
.Y(n_207)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_109),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_145),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_187),
.B(n_191),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_96),
.B(n_100),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_188),
.B(n_180),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_96),
.A2(n_120),
.B(n_102),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_189),
.A2(n_166),
.B(n_151),
.Y(n_213)
);

A2O1A1Ixp33_ASAP7_75t_SL g190 ( 
.A1(n_96),
.A2(n_120),
.B(n_146),
.C(n_82),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_113),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_101),
.B(n_95),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_192),
.B(n_183),
.Y(n_215)
);

INVx1_ASAP7_75t_SL g242 ( 
.A(n_193),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_173),
.A2(n_153),
.B1(n_170),
.B2(n_158),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_194),
.A2(n_198),
.B1(n_150),
.B2(n_156),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_153),
.A2(n_176),
.B1(n_164),
.B2(n_190),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_205),
.B(n_221),
.Y(n_239)
);

FAx1_ASAP7_75t_SL g210 ( 
.A(n_190),
.B(n_189),
.CI(n_172),
.CON(n_210),
.SN(n_210)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_210),
.B(n_226),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_182),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_212),
.B(n_224),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_213),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_215),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_217),
.B(n_225),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_222),
.B(n_185),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_169),
.B(n_162),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_190),
.B(n_150),
.C(n_163),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_149),
.B(n_177),
.Y(n_226)
);

INVx13_ASAP7_75t_L g228 ( 
.A(n_208),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_228),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_229),
.B(n_247),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_220),
.A2(n_150),
.B1(n_154),
.B2(n_168),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_231),
.A2(n_240),
.B1(n_222),
.B2(n_203),
.Y(n_267)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_218),
.Y(n_232)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_232),
.Y(n_252)
);

BUFx4f_ASAP7_75t_L g233 ( 
.A(n_200),
.Y(n_233)
);

INVx4_ASAP7_75t_L g257 ( 
.A(n_233),
.Y(n_257)
);

INVx13_ASAP7_75t_L g234 ( 
.A(n_208),
.Y(n_234)
);

CKINVDCx16_ASAP7_75t_R g261 ( 
.A(n_234),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_207),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_235),
.B(n_238),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_237),
.A2(n_244),
.B(n_231),
.Y(n_269)
);

INVx8_ASAP7_75t_L g238 ( 
.A(n_199),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_239),
.B(n_249),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_194),
.A2(n_225),
.B1(n_198),
.B2(n_195),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_214),
.B(n_206),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_243),
.B(n_245),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_223),
.A2(n_201),
.B(n_206),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_204),
.B(n_216),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_214),
.B(n_206),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_246),
.B(n_248),
.Y(n_259)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_218),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_196),
.B(n_217),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_209),
.B(n_202),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_219),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_250),
.B(n_219),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_241),
.Y(n_253)
);

BUFx4f_ASAP7_75t_SL g283 ( 
.A(n_253),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_236),
.B(n_213),
.C(n_201),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_260),
.B(n_265),
.C(n_266),
.Y(n_276)
);

OR2x2_ASAP7_75t_L g262 ( 
.A(n_244),
.B(n_220),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_262),
.A2(n_222),
.B(n_242),
.Y(n_284)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_263),
.Y(n_272)
);

AOI322xp5_ASAP7_75t_L g264 ( 
.A1(n_236),
.A2(n_210),
.A3(n_222),
.B1(n_223),
.B2(n_193),
.C1(n_199),
.C2(n_203),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_264),
.B(n_230),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_248),
.B(n_210),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_240),
.B(n_227),
.C(n_246),
.Y(n_266)
);

AND2x2_ASAP7_75t_L g282 ( 
.A(n_267),
.B(n_242),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_269),
.A2(n_237),
.B(n_239),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_270),
.B(n_230),
.Y(n_287)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_263),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_271),
.B(n_274),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_258),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_273),
.B(n_284),
.Y(n_289)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_252),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_254),
.B(n_243),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_275),
.B(n_278),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_260),
.B(n_229),
.C(n_235),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_277),
.B(n_266),
.Y(n_290)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_252),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_255),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_279),
.B(n_280),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_254),
.B(n_232),
.Y(n_280)
);

OA21x2_ASAP7_75t_SL g286 ( 
.A1(n_281),
.A2(n_268),
.B(n_259),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_282),
.A2(n_262),
.B1(n_256),
.B2(n_267),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_286),
.B(n_249),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_L g297 ( 
.A1(n_287),
.A2(n_288),
.B(n_280),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_290),
.B(n_282),
.C(n_247),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_283),
.B(n_251),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_292),
.B(n_296),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_SL g294 ( 
.A(n_276),
.B(n_265),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_294),
.B(n_295),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_276),
.B(n_259),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_283),
.B(n_253),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_297),
.A2(n_298),
.B1(n_303),
.B2(n_288),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_L g300 ( 
.A1(n_289),
.A2(n_270),
.B(n_284),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_300),
.B(n_289),
.Y(n_306)
);

AOI321xp33_ASAP7_75t_L g301 ( 
.A1(n_294),
.A2(n_245),
.A3(n_272),
.B1(n_275),
.B2(n_278),
.C(n_269),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_SL g308 ( 
.A(n_301),
.B(n_290),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_285),
.A2(n_256),
.B1(n_273),
.B2(n_293),
.Y(n_303)
);

AOI322xp5_ASAP7_75t_L g304 ( 
.A1(n_291),
.A2(n_282),
.A3(n_272),
.B1(n_283),
.B2(n_277),
.C1(n_262),
.C2(n_222),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_304),
.B(n_257),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_305),
.B(n_261),
.C(n_250),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_306),
.B(n_307),
.Y(n_312)
);

OAI21x1_ASAP7_75t_L g314 ( 
.A1(n_308),
.A2(n_299),
.B(n_300),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_302),
.A2(n_255),
.B1(n_295),
.B2(n_261),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_309),
.B(n_305),
.C(n_299),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_310),
.B(n_311),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_SL g313 ( 
.A(n_310),
.B(n_297),
.Y(n_313)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_313),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_314),
.B(n_306),
.C(n_211),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_315),
.B(n_309),
.Y(n_318)
);

HB1xp67_ASAP7_75t_L g317 ( 
.A(n_312),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_317),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_318),
.B(n_320),
.Y(n_321)
);

A2O1A1Ixp33_ASAP7_75t_L g322 ( 
.A1(n_319),
.A2(n_316),
.B(n_315),
.C(n_197),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_L g324 ( 
.A1(n_322),
.A2(n_317),
.B(n_257),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_L g326 ( 
.A1(n_324),
.A2(n_325),
.B(n_323),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_321),
.B(n_197),
.C(n_211),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_326),
.B(n_238),
.Y(n_327)
);


endmodule