module fake_jpeg_4709_n_53 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_53);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_53;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_37;
wire n_29;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx4_ASAP7_75t_L g7 ( 
.A(n_5),
.Y(n_7)
);

BUFx3_ASAP7_75t_L g8 ( 
.A(n_2),
.Y(n_8)
);

INVx2_ASAP7_75t_L g9 ( 
.A(n_0),
.Y(n_9)
);

INVx4_ASAP7_75t_L g10 ( 
.A(n_1),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_3),
.Y(n_11)
);

INVx6_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

INVx3_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

INVx8_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_17),
.B(n_18),
.Y(n_33)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

HB1xp67_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_19),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_14),
.B(n_0),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_20),
.B(n_21),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_16),
.B(n_2),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_7),
.B(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_7),
.B(n_3),
.Y(n_24)
);

INVx13_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

OAI22xp33_ASAP7_75t_SL g25 ( 
.A1(n_13),
.A2(n_4),
.B1(n_6),
.B2(n_9),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g30 ( 
.A(n_25),
.B(n_26),
.C(n_27),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_13),
.B(n_4),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_10),
.B(n_4),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g35 ( 
.A(n_27),
.B(n_10),
.C(n_11),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_35),
.B(n_22),
.Y(n_37)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_36),
.B(n_38),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_L g43 ( 
.A1(n_37),
.A2(n_39),
.B(n_30),
.Y(n_43)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_35),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_L g39 ( 
.A1(n_29),
.A2(n_23),
.B1(n_15),
.B2(n_18),
.Y(n_39)
);

XOR2xp5_ASAP7_75t_L g40 ( 
.A(n_38),
.B(n_30),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_40),
.B(n_28),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_37),
.B(n_17),
.C(n_28),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_41),
.B(n_43),
.Y(n_45)
);

XOR2xp5_ASAP7_75t_L g47 ( 
.A(n_44),
.B(n_46),
.Y(n_47)
);

OAI321xp33_ASAP7_75t_L g46 ( 
.A1(n_40),
.A2(n_31),
.A3(n_34),
.B1(n_29),
.B2(n_32),
.C(n_21),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_45),
.B(n_42),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_48),
.B(n_32),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_49),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_47),
.B(n_26),
.C(n_34),
.Y(n_50)
);

AO22x1_ASAP7_75t_L g52 ( 
.A1(n_51),
.A2(n_50),
.B1(n_47),
.B2(n_15),
.Y(n_52)
);

AOI21xp5_ASAP7_75t_L g53 ( 
.A1(n_52),
.A2(n_20),
.B(n_11),
.Y(n_53)
);


endmodule