module fake_jpeg_11233_n_186 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_186);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_186;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

BUFx10_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_7),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_4),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_10),
.B(n_8),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

INVx11_ASAP7_75t_SL g24 ( 
.A(n_5),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx4f_ASAP7_75t_SL g28 ( 
.A(n_1),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_12),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_9),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx12_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_8),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_35),
.B(n_36),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_17),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_37),
.B(n_40),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_17),
.B(n_11),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_38),
.B(n_43),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_39),
.Y(n_74)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_41),
.B(n_44),
.Y(n_97)
);

AOI21xp33_ASAP7_75t_L g42 ( 
.A1(n_14),
.A2(n_2),
.B(n_3),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_42),
.B(n_70),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_19),
.B(n_2),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_22),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_45),
.B(n_53),
.Y(n_102)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_13),
.Y(n_46)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_46),
.Y(n_77)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_13),
.Y(n_47)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_47),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_26),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_48),
.A2(n_61),
.B1(n_67),
.B2(n_25),
.Y(n_81)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_13),
.Y(n_49)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_49),
.Y(n_85)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_13),
.Y(n_50)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_50),
.Y(n_83)
);

BUFx2_ASAP7_75t_L g51 ( 
.A(n_13),
.Y(n_51)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_51),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_19),
.B(n_6),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_52),
.B(n_59),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_33),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_29),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_54),
.B(n_60),
.Y(n_103)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_21),
.Y(n_55)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_55),
.Y(n_90)
);

BUFx8_ASAP7_75t_L g56 ( 
.A(n_21),
.Y(n_56)
);

BUFx4f_ASAP7_75t_SL g94 ( 
.A(n_56),
.Y(n_94)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_21),
.Y(n_57)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_57),
.Y(n_93)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_29),
.Y(n_58)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_58),
.Y(n_96)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_21),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_28),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_26),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_61)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_28),
.Y(n_62)
);

CKINVDCx5p33_ASAP7_75t_R g89 ( 
.A(n_62),
.Y(n_89)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_24),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_63),
.A2(n_27),
.B1(n_32),
.B2(n_31),
.Y(n_80)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_28),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_64),
.B(n_66),
.Y(n_84)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_33),
.Y(n_65)
);

OR2x2_ASAP7_75t_SL g101 ( 
.A(n_65),
.B(n_69),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_20),
.B(n_30),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_14),
.A2(n_15),
.B1(n_32),
.B2(n_23),
.Y(n_67)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_33),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_68),
.B(n_56),
.Y(n_100)
);

NAND2xp33_ASAP7_75t_SL g69 ( 
.A(n_33),
.B(n_15),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_20),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_25),
.B(n_30),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_71),
.B(n_34),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_67),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_75),
.B(n_80),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_35),
.B(n_23),
.C(n_27),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_76),
.B(n_73),
.C(n_79),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_81),
.B(n_100),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_49),
.A2(n_31),
.B1(n_34),
.B2(n_51),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_82),
.A2(n_89),
.B1(n_96),
.B2(n_85),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_87),
.B(n_98),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_46),
.A2(n_50),
.B1(n_55),
.B2(n_64),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_88),
.B(n_94),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_65),
.A2(n_56),
.B(n_62),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_92),
.A2(n_89),
.B(n_100),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_39),
.A2(n_60),
.B1(n_68),
.B2(n_56),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_95),
.B(n_92),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_66),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_104),
.B(n_105),
.Y(n_133)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_99),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_108),
.B(n_110),
.Y(n_136)
);

MAJx2_ASAP7_75t_L g109 ( 
.A(n_101),
.B(n_84),
.C(n_91),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_109),
.A2(n_104),
.B(n_119),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_84),
.B(n_101),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_76),
.B(n_81),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_111),
.B(n_114),
.Y(n_138)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_74),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_112),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_113),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_86),
.Y(n_114)
);

INVx13_ASAP7_75t_L g115 ( 
.A(n_94),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_115),
.B(n_116),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_72),
.B(n_97),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_99),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_117),
.B(n_118),
.Y(n_142)
);

INVx13_ASAP7_75t_L g118 ( 
.A(n_94),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_120),
.A2(n_127),
.B1(n_119),
.B2(n_124),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_103),
.B(n_96),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_121),
.B(n_125),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_102),
.B(n_93),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_122),
.B(n_123),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_93),
.B(n_78),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_88),
.B(n_85),
.C(n_78),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_124),
.B(n_90),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_77),
.B(n_83),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_77),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_126),
.B(n_90),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_105),
.A2(n_74),
.B(n_83),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_131),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_132),
.B(n_140),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_135),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_111),
.A2(n_119),
.B1(n_110),
.B2(n_106),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_137),
.A2(n_127),
.B1(n_117),
.B2(n_126),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_114),
.B(n_107),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_141),
.B(n_108),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_143),
.A2(n_125),
.B(n_120),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_142),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_144),
.B(n_145),
.Y(n_161)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_135),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_140),
.B(n_109),
.C(n_121),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_146),
.B(n_133),
.C(n_138),
.Y(n_157)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_130),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_147),
.B(n_148),
.Y(n_156)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_128),
.Y(n_148)
);

NAND3xp33_ASAP7_75t_L g159 ( 
.A(n_149),
.B(n_139),
.C(n_136),
.Y(n_159)
);

MAJx2_ASAP7_75t_L g163 ( 
.A(n_150),
.B(n_133),
.C(n_134),
.Y(n_163)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_128),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_154),
.B(n_112),
.Y(n_164)
);

AOI221xp5_ASAP7_75t_L g162 ( 
.A1(n_155),
.A2(n_137),
.B1(n_134),
.B2(n_133),
.C(n_129),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_157),
.B(n_163),
.C(n_146),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_151),
.A2(n_131),
.B(n_143),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_158),
.A2(n_162),
.B(n_155),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_159),
.B(n_164),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_152),
.Y(n_160)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_160),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_166),
.B(n_170),
.C(n_158),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_168),
.B(n_150),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_161),
.A2(n_151),
.B1(n_156),
.B2(n_152),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_169),
.B(n_153),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_157),
.B(n_153),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_171),
.B(n_174),
.C(n_166),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_172),
.B(n_173),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_170),
.B(n_163),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_176),
.B(n_168),
.C(n_165),
.Y(n_179)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_174),
.Y(n_177)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_177),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_172),
.B(n_167),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_178),
.B(n_165),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_179),
.B(n_181),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_180),
.A2(n_175),
.B(n_176),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_182),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_184),
.A2(n_183),
.B(n_129),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_185),
.B(n_115),
.Y(n_186)
);


endmodule