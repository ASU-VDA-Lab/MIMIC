module real_aes_6590_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_369;
wire n_343;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_725;
wire n_310;
wire n_504;
wire n_455;
wire n_164;
wire n_671;
wire n_231;
wire n_659;
wire n_547;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_363;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_720;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND3xp33_ASAP7_75t_SL g111 ( .A(n_0), .B(n_112), .C(n_113), .Y(n_111) );
INVx1_ASAP7_75t_L g443 ( .A(n_0), .Y(n_443) );
A2O1A1Ixp33_ASAP7_75t_L g189 ( .A1(n_1), .A2(n_148), .B(n_153), .C(n_190), .Y(n_189) );
AOI21xp5_ASAP7_75t_L g212 ( .A1(n_2), .A2(n_143), .B(n_213), .Y(n_212) );
INVx1_ASAP7_75t_L g461 ( .A(n_3), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_4), .B(n_167), .Y(n_220) );
AOI22xp5_ASAP7_75t_L g722 ( .A1(n_5), .A2(n_15), .B1(n_723), .B2(n_724), .Y(n_722) );
CKINVDCx20_ASAP7_75t_R g724 ( .A(n_5), .Y(n_724) );
AOI21xp33_ASAP7_75t_L g478 ( .A1(n_6), .A2(n_143), .B(n_479), .Y(n_478) );
AND2x6_ASAP7_75t_L g148 ( .A(n_7), .B(n_149), .Y(n_148) );
INVx1_ASAP7_75t_L g177 ( .A(n_8), .Y(n_177) );
INVx1_ASAP7_75t_L g109 ( .A(n_9), .Y(n_109) );
NOR2xp33_ASAP7_75t_L g444 ( .A(n_9), .B(n_43), .Y(n_444) );
AOI21xp5_ASAP7_75t_L g538 ( .A1(n_10), .A2(n_255), .B(n_539), .Y(n_538) );
NAND2xp5_ASAP7_75t_SL g194 ( .A(n_11), .B(n_158), .Y(n_194) );
INVx1_ASAP7_75t_L g483 ( .A(n_12), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_13), .B(n_157), .Y(n_531) );
INVx1_ASAP7_75t_L g141 ( .A(n_14), .Y(n_141) );
CKINVDCx20_ASAP7_75t_R g723 ( .A(n_15), .Y(n_723) );
INVx1_ASAP7_75t_L g543 ( .A(n_16), .Y(n_543) );
A2O1A1Ixp33_ASAP7_75t_L g202 ( .A1(n_17), .A2(n_178), .B(n_203), .C(n_205), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_18), .B(n_167), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_19), .B(n_472), .Y(n_522) );
NAND2xp5_ASAP7_75t_SL g509 ( .A(n_20), .B(n_143), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_21), .B(n_263), .Y(n_262) );
A2O1A1Ixp33_ASAP7_75t_L g156 ( .A1(n_22), .A2(n_157), .B(n_159), .C(n_163), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_23), .B(n_167), .Y(n_475) );
NAND2xp5_ASAP7_75t_SL g227 ( .A(n_24), .B(n_158), .Y(n_227) );
A2O1A1Ixp33_ASAP7_75t_L g541 ( .A1(n_25), .A2(n_161), .B(n_205), .C(n_542), .Y(n_541) );
NAND2xp5_ASAP7_75t_SL g239 ( .A(n_26), .B(n_158), .Y(n_239) );
CKINVDCx16_ASAP7_75t_R g223 ( .A(n_27), .Y(n_223) );
INVx1_ASAP7_75t_L g237 ( .A(n_28), .Y(n_237) );
BUFx6f_ASAP7_75t_L g147 ( .A(n_29), .Y(n_147) );
CKINVDCx20_ASAP7_75t_R g187 ( .A(n_30), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_31), .B(n_158), .Y(n_462) );
INVx1_ASAP7_75t_L g260 ( .A(n_32), .Y(n_260) );
INVx1_ASAP7_75t_L g496 ( .A(n_33), .Y(n_496) );
NAND2xp5_ASAP7_75t_SL g445 ( .A(n_34), .B(n_446), .Y(n_445) );
INVx2_ASAP7_75t_L g146 ( .A(n_35), .Y(n_146) );
CKINVDCx20_ASAP7_75t_R g197 ( .A(n_36), .Y(n_197) );
A2O1A1Ixp33_ASAP7_75t_L g215 ( .A1(n_37), .A2(n_157), .B(n_216), .C(n_218), .Y(n_215) );
INVxp67_ASAP7_75t_L g261 ( .A(n_38), .Y(n_261) );
CKINVDCx14_ASAP7_75t_R g214 ( .A(n_39), .Y(n_214) );
A2O1A1Ixp33_ASAP7_75t_L g235 ( .A1(n_40), .A2(n_153), .B(n_236), .C(n_242), .Y(n_235) );
A2O1A1Ixp33_ASAP7_75t_L g510 ( .A1(n_41), .A2(n_148), .B(n_153), .C(n_511), .Y(n_510) );
OAI22xp5_ASAP7_75t_SL g125 ( .A1(n_42), .A2(n_92), .B1(n_126), .B2(n_127), .Y(n_125) );
CKINVDCx20_ASAP7_75t_R g127 ( .A(n_42), .Y(n_127) );
NAND2xp5_ASAP7_75t_L g108 ( .A(n_43), .B(n_109), .Y(n_108) );
INVx1_ASAP7_75t_L g495 ( .A(n_44), .Y(n_495) );
A2O1A1Ixp33_ASAP7_75t_L g174 ( .A1(n_45), .A2(n_175), .B(n_176), .C(n_179), .Y(n_174) );
NAND2xp5_ASAP7_75t_SL g521 ( .A(n_46), .B(n_158), .Y(n_521) );
AOI22xp33_ASAP7_75t_L g103 ( .A1(n_47), .A2(n_104), .B1(n_116), .B2(n_735), .Y(n_103) );
AOI22xp33_ASAP7_75t_L g123 ( .A1(n_48), .A2(n_124), .B1(n_436), .B2(n_437), .Y(n_123) );
CKINVDCx20_ASAP7_75t_R g436 ( .A(n_48), .Y(n_436) );
CKINVDCx20_ASAP7_75t_R g244 ( .A(n_49), .Y(n_244) );
CKINVDCx20_ASAP7_75t_R g257 ( .A(n_50), .Y(n_257) );
INVx1_ASAP7_75t_L g151 ( .A(n_51), .Y(n_151) );
CKINVDCx16_ASAP7_75t_R g497 ( .A(n_52), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_53), .B(n_143), .Y(n_533) );
AOI22xp5_ASAP7_75t_L g493 ( .A1(n_54), .A2(n_153), .B1(n_163), .B2(n_494), .Y(n_493) );
CKINVDCx20_ASAP7_75t_R g515 ( .A(n_55), .Y(n_515) );
CKINVDCx16_ASAP7_75t_R g458 ( .A(n_56), .Y(n_458) );
CKINVDCx14_ASAP7_75t_R g173 ( .A(n_57), .Y(n_173) );
A2O1A1Ixp33_ASAP7_75t_L g481 ( .A1(n_58), .A2(n_175), .B(n_218), .C(n_482), .Y(n_481) );
CKINVDCx20_ASAP7_75t_R g524 ( .A(n_59), .Y(n_524) );
INVx1_ASAP7_75t_L g480 ( .A(n_60), .Y(n_480) );
INVx1_ASAP7_75t_L g149 ( .A(n_61), .Y(n_149) );
INVx1_ASAP7_75t_L g140 ( .A(n_62), .Y(n_140) );
INVx1_ASAP7_75t_SL g217 ( .A(n_63), .Y(n_217) );
CKINVDCx20_ASAP7_75t_R g121 ( .A(n_64), .Y(n_121) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_65), .B(n_167), .Y(n_166) );
INVx1_ASAP7_75t_L g226 ( .A(n_66), .Y(n_226) );
A2O1A1Ixp33_ASAP7_75t_SL g471 ( .A1(n_67), .A2(n_218), .B(n_472), .C(n_473), .Y(n_471) );
INVxp67_ASAP7_75t_L g474 ( .A(n_68), .Y(n_474) );
INVx1_ASAP7_75t_L g115 ( .A(n_69), .Y(n_115) );
AOI21xp5_ASAP7_75t_L g171 ( .A1(n_70), .A2(n_143), .B(n_172), .Y(n_171) );
CKINVDCx20_ASAP7_75t_R g230 ( .A(n_71), .Y(n_230) );
AOI21xp5_ASAP7_75t_L g199 ( .A1(n_72), .A2(n_143), .B(n_200), .Y(n_199) );
CKINVDCx20_ASAP7_75t_R g499 ( .A(n_73), .Y(n_499) );
INVx1_ASAP7_75t_L g518 ( .A(n_74), .Y(n_518) );
AOI21xp5_ASAP7_75t_L g254 ( .A1(n_75), .A2(n_255), .B(n_256), .Y(n_254) );
INVx1_ASAP7_75t_L g201 ( .A(n_76), .Y(n_201) );
CKINVDCx16_ASAP7_75t_R g234 ( .A(n_77), .Y(n_234) );
AOI222xp33_ASAP7_75t_L g448 ( .A1(n_78), .A2(n_449), .B1(n_720), .B2(n_726), .C1(n_730), .C2(n_731), .Y(n_448) );
A2O1A1Ixp33_ASAP7_75t_L g519 ( .A1(n_79), .A2(n_148), .B(n_153), .C(n_520), .Y(n_519) );
AOI21xp5_ASAP7_75t_L g142 ( .A1(n_80), .A2(n_143), .B(n_150), .Y(n_142) );
INVx1_ASAP7_75t_L g204 ( .A(n_81), .Y(n_204) );
NAND2xp5_ASAP7_75t_SL g512 ( .A(n_82), .B(n_238), .Y(n_512) );
INVx2_ASAP7_75t_L g138 ( .A(n_83), .Y(n_138) );
INVx1_ASAP7_75t_L g191 ( .A(n_84), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_85), .B(n_472), .Y(n_513) );
A2O1A1Ixp33_ASAP7_75t_L g459 ( .A1(n_86), .A2(n_148), .B(n_153), .C(n_460), .Y(n_459) );
INVx2_ASAP7_75t_L g112 ( .A(n_87), .Y(n_112) );
OR2x2_ASAP7_75t_L g440 ( .A(n_87), .B(n_441), .Y(n_440) );
OR2x2_ASAP7_75t_L g719 ( .A(n_87), .B(n_442), .Y(n_719) );
A2O1A1Ixp33_ASAP7_75t_L g224 ( .A1(n_88), .A2(n_153), .B(n_225), .C(n_228), .Y(n_224) );
OAI22xp5_ASAP7_75t_SL g720 ( .A1(n_89), .A2(n_721), .B1(n_722), .B2(n_725), .Y(n_720) );
CKINVDCx20_ASAP7_75t_R g725 ( .A(n_89), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_90), .B(n_170), .Y(n_484) );
CKINVDCx20_ASAP7_75t_R g465 ( .A(n_91), .Y(n_465) );
CKINVDCx20_ASAP7_75t_R g126 ( .A(n_92), .Y(n_126) );
A2O1A1Ixp33_ASAP7_75t_L g528 ( .A1(n_93), .A2(n_148), .B(n_153), .C(n_529), .Y(n_528) );
CKINVDCx20_ASAP7_75t_R g535 ( .A(n_94), .Y(n_535) );
INVx1_ASAP7_75t_L g470 ( .A(n_95), .Y(n_470) );
CKINVDCx16_ASAP7_75t_R g540 ( .A(n_96), .Y(n_540) );
NAND2xp5_ASAP7_75t_SL g530 ( .A(n_97), .B(n_238), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_98), .B(n_136), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_99), .B(n_136), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g114 ( .A(n_100), .B(n_115), .Y(n_114) );
INVx2_ASAP7_75t_L g160 ( .A(n_101), .Y(n_160) );
AOI21xp5_ASAP7_75t_L g468 ( .A1(n_102), .A2(n_143), .B(n_469), .Y(n_468) );
INVx1_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
INVx2_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
INVx2_ASAP7_75t_SL g735 ( .A(n_106), .Y(n_735) );
AND2x2_ASAP7_75t_L g106 ( .A(n_107), .B(n_110), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
INVx1_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
OR2x2_ASAP7_75t_L g718 ( .A(n_112), .B(n_442), .Y(n_718) );
NOR2x2_ASAP7_75t_L g733 ( .A(n_112), .B(n_441), .Y(n_733) );
INVx1_ASAP7_75t_SL g113 ( .A(n_114), .Y(n_113) );
AO21x1_ASAP7_75t_L g116 ( .A1(n_117), .A2(n_122), .B(n_447), .Y(n_116) );
INVx1_ASAP7_75t_SL g117 ( .A(n_118), .Y(n_117) );
BUFx2_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVx2_ASAP7_75t_SL g734 ( .A(n_119), .Y(n_734) );
BUFx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx2_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
OAI21xp5_ASAP7_75t_SL g122 ( .A1(n_123), .A2(n_438), .B(n_445), .Y(n_122) );
INVx1_ASAP7_75t_L g437 ( .A(n_124), .Y(n_437) );
AOI22xp5_ASAP7_75t_L g124 ( .A1(n_125), .A2(n_128), .B1(n_434), .B2(n_435), .Y(n_124) );
CKINVDCx20_ASAP7_75t_R g434 ( .A(n_125), .Y(n_434) );
OAI22xp5_ASAP7_75t_L g726 ( .A1(n_128), .A2(n_718), .B1(n_727), .B2(n_728), .Y(n_726) );
BUFx2_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
INVx1_ASAP7_75t_L g435 ( .A(n_129), .Y(n_435) );
AND2x2_ASAP7_75t_L g129 ( .A(n_130), .B(n_360), .Y(n_129) );
NOR4xp25_ASAP7_75t_L g130 ( .A(n_131), .B(n_302), .C(n_332), .D(n_342), .Y(n_130) );
OAI211xp5_ASAP7_75t_L g131 ( .A1(n_132), .A2(n_207), .B(n_265), .C(n_292), .Y(n_131) );
OAI222xp33_ASAP7_75t_L g387 ( .A1(n_132), .A2(n_307), .B1(n_388), .B2(n_389), .C1(n_390), .C2(n_391), .Y(n_387) );
OR2x2_ASAP7_75t_L g132 ( .A(n_133), .B(n_182), .Y(n_132) );
AOI33xp33_ASAP7_75t_L g313 ( .A1(n_133), .A2(n_300), .A3(n_301), .B1(n_314), .B2(n_319), .B3(n_321), .Y(n_313) );
OAI211xp5_ASAP7_75t_SL g370 ( .A1(n_133), .A2(n_371), .B(n_373), .C(n_375), .Y(n_370) );
OR2x2_ASAP7_75t_L g386 ( .A(n_133), .B(n_372), .Y(n_386) );
INVx1_ASAP7_75t_L g419 ( .A(n_133), .Y(n_419) );
OR2x2_ASAP7_75t_L g133 ( .A(n_134), .B(n_169), .Y(n_133) );
INVx2_ASAP7_75t_L g296 ( .A(n_134), .Y(n_296) );
AND2x2_ASAP7_75t_L g312 ( .A(n_134), .B(n_198), .Y(n_312) );
HB1xp67_ASAP7_75t_L g347 ( .A(n_134), .Y(n_347) );
AND2x2_ASAP7_75t_L g376 ( .A(n_134), .B(n_169), .Y(n_376) );
OA21x2_ASAP7_75t_L g134 ( .A1(n_135), .A2(n_142), .B(n_166), .Y(n_134) );
OA21x2_ASAP7_75t_L g198 ( .A1(n_135), .A2(n_199), .B(n_206), .Y(n_198) );
OA21x2_ASAP7_75t_L g211 ( .A1(n_135), .A2(n_212), .B(n_220), .Y(n_211) );
HB1xp67_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
INVx4_ASAP7_75t_L g168 ( .A(n_136), .Y(n_168) );
OA21x2_ASAP7_75t_L g467 ( .A1(n_136), .A2(n_468), .B(n_475), .Y(n_467) );
BUFx6f_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
INVx1_ASAP7_75t_L g253 ( .A(n_137), .Y(n_253) );
AND2x2_ASAP7_75t_L g137 ( .A(n_138), .B(n_139), .Y(n_137) );
AND2x2_ASAP7_75t_SL g170 ( .A(n_138), .B(n_139), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g139 ( .A(n_140), .B(n_141), .Y(n_139) );
BUFx2_ASAP7_75t_L g255 ( .A(n_143), .Y(n_255) );
AND2x4_ASAP7_75t_L g143 ( .A(n_144), .B(n_148), .Y(n_143) );
NAND2x1p5_ASAP7_75t_L g188 ( .A(n_144), .B(n_148), .Y(n_188) );
AND2x2_ASAP7_75t_L g144 ( .A(n_145), .B(n_147), .Y(n_144) );
INVx1_ASAP7_75t_L g241 ( .A(n_145), .Y(n_241) );
INVx1_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx2_ASAP7_75t_L g154 ( .A(n_146), .Y(n_154) );
INVx1_ASAP7_75t_L g164 ( .A(n_146), .Y(n_164) );
INVx1_ASAP7_75t_L g155 ( .A(n_147), .Y(n_155) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_147), .Y(n_158) );
BUFx6f_ASAP7_75t_L g162 ( .A(n_147), .Y(n_162) );
INVx3_ASAP7_75t_L g178 ( .A(n_147), .Y(n_178) );
INVx1_ASAP7_75t_L g472 ( .A(n_147), .Y(n_472) );
INVx4_ASAP7_75t_SL g165 ( .A(n_148), .Y(n_165) );
BUFx3_ASAP7_75t_L g242 ( .A(n_148), .Y(n_242) );
O2A1O1Ixp33_ASAP7_75t_SL g150 ( .A1(n_151), .A2(n_152), .B(n_156), .C(n_165), .Y(n_150) );
O2A1O1Ixp33_ASAP7_75t_SL g172 ( .A1(n_152), .A2(n_165), .B(n_173), .C(n_174), .Y(n_172) );
O2A1O1Ixp33_ASAP7_75t_SL g200 ( .A1(n_152), .A2(n_165), .B(n_201), .C(n_202), .Y(n_200) );
O2A1O1Ixp33_ASAP7_75t_L g213 ( .A1(n_152), .A2(n_165), .B(n_214), .C(n_215), .Y(n_213) );
O2A1O1Ixp33_ASAP7_75t_SL g256 ( .A1(n_152), .A2(n_165), .B(n_257), .C(n_258), .Y(n_256) );
O2A1O1Ixp33_ASAP7_75t_L g469 ( .A1(n_152), .A2(n_165), .B(n_470), .C(n_471), .Y(n_469) );
O2A1O1Ixp33_ASAP7_75t_L g479 ( .A1(n_152), .A2(n_165), .B(n_480), .C(n_481), .Y(n_479) );
O2A1O1Ixp33_ASAP7_75t_L g539 ( .A1(n_152), .A2(n_165), .B(n_540), .C(n_541), .Y(n_539) );
INVx5_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
AND2x6_ASAP7_75t_L g153 ( .A(n_154), .B(n_155), .Y(n_153) );
BUFx3_ASAP7_75t_L g180 ( .A(n_154), .Y(n_180) );
BUFx6f_ASAP7_75t_L g219 ( .A(n_154), .Y(n_219) );
NOR2xp33_ASAP7_75t_L g216 ( .A(n_157), .B(n_217), .Y(n_216) );
INVx4_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx2_ASAP7_75t_L g175 ( .A(n_158), .Y(n_175) );
NOR2xp33_ASAP7_75t_L g159 ( .A(n_160), .B(n_161), .Y(n_159) );
NOR2xp33_ASAP7_75t_L g203 ( .A(n_161), .B(n_204), .Y(n_203) );
OAI22xp33_ASAP7_75t_L g259 ( .A1(n_161), .A2(n_238), .B1(n_260), .B2(n_261), .Y(n_259) );
NOR2xp33_ASAP7_75t_L g542 ( .A(n_161), .B(n_543), .Y(n_542) );
INVx4_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
INVx2_ASAP7_75t_L g193 ( .A(n_162), .Y(n_193) );
OAI22xp5_ASAP7_75t_SL g494 ( .A1(n_162), .A2(n_193), .B1(n_495), .B2(n_496), .Y(n_494) );
INVx2_ASAP7_75t_L g463 ( .A(n_163), .Y(n_463) );
INVx3_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVx1_ASAP7_75t_L g228 ( .A(n_165), .Y(n_228) );
OAI22xp33_ASAP7_75t_L g492 ( .A1(n_165), .A2(n_188), .B1(n_493), .B2(n_497), .Y(n_492) );
OA21x2_ASAP7_75t_L g477 ( .A1(n_167), .A2(n_478), .B(n_484), .Y(n_477) );
INVx3_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
NOR2xp33_ASAP7_75t_L g196 ( .A(n_168), .B(n_197), .Y(n_196) );
AO21x2_ASAP7_75t_L g221 ( .A1(n_168), .A2(n_222), .B(n_229), .Y(n_221) );
NOR2xp33_ASAP7_75t_L g243 ( .A(n_168), .B(n_244), .Y(n_243) );
NOR2xp33_ASAP7_75t_SL g514 ( .A(n_168), .B(n_515), .Y(n_514) );
INVx2_ASAP7_75t_L g276 ( .A(n_169), .Y(n_276) );
BUFx3_ASAP7_75t_L g284 ( .A(n_169), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_169), .B(n_287), .Y(n_286) );
AND2x2_ASAP7_75t_L g295 ( .A(n_169), .B(n_296), .Y(n_295) );
NOR2xp33_ASAP7_75t_L g324 ( .A(n_169), .B(n_183), .Y(n_324) );
AND2x2_ASAP7_75t_L g393 ( .A(n_169), .B(n_327), .Y(n_393) );
OA21x2_ASAP7_75t_L g169 ( .A1(n_170), .A2(n_171), .B(n_181), .Y(n_169) );
INVx1_ASAP7_75t_L g185 ( .A(n_170), .Y(n_185) );
INVx2_ASAP7_75t_L g231 ( .A(n_170), .Y(n_231) );
O2A1O1Ixp33_ASAP7_75t_L g233 ( .A1(n_170), .A2(n_188), .B(n_234), .C(n_235), .Y(n_233) );
OA21x2_ASAP7_75t_L g537 ( .A1(n_170), .A2(n_538), .B(n_544), .Y(n_537) );
NOR2xp33_ASAP7_75t_L g176 ( .A(n_177), .B(n_178), .Y(n_176) );
INVx5_ASAP7_75t_L g238 ( .A(n_178), .Y(n_238) );
NOR2xp33_ASAP7_75t_L g473 ( .A(n_178), .B(n_474), .Y(n_473) );
NOR2xp33_ASAP7_75t_L g482 ( .A(n_178), .B(n_483), .Y(n_482) );
INVx2_ASAP7_75t_L g195 ( .A(n_179), .Y(n_195) );
INVx2_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
INVx1_ASAP7_75t_L g205 ( .A(n_180), .Y(n_205) );
INVx2_ASAP7_75t_SL g287 ( .A(n_182), .Y(n_287) );
OR2x2_ASAP7_75t_L g182 ( .A(n_183), .B(n_198), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_183), .B(n_276), .Y(n_275) );
INVx1_ASAP7_75t_L g329 ( .A(n_183), .Y(n_329) );
AND2x2_ASAP7_75t_L g340 ( .A(n_183), .B(n_296), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_183), .B(n_325), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_183), .B(n_327), .Y(n_372) );
AND2x2_ASAP7_75t_L g431 ( .A(n_183), .B(n_376), .Y(n_431) );
INVx4_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
AND2x2_ASAP7_75t_L g301 ( .A(n_184), .B(n_198), .Y(n_301) );
AND2x2_ASAP7_75t_L g311 ( .A(n_184), .B(n_312), .Y(n_311) );
BUFx3_ASAP7_75t_L g333 ( .A(n_184), .Y(n_333) );
AND3x2_ASAP7_75t_L g392 ( .A(n_184), .B(n_393), .C(n_394), .Y(n_392) );
AO21x2_ASAP7_75t_L g184 ( .A1(n_185), .A2(n_186), .B(n_196), .Y(n_184) );
NOR2xp33_ASAP7_75t_L g464 ( .A(n_185), .B(n_465), .Y(n_464) );
NOR2xp33_ASAP7_75t_L g523 ( .A(n_185), .B(n_524), .Y(n_523) );
NOR2xp33_ASAP7_75t_L g534 ( .A(n_185), .B(n_535), .Y(n_534) );
OAI21xp5_ASAP7_75t_L g186 ( .A1(n_187), .A2(n_188), .B(n_189), .Y(n_186) );
OAI21xp5_ASAP7_75t_L g222 ( .A1(n_188), .A2(n_223), .B(n_224), .Y(n_222) );
OAI21xp5_ASAP7_75t_L g457 ( .A1(n_188), .A2(n_458), .B(n_459), .Y(n_457) );
OAI21xp5_ASAP7_75t_L g517 ( .A1(n_188), .A2(n_518), .B(n_519), .Y(n_517) );
O2A1O1Ixp5_ASAP7_75t_L g190 ( .A1(n_191), .A2(n_192), .B(n_194), .C(n_195), .Y(n_190) );
O2A1O1Ixp33_ASAP7_75t_L g225 ( .A1(n_192), .A2(n_195), .B(n_226), .C(n_227), .Y(n_225) );
INVx2_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
AOI21xp5_ASAP7_75t_L g511 ( .A1(n_195), .A2(n_512), .B(n_513), .Y(n_511) );
AOI21xp5_ASAP7_75t_L g520 ( .A1(n_195), .A2(n_521), .B(n_522), .Y(n_520) );
HB1xp67_ASAP7_75t_L g283 ( .A(n_198), .Y(n_283) );
INVx1_ASAP7_75t_SL g327 ( .A(n_198), .Y(n_327) );
NAND3xp33_ASAP7_75t_L g339 ( .A(n_198), .B(n_276), .C(n_340), .Y(n_339) );
NOR2xp33_ASAP7_75t_L g207 ( .A(n_208), .B(n_245), .Y(n_207) );
A2O1A1Ixp33_ASAP7_75t_L g362 ( .A1(n_208), .A2(n_311), .B(n_363), .C(n_365), .Y(n_362) );
INVx1_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
NAND2xp5_ASAP7_75t_SL g209 ( .A(n_210), .B(n_232), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_210), .B(n_369), .Y(n_368) );
INVx2_ASAP7_75t_SL g379 ( .A(n_210), .Y(n_379) );
AND2x2_ASAP7_75t_L g400 ( .A(n_210), .B(n_247), .Y(n_400) );
NOR2xp33_ASAP7_75t_L g428 ( .A(n_210), .B(n_309), .Y(n_428) );
AND2x2_ASAP7_75t_L g210 ( .A(n_211), .B(n_221), .Y(n_210) );
AND2x2_ASAP7_75t_L g273 ( .A(n_211), .B(n_264), .Y(n_273) );
INVx2_ASAP7_75t_L g280 ( .A(n_211), .Y(n_280) );
AND2x2_ASAP7_75t_L g300 ( .A(n_211), .B(n_247), .Y(n_300) );
AND2x2_ASAP7_75t_L g350 ( .A(n_211), .B(n_232), .Y(n_350) );
INVx1_ASAP7_75t_L g354 ( .A(n_211), .Y(n_354) );
INVx3_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
HB1xp67_ASAP7_75t_L g532 ( .A(n_219), .Y(n_532) );
INVx2_ASAP7_75t_SL g264 ( .A(n_221), .Y(n_264) );
BUFx2_ASAP7_75t_L g290 ( .A(n_221), .Y(n_290) );
AND2x2_ASAP7_75t_L g417 ( .A(n_221), .B(n_232), .Y(n_417) );
NOR2xp33_ASAP7_75t_L g229 ( .A(n_230), .B(n_231), .Y(n_229) );
INVx1_ASAP7_75t_L g263 ( .A(n_231), .Y(n_263) );
AO21x2_ASAP7_75t_L g526 ( .A1(n_231), .A2(n_527), .B(n_534), .Y(n_526) );
INVx3_ASAP7_75t_SL g247 ( .A(n_232), .Y(n_247) );
AND2x2_ASAP7_75t_L g272 ( .A(n_232), .B(n_273), .Y(n_272) );
AND2x4_ASAP7_75t_L g279 ( .A(n_232), .B(n_280), .Y(n_279) );
OR2x2_ASAP7_75t_L g309 ( .A(n_232), .B(n_269), .Y(n_309) );
OR2x2_ASAP7_75t_L g318 ( .A(n_232), .B(n_264), .Y(n_318) );
HB1xp67_ASAP7_75t_L g336 ( .A(n_232), .Y(n_336) );
AND2x2_ASAP7_75t_L g341 ( .A(n_232), .B(n_294), .Y(n_341) );
AND2x2_ASAP7_75t_L g369 ( .A(n_232), .B(n_249), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_232), .B(n_405), .Y(n_404) );
OR2x2_ASAP7_75t_L g407 ( .A(n_232), .B(n_248), .Y(n_407) );
OR2x6_ASAP7_75t_L g232 ( .A(n_233), .B(n_243), .Y(n_232) );
O2A1O1Ixp33_ASAP7_75t_L g236 ( .A1(n_237), .A2(n_238), .B(n_239), .C(n_240), .Y(n_236) );
O2A1O1Ixp33_ASAP7_75t_L g460 ( .A1(n_238), .A2(n_461), .B(n_462), .C(n_463), .Y(n_460) );
INVx2_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
NAND2xp5_ASAP7_75t_SL g258 ( .A(n_241), .B(n_259), .Y(n_258) );
INVx1_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
OR2x2_ASAP7_75t_L g246 ( .A(n_247), .B(n_248), .Y(n_246) );
AND2x2_ASAP7_75t_L g331 ( .A(n_247), .B(n_280), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_247), .B(n_273), .Y(n_359) );
AND2x2_ASAP7_75t_L g377 ( .A(n_247), .B(n_294), .Y(n_377) );
OR2x2_ASAP7_75t_L g248 ( .A(n_249), .B(n_264), .Y(n_248) );
AND2x2_ASAP7_75t_L g278 ( .A(n_249), .B(n_264), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_249), .B(n_307), .Y(n_306) );
BUFx3_ASAP7_75t_L g316 ( .A(n_249), .Y(n_316) );
OR2x2_ASAP7_75t_L g364 ( .A(n_249), .B(n_284), .Y(n_364) );
OA21x2_ASAP7_75t_L g249 ( .A1(n_250), .A2(n_254), .B(n_262), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
AO21x2_ASAP7_75t_L g269 ( .A1(n_251), .A2(n_270), .B(n_271), .Y(n_269) );
AO21x2_ASAP7_75t_L g516 ( .A1(n_251), .A2(n_517), .B(n_523), .Y(n_516) );
INVx1_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
AOI21xp5_ASAP7_75t_SL g508 ( .A1(n_252), .A2(n_509), .B(n_510), .Y(n_508) );
INVx2_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
AO21x2_ASAP7_75t_L g456 ( .A1(n_253), .A2(n_457), .B(n_464), .Y(n_456) );
AO21x2_ASAP7_75t_L g491 ( .A1(n_253), .A2(n_492), .B(n_498), .Y(n_491) );
NOR2xp33_ASAP7_75t_L g498 ( .A(n_253), .B(n_499), .Y(n_498) );
INVx1_ASAP7_75t_L g270 ( .A(n_254), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_262), .Y(n_271) );
AND2x2_ASAP7_75t_L g299 ( .A(n_264), .B(n_269), .Y(n_299) );
INVx1_ASAP7_75t_L g307 ( .A(n_264), .Y(n_307) );
AND2x2_ASAP7_75t_L g402 ( .A(n_264), .B(n_280), .Y(n_402) );
AOI222xp33_ASAP7_75t_L g265 ( .A1(n_266), .A2(n_274), .B1(n_277), .B2(n_281), .C1(n_285), .C2(n_288), .Y(n_265) );
INVx1_ASAP7_75t_L g397 ( .A(n_266), .Y(n_397) );
AND2x2_ASAP7_75t_L g266 ( .A(n_267), .B(n_272), .Y(n_266) );
AND2x2_ASAP7_75t_L g293 ( .A(n_267), .B(n_294), .Y(n_293) );
AND2x2_ASAP7_75t_L g304 ( .A(n_267), .B(n_273), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_267), .B(n_295), .Y(n_320) );
OAI222xp33_ASAP7_75t_L g342 ( .A1(n_267), .A2(n_343), .B1(n_348), .B2(n_349), .C1(n_357), .C2(n_359), .Y(n_342) );
INVx2_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
INVx1_ASAP7_75t_SL g268 ( .A(n_269), .Y(n_268) );
AND2x2_ASAP7_75t_L g330 ( .A(n_269), .B(n_331), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_269), .B(n_350), .Y(n_390) );
AND2x2_ASAP7_75t_L g401 ( .A(n_269), .B(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g409 ( .A(n_272), .Y(n_409) );
NAND2xp5_ASAP7_75t_SL g388 ( .A(n_274), .B(n_325), .Y(n_388) );
INVx1_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
NOR2xp33_ASAP7_75t_L g328 ( .A(n_276), .B(n_329), .Y(n_328) );
AND2x2_ASAP7_75t_L g346 ( .A(n_276), .B(n_347), .Y(n_346) );
AND2x2_ASAP7_75t_L g277 ( .A(n_278), .B(n_279), .Y(n_277) );
INVx3_ASAP7_75t_L g291 ( .A(n_279), .Y(n_291) );
O2A1O1Ixp33_ASAP7_75t_L g381 ( .A1(n_279), .A2(n_382), .B(n_385), .C(n_387), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_279), .B(n_316), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_279), .B(n_299), .Y(n_421) );
AND2x2_ASAP7_75t_L g294 ( .A(n_280), .B(n_290), .Y(n_294) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_283), .B(n_284), .Y(n_282) );
INVx1_ASAP7_75t_L g321 ( .A(n_283), .Y(n_321) );
NAND2xp5_ASAP7_75t_SL g310 ( .A(n_284), .B(n_311), .Y(n_310) );
OR2x2_ASAP7_75t_L g373 ( .A(n_284), .B(n_374), .Y(n_373) );
AND2x2_ASAP7_75t_L g412 ( .A(n_284), .B(n_312), .Y(n_412) );
INVx1_ASAP7_75t_L g424 ( .A(n_284), .Y(n_424) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_287), .B(n_426), .Y(n_425) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
OR2x2_ASAP7_75t_L g289 ( .A(n_290), .B(n_291), .Y(n_289) );
INVx1_ASAP7_75t_L g405 ( .A(n_290), .Y(n_405) );
A2O1A1Ixp33_ASAP7_75t_SL g292 ( .A1(n_293), .A2(n_295), .B(n_297), .C(n_301), .Y(n_292) );
AOI22xp33_ASAP7_75t_L g337 ( .A1(n_293), .A2(n_323), .B1(n_338), .B2(n_341), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_294), .B(n_308), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_294), .B(n_316), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_295), .B(n_353), .Y(n_352) );
INVx1_ASAP7_75t_SL g358 ( .A(n_295), .Y(n_358) );
AND2x2_ASAP7_75t_L g365 ( .A(n_295), .B(n_345), .Y(n_365) );
INVx2_ASAP7_75t_L g326 ( .A(n_296), .Y(n_326) );
INVxp67_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_299), .B(n_300), .Y(n_298) );
NOR4xp25_ASAP7_75t_L g303 ( .A(n_300), .B(n_304), .C(n_305), .D(n_308), .Y(n_303) );
INVx1_ASAP7_75t_SL g374 ( .A(n_301), .Y(n_374) );
AND2x2_ASAP7_75t_L g418 ( .A(n_301), .B(n_419), .Y(n_418) );
OAI211xp5_ASAP7_75t_SL g302 ( .A1(n_303), .A2(n_310), .B(n_313), .C(n_322), .Y(n_302) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
INVx1_ASAP7_75t_SL g308 ( .A(n_309), .Y(n_308) );
NOR2xp33_ASAP7_75t_L g430 ( .A(n_309), .B(n_379), .Y(n_430) );
AOI22xp5_ASAP7_75t_L g429 ( .A1(n_311), .A2(n_430), .B1(n_431), .B2(n_432), .Y(n_429) );
INVx1_ASAP7_75t_SL g384 ( .A(n_312), .Y(n_384) );
AND2x2_ASAP7_75t_L g423 ( .A(n_312), .B(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_316), .B(n_317), .Y(n_315) );
NAND2xp5_ASAP7_75t_SL g416 ( .A(n_316), .B(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
NOR2xp33_ASAP7_75t_L g335 ( .A(n_320), .B(n_336), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_321), .B(n_346), .Y(n_406) );
OAI21xp5_ASAP7_75t_SL g322 ( .A1(n_323), .A2(n_328), .B(n_330), .Y(n_322) );
AND2x2_ASAP7_75t_L g323 ( .A(n_324), .B(n_325), .Y(n_323) );
INVx1_ASAP7_75t_L g398 ( .A(n_325), .Y(n_398) );
AND2x2_ASAP7_75t_L g325 ( .A(n_326), .B(n_327), .Y(n_325) );
INVx2_ASAP7_75t_L g426 ( .A(n_326), .Y(n_426) );
HB1xp67_ASAP7_75t_L g353 ( .A(n_327), .Y(n_353) );
OAI21xp33_ASAP7_75t_L g332 ( .A1(n_333), .A2(n_334), .B(n_337), .Y(n_332) );
CKINVDCx16_ASAP7_75t_R g345 ( .A(n_333), .Y(n_345) );
OR2x2_ASAP7_75t_L g383 ( .A(n_333), .B(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
AOI21xp33_ASAP7_75t_SL g378 ( .A1(n_336), .A2(n_379), .B(n_380), .Y(n_378) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
AOI221xp5_ASAP7_75t_L g366 ( .A1(n_340), .A2(n_367), .B1(n_370), .B2(n_377), .C(n_378), .Y(n_366) );
INVx1_ASAP7_75t_SL g410 ( .A(n_341), .Y(n_410) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
AND2x2_ASAP7_75t_L g344 ( .A(n_345), .B(n_346), .Y(n_344) );
OR2x2_ASAP7_75t_L g357 ( .A(n_345), .B(n_358), .Y(n_357) );
INVxp67_ASAP7_75t_L g394 ( .A(n_347), .Y(n_394) );
AOI22xp5_ASAP7_75t_L g349 ( .A1(n_350), .A2(n_351), .B1(n_354), .B2(n_355), .Y(n_349) );
INVx1_ASAP7_75t_L g389 ( .A(n_350), .Y(n_389) );
INVxp67_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_353), .B(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
NOR4xp25_ASAP7_75t_L g360 ( .A(n_361), .B(n_395), .C(n_408), .D(n_420), .Y(n_360) );
NAND3xp33_ASAP7_75t_SL g361 ( .A(n_362), .B(n_366), .C(n_381), .Y(n_361) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
NOR2xp33_ASAP7_75t_L g382 ( .A(n_364), .B(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_371), .B(n_376), .Y(n_380) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
OAI221xp5_ASAP7_75t_SL g408 ( .A1(n_383), .A2(n_409), .B1(n_410), .B2(n_411), .C(n_413), .Y(n_408) );
O2A1O1Ixp33_ASAP7_75t_L g399 ( .A1(n_385), .A2(n_400), .B(n_401), .C(n_403), .Y(n_399) );
INVx2_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
OAI22xp5_ASAP7_75t_L g403 ( .A1(n_386), .A2(n_404), .B1(n_406), .B2(n_407), .Y(n_403) );
INVx2_ASAP7_75t_SL g391 ( .A(n_392), .Y(n_391) );
A2O1A1Ixp33_ASAP7_75t_L g395 ( .A1(n_396), .A2(n_397), .B(n_398), .C(n_399), .Y(n_395) );
INVx1_ASAP7_75t_L g414 ( .A(n_407), .Y(n_414) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
OAI21xp5_ASAP7_75t_SL g413 ( .A1(n_414), .A2(n_415), .B(n_418), .Y(n_413) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
OAI221xp5_ASAP7_75t_SL g420 ( .A1(n_421), .A2(n_422), .B1(n_425), .B2(n_427), .C(n_429), .Y(n_420) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVxp67_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
OAI22xp5_ASAP7_75t_SL g449 ( .A1(n_435), .A2(n_450), .B1(n_718), .B2(n_719), .Y(n_449) );
INVx1_ASAP7_75t_SL g438 ( .A(n_439), .Y(n_438) );
HB1xp67_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx1_ASAP7_75t_SL g446 ( .A(n_440), .Y(n_446) );
INVx2_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_443), .B(n_444), .Y(n_442) );
AOI21xp33_ASAP7_75t_SL g447 ( .A1(n_445), .A2(n_448), .B(n_734), .Y(n_447) );
INVx1_ASAP7_75t_L g727 ( .A(n_450), .Y(n_727) );
NAND2x1_ASAP7_75t_L g450 ( .A(n_451), .B(n_634), .Y(n_450) );
NOR5xp2_ASAP7_75t_L g451 ( .A(n_452), .B(n_557), .C(n_589), .D(n_604), .E(n_621), .Y(n_451) );
A2O1A1Ixp33_ASAP7_75t_L g452 ( .A1(n_453), .A2(n_485), .B(n_504), .C(n_545), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_454), .B(n_466), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_454), .B(n_657), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_454), .B(n_609), .Y(n_672) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_455), .B(n_554), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_455), .B(n_501), .Y(n_558) );
AND2x2_ASAP7_75t_L g599 ( .A(n_455), .B(n_600), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_455), .B(n_568), .Y(n_603) );
OR2x2_ASAP7_75t_L g640 ( .A(n_455), .B(n_491), .Y(n_640) );
INVx3_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
AND2x2_ASAP7_75t_L g490 ( .A(n_456), .B(n_491), .Y(n_490) );
INVx3_ASAP7_75t_L g548 ( .A(n_456), .Y(n_548) );
OR2x2_ASAP7_75t_L g711 ( .A(n_456), .B(n_551), .Y(n_711) );
AOI22xp5_ASAP7_75t_L g613 ( .A1(n_466), .A2(n_614), .B1(n_615), .B2(n_618), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_466), .B(n_548), .Y(n_697) );
AND2x2_ASAP7_75t_L g466 ( .A(n_467), .B(n_476), .Y(n_466) );
AND2x2_ASAP7_75t_L g503 ( .A(n_467), .B(n_491), .Y(n_503) );
AND2x2_ASAP7_75t_L g550 ( .A(n_467), .B(n_551), .Y(n_550) );
INVx1_ASAP7_75t_L g555 ( .A(n_467), .Y(n_555) );
INVx3_ASAP7_75t_L g568 ( .A(n_467), .Y(n_568) );
OR2x2_ASAP7_75t_L g588 ( .A(n_467), .B(n_551), .Y(n_588) );
AND2x2_ASAP7_75t_L g607 ( .A(n_467), .B(n_477), .Y(n_607) );
BUFx2_ASAP7_75t_L g639 ( .A(n_467), .Y(n_639) );
AND2x4_ASAP7_75t_L g554 ( .A(n_476), .B(n_555), .Y(n_554) );
INVx1_ASAP7_75t_SL g476 ( .A(n_477), .Y(n_476) );
BUFx2_ASAP7_75t_L g489 ( .A(n_477), .Y(n_489) );
INVx2_ASAP7_75t_L g502 ( .A(n_477), .Y(n_502) );
OR2x2_ASAP7_75t_L g570 ( .A(n_477), .B(n_551), .Y(n_570) );
AND2x2_ASAP7_75t_L g600 ( .A(n_477), .B(n_491), .Y(n_600) );
AND2x2_ASAP7_75t_L g617 ( .A(n_477), .B(n_548), .Y(n_617) );
AND2x2_ASAP7_75t_L g657 ( .A(n_477), .B(n_568), .Y(n_657) );
AND2x2_ASAP7_75t_SL g693 ( .A(n_477), .B(n_503), .Y(n_693) );
INVx1_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
NAND2xp33_ASAP7_75t_SL g486 ( .A(n_487), .B(n_500), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_488), .B(n_490), .Y(n_487) );
NOR2xp33_ASAP7_75t_L g671 ( .A(n_488), .B(n_672), .Y(n_671) );
INVx1_ASAP7_75t_SL g488 ( .A(n_489), .Y(n_488) );
OAI21xp33_ASAP7_75t_L g631 ( .A1(n_489), .A2(n_503), .B(n_632), .Y(n_631) );
NOR2xp33_ASAP7_75t_L g687 ( .A(n_489), .B(n_491), .Y(n_687) );
AND2x2_ASAP7_75t_L g623 ( .A(n_490), .B(n_624), .Y(n_623) );
INVx3_ASAP7_75t_L g551 ( .A(n_491), .Y(n_551) );
HB1xp67_ASAP7_75t_L g649 ( .A(n_491), .Y(n_649) );
NOR2xp33_ASAP7_75t_L g716 ( .A(n_500), .B(n_548), .Y(n_716) );
INVx2_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
AOI22xp33_ASAP7_75t_L g658 ( .A1(n_501), .A2(n_659), .B1(n_660), .B2(n_665), .Y(n_658) );
AND2x2_ASAP7_75t_L g501 ( .A(n_502), .B(n_503), .Y(n_501) );
AND2x2_ASAP7_75t_L g549 ( .A(n_502), .B(n_550), .Y(n_549) );
OR2x2_ASAP7_75t_L g587 ( .A(n_502), .B(n_588), .Y(n_587) );
INVx1_ASAP7_75t_SL g624 ( .A(n_502), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_503), .B(n_617), .Y(n_616) );
INVx1_ASAP7_75t_L g678 ( .A(n_503), .Y(n_678) );
CKINVDCx16_ASAP7_75t_R g504 ( .A(n_505), .Y(n_504) );
AND2x2_ASAP7_75t_L g505 ( .A(n_506), .B(n_525), .Y(n_505) );
INVx4_ASAP7_75t_L g564 ( .A(n_506), .Y(n_564) );
AND2x2_ASAP7_75t_L g642 ( .A(n_506), .B(n_609), .Y(n_642) );
AND2x2_ASAP7_75t_L g506 ( .A(n_507), .B(n_516), .Y(n_506) );
INVx3_ASAP7_75t_L g561 ( .A(n_507), .Y(n_561) );
AND2x2_ASAP7_75t_L g575 ( .A(n_507), .B(n_576), .Y(n_575) );
INVx1_ASAP7_75t_L g579 ( .A(n_507), .Y(n_579) );
INVx2_ASAP7_75t_L g593 ( .A(n_507), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_507), .B(n_609), .Y(n_608) );
AND2x2_ASAP7_75t_L g650 ( .A(n_507), .B(n_645), .Y(n_650) );
AND2x2_ASAP7_75t_L g715 ( .A(n_507), .B(n_685), .Y(n_715) );
OR2x6_ASAP7_75t_L g507 ( .A(n_508), .B(n_514), .Y(n_507) );
AND2x2_ASAP7_75t_L g556 ( .A(n_516), .B(n_537), .Y(n_556) );
INVx2_ASAP7_75t_L g576 ( .A(n_516), .Y(n_576) );
INVx1_ASAP7_75t_L g581 ( .A(n_525), .Y(n_581) );
AND2x2_ASAP7_75t_L g627 ( .A(n_525), .B(n_575), .Y(n_627) );
AND2x2_ASAP7_75t_L g525 ( .A(n_526), .B(n_536), .Y(n_525) );
INVx2_ASAP7_75t_L g566 ( .A(n_526), .Y(n_566) );
INVx1_ASAP7_75t_L g574 ( .A(n_526), .Y(n_574) );
AND2x2_ASAP7_75t_L g592 ( .A(n_526), .B(n_593), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_526), .B(n_576), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_528), .B(n_533), .Y(n_527) );
AOI21xp5_ASAP7_75t_L g529 ( .A1(n_530), .A2(n_531), .B(n_532), .Y(n_529) );
AND2x2_ASAP7_75t_L g609 ( .A(n_536), .B(n_566), .Y(n_609) );
INVx1_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
INVx2_ASAP7_75t_L g562 ( .A(n_537), .Y(n_562) );
AND2x2_ASAP7_75t_L g645 ( .A(n_537), .B(n_576), .Y(n_645) );
OAI21xp5_ASAP7_75t_SL g545 ( .A1(n_546), .A2(n_552), .B(n_556), .Y(n_545) );
INVx1_ASAP7_75t_SL g590 ( .A(n_546), .Y(n_590) );
AND2x2_ASAP7_75t_L g546 ( .A(n_547), .B(n_549), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_547), .B(n_554), .Y(n_647) );
INVx1_ASAP7_75t_SL g547 ( .A(n_548), .Y(n_547) );
AND2x2_ASAP7_75t_L g596 ( .A(n_548), .B(n_551), .Y(n_596) );
AND2x2_ASAP7_75t_L g625 ( .A(n_548), .B(n_569), .Y(n_625) );
OR2x2_ASAP7_75t_L g628 ( .A(n_548), .B(n_588), .Y(n_628) );
AOI222xp33_ASAP7_75t_L g692 ( .A1(n_549), .A2(n_641), .B1(n_693), .B2(n_694), .C1(n_696), .C2(n_698), .Y(n_692) );
BUFx2_ASAP7_75t_L g606 ( .A(n_551), .Y(n_606) );
INVx1_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
AND2x2_ASAP7_75t_L g595 ( .A(n_554), .B(n_596), .Y(n_595) );
INVx3_ASAP7_75t_SL g612 ( .A(n_554), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_554), .B(n_606), .Y(n_666) );
AND2x2_ASAP7_75t_L g601 ( .A(n_556), .B(n_561), .Y(n_601) );
INVx1_ASAP7_75t_L g620 ( .A(n_556), .Y(n_620) );
OAI221xp5_ASAP7_75t_SL g557 ( .A1(n_558), .A2(n_559), .B1(n_563), .B2(n_567), .C(n_571), .Y(n_557) );
OR2x2_ASAP7_75t_L g629 ( .A(n_559), .B(n_630), .Y(n_629) );
INVx1_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
AND2x2_ASAP7_75t_L g560 ( .A(n_561), .B(n_562), .Y(n_560) );
AND2x2_ASAP7_75t_L g614 ( .A(n_561), .B(n_584), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_561), .B(n_574), .Y(n_654) );
AND2x2_ASAP7_75t_L g659 ( .A(n_561), .B(n_609), .Y(n_659) );
HB1xp67_ASAP7_75t_L g669 ( .A(n_561), .Y(n_669) );
NAND2x1_ASAP7_75t_SL g680 ( .A(n_561), .B(n_681), .Y(n_680) );
OR2x2_ASAP7_75t_L g565 ( .A(n_562), .B(n_566), .Y(n_565) );
INVx2_ASAP7_75t_L g585 ( .A(n_562), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_562), .B(n_580), .Y(n_611) );
INVx1_ASAP7_75t_L g677 ( .A(n_562), .Y(n_677) );
INVx1_ASAP7_75t_L g652 ( .A(n_563), .Y(n_652) );
OR2x2_ASAP7_75t_L g563 ( .A(n_564), .B(n_565), .Y(n_563) );
INVx1_ASAP7_75t_L g664 ( .A(n_564), .Y(n_664) );
NOR2xp67_ASAP7_75t_L g676 ( .A(n_564), .B(n_677), .Y(n_676) );
INVx2_ASAP7_75t_L g681 ( .A(n_565), .Y(n_681) );
NOR2xp33_ASAP7_75t_L g688 ( .A(n_565), .B(n_689), .Y(n_688) );
AND2x2_ASAP7_75t_L g584 ( .A(n_566), .B(n_585), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_566), .B(n_576), .Y(n_597) );
INVx1_ASAP7_75t_L g663 ( .A(n_566), .Y(n_663) );
INVx1_ASAP7_75t_L g684 ( .A(n_567), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_568), .B(n_569), .Y(n_567) );
INVx1_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
OAI21xp5_ASAP7_75t_SL g571 ( .A1(n_572), .A2(n_577), .B(n_586), .Y(n_571) );
AND2x2_ASAP7_75t_L g572 ( .A(n_573), .B(n_575), .Y(n_572) );
AND2x2_ASAP7_75t_L g717 ( .A(n_573), .B(n_650), .Y(n_717) );
INVx1_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
AND2x2_ASAP7_75t_L g685 ( .A(n_574), .B(n_645), .Y(n_685) );
AOI32xp33_ASAP7_75t_L g598 ( .A1(n_575), .A2(n_581), .A3(n_599), .B1(n_601), .B2(n_602), .Y(n_598) );
AOI322xp5_ASAP7_75t_L g700 ( .A1(n_575), .A2(n_607), .A3(n_690), .B1(n_701), .B2(n_702), .C1(n_703), .C2(n_705), .Y(n_700) );
INVx2_ASAP7_75t_L g580 ( .A(n_576), .Y(n_580) );
INVx1_ASAP7_75t_L g690 ( .A(n_576), .Y(n_690) );
OAI22xp5_ASAP7_75t_L g577 ( .A1(n_578), .A2(n_581), .B1(n_582), .B2(n_583), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_578), .B(n_584), .Y(n_633) );
AND2x2_ASAP7_75t_L g578 ( .A(n_579), .B(n_580), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_579), .B(n_645), .Y(n_695) );
INVx1_ASAP7_75t_L g582 ( .A(n_580), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_580), .B(n_609), .Y(n_699) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
INVx1_ASAP7_75t_SL g586 ( .A(n_587), .Y(n_586) );
NOR2xp33_ASAP7_75t_L g682 ( .A(n_588), .B(n_683), .Y(n_682) );
OAI221xp5_ASAP7_75t_SL g589 ( .A1(n_590), .A2(n_591), .B1(n_594), .B2(n_597), .C(n_598), .Y(n_589) );
OR2x2_ASAP7_75t_L g610 ( .A(n_591), .B(n_611), .Y(n_610) );
OR2x2_ASAP7_75t_L g619 ( .A(n_591), .B(n_620), .Y(n_619) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
AND2x2_ASAP7_75t_L g644 ( .A(n_592), .B(n_645), .Y(n_644) );
INVx2_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
AND2x2_ASAP7_75t_L g648 ( .A(n_602), .B(n_649), .Y(n_648) );
INVx1_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
OAI221xp5_ASAP7_75t_L g604 ( .A1(n_605), .A2(n_608), .B1(n_610), .B2(n_612), .C(n_613), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_606), .B(n_607), .Y(n_605) );
AOI22xp5_ASAP7_75t_L g636 ( .A1(n_606), .A2(n_637), .B1(n_641), .B2(n_642), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_607), .B(n_708), .Y(n_707) );
INVx1_ASAP7_75t_L g712 ( .A(n_607), .Y(n_712) );
INVx1_ASAP7_75t_L g706 ( .A(n_609), .Y(n_706) );
INVx1_ASAP7_75t_SL g641 ( .A(n_610), .Y(n_641) );
NOR2xp33_ASAP7_75t_L g702 ( .A(n_612), .B(n_640), .Y(n_702) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_617), .B(n_676), .Y(n_675) );
INVx1_ASAP7_75t_SL g683 ( .A(n_617), .Y(n_683) );
INVx1_ASAP7_75t_SL g618 ( .A(n_619), .Y(n_618) );
OAI221xp5_ASAP7_75t_SL g621 ( .A1(n_622), .A2(n_626), .B1(n_628), .B2(n_629), .C(n_631), .Y(n_621) );
NOR2xp33_ASAP7_75t_SL g622 ( .A(n_623), .B(n_625), .Y(n_622) );
AOI22xp5_ASAP7_75t_L g686 ( .A1(n_623), .A2(n_641), .B1(n_687), .B2(n_688), .Y(n_686) );
CKINVDCx14_ASAP7_75t_R g626 ( .A(n_627), .Y(n_626) );
OAI21xp33_ASAP7_75t_L g705 ( .A1(n_628), .A2(n_706), .B(n_707), .Y(n_705) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
NOR3xp33_ASAP7_75t_SL g634 ( .A(n_635), .B(n_667), .C(n_691), .Y(n_634) );
NAND4xp25_ASAP7_75t_L g635 ( .A(n_636), .B(n_643), .C(n_651), .D(n_658), .Y(n_635) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
OR2x2_ASAP7_75t_L g638 ( .A(n_639), .B(n_640), .Y(n_638) );
INVx1_ASAP7_75t_L g714 ( .A(n_639), .Y(n_714) );
INVx3_ASAP7_75t_SL g708 ( .A(n_640), .Y(n_708) );
OR2x2_ASAP7_75t_L g713 ( .A(n_640), .B(n_714), .Y(n_713) );
AOI22xp5_ASAP7_75t_L g643 ( .A1(n_644), .A2(n_646), .B1(n_648), .B2(n_650), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_645), .B(n_663), .Y(n_704) );
INVxp67_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
OAI21xp5_ASAP7_75t_SL g651 ( .A1(n_652), .A2(n_653), .B(n_655), .Y(n_651) );
INVxp67_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_662), .B(n_664), .Y(n_661) );
INVxp67_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
OAI211xp5_ASAP7_75t_SL g667 ( .A1(n_668), .A2(n_670), .B(n_673), .C(n_686), .Y(n_667) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
INVx1_ASAP7_75t_L g701 ( .A(n_672), .Y(n_701) );
AOI222xp33_ASAP7_75t_L g673 ( .A1(n_674), .A2(n_678), .B1(n_679), .B2(n_682), .C1(n_684), .C2(n_685), .Y(n_673) );
INVxp67_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
NAND4xp25_ASAP7_75t_SL g710 ( .A(n_683), .B(n_711), .C(n_712), .D(n_713), .Y(n_710) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
NAND3xp33_ASAP7_75t_SL g691 ( .A(n_692), .B(n_700), .C(n_709), .Y(n_691) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
AOI22xp33_ASAP7_75t_L g709 ( .A1(n_710), .A2(n_715), .B1(n_716), .B2(n_717), .Y(n_709) );
INVx1_ASAP7_75t_L g729 ( .A(n_719), .Y(n_729) );
INVx1_ASAP7_75t_L g730 ( .A(n_720), .Y(n_730) );
INVx1_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
INVx2_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
INVx1_ASAP7_75t_SL g731 ( .A(n_732), .Y(n_731) );
INVx2_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
endmodule