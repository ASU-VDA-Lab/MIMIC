module fake_jpeg_15781_n_144 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_144);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_144;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_9),
.Y(n_13)
);

INVx11_ASAP7_75t_SL g14 ( 
.A(n_5),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_2),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_26),
.B(n_1),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_28),
.B(n_30),
.Y(n_38)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_26),
.Y(n_29)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_13),
.B(n_15),
.Y(n_30)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx2_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_33),
.B(n_34),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_13),
.B(n_15),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_17),
.B(n_1),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_35),
.B(n_36),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_29),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_37)
);

OAI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_37),
.A2(n_42),
.B1(n_46),
.B2(n_20),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g42 ( 
.A1(n_29),
.A2(n_20),
.B1(n_25),
.B2(n_27),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_30),
.B(n_21),
.Y(n_43)
);

CKINVDCx14_ASAP7_75t_R g53 ( 
.A(n_43),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_28),
.B(n_23),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_44),
.B(n_50),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_16),
.Y(n_45)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_L g46 ( 
.A1(n_36),
.A2(n_20),
.B1(n_25),
.B2(n_27),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_33),
.A2(n_24),
.B1(n_21),
.B2(n_19),
.Y(n_48)
);

AO22x2_ASAP7_75t_L g64 ( 
.A1(n_48),
.A2(n_17),
.B1(n_24),
.B2(n_18),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_32),
.B(n_23),
.Y(n_50)
);

INVx3_ASAP7_75t_SL g51 ( 
.A(n_47),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_51),
.B(n_57),
.Y(n_77)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_54),
.Y(n_68)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_49),
.Y(n_56)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_56),
.Y(n_76)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_49),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_58),
.Y(n_81)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_59),
.Y(n_69)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_60),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_47),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_61),
.B(n_63),
.Y(n_80)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_62),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_45),
.B(n_35),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_64),
.A2(n_22),
.B1(n_16),
.B2(n_48),
.Y(n_82)
);

AO22x2_ASAP7_75t_L g65 ( 
.A1(n_37),
.A2(n_36),
.B1(n_32),
.B2(n_27),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_65),
.A2(n_66),
.B1(n_62),
.B2(n_56),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_66),
.A2(n_46),
.B1(n_42),
.B2(n_41),
.Y(n_73)
);

XNOR2xp5_ASAP7_75t_SL g67 ( 
.A(n_64),
.B(n_44),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_67),
.A2(n_71),
.B1(n_33),
.B2(n_54),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_65),
.B(n_50),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_64),
.A2(n_31),
.B1(n_19),
.B2(n_18),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_72),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_73),
.A2(n_65),
.B1(n_51),
.B2(n_36),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_53),
.B(n_38),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_74),
.B(n_82),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_55),
.B(n_41),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_78),
.B(n_83),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_79),
.B(n_65),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_64),
.B(n_38),
.Y(n_83)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_68),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_85),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_80),
.B(n_52),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_86),
.B(n_87),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_77),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_68),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_88),
.B(n_89),
.Y(n_98)
);

CKINVDCx14_ASAP7_75t_R g89 ( 
.A(n_82),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_76),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_91),
.B(n_76),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_92),
.A2(n_93),
.B1(n_97),
.B2(n_71),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_95),
.B(n_81),
.Y(n_106)
);

INVx1_ASAP7_75t_SL g96 ( 
.A(n_70),
.Y(n_96)
);

CKINVDCx14_ASAP7_75t_R g109 ( 
.A(n_96),
.Y(n_109)
);

NOR2x1_ASAP7_75t_L g97 ( 
.A(n_83),
.B(n_43),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_95),
.B(n_67),
.C(n_78),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_99),
.B(n_106),
.C(n_84),
.Y(n_110)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_101),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_91),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_103),
.B(n_107),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_104),
.A2(n_93),
.B(n_94),
.Y(n_112)
);

OAI22xp33_ASAP7_75t_L g105 ( 
.A1(n_90),
.A2(n_79),
.B1(n_71),
.B2(n_75),
.Y(n_105)
);

AOI322xp5_ASAP7_75t_L g116 ( 
.A1(n_105),
.A2(n_108),
.A3(n_93),
.B1(n_85),
.B2(n_96),
.C1(n_70),
.C2(n_32),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_106),
.B(n_3),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_84),
.B(n_97),
.Y(n_107)
);

AOI322xp5_ASAP7_75t_L g108 ( 
.A1(n_94),
.A2(n_81),
.A3(n_69),
.B1(n_22),
.B2(n_31),
.C1(n_32),
.C2(n_75),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_110),
.B(n_117),
.C(n_104),
.Y(n_121)
);

XNOR2x1_ASAP7_75t_L g111 ( 
.A(n_99),
.B(n_90),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_111),
.B(n_118),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g120 ( 
.A1(n_112),
.A2(n_116),
.B1(n_98),
.B2(n_109),
.Y(n_120)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_100),
.Y(n_113)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_113),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_102),
.B(n_88),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_114),
.A2(n_4),
.B(n_6),
.Y(n_126)
);

AOI322xp5_ASAP7_75t_L g117 ( 
.A1(n_105),
.A2(n_32),
.A3(n_12),
.B1(n_11),
.B2(n_5),
.C1(n_6),
.C2(n_2),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_120),
.B(n_123),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_121),
.B(n_124),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_115),
.A2(n_107),
.B1(n_101),
.B2(n_100),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_110),
.B(n_12),
.C(n_5),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_126),
.B(n_6),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_121),
.A2(n_119),
.B(n_112),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_129),
.B(n_130),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_123),
.B(n_115),
.Y(n_131)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_131),
.Y(n_133)
);

OR2x2_ASAP7_75t_L g132 ( 
.A(n_124),
.B(n_113),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_132),
.B(n_118),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_128),
.A2(n_111),
.B1(n_122),
.B2(n_125),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_134),
.B(n_135),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_136),
.B(n_127),
.C(n_128),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_137),
.B(n_138),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_133),
.A2(n_125),
.B1(n_8),
.B2(n_9),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_139),
.B(n_134),
.Y(n_141)
);

BUFx24_ASAP7_75t_SL g142 ( 
.A(n_141),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_142),
.A2(n_140),
.B(n_7),
.Y(n_143)
);

MAJx2_ASAP7_75t_L g144 ( 
.A(n_143),
.B(n_7),
.C(n_142),
.Y(n_144)
);


endmodule