module fake_netlist_5_1081_n_324 (n_82, n_10, n_24, n_83, n_61, n_75, n_65, n_78, n_74, n_57, n_37, n_31, n_13, n_66, n_60, n_16, n_43, n_0, n_58, n_9, n_69, n_18, n_42, n_22, n_1, n_45, n_46, n_21, n_38, n_80, n_4, n_35, n_73, n_17, n_19, n_30, n_5, n_33, n_14, n_23, n_29, n_79, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_62, n_71, n_59, n_26, n_55, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_12, n_67, n_36, n_76, n_27, n_64, n_77, n_81, n_28, n_70, n_68, n_72, n_32, n_41, n_56, n_51, n_63, n_11, n_7, n_15, n_48, n_50, n_52, n_324);

input n_82;
input n_10;
input n_24;
input n_83;
input n_61;
input n_75;
input n_65;
input n_78;
input n_74;
input n_57;
input n_37;
input n_31;
input n_13;
input n_66;
input n_60;
input n_16;
input n_43;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_42;
input n_22;
input n_1;
input n_45;
input n_46;
input n_21;
input n_38;
input n_80;
input n_4;
input n_35;
input n_73;
input n_17;
input n_19;
input n_30;
input n_5;
input n_33;
input n_14;
input n_23;
input n_29;
input n_79;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_62;
input n_71;
input n_59;
input n_26;
input n_55;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_12;
input n_67;
input n_36;
input n_76;
input n_27;
input n_64;
input n_77;
input n_81;
input n_28;
input n_70;
input n_68;
input n_72;
input n_32;
input n_41;
input n_56;
input n_51;
input n_63;
input n_11;
input n_7;
input n_15;
input n_48;
input n_50;
input n_52;

output n_324;

wire n_137;
wire n_294;
wire n_318;
wire n_194;
wire n_316;
wire n_248;
wire n_136;
wire n_86;
wire n_146;
wire n_124;
wire n_315;
wire n_268;
wire n_127;
wire n_235;
wire n_226;
wire n_111;
wire n_155;
wire n_116;
wire n_284;
wire n_245;
wire n_139;
wire n_105;
wire n_280;
wire n_254;
wire n_302;
wire n_265;
wire n_293;
wire n_244;
wire n_173;
wire n_198;
wire n_247;
wire n_314;
wire n_321;
wire n_292;
wire n_100;
wire n_212;
wire n_119;
wire n_275;
wire n_252;
wire n_295;
wire n_133;
wire n_147;
wire n_307;
wire n_87;
wire n_150;
wire n_106;
wire n_209;
wire n_259;
wire n_301;
wire n_93;
wire n_186;
wire n_134;
wire n_191;
wire n_171;
wire n_153;
wire n_204;
wire n_250;
wire n_260;
wire n_298;
wire n_320;
wire n_286;
wire n_122;
wire n_282;
wire n_132;
wire n_90;
wire n_101;
wire n_281;
wire n_240;
wire n_189;
wire n_220;
wire n_291;
wire n_231;
wire n_257;
wire n_152;
wire n_317;
wire n_323;
wire n_195;
wire n_227;
wire n_271;
wire n_94;
wire n_123;
wire n_167;
wire n_234;
wire n_308;
wire n_267;
wire n_297;
wire n_156;
wire n_225;
wire n_219;
wire n_157;
wire n_131;
wire n_192;
wire n_223;
wire n_158;
wire n_138;
wire n_264;
wire n_109;
wire n_163;
wire n_276;
wire n_95;
wire n_183;
wire n_185;
wire n_243;
wire n_169;
wire n_255;
wire n_215;
wire n_196;
wire n_211;
wire n_218;
wire n_181;
wire n_290;
wire n_221;
wire n_178;
wire n_287;
wire n_104;
wire n_141;
wire n_145;
wire n_313;
wire n_88;
wire n_216;
wire n_168;
wire n_164;
wire n_311;
wire n_208;
wire n_142;
wire n_214;
wire n_140;
wire n_299;
wire n_303;
wire n_296;
wire n_241;
wire n_184;
wire n_144;
wire n_114;
wire n_96;
wire n_165;
wire n_213;
wire n_129;
wire n_98;
wire n_197;
wire n_107;
wire n_236;
wire n_249;
wire n_304;
wire n_203;
wire n_274;
wire n_277;
wire n_92;
wire n_149;
wire n_309;
wire n_84;
wire n_130;
wire n_322;
wire n_258;
wire n_151;
wire n_306;
wire n_288;
wire n_188;
wire n_190;
wire n_201;
wire n_263;
wire n_224;
wire n_228;
wire n_283;
wire n_112;
wire n_85;
wire n_239;
wire n_310;
wire n_170;
wire n_102;
wire n_161;
wire n_273;
wire n_270;
wire n_230;
wire n_118;
wire n_279;
wire n_253;
wire n_261;
wire n_174;
wire n_289;
wire n_172;
wire n_206;
wire n_217;
wire n_312;
wire n_210;
wire n_91;
wire n_176;
wire n_182;
wire n_143;
wire n_237;
wire n_180;
wire n_207;
wire n_229;
wire n_108;
wire n_177;
wire n_117;
wire n_233;
wire n_205;
wire n_113;
wire n_246;
wire n_179;
wire n_125;
wire n_269;
wire n_128;
wire n_285;
wire n_120;
wire n_232;
wire n_135;
wire n_126;
wire n_202;
wire n_266;
wire n_272;
wire n_193;
wire n_251;
wire n_160;
wire n_154;
wire n_148;
wire n_300;
wire n_159;
wire n_175;
wire n_262;
wire n_238;
wire n_99;
wire n_319;
wire n_121;
wire n_242;
wire n_200;
wire n_162;
wire n_222;
wire n_89;
wire n_115;
wire n_199;
wire n_187;
wire n_103;
wire n_97;
wire n_166;
wire n_256;
wire n_305;
wire n_278;
wire n_110;

INVx1_ASAP7_75t_L g84 ( 
.A(n_43),
.Y(n_84)
);

INVxp67_ASAP7_75t_SL g85 ( 
.A(n_58),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_81),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_7),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_29),
.Y(n_88)
);

INVxp33_ASAP7_75t_L g89 ( 
.A(n_80),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_64),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_14),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_51),
.Y(n_92)
);

CKINVDCx5p33_ASAP7_75t_R g93 ( 
.A(n_56),
.Y(n_93)
);

INVxp33_ASAP7_75t_L g94 ( 
.A(n_13),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_63),
.Y(n_95)
);

INVxp33_ASAP7_75t_L g96 ( 
.A(n_49),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_16),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_44),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_48),
.Y(n_99)
);

INVxp33_ASAP7_75t_SL g100 ( 
.A(n_83),
.Y(n_100)
);

INVxp67_ASAP7_75t_SL g101 ( 
.A(n_30),
.Y(n_101)
);

INVxp33_ASAP7_75t_L g102 ( 
.A(n_35),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_32),
.Y(n_103)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_5),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_2),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_1),
.Y(n_106)
);

INVxp33_ASAP7_75t_L g107 ( 
.A(n_60),
.Y(n_107)
);

BUFx2_ASAP7_75t_L g108 ( 
.A(n_55),
.Y(n_108)
);

INVxp67_ASAP7_75t_SL g109 ( 
.A(n_76),
.Y(n_109)
);

NOR2xp67_ASAP7_75t_L g110 ( 
.A(n_40),
.B(n_65),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_46),
.Y(n_111)
);

CKINVDCx5p33_ASAP7_75t_R g112 ( 
.A(n_38),
.Y(n_112)
);

INVx2_ASAP7_75t_SL g113 ( 
.A(n_23),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_6),
.Y(n_114)
);

INVx1_ASAP7_75t_SL g115 ( 
.A(n_18),
.Y(n_115)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_71),
.Y(n_116)
);

INVxp67_ASAP7_75t_SL g117 ( 
.A(n_54),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_73),
.Y(n_118)
);

INVx1_ASAP7_75t_SL g119 ( 
.A(n_42),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_82),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_1),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_10),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_52),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_68),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_17),
.Y(n_125)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_45),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_20),
.Y(n_127)
);

INVxp33_ASAP7_75t_L g128 ( 
.A(n_78),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_6),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_19),
.Y(n_130)
);

INVxp67_ASAP7_75t_SL g131 ( 
.A(n_57),
.Y(n_131)
);

INVx1_ASAP7_75t_SL g132 ( 
.A(n_70),
.Y(n_132)
);

INVxp33_ASAP7_75t_L g133 ( 
.A(n_7),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_33),
.Y(n_134)
);

INVxp33_ASAP7_75t_L g135 ( 
.A(n_66),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_41),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_31),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_50),
.Y(n_138)
);

INVxp33_ASAP7_75t_SL g139 ( 
.A(n_15),
.Y(n_139)
);

INVxp67_ASAP7_75t_SL g140 ( 
.A(n_67),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_22),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_8),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_105),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_87),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_106),
.Y(n_145)
);

CKINVDCx5p33_ASAP7_75t_R g146 ( 
.A(n_93),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_114),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_108),
.B(n_0),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_121),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_122),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_95),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_129),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_112),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_94),
.B(n_2),
.Y(n_154)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_95),
.Y(n_155)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_104),
.Y(n_156)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_116),
.Y(n_157)
);

BUFx12f_ASAP7_75t_L g158 ( 
.A(n_113),
.Y(n_158)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_104),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_88),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_142),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_138),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_94),
.B(n_3),
.Y(n_163)
);

BUFx10_ASAP7_75t_L g164 ( 
.A(n_84),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_116),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_138),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_111),
.B(n_3),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_89),
.B(n_4),
.Y(n_168)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_126),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_86),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_97),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_90),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_151),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_151),
.B(n_125),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_171),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_151),
.B(n_115),
.Y(n_176)
);

INVx5_ASAP7_75t_L g177 ( 
.A(n_151),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_146),
.B(n_96),
.Y(n_178)
);

BUFx10_ASAP7_75t_L g179 ( 
.A(n_153),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_L g180 ( 
.A1(n_154),
.A2(n_133),
.B1(n_128),
.B2(n_107),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_165),
.Y(n_181)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_165),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_165),
.B(n_119),
.Y(n_183)
);

NAND2x1p5_ASAP7_75t_L g184 ( 
.A(n_167),
.B(n_132),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_169),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_156),
.Y(n_186)
);

NOR3xp33_ASAP7_75t_L g187 ( 
.A(n_167),
.B(n_168),
.C(n_148),
.Y(n_187)
);

AND2x4_ASAP7_75t_L g188 ( 
.A(n_163),
.B(n_127),
.Y(n_188)
);

NAND3xp33_ASAP7_75t_L g189 ( 
.A(n_150),
.B(n_133),
.C(n_107),
.Y(n_189)
);

INVx1_ASAP7_75t_SL g190 ( 
.A(n_162),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_158),
.B(n_96),
.Y(n_191)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_158),
.Y(n_192)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_156),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_169),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_159),
.Y(n_195)
);

INVx3_ASAP7_75t_R g196 ( 
.A(n_159),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_143),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_144),
.A2(n_102),
.B1(n_135),
.B2(n_128),
.Y(n_198)
);

INVx2_ASAP7_75t_SL g199 ( 
.A(n_164),
.Y(n_199)
);

INVxp33_ASAP7_75t_L g200 ( 
.A(n_170),
.Y(n_200)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_155),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_164),
.B(n_135),
.Y(n_202)
);

AND2x6_ASAP7_75t_L g203 ( 
.A(n_155),
.B(n_126),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_145),
.Y(n_204)
);

INVx4_ASAP7_75t_L g205 ( 
.A(n_181),
.Y(n_205)
);

INVx3_ASAP7_75t_SL g206 ( 
.A(n_175),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_204),
.Y(n_207)
);

AND2x4_ASAP7_75t_SL g208 ( 
.A(n_179),
.B(n_171),
.Y(n_208)
);

NOR3xp33_ASAP7_75t_SL g209 ( 
.A(n_198),
.B(n_160),
.C(n_149),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_174),
.B(n_172),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_204),
.Y(n_211)
);

NOR2xp67_ASAP7_75t_L g212 ( 
.A(n_177),
.B(n_155),
.Y(n_212)
);

NOR3xp33_ASAP7_75t_SL g213 ( 
.A(n_198),
.B(n_147),
.C(n_152),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_174),
.A2(n_85),
.B(n_131),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_184),
.A2(n_166),
.B1(n_162),
.B2(n_98),
.Y(n_215)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_181),
.Y(n_216)
);

AOI211xp5_ASAP7_75t_L g217 ( 
.A1(n_187),
.A2(n_189),
.B(n_202),
.C(n_178),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g218 ( 
.A(n_200),
.B(n_161),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_180),
.B(n_100),
.Y(n_219)
);

AND3x1_ASAP7_75t_SL g220 ( 
.A(n_184),
.B(n_120),
.C(n_92),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_197),
.Y(n_221)
);

NOR3xp33_ASAP7_75t_SL g222 ( 
.A(n_189),
.B(n_118),
.C(n_141),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_186),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_199),
.B(n_139),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_186),
.Y(n_225)
);

AO22x1_ASAP7_75t_L g226 ( 
.A1(n_191),
.A2(n_101),
.B1(n_109),
.B2(n_117),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_188),
.B(n_157),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_186),
.Y(n_228)
);

AND2x6_ASAP7_75t_L g229 ( 
.A(n_173),
.B(n_91),
.Y(n_229)
);

INVx1_ASAP7_75t_SL g230 ( 
.A(n_190),
.Y(n_230)
);

AND2x4_ASAP7_75t_L g231 ( 
.A(n_176),
.B(n_123),
.Y(n_231)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_182),
.Y(n_232)
);

NAND2x1p5_ASAP7_75t_L g233 ( 
.A(n_192),
.B(n_110),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_223),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_210),
.A2(n_183),
.B(n_177),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_206),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_221),
.Y(n_237)
);

AOI221xp5_ASAP7_75t_L g238 ( 
.A1(n_219),
.A2(n_166),
.B1(n_190),
.B2(n_99),
.C(n_136),
.Y(n_238)
);

INVx4_ASAP7_75t_L g239 ( 
.A(n_228),
.Y(n_239)
);

INVx4_ASAP7_75t_L g240 ( 
.A(n_228),
.Y(n_240)
);

INVx3_ASAP7_75t_L g241 ( 
.A(n_228),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_217),
.A2(n_231),
.B1(n_213),
.B2(n_227),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_214),
.A2(n_140),
.B(n_103),
.Y(n_243)
);

INVx1_ASAP7_75t_SL g244 ( 
.A(n_230),
.Y(n_244)
);

AND2x4_ASAP7_75t_L g245 ( 
.A(n_207),
.B(n_193),
.Y(n_245)
);

INVx3_ASAP7_75t_L g246 ( 
.A(n_232),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_218),
.Y(n_247)
);

A2O1A1Ixp33_ASAP7_75t_L g248 ( 
.A1(n_222),
.A2(n_124),
.B(n_130),
.C(n_134),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_225),
.B(n_201),
.Y(n_249)
);

O2A1O1Ixp33_ASAP7_75t_SL g250 ( 
.A1(n_224),
.A2(n_137),
.B(n_194),
.C(n_185),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_L g251 ( 
.A1(n_211),
.A2(n_203),
.B1(n_195),
.B2(n_201),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g252 ( 
.A(n_229),
.Y(n_252)
);

OR2x2_ASAP7_75t_L g253 ( 
.A(n_226),
.B(n_8),
.Y(n_253)
);

OA21x2_ASAP7_75t_L g254 ( 
.A1(n_243),
.A2(n_212),
.B(n_209),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_237),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_242),
.A2(n_215),
.B1(n_233),
.B2(n_208),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_236),
.Y(n_257)
);

OAI22xp33_ASAP7_75t_L g258 ( 
.A1(n_253),
.A2(n_220),
.B1(n_216),
.B2(n_205),
.Y(n_258)
);

AOI221xp5_ASAP7_75t_L g259 ( 
.A1(n_238),
.A2(n_205),
.B1(n_10),
.B2(n_11),
.C(n_12),
.Y(n_259)
);

AND2x2_ASAP7_75t_L g260 ( 
.A(n_244),
.B(n_247),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_245),
.Y(n_261)
);

OAI21x1_ASAP7_75t_SL g262 ( 
.A1(n_243),
.A2(n_229),
.B(n_47),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_246),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_249),
.Y(n_264)
);

A2O1A1Ixp33_ASAP7_75t_L g265 ( 
.A1(n_235),
.A2(n_196),
.B(n_203),
.C(n_9),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_246),
.Y(n_266)
);

INVx4_ASAP7_75t_L g267 ( 
.A(n_234),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g268 ( 
.A(n_260),
.B(n_248),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_257),
.Y(n_269)
);

OA21x2_ASAP7_75t_L g270 ( 
.A1(n_262),
.A2(n_251),
.B(n_250),
.Y(n_270)
);

AO21x2_ASAP7_75t_L g271 ( 
.A1(n_258),
.A2(n_241),
.B(n_240),
.Y(n_271)
);

AND2x2_ASAP7_75t_L g272 ( 
.A(n_264),
.B(n_252),
.Y(n_272)
);

AOI33xp33_ASAP7_75t_L g273 ( 
.A1(n_259),
.A2(n_239),
.A3(n_234),
.B1(n_21),
.B2(n_24),
.B3(n_25),
.Y(n_273)
);

AOI22xp33_ASAP7_75t_L g274 ( 
.A1(n_256),
.A2(n_26),
.B1(n_27),
.B2(n_28),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_255),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_261),
.Y(n_276)
);

AND2x2_ASAP7_75t_L g277 ( 
.A(n_263),
.B(n_34),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_266),
.Y(n_278)
);

OA21x2_ASAP7_75t_L g279 ( 
.A1(n_265),
.A2(n_36),
.B(n_37),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_275),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_269),
.B(n_254),
.Y(n_281)
);

AND2x2_ASAP7_75t_L g282 ( 
.A(n_268),
.B(n_276),
.Y(n_282)
);

NAND4xp25_ASAP7_75t_L g283 ( 
.A(n_275),
.B(n_273),
.C(n_278),
.D(n_274),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_272),
.B(n_267),
.Y(n_284)
);

AND2x4_ASAP7_75t_SL g285 ( 
.A(n_269),
.B(n_39),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_278),
.Y(n_286)
);

INVx3_ASAP7_75t_L g287 ( 
.A(n_271),
.Y(n_287)
);

BUFx2_ASAP7_75t_L g288 ( 
.A(n_277),
.Y(n_288)
);

INVx1_ASAP7_75t_SL g289 ( 
.A(n_277),
.Y(n_289)
);

BUFx3_ASAP7_75t_L g290 ( 
.A(n_282),
.Y(n_290)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_281),
.B(n_288),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_280),
.Y(n_292)
);

OR2x2_ASAP7_75t_L g293 ( 
.A(n_289),
.B(n_271),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_286),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_284),
.Y(n_295)
);

HB1xp67_ASAP7_75t_L g296 ( 
.A(n_289),
.Y(n_296)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_287),
.B(n_279),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_287),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_283),
.Y(n_299)
);

AND2x2_ASAP7_75t_L g300 ( 
.A(n_291),
.B(n_285),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_294),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_295),
.B(n_270),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_299),
.B(n_270),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_296),
.Y(n_304)
);

HB1xp67_ASAP7_75t_L g305 ( 
.A(n_293),
.Y(n_305)
);

AND2x2_ASAP7_75t_L g306 ( 
.A(n_290),
.B(n_53),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_292),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_298),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_304),
.Y(n_309)
);

NOR2x1_ASAP7_75t_L g310 ( 
.A(n_303),
.B(n_297),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g311 ( 
.A(n_300),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_301),
.Y(n_312)
);

AND2x2_ASAP7_75t_L g313 ( 
.A(n_310),
.B(n_305),
.Y(n_313)
);

NOR4xp25_ASAP7_75t_SL g314 ( 
.A(n_309),
.B(n_308),
.C(n_307),
.D(n_305),
.Y(n_314)
);

AND2x2_ASAP7_75t_L g315 ( 
.A(n_311),
.B(n_297),
.Y(n_315)
);

NAND4xp75_ASAP7_75t_L g316 ( 
.A(n_313),
.B(n_306),
.C(n_312),
.D(n_301),
.Y(n_316)
);

INVx1_ASAP7_75t_SL g317 ( 
.A(n_316),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_317),
.A2(n_314),
.B1(n_315),
.B2(n_302),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_318),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_L g320 ( 
.A1(n_319),
.A2(n_59),
.B(n_61),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_320),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_321),
.Y(n_322)
);

AOI22xp33_ASAP7_75t_L g323 ( 
.A1(n_322),
.A2(n_62),
.B1(n_69),
.B2(n_72),
.Y(n_323)
);

AOI221xp5_ASAP7_75t_L g324 ( 
.A1(n_323),
.A2(n_74),
.B1(n_75),
.B2(n_77),
.C(n_79),
.Y(n_324)
);


endmodule