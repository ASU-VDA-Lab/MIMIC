module real_jpeg_22720_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_320, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_320;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_13;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_14;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_0),
.A2(n_37),
.B1(n_38),
.B2(n_50),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_0),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_0),
.A2(n_41),
.B1(n_42),
.B2(n_50),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_0),
.A2(n_27),
.B1(n_28),
.B2(n_50),
.Y(n_97)
);

OAI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_0),
.A2(n_21),
.B1(n_22),
.B2(n_50),
.Y(n_100)
);

OAI22xp33_ASAP7_75t_SL g32 ( 
.A1(n_1),
.A2(n_21),
.B1(n_22),
.B2(n_33),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_1),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_1),
.A2(n_33),
.B1(n_41),
.B2(n_42),
.Y(n_59)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_1),
.A2(n_37),
.B(n_80),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_1),
.B(n_37),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_1),
.B(n_73),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_1),
.A2(n_27),
.B1(n_28),
.B2(n_33),
.Y(n_145)
);

AOI21xp33_ASAP7_75t_L g159 ( 
.A1(n_1),
.A2(n_10),
.B(n_27),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_1),
.B(n_54),
.Y(n_180)
);

O2A1O1Ixp33_ASAP7_75t_L g193 ( 
.A1(n_1),
.A2(n_41),
.B(n_56),
.C(n_194),
.Y(n_193)
);

BUFx16f_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_3),
.A2(n_37),
.B1(n_38),
.B2(n_39),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_3),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_3),
.A2(n_27),
.B1(n_28),
.B2(n_39),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_3),
.A2(n_21),
.B1(n_22),
.B2(n_39),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_L g273 ( 
.A1(n_3),
.A2(n_39),
.B1(n_41),
.B2(n_42),
.Y(n_273)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_4),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_4),
.B(n_97),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_4),
.B(n_155),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_4),
.B(n_144),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_5),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_6),
.A2(n_37),
.B1(n_38),
.B2(n_106),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_6),
.Y(n_106)
);

OAI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_6),
.A2(n_41),
.B1(n_42),
.B2(n_106),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_6),
.A2(n_27),
.B1(n_28),
.B2(n_106),
.Y(n_155)
);

OAI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_6),
.A2(n_21),
.B1(n_22),
.B2(n_106),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

INVx13_ASAP7_75t_L g57 ( 
.A(n_8),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_9),
.A2(n_41),
.B1(n_42),
.B2(n_43),
.Y(n_40)
);

INVx13_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_9),
.B(n_37),
.Y(n_48)
);

O2A1O1Ixp33_ASAP7_75t_L g20 ( 
.A1(n_10),
.A2(n_21),
.B(n_25),
.C(n_26),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_10),
.B(n_21),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_10),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_26)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

INVx11_ASAP7_75t_SL g24 ( 
.A(n_11),
.Y(n_24)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_83),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_81),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_SL g14 ( 
.A(n_15),
.B(n_75),
.Y(n_14)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_15),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_66),
.C(n_68),
.Y(n_15)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_16),
.A2(n_17),
.B1(n_314),
.B2(n_316),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_17),
.Y(n_16)
);

MAJIxp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_34),
.C(n_51),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_18),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_18),
.A2(n_108),
.B1(n_109),
.B2(n_110),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_18),
.A2(n_108),
.B1(n_295),
.B2(n_296),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_18),
.A2(n_51),
.B1(n_52),
.B2(n_108),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_SL g18 ( 
.A1(n_19),
.A2(n_30),
.B(n_31),
.Y(n_18)
);

OAI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_19),
.A2(n_99),
.B(n_236),
.Y(n_261)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_20),
.B(n_32),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_20),
.B(n_163),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_20),
.B(n_100),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_21),
.A2(n_22),
.B1(n_56),
.B2(n_58),
.Y(n_55)
);

OAI21xp33_ASAP7_75t_L g194 ( 
.A1(n_21),
.A2(n_33),
.B(n_58),
.Y(n_194)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

A2O1A1Ixp33_ASAP7_75t_L g158 ( 
.A1(n_22),
.A2(n_29),
.B(n_33),
.C(n_159),
.Y(n_158)
);

BUFx10_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_26),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_26),
.B(n_100),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_26),
.B(n_163),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_26),
.B(n_32),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_27),
.B(n_94),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_28),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_28),
.B(n_172),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_30),
.B(n_33),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_30),
.A2(n_199),
.B(n_236),
.Y(n_235)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_33),
.B(n_94),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_34),
.A2(n_35),
.B1(n_303),
.B2(n_304),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_35),
.Y(n_34)
);

OAI21xp5_ASAP7_75t_L g35 ( 
.A1(n_36),
.A2(n_40),
.B(n_44),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_36),
.Y(n_70)
);

A2O1A1Ixp33_ASAP7_75t_L g46 ( 
.A1(n_37),
.A2(n_40),
.B(n_47),
.C(n_48),
.Y(n_46)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_40),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_40),
.B(n_105),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_40),
.A2(n_46),
.B(n_79),
.Y(n_279)
);

A2O1A1Ixp33_ASAP7_75t_L g62 ( 
.A1(n_41),
.A2(n_55),
.B(n_56),
.C(n_63),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_41),
.B(n_56),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_41),
.B(n_43),
.Y(n_129)
);

INVx4_ASAP7_75t_SL g41 ( 
.A(n_42),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_42),
.A2(n_129),
.B1(n_130),
.B2(n_131),
.Y(n_128)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_44),
.B(n_77),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g44 ( 
.A(n_45),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_45),
.B(n_104),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_49),
.Y(n_45)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_46),
.B(n_79),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_48),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_60),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_53),
.B(n_119),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_59),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_54),
.B(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g66 ( 
.A1(n_55),
.A2(n_62),
.B(n_67),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_55),
.B(n_65),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_55),
.A2(n_60),
.B(n_273),
.Y(n_272)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_56),
.Y(n_58)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_59),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_59),
.B(n_61),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_60),
.B(n_111),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_61),
.B(n_64),
.Y(n_60)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_61),
.A2(n_139),
.B(n_297),
.Y(n_296)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_62),
.B(n_121),
.Y(n_120)
);

CKINVDCx14_ASAP7_75t_R g64 ( 
.A(n_65),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_66),
.A2(n_240),
.B1(n_241),
.B2(n_242),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_66),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_66),
.A2(n_68),
.B1(n_242),
.B2(n_315),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_68),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_70),
.B(n_71),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_69),
.B(n_117),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_72),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_72),
.B(n_116),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_72),
.B(n_292),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_74),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_73),
.B(n_78),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_76),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_76),
.B(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_77),
.B(n_116),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_80),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_311),
.B(n_317),
.Y(n_83)
);

OAI321xp33_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_287),
.A3(n_306),
.B1(n_309),
.B2(n_310),
.C(n_320),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_265),
.B(n_286),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_87),
.A2(n_246),
.B(n_264),
.Y(n_86)
);

O2A1O1Ixp33_ASAP7_75t_SL g87 ( 
.A1(n_88),
.A2(n_146),
.B(n_228),
.C(n_245),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_132),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_89),
.B(n_132),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_113),
.Y(n_89)
);

XOR2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_102),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_91),
.B(n_102),
.C(n_113),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_98),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_92),
.B(n_98),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_93),
.A2(n_95),
.B(n_96),
.Y(n_92)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_93),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_93),
.A2(n_94),
.B(n_145),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_94),
.A2(n_95),
.B(n_125),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_96),
.B(n_143),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_96),
.B(n_168),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_97),
.B(n_126),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_101),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_99),
.B(n_183),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_101),
.B(n_162),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_108),
.C(n_109),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_103),
.B(n_134),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_107),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_105),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g292 ( 
.A(n_107),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_108),
.B(n_291),
.C(n_296),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_110),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_111),
.B(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_112),
.Y(n_121)
);

CKINVDCx5p33_ASAP7_75t_R g113 ( 
.A(n_114),
.Y(n_113)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_114),
.Y(n_243)
);

FAx1_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_118),
.CI(n_122),
.CON(n_114),
.SN(n_114)
);

CKINVDCx14_ASAP7_75t_R g119 ( 
.A(n_120),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_120),
.B(n_139),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_123),
.B(n_127),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_123),
.A2(n_124),
.B1(n_127),
.B2(n_128),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_124),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_125),
.B(n_154),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_125),
.B(n_185),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_126),
.B(n_144),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_126),
.B(n_155),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_128),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_135),
.C(n_136),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_133),
.B(n_224),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_135),
.A2(n_136),
.B1(n_137),
.B2(n_225),
.Y(n_224)
);

CKINVDCx14_ASAP7_75t_R g225 ( 
.A(n_135),
.Y(n_225)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_140),
.C(n_141),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_SL g210 ( 
.A(n_138),
.B(n_211),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_139),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_140),
.A2(n_141),
.B1(n_142),
.B2(n_212),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_140),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_142),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_143),
.B(n_154),
.Y(n_170)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_147),
.B(n_227),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_148),
.A2(n_221),
.B(n_226),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_149),
.A2(n_206),
.B(n_220),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_150),
.A2(n_187),
.B(n_205),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_151),
.A2(n_175),
.B(n_186),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_164),
.B(n_174),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_156),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_153),
.B(n_156),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_158),
.B1(n_160),
.B2(n_161),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_158),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_158),
.B(n_160),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_161),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_162),
.B(n_199),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_165),
.A2(n_169),
.B(n_173),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_167),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_166),
.B(n_167),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_168),
.B(n_185),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_170),
.B(n_171),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_177),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_176),
.B(n_177),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_184),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_179),
.A2(n_180),
.B1(n_181),
.B2(n_182),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_179),
.B(n_182),
.C(n_184),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_180),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_182),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_183),
.B(n_216),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_189),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_188),
.B(n_189),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_190),
.A2(n_196),
.B1(n_197),
.B2(n_204),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_190),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_191),
.A2(n_192),
.B1(n_193),
.B2(n_195),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_191),
.A2(n_192),
.B1(n_261),
.B2(n_262),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_191),
.A2(n_192),
.B1(n_278),
.B2(n_279),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_L g298 ( 
.A1(n_191),
.A2(n_279),
.B(n_281),
.Y(n_298)
);

CKINVDCx16_ASAP7_75t_R g191 ( 
.A(n_192),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_192),
.B(n_193),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_192),
.B(n_261),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_193),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_198),
.A2(n_200),
.B1(n_201),
.B2(n_203),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_198),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_199),
.B(n_216),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_200),
.B(n_203),
.C(n_204),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_201),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_202),
.B(n_257),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_208),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_207),
.B(n_208),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_209),
.A2(n_210),
.B1(n_213),
.B2(n_214),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_209),
.B(n_215),
.C(n_219),
.Y(n_222)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_215),
.A2(n_217),
.B1(n_218),
.B2(n_219),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_215),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_217),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_223),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_222),
.B(n_223),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_230),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_229),
.B(n_230),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_231),
.A2(n_232),
.B1(n_243),
.B2(n_244),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_237),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_233),
.B(n_237),
.C(n_244),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_235),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_234),
.B(n_235),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_239),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_238),
.B(n_241),
.C(n_242),
.Y(n_263)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

CKINVDCx16_ASAP7_75t_R g244 ( 
.A(n_243),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_248),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_247),
.B(n_248),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_263),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_250),
.A2(n_251),
.B1(n_259),
.B2(n_260),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_250),
.B(n_260),
.C(n_263),
.Y(n_266)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_253),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_252),
.B(n_254),
.C(n_258),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_254),
.A2(n_255),
.B1(n_256),
.B2(n_258),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_255),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_256),
.Y(n_258)
);

CKINVDCx16_ASAP7_75t_R g259 ( 
.A(n_260),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_261),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_267),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_266),
.B(n_267),
.Y(n_286)
);

AOI22xp33_ASAP7_75t_SL g267 ( 
.A1(n_268),
.A2(n_269),
.B1(n_284),
.B2(n_285),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_270),
.A2(n_275),
.B1(n_282),
.B2(n_283),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_270),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_270),
.B(n_283),
.C(n_285),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_271),
.A2(n_272),
.B(n_274),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_271),
.B(n_272),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_273),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_274),
.B(n_289),
.C(n_298),
.Y(n_288)
);

FAx1_ASAP7_75t_SL g308 ( 
.A(n_274),
.B(n_289),
.CI(n_298),
.CON(n_308),
.SN(n_308)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_275),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_276),
.A2(n_277),
.B1(n_280),
.B2(n_281),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_276),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_277),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_279),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_284),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_299),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_288),
.B(n_299),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_290),
.A2(n_291),
.B1(n_293),
.B2(n_294),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_290),
.A2(n_291),
.B1(n_301),
.B2(n_302),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_291),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_291),
.B(n_301),
.C(n_305),
.Y(n_312)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_296),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_305),
.Y(n_299)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_304),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_308),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_307),
.B(n_308),
.Y(n_309)
);

BUFx24_ASAP7_75t_SL g318 ( 
.A(n_308),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_312),
.B(n_313),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_312),
.B(n_313),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_314),
.Y(n_316)
);


endmodule