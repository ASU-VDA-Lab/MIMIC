module fake_jpeg_14711_n_333 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_333);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_333;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_3),
.Y(n_16)
);

INVx6_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx14_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

CKINVDCx14_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

INVx2_ASAP7_75t_SL g35 ( 
.A(n_7),
.Y(n_35)
);

CKINVDCx16_ASAP7_75t_R g36 ( 
.A(n_19),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_36),
.B(n_38),
.Y(n_51)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_34),
.B(n_8),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

HAxp5_ASAP7_75t_SL g40 ( 
.A(n_16),
.B(n_0),
.CON(n_40),
.SN(n_40)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_40),
.B(n_42),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_43),
.Y(n_46)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

BUFx4f_ASAP7_75t_L g45 ( 
.A(n_26),
.Y(n_45)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_45),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_39),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_48),
.B(n_50),
.Y(n_68)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_45),
.Y(n_49)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_39),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_45),
.B(n_0),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_53),
.A2(n_28),
.B(n_18),
.Y(n_103)
);

HB1xp67_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_54),
.Y(n_94)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_55),
.Y(n_71)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_56),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_38),
.B(n_40),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_58),
.B(n_18),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_37),
.A2(n_17),
.B1(n_35),
.B2(n_34),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_60),
.A2(n_35),
.B1(n_17),
.B2(n_30),
.Y(n_75)
);

OAI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_42),
.A2(n_17),
.B1(n_31),
.B2(n_30),
.Y(n_63)
);

OAI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_63),
.A2(n_42),
.B1(n_17),
.B2(n_30),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_38),
.B(n_24),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_64),
.B(n_66),
.Y(n_95)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_65),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_36),
.B(n_20),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_36),
.B(n_20),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_67),
.B(n_18),
.Y(n_100)
);

AND2x2_ASAP7_75t_SL g69 ( 
.A(n_58),
.B(n_45),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_69),
.B(n_96),
.C(n_39),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_64),
.B(n_24),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_70),
.B(n_83),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_57),
.B(n_51),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_72),
.B(n_101),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_74),
.A2(n_99),
.B1(n_28),
.B2(n_37),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_75),
.A2(n_56),
.B1(n_49),
.B2(n_65),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_57),
.A2(n_44),
.B1(n_42),
.B2(n_34),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_76),
.A2(n_85),
.B1(n_93),
.B2(n_37),
.Y(n_108)
);

HB1xp67_ASAP7_75t_L g77 ( 
.A(n_62),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_77),
.B(n_80),
.Y(n_116)
);

HB1xp67_ASAP7_75t_L g80 ( 
.A(n_62),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_52),
.Y(n_81)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_81),
.Y(n_114)
);

INVx2_ASAP7_75t_SL g82 ( 
.A(n_59),
.Y(n_82)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_82),
.Y(n_118)
);

INVx1_ASAP7_75t_SL g83 ( 
.A(n_61),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_52),
.Y(n_84)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_84),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_51),
.A2(n_31),
.B1(n_44),
.B2(n_27),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_46),
.Y(n_86)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_86),
.Y(n_132)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_46),
.Y(n_87)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_87),
.Y(n_111)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_66),
.Y(n_88)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_88),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_67),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_89),
.B(n_90),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_59),
.B(n_31),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_59),
.B(n_35),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_91),
.B(n_92),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_48),
.B(n_35),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_47),
.A2(n_44),
.B1(n_27),
.B2(n_42),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_53),
.B(n_27),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_55),
.Y(n_97)
);

INVx11_ASAP7_75t_L g135 ( 
.A(n_97),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_53),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_98),
.Y(n_137)
);

OAI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_53),
.A2(n_37),
.B1(n_22),
.B2(n_16),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_SL g117 ( 
.A(n_100),
.B(n_103),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_50),
.B(n_19),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_55),
.B(n_19),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_102),
.B(n_56),
.Y(n_113)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_61),
.Y(n_104)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_104),
.Y(n_136)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_61),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_105),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_54),
.B(n_22),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_106),
.Y(n_130)
);

XNOR2x1_ASAP7_75t_L g129 ( 
.A(n_107),
.B(n_33),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_108),
.B(n_76),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_110),
.A2(n_124),
.B1(n_23),
.B2(n_82),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_113),
.B(n_119),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_72),
.B(n_96),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_115),
.B(n_127),
.C(n_103),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_69),
.B(n_65),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_69),
.A2(n_0),
.B(n_1),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_120),
.A2(n_100),
.B(n_95),
.Y(n_154)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_81),
.Y(n_126)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_126),
.Y(n_145)
);

INVx2_ASAP7_75t_SL g128 ( 
.A(n_82),
.Y(n_128)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_128),
.Y(n_139)
);

NAND2xp33_ASAP7_75t_SL g153 ( 
.A(n_129),
.B(n_102),
.Y(n_153)
);

A2O1A1Ixp33_ASAP7_75t_L g131 ( 
.A1(n_98),
.A2(n_23),
.B(n_16),
.C(n_8),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_131),
.B(n_134),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_101),
.B(n_47),
.Y(n_134)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_135),
.Y(n_138)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_138),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_141),
.B(n_25),
.C(n_29),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_137),
.A2(n_107),
.B(n_68),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_142),
.A2(n_153),
.B(n_154),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_143),
.A2(n_148),
.B1(n_149),
.B2(n_157),
.Y(n_170)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_134),
.Y(n_144)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_144),
.Y(n_176)
);

BUFx2_ASAP7_75t_L g146 ( 
.A(n_136),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_146),
.B(n_155),
.Y(n_173)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_128),
.Y(n_147)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_147),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_119),
.A2(n_47),
.B1(n_68),
.B2(n_49),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_127),
.A2(n_107),
.B1(n_89),
.B2(n_88),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_128),
.Y(n_150)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_150),
.Y(n_186)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_123),
.Y(n_151)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_151),
.Y(n_193)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_123),
.Y(n_152)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_152),
.Y(n_194)
);

HB1xp67_ASAP7_75t_L g155 ( 
.A(n_118),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_130),
.B(n_95),
.Y(n_156)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_156),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_113),
.A2(n_94),
.B1(n_84),
.B2(n_79),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_114),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_158),
.B(n_167),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_137),
.A2(n_117),
.B1(n_129),
.B2(n_133),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_159),
.Y(n_202)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_126),
.Y(n_160)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_160),
.Y(n_195)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_111),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_161),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_162),
.A2(n_163),
.B1(n_165),
.B2(n_132),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_109),
.A2(n_94),
.B1(n_79),
.B2(n_73),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_130),
.B(n_121),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g198 ( 
.A(n_164),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_109),
.A2(n_73),
.B1(n_78),
.B2(n_87),
.Y(n_165)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_112),
.Y(n_166)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_166),
.Y(n_203)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_112),
.Y(n_167)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_111),
.Y(n_169)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_169),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_144),
.B(n_120),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_172),
.B(n_174),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_140),
.B(n_115),
.Y(n_174)
);

AND2x6_ASAP7_75t_L g175 ( 
.A(n_141),
.B(n_117),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_175),
.Y(n_204)
);

NOR2x1_ASAP7_75t_L g177 ( 
.A(n_168),
.B(n_131),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_177),
.B(n_149),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_140),
.B(n_125),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_178),
.B(n_184),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_159),
.A2(n_133),
.B1(n_108),
.B2(n_122),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_181),
.A2(n_187),
.B(n_23),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_165),
.B(n_121),
.Y(n_182)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_182),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_157),
.B(n_154),
.Y(n_184)
);

OA21x2_ASAP7_75t_L g187 ( 
.A1(n_148),
.A2(n_116),
.B(n_163),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_145),
.B(n_118),
.Y(n_188)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_188),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_138),
.B(n_135),
.Y(n_189)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_189),
.Y(n_219)
);

OAI22xp33_ASAP7_75t_L g191 ( 
.A1(n_151),
.A2(n_105),
.B1(n_78),
.B2(n_83),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_191),
.A2(n_104),
.B1(n_41),
.B2(n_43),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_160),
.B(n_114),
.Y(n_196)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_196),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_152),
.B(n_132),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_197),
.B(n_200),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_199),
.A2(n_43),
.B1(n_33),
.B2(n_32),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_167),
.B(n_112),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_201),
.B(n_142),
.C(n_150),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_206),
.A2(n_177),
.B(n_187),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_209),
.B(n_210),
.C(n_211),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_174),
.B(n_139),
.C(n_147),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_201),
.B(n_139),
.C(n_169),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_171),
.B(n_97),
.C(n_71),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_212),
.B(n_213),
.C(n_216),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_171),
.B(n_71),
.C(n_41),
.Y(n_213)
);

AO21x1_ASAP7_75t_L g250 ( 
.A1(n_214),
.A2(n_179),
.B(n_186),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_202),
.A2(n_166),
.B1(n_86),
.B2(n_136),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_215),
.A2(n_183),
.B1(n_203),
.B2(n_199),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_184),
.B(n_146),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_178),
.B(n_41),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_217),
.B(n_221),
.Y(n_241)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_218),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_175),
.B(n_41),
.C(n_43),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_190),
.B(n_2),
.Y(n_222)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_222),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_195),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_223),
.B(n_232),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_172),
.B(n_43),
.C(n_39),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_225),
.B(n_231),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_226),
.A2(n_193),
.B1(n_194),
.B2(n_203),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_198),
.B(n_2),
.Y(n_228)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_228),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_181),
.B(n_25),
.Y(n_229)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_229),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_SL g230 ( 
.A(n_170),
.B(n_25),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_230),
.A2(n_183),
.B1(n_194),
.B2(n_193),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_170),
.B(n_43),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_202),
.B(n_33),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_233),
.A2(n_243),
.B1(n_246),
.B2(n_192),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_215),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_234),
.B(n_252),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_205),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_235),
.B(n_252),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_214),
.A2(n_187),
.B(n_197),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_236),
.A2(n_250),
.B(n_173),
.Y(n_260)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_238),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_242),
.B(n_212),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_207),
.A2(n_227),
.B1(n_221),
.B2(n_204),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_208),
.B(n_224),
.Y(n_251)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_251),
.Y(n_263)
);

OR2x2_ASAP7_75t_L g252 ( 
.A(n_227),
.B(n_176),
.Y(n_252)
);

INVx1_ASAP7_75t_SL g253 ( 
.A(n_219),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_253),
.B(n_192),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_231),
.A2(n_176),
.B1(n_185),
.B2(n_186),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_254),
.A2(n_225),
.B1(n_213),
.B2(n_220),
.Y(n_257)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_216),
.Y(n_255)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_255),
.Y(n_264)
);

A2O1A1Ixp33_ASAP7_75t_SL g256 ( 
.A1(n_229),
.A2(n_185),
.B(n_195),
.C(n_191),
.Y(n_256)
);

AOI22x1_ASAP7_75t_L g267 ( 
.A1(n_256),
.A2(n_250),
.B1(n_238),
.B2(n_242),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_257),
.B(n_275),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_258),
.B(n_241),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_240),
.B(n_211),
.C(n_245),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_259),
.B(n_265),
.C(n_276),
.Y(n_280)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_260),
.Y(n_279)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_261),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_240),
.B(n_210),
.C(n_209),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_234),
.A2(n_220),
.B1(n_230),
.B2(n_232),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_266),
.A2(n_267),
.B1(n_256),
.B2(n_239),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_269),
.A2(n_239),
.B1(n_256),
.B2(n_243),
.Y(n_286)
);

HB1xp67_ASAP7_75t_L g270 ( 
.A(n_248),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_270),
.B(n_272),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_253),
.B(n_180),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_271),
.B(n_272),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_237),
.B(n_217),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_273),
.B(n_274),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_254),
.B(n_218),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_249),
.B(n_11),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_245),
.B(n_33),
.C(n_32),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_277),
.B(n_290),
.Y(n_303)
);

NOR2xp67_ASAP7_75t_L g278 ( 
.A(n_267),
.B(n_233),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g300 ( 
.A1(n_278),
.A2(n_286),
.B1(n_32),
.B2(n_29),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_259),
.B(n_241),
.C(n_248),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_281),
.B(n_283),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_265),
.B(n_244),
.C(n_247),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_258),
.B(n_247),
.C(n_236),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_284),
.B(n_289),
.Y(n_298)
);

AOI221xp5_ASAP7_75t_L g304 ( 
.A1(n_285),
.A2(n_32),
.B1(n_29),
.B2(n_26),
.C(n_5),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_287),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_276),
.B(n_257),
.C(n_264),
.Y(n_289)
);

A2O1A1Ixp33_ASAP7_75t_L g290 ( 
.A1(n_260),
.A2(n_256),
.B(n_10),
.C(n_12),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_279),
.A2(n_267),
.B1(n_262),
.B2(n_268),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_293),
.B(n_296),
.C(n_295),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_291),
.A2(n_268),
.B(n_262),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_294),
.A2(n_300),
.B1(n_304),
.B2(n_2),
.Y(n_309)
);

A2O1A1Ixp33_ASAP7_75t_SL g295 ( 
.A1(n_290),
.A2(n_266),
.B(n_264),
.C(n_263),
.Y(n_295)
);

AND2x2_ASAP7_75t_L g311 ( 
.A(n_295),
.B(n_277),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_288),
.A2(n_9),
.B1(n_15),
.B2(n_14),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_292),
.B(n_10),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_297),
.B(n_302),
.Y(n_308)
);

NAND2xp33_ASAP7_75t_SL g299 ( 
.A(n_282),
.B(n_8),
.Y(n_299)
);

OR2x2_ASAP7_75t_L g310 ( 
.A(n_299),
.B(n_306),
.Y(n_310)
);

BUFx3_ASAP7_75t_L g302 ( 
.A(n_289),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_283),
.B(n_7),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_SL g307 ( 
.A1(n_298),
.A2(n_280),
.B(n_284),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_SL g321 ( 
.A1(n_307),
.A2(n_6),
.B(n_14),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_309),
.B(n_314),
.Y(n_317)
);

AOI322xp5_ASAP7_75t_L g319 ( 
.A1(n_311),
.A2(n_313),
.A3(n_315),
.B1(n_294),
.B2(n_295),
.C1(n_304),
.C2(n_310),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_305),
.B(n_280),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_312),
.B(n_13),
.Y(n_323)
);

NOR2xp67_ASAP7_75t_SL g313 ( 
.A(n_302),
.B(n_281),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_L g314 ( 
.A1(n_301),
.A2(n_7),
.B(n_15),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_303),
.B(n_6),
.Y(n_315)
);

AND2x2_ASAP7_75t_L g318 ( 
.A(n_315),
.B(n_308),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_316),
.B(n_29),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_318),
.A2(n_319),
.B1(n_13),
.B2(n_14),
.Y(n_324)
);

NOR2x1_ASAP7_75t_L g320 ( 
.A(n_311),
.B(n_6),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_L g327 ( 
.A1(n_320),
.A2(n_322),
.B1(n_323),
.B2(n_2),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_321),
.B(n_26),
.C(n_3),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_324),
.B(n_325),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_323),
.B(n_318),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_SL g329 ( 
.A1(n_326),
.A2(n_327),
.B(n_317),
.Y(n_329)
);

AOI31xp33_ASAP7_75t_L g330 ( 
.A1(n_329),
.A2(n_326),
.A3(n_325),
.B(n_5),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_330),
.B(n_328),
.Y(n_331)
);

MAJx2_ASAP7_75t_L g332 ( 
.A(n_331),
.B(n_4),
.C(n_5),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_R g333 ( 
.A(n_332),
.B(n_4),
.Y(n_333)
);


endmodule