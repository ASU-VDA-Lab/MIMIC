module real_jpeg_5725_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_13;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_176;
wire n_166;
wire n_312;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_14;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx8_ASAP7_75t_L g48 ( 
.A(n_0),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_1),
.A2(n_37),
.B1(n_38),
.B2(n_41),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_1),
.A2(n_37),
.B1(n_45),
.B2(n_49),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_1),
.A2(n_83),
.B1(n_86),
.B2(n_87),
.Y(n_82)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_1),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_1),
.A2(n_114),
.B1(n_116),
.B2(n_117),
.Y(n_113)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_1),
.Y(n_116)
);

O2A1O1Ixp33_ASAP7_75t_L g199 ( 
.A1(n_1),
.A2(n_200),
.B(n_203),
.C(n_206),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_1),
.B(n_214),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_1),
.B(n_73),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_1),
.B(n_57),
.C(n_243),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_1),
.B(n_251),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_1),
.B(n_108),
.C(n_263),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_1),
.B(n_119),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_2),
.A2(n_152),
.B1(n_154),
.B2(n_155),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_2),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g20 ( 
.A1(n_3),
.A2(n_21),
.B1(n_22),
.B2(n_25),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_3),
.A2(n_21),
.B1(n_177),
.B2(n_181),
.Y(n_176)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_4),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_4),
.Y(n_153)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_5),
.Y(n_95)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g186 ( 
.A(n_6),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_6),
.Y(n_214)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_7),
.Y(n_123)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_7),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_7),
.Y(n_202)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_8),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_9),
.A2(n_75),
.B1(n_78),
.B2(n_79),
.Y(n_74)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_9),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g134 ( 
.A1(n_9),
.A2(n_78),
.B1(n_114),
.B2(n_135),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_9),
.A2(n_78),
.B1(n_164),
.B2(n_169),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_9),
.A2(n_31),
.B1(n_78),
.B2(n_212),
.Y(n_211)
);

BUFx5_ASAP7_75t_L g115 ( 
.A(n_10),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_10),
.Y(n_117)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_10),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_10),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_10),
.Y(n_137)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_10),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_11),
.Y(n_57)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_11),
.Y(n_59)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_11),
.Y(n_64)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_217),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_215),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_SL g14 ( 
.A(n_15),
.B(n_188),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_15),
.B(n_188),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_139),
.Y(n_15)
);

MAJIxp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_80),
.C(n_112),
.Y(n_16)
);

INVxp67_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_18),
.B(n_191),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_42),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_19),
.A2(n_42),
.B1(n_239),
.B2(n_306),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_19),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_26),
.B(n_28),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_20),
.Y(n_149)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_22),
.Y(n_25)
);

BUFx2_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

BUFx8_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_27),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_35),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_29),
.A2(n_149),
.B1(n_150),
.B2(n_157),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_29),
.B(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_30),
.A2(n_36),
.B1(n_211),
.B2(n_214),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_30),
.A2(n_36),
.B1(n_211),
.B2(n_232),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_34),
.Y(n_30)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_31),
.Y(n_229)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_33),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_36),
.B(n_184),
.Y(n_264)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_40),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_42),
.A2(n_239),
.B1(n_240),
.B2(n_244),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_42),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_42),
.A2(n_161),
.B1(n_162),
.B2(n_239),
.Y(n_266)
);

AND2x2_ASAP7_75t_SL g42 ( 
.A(n_43),
.B(n_72),
.Y(n_42)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_43),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_53),
.Y(n_43)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_44),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_44),
.B(n_290),
.Y(n_289)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_47),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_47),
.Y(n_79)
);

INVx6_ASAP7_75t_L g180 ( 
.A(n_47),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_47),
.Y(n_241)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_48),
.Y(n_52)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_48),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_48),
.Y(n_109)
);

INVx5_ASAP7_75t_SL g49 ( 
.A(n_50),
.Y(n_49)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_53),
.Y(n_145)
);

NOR2x1_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_62),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_56),
.B1(n_58),
.B2(n_60),
.Y(n_54)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_62),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_63),
.A2(n_65),
.B1(n_66),
.B2(n_70),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_64),
.Y(n_71)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_69),
.Y(n_156)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_74),
.Y(n_72)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_73),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_73),
.A2(n_176),
.B(n_182),
.Y(n_175)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_74),
.Y(n_144)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_80),
.A2(n_112),
.B1(n_192),
.B2(n_193),
.Y(n_191)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_80),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_89),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

OA22x2_ASAP7_75t_L g162 ( 
.A1(n_82),
.A2(n_90),
.B1(n_101),
.B2(n_163),
.Y(n_162)
);

OA22x2_ASAP7_75t_L g197 ( 
.A1(n_82),
.A2(n_90),
.B1(n_101),
.B2(n_163),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_83),
.A2(n_120),
.B1(n_121),
.B2(n_122),
.Y(n_119)
);

INVx5_ASAP7_75t_L g205 ( 
.A(n_83),
.Y(n_205)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_85),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_85),
.Y(n_168)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_85),
.Y(n_171)
);

OAI21xp33_ASAP7_75t_L g203 ( 
.A1(n_86),
.A2(n_201),
.B(n_204),
.Y(n_203)
);

BUFx5_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_88),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_88),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_88),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_90),
.B(n_101),
.Y(n_89)
);

NAND2x1_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_101),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_92),
.A2(n_96),
.B1(n_98),
.B2(n_100),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_94),
.Y(n_111)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_95),
.Y(n_99)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_95),
.Y(n_107)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_97),
.Y(n_261)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_101),
.Y(n_251)
);

AOI22x1_ASAP7_75t_L g101 ( 
.A1(n_102),
.A2(n_105),
.B1(n_108),
.B2(n_110),
.Y(n_101)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_104),
.Y(n_181)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx8_ASAP7_75t_L g263 ( 
.A(n_106),
.Y(n_263)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx2_ASAP7_75t_SL g192 ( 
.A(n_112),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_112),
.A2(n_192),
.B1(n_287),
.B2(n_288),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_112),
.B(n_162),
.C(n_289),
.Y(n_307)
);

OA22x2_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_118),
.B1(n_134),
.B2(n_138),
.Y(n_112)
);

OA22x2_ASAP7_75t_L g160 ( 
.A1(n_113),
.A2(n_118),
.B1(n_134),
.B2(n_138),
.Y(n_160)
);

INVx8_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

OR2x2_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_124),
.Y(n_118)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_119),
.Y(n_138)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_123),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_L g124 ( 
.A1(n_125),
.A2(n_127),
.B1(n_130),
.B2(n_132),
.Y(n_124)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx8_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_173),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_159),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_142),
.B(n_148),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_142),
.A2(n_143),
.B1(n_148),
.B2(n_195),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_142),
.A2(n_143),
.B1(n_250),
.B2(n_252),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_142),
.A2(n_143),
.B1(n_271),
.B2(n_272),
.Y(n_270)
);

INVx2_ASAP7_75t_SL g142 ( 
.A(n_143),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_143),
.B(n_210),
.C(n_250),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_143),
.B(n_271),
.C(n_273),
.Y(n_284)
);

OA22x2_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_145),
.B1(n_146),
.B2(n_147),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_145),
.B(n_146),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_148),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_151),
.B(n_184),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_153),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_153),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_160),
.A2(n_161),
.B1(n_162),
.B2(n_172),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_160),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_160),
.B(n_197),
.C(n_198),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_160),
.A2(n_172),
.B1(n_197),
.B2(n_279),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_161),
.B(n_239),
.C(n_258),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_161),
.A2(n_162),
.B1(n_289),
.B2(n_291),
.Y(n_288)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_162),
.Y(n_161)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_174),
.A2(n_175),
.B1(n_183),
.B2(n_187),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx6_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_183),
.Y(n_187)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_185),
.Y(n_232)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_194),
.C(n_196),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_190),
.B(n_194),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_196),
.B(n_313),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_197),
.A2(n_275),
.B1(n_276),
.B2(n_279),
.Y(n_274)
);

CKINVDCx16_ASAP7_75t_R g279 ( 
.A(n_197),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_198),
.B(n_303),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_209),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_199),
.A2(n_209),
.B1(n_210),
.B2(n_297),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_199),
.Y(n_297)
);

INVx6_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx4_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx2_ASAP7_75t_SL g206 ( 
.A(n_207),
.Y(n_206)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_209),
.A2(n_210),
.B1(n_248),
.B2(n_249),
.Y(n_247)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_210),
.B(n_234),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_210),
.B(n_234),
.Y(n_235)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_218),
.A2(n_299),
.B(n_314),
.Y(n_217)
);

HB1xp67_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_220),
.A2(n_283),
.B(n_298),
.Y(n_219)
);

AOI21x1_ASAP7_75t_L g220 ( 
.A1(n_221),
.A2(n_268),
.B(n_282),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_222),
.A2(n_255),
.B(n_267),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_223),
.A2(n_246),
.B(n_254),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_224),
.A2(n_236),
.B(n_245),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_225),
.A2(n_233),
.B(n_235),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_231),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_230),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx1_ASAP7_75t_SL g228 ( 
.A(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_231),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_231),
.A2(n_237),
.B1(n_277),
.B2(n_278),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_238),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_237),
.B(n_238),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_237),
.B(n_277),
.C(n_279),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_239),
.B(n_244),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g244 ( 
.A(n_240),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_242),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_247),
.B(n_253),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_247),
.B(n_253),
.Y(n_254)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_250),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_257),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_256),
.B(n_257),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_266),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_259),
.A2(n_260),
.B1(n_264),
.B2(n_265),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_259),
.B(n_265),
.Y(n_271)
);

CKINVDCx16_ASAP7_75t_R g259 ( 
.A(n_260),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_262),
.Y(n_260)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_264),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_269),
.B(n_281),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_269),
.B(n_281),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_270),
.A2(n_273),
.B1(n_274),
.B2(n_280),
.Y(n_269)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_270),
.Y(n_280)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_271),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

CKINVDCx14_ASAP7_75t_R g277 ( 
.A(n_278),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_285),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_284),
.B(n_285),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_292),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_286),
.B(n_294),
.C(n_295),
.Y(n_308)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_289),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_293),
.A2(n_294),
.B1(n_295),
.B2(n_296),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

NOR2x1_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_309),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_301),
.B(n_308),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_301),
.B(n_308),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_304),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g311 ( 
.A(n_302),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_307),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_305),
.B(n_307),
.C(n_311),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_L g314 ( 
.A1(n_309),
.A2(n_315),
.B(n_316),
.Y(n_314)
);

AND2x2_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_312),
.Y(n_309)
);

OR2x2_ASAP7_75t_L g316 ( 
.A(n_310),
.B(n_312),
.Y(n_316)
);


endmodule