module fake_jpeg_18861_n_319 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_319);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_319;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx16f_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx16f_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_0),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_18),
.B(n_1),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_37),
.B(n_38),
.Y(n_46)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_18),
.B(n_1),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_32),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_39),
.B(n_17),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_43),
.B(n_44),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_35),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_35),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_45),
.B(n_51),
.Y(n_79)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_47),
.Y(n_75)
);

HB1xp67_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_48),
.Y(n_68)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_37),
.B(n_17),
.Y(n_52)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_52),
.Y(n_87)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_55),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_37),
.B(n_32),
.Y(n_59)
);

XOR2xp5_ASAP7_75t_L g74 ( 
.A(n_59),
.B(n_63),
.Y(n_74)
);

HB1xp67_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_60),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_36),
.B(n_26),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_61),
.Y(n_93)
);

AND2x2_ASAP7_75t_SL g62 ( 
.A(n_40),
.B(n_21),
.Y(n_62)
);

OR2x4_ASAP7_75t_L g64 ( 
.A(n_62),
.B(n_36),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_40),
.B(n_32),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_64),
.B(n_32),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_52),
.A2(n_30),
.B1(n_24),
.B2(n_31),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_65),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_51),
.A2(n_42),
.B1(n_30),
.B2(n_22),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_67),
.A2(n_83),
.B1(n_84),
.B2(n_58),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_47),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_69),
.B(n_85),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_43),
.A2(n_30),
.B1(n_24),
.B2(n_42),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_70),
.A2(n_82),
.B1(n_86),
.B2(n_89),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_53),
.Y(n_72)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_72),
.Y(n_103)
);

BUFx2_ASAP7_75t_SL g73 ( 
.A(n_53),
.Y(n_73)
);

INVx1_ASAP7_75t_SL g109 ( 
.A(n_73),
.Y(n_109)
);

A2O1A1Ixp33_ASAP7_75t_L g77 ( 
.A1(n_46),
.A2(n_31),
.B(n_28),
.C(n_24),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_77),
.B(n_32),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_56),
.A2(n_17),
.B1(n_26),
.B2(n_22),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_78),
.Y(n_100)
);

AO22x2_ASAP7_75t_L g81 ( 
.A1(n_62),
.A2(n_56),
.B1(n_63),
.B2(n_46),
.Y(n_81)
);

OA22x2_ASAP7_75t_L g98 ( 
.A1(n_81),
.A2(n_45),
.B1(n_54),
.B2(n_49),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_56),
.A2(n_26),
.B1(n_22),
.B2(n_31),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_59),
.A2(n_28),
.B1(n_20),
.B2(n_25),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_61),
.A2(n_28),
.B1(n_20),
.B2(n_25),
.Y(n_84)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_58),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_62),
.A2(n_33),
.B1(n_23),
.B2(n_25),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_62),
.A2(n_20),
.B1(n_33),
.B2(n_23),
.Y(n_88)
);

INVx1_ASAP7_75t_SL g112 ( 
.A(n_88),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_58),
.A2(n_33),
.B1(n_23),
.B2(n_29),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_55),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_90),
.B(n_91),
.Y(n_121)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_54),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g92 ( 
.A(n_44),
.B(n_29),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_92),
.B(n_32),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_95),
.A2(n_108),
.B1(n_110),
.B2(n_94),
.Y(n_128)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_75),
.Y(n_96)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_96),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_97),
.B(n_98),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_93),
.B(n_57),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_99),
.B(n_104),
.Y(n_133)
);

AO21x2_ASAP7_75t_SL g101 ( 
.A1(n_64),
.A2(n_53),
.B(n_50),
.Y(n_101)
);

AO21x1_ASAP7_75t_L g124 ( 
.A1(n_101),
.A2(n_106),
.B(n_107),
.Y(n_124)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_75),
.Y(n_102)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_102),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_93),
.B(n_87),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_79),
.Y(n_105)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_105),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_84),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_110),
.B(n_114),
.Y(n_140)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_79),
.Y(n_113)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_113),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_88),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_66),
.Y(n_115)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_115),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_74),
.B(n_54),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_116),
.B(n_119),
.Y(n_135)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_66),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_117),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_68),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_118),
.B(n_90),
.Y(n_138)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_72),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_67),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_120),
.B(n_71),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_120),
.A2(n_81),
.B1(n_65),
.B2(n_87),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_122),
.A2(n_134),
.B1(n_142),
.B2(n_146),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_116),
.B(n_74),
.C(n_92),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_123),
.B(n_126),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_114),
.A2(n_81),
.B(n_77),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_126),
.A2(n_139),
.B(n_1),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_128),
.A2(n_132),
.B1(n_143),
.B2(n_145),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_121),
.Y(n_129)
);

INVx13_ASAP7_75t_L g168 ( 
.A(n_129),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_95),
.A2(n_81),
.B1(n_83),
.B2(n_68),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_L g134 ( 
.A1(n_112),
.A2(n_81),
.B1(n_85),
.B2(n_71),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_136),
.B(n_141),
.Y(n_167)
);

CKINVDCx14_ASAP7_75t_R g182 ( 
.A(n_138),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_94),
.A2(n_21),
.B(n_19),
.Y(n_139)
);

OAI32xp33_ASAP7_75t_L g141 ( 
.A1(n_105),
.A2(n_57),
.A3(n_76),
.B1(n_27),
.B2(n_29),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_113),
.A2(n_112),
.B1(n_117),
.B2(n_115),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_106),
.A2(n_80),
.B1(n_91),
.B2(n_76),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_106),
.A2(n_100),
.B1(n_107),
.B2(n_101),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_100),
.A2(n_80),
.B1(n_27),
.B2(n_29),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_111),
.B(n_19),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_147),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_97),
.B(n_32),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_148),
.B(n_151),
.Y(n_170)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_98),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_149),
.B(n_98),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_101),
.A2(n_11),
.B1(n_15),
.B2(n_3),
.Y(n_151)
);

INVx1_ASAP7_75t_SL g152 ( 
.A(n_125),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_152),
.B(n_161),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_153),
.B(n_154),
.Y(n_188)
);

AND2x2_ASAP7_75t_SL g154 ( 
.A(n_127),
.B(n_98),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_150),
.B(n_96),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_155),
.B(n_156),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_150),
.B(n_102),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_133),
.B(n_119),
.Y(n_158)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_158),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_133),
.B(n_103),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_159),
.B(n_171),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_149),
.B(n_145),
.Y(n_160)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_160),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_136),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_125),
.Y(n_162)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_162),
.Y(n_193)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_130),
.Y(n_164)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_164),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_140),
.B(n_101),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_165),
.B(n_178),
.Y(n_199)
);

INVxp67_ASAP7_75t_SL g166 ( 
.A(n_129),
.Y(n_166)
);

INVxp67_ASAP7_75t_SL g194 ( 
.A(n_166),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_140),
.A2(n_109),
.B(n_103),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_169),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_142),
.B(n_109),
.Y(n_171)
);

AND2x6_ASAP7_75t_L g173 ( 
.A(n_124),
.B(n_50),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_173),
.B(n_174),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_130),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_131),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_175),
.B(n_176),
.Y(n_210)
);

INVx2_ASAP7_75t_SL g176 ( 
.A(n_141),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_177),
.B(n_148),
.C(n_122),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_135),
.B(n_27),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_179),
.A2(n_165),
.B1(n_170),
.B2(n_161),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_132),
.B(n_19),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_180),
.B(n_181),
.Y(n_197)
);

AND2x6_ASAP7_75t_L g181 ( 
.A(n_124),
.B(n_50),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_124),
.A2(n_127),
.B(n_143),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_183),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_135),
.B(n_1),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_184),
.B(n_2),
.Y(n_202)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_131),
.Y(n_185)
);

CKINVDCx16_ASAP7_75t_R g201 ( 
.A(n_185),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_SL g187 ( 
.A(n_177),
.B(n_123),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_187),
.B(n_203),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_176),
.A2(n_128),
.B1(n_137),
.B2(n_144),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_189),
.A2(n_208),
.B1(n_213),
.B2(n_155),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_190),
.B(n_204),
.C(n_206),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_157),
.A2(n_144),
.B1(n_137),
.B2(n_151),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_192),
.A2(n_205),
.B1(n_175),
.B2(n_174),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_202),
.B(n_184),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_183),
.B(n_139),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_154),
.B(n_19),
.C(n_16),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_157),
.A2(n_160),
.B1(n_176),
.B2(n_154),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_178),
.B(n_19),
.C(n_16),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_167),
.A2(n_16),
.B1(n_21),
.B2(n_2),
.Y(n_208)
);

HB1xp67_ASAP7_75t_L g209 ( 
.A(n_173),
.Y(n_209)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_209),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_167),
.B(n_16),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_211),
.B(n_3),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_186),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_215),
.B(n_217),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_214),
.A2(n_181),
.B(n_160),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_216),
.B(n_235),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_218),
.A2(n_234),
.B1(n_239),
.B2(n_199),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_187),
.B(n_179),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_219),
.B(n_211),
.Y(n_242)
);

AND2x6_ASAP7_75t_L g220 ( 
.A(n_207),
.B(n_169),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_220),
.B(n_237),
.Y(n_256)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_193),
.Y(n_221)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_221),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_193),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_222),
.B(n_227),
.Y(n_243)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_212),
.Y(n_223)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_223),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_190),
.B(n_172),
.C(n_185),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_225),
.B(n_236),
.C(n_206),
.Y(n_251)
);

AO22x1_ASAP7_75t_L g226 ( 
.A1(n_188),
.A2(n_170),
.B1(n_172),
.B2(n_156),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_226),
.B(n_232),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_195),
.B(n_182),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_196),
.B(n_168),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_228),
.B(n_233),
.Y(n_244)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_212),
.Y(n_231)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_231),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_198),
.B(n_163),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_197),
.A2(n_163),
.B1(n_152),
.B2(n_162),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_202),
.B(n_168),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_203),
.B(n_164),
.C(n_4),
.Y(n_236)
);

INVx1_ASAP7_75t_SL g237 ( 
.A(n_194),
.Y(n_237)
);

FAx1_ASAP7_75t_SL g255 ( 
.A(n_238),
.B(n_208),
.CI(n_192),
.CON(n_255),
.SN(n_255)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_198),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_240),
.A2(n_232),
.B1(n_210),
.B2(n_214),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_242),
.B(n_251),
.Y(n_273)
);

HB1xp67_ASAP7_75t_L g245 ( 
.A(n_220),
.Y(n_245)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_245),
.Y(n_267)
);

HB1xp67_ASAP7_75t_L g249 ( 
.A(n_216),
.Y(n_249)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_249),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_236),
.A2(n_200),
.B1(n_204),
.B2(n_191),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_252),
.A2(n_224),
.B(n_229),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_230),
.B(n_189),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_253),
.B(n_254),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_230),
.B(n_205),
.Y(n_254)
);

MAJx2_ASAP7_75t_L g266 ( 
.A(n_255),
.B(n_238),
.C(n_225),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_219),
.B(n_199),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_257),
.B(n_218),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_224),
.B(n_191),
.C(n_188),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_258),
.B(n_226),
.C(n_237),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_260),
.B(n_262),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_244),
.B(n_217),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_243),
.B(n_201),
.Y(n_263)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_263),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_241),
.B(n_221),
.Y(n_264)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_264),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_259),
.B(n_223),
.Y(n_265)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_265),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_L g285 ( 
.A1(n_266),
.A2(n_271),
.B(n_252),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_268),
.A2(n_258),
.B1(n_266),
.B2(n_267),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_269),
.B(n_270),
.Y(n_279)
);

A2O1A1Ixp33_ASAP7_75t_SL g271 ( 
.A1(n_255),
.A2(n_3),
.B(n_5),
.C(n_6),
.Y(n_271)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_246),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_274),
.B(n_275),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_251),
.B(n_5),
.C(n_7),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_SL g277 ( 
.A(n_270),
.B(n_242),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_277),
.B(n_278),
.Y(n_298)
);

OAI21x1_ASAP7_75t_L g278 ( 
.A1(n_271),
.A2(n_250),
.B(n_256),
.Y(n_278)
);

FAx1_ASAP7_75t_SL g280 ( 
.A(n_261),
.B(n_253),
.CI(n_254),
.CON(n_280),
.SN(n_280)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_280),
.B(n_284),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_282),
.A2(n_9),
.B(n_11),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_272),
.B(n_247),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_285),
.A2(n_271),
.B(n_247),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_275),
.B(n_257),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_288),
.B(n_286),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_290),
.B(n_280),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_281),
.A2(n_248),
.B1(n_271),
.B2(n_255),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_291),
.B(n_292),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_285),
.A2(n_273),
.B(n_8),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_283),
.B(n_273),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_293),
.B(n_294),
.Y(n_305)
);

NAND3xp33_ASAP7_75t_SL g294 ( 
.A(n_287),
.B(n_5),
.C(n_8),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_295),
.A2(n_296),
.B(n_297),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_L g297 ( 
.A1(n_282),
.A2(n_9),
.B(n_12),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_279),
.B(n_9),
.C(n_12),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_299),
.B(n_13),
.Y(n_306)
);

NOR2xp67_ASAP7_75t_L g300 ( 
.A(n_289),
.B(n_276),
.Y(n_300)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_300),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_293),
.B(n_277),
.C(n_280),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_303),
.B(n_306),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_304),
.B(n_13),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_SL g307 ( 
.A1(n_298),
.A2(n_13),
.B(n_14),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_SL g312 ( 
.A1(n_307),
.A2(n_14),
.B(n_15),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_305),
.B(n_294),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_309),
.B(n_312),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_311),
.B(n_302),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_L g316 ( 
.A1(n_313),
.A2(n_315),
.B(n_310),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_308),
.B(n_301),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_316),
.B(n_311),
.C(n_314),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_317),
.A2(n_303),
.B1(n_304),
.B2(n_14),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_318),
.B(n_15),
.Y(n_319)
);


endmodule