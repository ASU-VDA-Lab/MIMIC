module fake_jpeg_1181_n_329 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_329);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_329;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_260;
wire n_199;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx5_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_11),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_10),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_12),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_13),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_4),
.Y(n_37)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_6),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_5),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

INVx4_ASAP7_75t_SL g99 ( 
.A(n_42),
.Y(n_99)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_43),
.Y(n_78)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_44),
.Y(n_87)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

INVx11_ASAP7_75t_L g109 ( 
.A(n_45),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_20),
.B(n_22),
.Y(n_46)
);

OR2x2_ASAP7_75t_L g68 ( 
.A(n_46),
.B(n_48),
.Y(n_68)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_47),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_20),
.B(n_8),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_22),
.B(n_9),
.Y(n_49)
);

OR2x2_ASAP7_75t_L g97 ( 
.A(n_49),
.B(n_52),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_17),
.Y(n_51)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_28),
.B(n_7),
.Y(n_52)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_53),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_18),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_54),
.Y(n_81)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

HB1xp67_ASAP7_75t_L g82 ( 
.A(n_55),
.Y(n_82)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_19),
.Y(n_56)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_56),
.Y(n_84)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_18),
.Y(n_57)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_57),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_28),
.B(n_7),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_58),
.B(n_31),
.Y(n_93)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_27),
.Y(n_59)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_59),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_19),
.B(n_0),
.Y(n_60)
);

AND2x2_ASAP7_75t_SL g69 ( 
.A(n_60),
.B(n_32),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_18),
.Y(n_61)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_61),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_46),
.B(n_41),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_62),
.B(n_70),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_48),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_63),
.B(n_71),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_60),
.B(n_29),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_67),
.B(n_95),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_69),
.B(n_76),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_49),
.B(n_52),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_58),
.Y(n_71)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_73),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_54),
.A2(n_35),
.B1(n_25),
.B2(n_30),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_74),
.A2(n_77),
.B1(n_106),
.B2(n_32),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_42),
.B(n_41),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_75),
.B(n_83),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_60),
.B(n_32),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_61),
.A2(n_25),
.B1(n_30),
.B2(n_35),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_44),
.A2(n_39),
.B1(n_38),
.B2(n_24),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_80),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_50),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_45),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_85),
.B(n_91),
.Y(n_127)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_47),
.Y(n_88)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_88),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_59),
.A2(n_39),
.B1(n_38),
.B2(n_24),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_89),
.Y(n_123)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_50),
.Y(n_90)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_90),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_42),
.B(n_40),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_42),
.B(n_36),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_92),
.B(n_93),
.Y(n_141)
);

BUFx12f_ASAP7_75t_L g94 ( 
.A(n_54),
.Y(n_94)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_94),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_55),
.B(n_36),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_56),
.B(n_40),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_96),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_43),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_98),
.B(n_100),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_53),
.B(n_31),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_57),
.Y(n_101)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_101),
.Y(n_133)
);

A2O1A1Ixp33_ASAP7_75t_L g102 ( 
.A1(n_57),
.A2(n_37),
.B(n_33),
.C(n_17),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_102),
.B(n_108),
.Y(n_142)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_61),
.Y(n_103)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_103),
.Y(n_110)
);

BUFx12f_ASAP7_75t_L g104 ( 
.A(n_50),
.Y(n_104)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_104),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_57),
.A2(n_35),
.B1(n_25),
.B2(n_30),
.Y(n_106)
);

OA22x2_ASAP7_75t_L g107 ( 
.A1(n_57),
.A2(n_38),
.B1(n_24),
.B2(n_39),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_107),
.A2(n_23),
.B1(n_26),
.B2(n_21),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_46),
.B(n_37),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_111),
.A2(n_112),
.B1(n_123),
.B2(n_140),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_82),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_114),
.B(n_134),
.Y(n_175)
);

BUFx12_ASAP7_75t_L g115 ( 
.A(n_99),
.Y(n_115)
);

BUFx12f_ASAP7_75t_L g153 ( 
.A(n_115),
.Y(n_153)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_86),
.Y(n_116)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_116),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_63),
.A2(n_33),
.B1(n_23),
.B2(n_32),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_118),
.A2(n_135),
.B1(n_99),
.B2(n_106),
.Y(n_146)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_86),
.Y(n_119)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_119),
.Y(n_155)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_101),
.Y(n_122)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_122),
.Y(n_166)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_65),
.Y(n_125)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_125),
.Y(n_167)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_65),
.Y(n_126)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_126),
.Y(n_168)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_73),
.Y(n_130)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_130),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_64),
.Y(n_134)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_105),
.Y(n_137)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_137),
.Y(n_165)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_88),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_138),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_64),
.Y(n_139)
);

OAI21xp33_ASAP7_75t_L g177 ( 
.A1(n_139),
.A2(n_144),
.B(n_81),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_69),
.B(n_26),
.C(n_21),
.Y(n_140)
);

MAJx2_ASAP7_75t_L g154 ( 
.A(n_140),
.B(n_69),
.C(n_76),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_72),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_146),
.B(n_159),
.Y(n_210)
);

AOI21xp33_ASAP7_75t_L g147 ( 
.A1(n_113),
.A2(n_67),
.B(n_102),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_147),
.B(n_172),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_142),
.A2(n_107),
.B1(n_76),
.B2(n_71),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_148),
.A2(n_149),
.B1(n_156),
.B2(n_161),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_142),
.A2(n_97),
.B1(n_68),
.B2(n_107),
.Y(n_149)
);

INVx5_ASAP7_75t_L g151 ( 
.A(n_120),
.Y(n_151)
);

HB1xp67_ASAP7_75t_L g189 ( 
.A(n_151),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_154),
.B(n_84),
.C(n_143),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_L g156 ( 
.A1(n_112),
.A2(n_83),
.B1(n_107),
.B2(n_87),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_127),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_157),
.B(n_176),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_137),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_158),
.B(n_162),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_123),
.A2(n_98),
.B1(n_105),
.B2(n_78),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_110),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_160),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_135),
.A2(n_97),
.B1(n_68),
.B2(n_103),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_113),
.B(n_136),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_124),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_163),
.B(n_164),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_136),
.B(n_79),
.Y(n_164)
);

AND2x2_ASAP7_75t_SL g169 ( 
.A(n_132),
.B(n_79),
.Y(n_169)
);

CKINVDCx14_ASAP7_75t_R g213 ( 
.A(n_169),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_170),
.A2(n_179),
.B1(n_181),
.B2(n_109),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_129),
.B(n_66),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_171),
.B(n_116),
.Y(n_185)
);

NOR2xp67_ASAP7_75t_L g172 ( 
.A(n_117),
.B(n_141),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_132),
.A2(n_78),
.B(n_66),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_173),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_115),
.Y(n_176)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_177),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_132),
.A2(n_129),
.B(n_145),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_178),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_128),
.A2(n_125),
.B1(n_130),
.B2(n_126),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_128),
.A2(n_72),
.B1(n_81),
.B2(n_87),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_180),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_133),
.A2(n_90),
.B1(n_84),
.B2(n_94),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_148),
.A2(n_133),
.B1(n_110),
.B2(n_131),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_182),
.A2(n_184),
.B1(n_150),
.B2(n_174),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_162),
.A2(n_138),
.B1(n_131),
.B2(n_122),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_185),
.B(n_192),
.Y(n_222)
);

AO22x1_ASAP7_75t_SL g187 ( 
.A1(n_169),
.A2(n_119),
.B1(n_94),
.B2(n_104),
.Y(n_187)
);

AND2x2_ASAP7_75t_L g218 ( 
.A(n_187),
.B(n_197),
.Y(n_218)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_160),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_190),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_164),
.B(n_163),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_175),
.B(n_120),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_193),
.B(n_202),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_180),
.A2(n_121),
.B1(n_143),
.B2(n_109),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_195),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_171),
.B(n_121),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_198),
.B(n_158),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_200),
.B(n_155),
.Y(n_227)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_168),
.Y(n_201)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_201),
.Y(n_216)
);

A2O1A1Ixp33_ASAP7_75t_L g202 ( 
.A1(n_178),
.A2(n_115),
.B(n_11),
.C(n_13),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_173),
.Y(n_203)
);

BUFx3_ASAP7_75t_L g229 ( 
.A(n_203),
.Y(n_229)
);

O2A1O1Ixp33_ASAP7_75t_L g204 ( 
.A1(n_159),
.A2(n_104),
.B(n_94),
.C(n_2),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_204),
.A2(n_165),
.B(n_1),
.Y(n_232)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_168),
.Y(n_205)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_205),
.Y(n_217)
);

BUFx12f_ASAP7_75t_L g206 ( 
.A(n_153),
.Y(n_206)
);

INVx13_ASAP7_75t_L g239 ( 
.A(n_206),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_L g207 ( 
.A1(n_174),
.A2(n_104),
.B1(n_1),
.B2(n_2),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_207),
.A2(n_212),
.B1(n_0),
.B2(n_1),
.Y(n_237)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_166),
.Y(n_209)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_209),
.Y(n_221)
);

NAND3xp33_ASAP7_75t_L g214 ( 
.A(n_186),
.B(n_179),
.C(n_154),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_214),
.B(n_215),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_188),
.B(n_153),
.Y(n_215)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_219),
.Y(n_251)
);

OR2x2_ASAP7_75t_L g223 ( 
.A(n_191),
.B(n_150),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_223),
.B(n_226),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_210),
.A2(n_169),
.B1(n_181),
.B2(n_167),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_224),
.A2(n_225),
.B1(n_231),
.B2(n_233),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_210),
.A2(n_151),
.B1(n_155),
.B2(n_152),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g226 ( 
.A(n_189),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_227),
.B(n_187),
.Y(n_253)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_228),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_211),
.B(n_153),
.Y(n_230)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_230),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_210),
.A2(n_152),
.B1(n_165),
.B2(n_153),
.Y(n_231)
);

AND2x2_ASAP7_75t_L g257 ( 
.A(n_232),
.B(n_206),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_192),
.A2(n_10),
.B1(n_16),
.B2(n_3),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_196),
.A2(n_10),
.B1(n_16),
.B2(n_5),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_235),
.A2(n_237),
.B1(n_238),
.B2(n_212),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_182),
.A2(n_5),
.B1(n_6),
.B2(n_13),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_L g263 ( 
.A1(n_240),
.A2(n_244),
.B1(n_232),
.B2(n_236),
.Y(n_263)
);

FAx1_ASAP7_75t_SL g241 ( 
.A(n_222),
.B(n_191),
.CI(n_200),
.CON(n_241),
.SN(n_241)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_241),
.B(n_260),
.Y(n_270)
);

HB1xp67_ASAP7_75t_L g242 ( 
.A(n_221),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_242),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_227),
.B(n_208),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_243),
.B(n_255),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_235),
.A2(n_199),
.B1(n_183),
.B2(n_203),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_218),
.A2(n_213),
.B1(n_183),
.B2(n_185),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_245),
.B(n_249),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_222),
.B(n_184),
.C(n_198),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_246),
.B(n_247),
.C(n_253),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_223),
.B(n_228),
.C(n_218),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_218),
.A2(n_187),
.B1(n_204),
.B2(n_205),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_SL g254 ( 
.A1(n_234),
.A2(n_202),
.B(n_201),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_254),
.A2(n_231),
.B(n_233),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_219),
.B(n_190),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_224),
.B(n_194),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_256),
.B(n_220),
.Y(n_275)
);

OAI22x1_ASAP7_75t_L g276 ( 
.A1(n_257),
.A2(n_206),
.B1(n_239),
.B2(n_194),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_220),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_263),
.A2(n_264),
.B1(n_271),
.B2(n_252),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_248),
.B(n_217),
.Y(n_265)
);

HB1xp67_ASAP7_75t_L g285 ( 
.A(n_265),
.Y(n_285)
);

OA21x2_ASAP7_75t_SL g266 ( 
.A1(n_241),
.A2(n_229),
.B(n_221),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_266),
.B(n_259),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_258),
.B(n_217),
.Y(n_268)
);

CKINVDCx16_ASAP7_75t_R g280 ( 
.A(n_268),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_243),
.B(n_229),
.C(n_216),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_269),
.B(n_253),
.C(n_247),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_251),
.A2(n_236),
.B1(n_238),
.B2(n_216),
.Y(n_271)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_255),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_273),
.A2(n_274),
.B1(n_276),
.B2(n_277),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_246),
.B(n_225),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_275),
.B(n_250),
.Y(n_283)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_251),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_278),
.B(n_290),
.Y(n_295)
);

NOR2xp67_ASAP7_75t_SL g294 ( 
.A(n_279),
.B(n_287),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_262),
.B(n_256),
.C(n_245),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_281),
.B(n_289),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_282),
.A2(n_261),
.B1(n_271),
.B2(n_288),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_283),
.B(n_286),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_264),
.A2(n_252),
.B1(n_257),
.B2(n_254),
.Y(n_284)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_284),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_262),
.B(n_241),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_SL g287 ( 
.A(n_272),
.B(n_249),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_272),
.B(n_257),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_269),
.B(n_239),
.C(n_6),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_SL g291 ( 
.A(n_270),
.B(n_15),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_291),
.B(n_268),
.Y(n_298)
);

CKINVDCx16_ASAP7_75t_R g293 ( 
.A(n_285),
.Y(n_293)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_293),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_280),
.A2(n_261),
.B1(n_277),
.B2(n_274),
.Y(n_297)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_297),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_298),
.B(n_301),
.Y(n_304)
);

HB1xp67_ASAP7_75t_L g308 ( 
.A(n_300),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_278),
.B(n_266),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_290),
.Y(n_302)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_302),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_L g303 ( 
.A1(n_294),
.A2(n_281),
.B(n_286),
.Y(n_303)
);

AOI21xp33_ASAP7_75t_L g313 ( 
.A1(n_303),
.A2(n_306),
.B(n_307),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_L g306 ( 
.A1(n_301),
.A2(n_283),
.B(n_265),
.Y(n_306)
);

AOI221xp5_ASAP7_75t_L g307 ( 
.A1(n_299),
.A2(n_287),
.B1(n_273),
.B2(n_267),
.C(n_291),
.Y(n_307)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_300),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_310),
.B(n_298),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_312),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_309),
.A2(n_296),
.B1(n_267),
.B2(n_276),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_314),
.B(n_315),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_308),
.A2(n_311),
.B1(n_307),
.B2(n_305),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_L g316 ( 
.A1(n_308),
.A2(n_292),
.B(n_275),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_316),
.B(n_318),
.C(n_292),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_304),
.B(n_295),
.Y(n_317)
);

BUFx5_ASAP7_75t_L g320 ( 
.A(n_317),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_309),
.B(n_295),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_322),
.B(n_314),
.Y(n_323)
);

NAND4xp25_ASAP7_75t_SL g325 ( 
.A(n_323),
.B(n_324),
.C(n_320),
.D(n_313),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_321),
.B(n_315),
.C(n_316),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_325),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_326),
.B(n_320),
.C(n_322),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_327),
.B(n_319),
.Y(n_328)
);

HB1xp67_ASAP7_75t_L g329 ( 
.A(n_328),
.Y(n_329)
);


endmodule