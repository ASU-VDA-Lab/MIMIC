module real_jpeg_261_n_25 (n_17, n_8, n_0, n_21, n_141, n_2, n_139, n_142, n_143, n_10, n_137, n_9, n_12, n_135, n_24, n_6, n_136, n_23, n_11, n_14, n_138, n_7, n_22, n_18, n_3, n_145, n_144, n_5, n_4, n_1, n_20, n_19, n_140, n_16, n_15, n_13, n_25);

input n_17;
input n_8;
input n_0;
input n_21;
input n_141;
input n_2;
input n_139;
input n_142;
input n_143;
input n_10;
input n_137;
input n_9;
input n_12;
input n_135;
input n_24;
input n_6;
input n_136;
input n_23;
input n_11;
input n_14;
input n_138;
input n_7;
input n_22;
input n_18;
input n_3;
input n_145;
input n_144;
input n_5;
input n_4;
input n_1;
input n_20;
input n_19;
input n_140;
input n_16;
input n_15;
input n_13;

output n_25;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_78;
wire n_83;
wire n_104;
wire n_64;
wire n_47;
wire n_131;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_126;
wire n_120;
wire n_113;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_118;
wire n_123;
wire n_116;
wire n_50;
wire n_69;
wire n_31;
wire n_129;
wire n_72;
wire n_100;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_30;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;

INVx1_ASAP7_75t_L g85 ( 
.A(n_0),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_SL g64 ( 
.A1(n_1),
.A2(n_65),
.B(n_69),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_2),
.A2(n_56),
.B1(n_89),
.B2(n_92),
.Y(n_55)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_2),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_3),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_4),
.B(n_58),
.C(n_82),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_5),
.Y(n_121)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_6),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_7),
.B(n_66),
.Y(n_65)
);

AO22x1_ASAP7_75t_L g60 ( 
.A1(n_8),
.A2(n_61),
.B1(n_63),
.B2(n_74),
.Y(n_60)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_8),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_9),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_10),
.Y(n_131)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx16f_ASAP7_75t_L g68 ( 
.A(n_11),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_11),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_12),
.B(n_98),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_12),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_13),
.B(n_101),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_13),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_14),
.Y(n_29)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_15),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_16),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_17),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_18),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_18),
.B(n_38),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_19),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_20),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_20),
.B(n_52),
.Y(n_96)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_21),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_22),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_23),
.A2(n_27),
.B1(n_28),
.B2(n_32),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_23),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_24),
.B(n_60),
.C(n_75),
.Y(n_59)
);

XNOR2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_33),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_28),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_30),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_30),
.B(n_48),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_30),
.B(n_53),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_30),
.B(n_88),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_30),
.B(n_93),
.Y(n_92)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

INVx6_ASAP7_75t_SL g81 ( 
.A(n_31),
.Y(n_81)
);

INVx4_ASAP7_75t_SL g84 ( 
.A(n_31),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_SL g33 ( 
.A1(n_34),
.A2(n_126),
.B(n_132),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

A2O1A1Ixp33_ASAP7_75t_L g35 ( 
.A1(n_36),
.A2(n_37),
.B(n_43),
.C(n_125),
.Y(n_35)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_40),
.Y(n_38)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx13_ASAP7_75t_L g103 ( 
.A(n_41),
.Y(n_103)
);

CKINVDCx6p67_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_42),
.B(n_62),
.Y(n_61)
);

BUFx10_ASAP7_75t_L g109 ( 
.A(n_42),
.Y(n_109)
);

MAJx2_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_121),
.C(n_122),
.Y(n_43)
);

AOI21xp5_ASAP7_75t_L g44 ( 
.A1(n_45),
.A2(n_50),
.B(n_120),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_46),
.B(n_49),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_46),
.B(n_49),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g46 ( 
.A(n_47),
.Y(n_46)
);

OAI221xp5_ASAP7_75t_L g50 ( 
.A1(n_51),
.A2(n_54),
.B1(n_55),
.B2(n_94),
.C(n_110),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_85),
.C(n_86),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_77),
.C(n_78),
.Y(n_58)
);

NAND3xp33_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_72),
.C(n_73),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_64),
.B(n_72),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_65),
.B(n_69),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_68),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_68),
.B(n_76),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_68),
.B(n_99),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_71),
.Y(n_69)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_81),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_84),
.Y(n_82)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_91),
.Y(n_89)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_95),
.B(n_104),
.Y(n_94)
);

AOI322xp5_ASAP7_75t_L g110 ( 
.A1(n_95),
.A2(n_111),
.A3(n_112),
.B1(n_115),
.B2(n_116),
.C1(n_119),
.C2(n_145),
.Y(n_110)
);

NOR3xp33_ASAP7_75t_SL g95 ( 
.A(n_96),
.B(n_97),
.C(n_100),
.Y(n_95)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_96),
.Y(n_115)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_98),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_100),
.Y(n_111)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_101),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_103),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_103),
.B(n_124),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_103),
.B(n_130),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_106),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_105),
.B(n_106),
.Y(n_119)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_109),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_114),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_118),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_123),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_128),
.B(n_131),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_128),
.B(n_131),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_129),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_135),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_136),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_137),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_138),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_139),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_140),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_141),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_142),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_143),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_144),
.Y(n_108)
);


endmodule