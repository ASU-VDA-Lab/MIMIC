module real_jpeg_3438_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_320, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_320;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_176;
wire n_166;
wire n_312;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_1),
.A2(n_26),
.B1(n_27),
.B2(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_1),
.A2(n_35),
.B1(n_49),
.B2(n_50),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_1),
.A2(n_35),
.B1(n_42),
.B2(n_46),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_1),
.A2(n_32),
.B1(n_33),
.B2(n_35),
.Y(n_164)
);

BUFx5_ASAP7_75t_L g104 ( 
.A(n_2),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_3),
.A2(n_26),
.B1(n_27),
.B2(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_3),
.A2(n_32),
.B1(n_33),
.B2(n_37),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_3),
.A2(n_37),
.B1(n_42),
.B2(n_46),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_3),
.A2(n_37),
.B1(n_49),
.B2(n_50),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_4),
.A2(n_49),
.B1(n_50),
.B2(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_4),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_4),
.A2(n_32),
.B1(n_33),
.B2(n_54),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_4),
.A2(n_42),
.B1(n_46),
.B2(n_54),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_4),
.A2(n_26),
.B1(n_27),
.B2(n_54),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_5),
.A2(n_26),
.B1(n_27),
.B2(n_146),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_5),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_5),
.A2(n_49),
.B1(n_50),
.B2(n_146),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_5),
.A2(n_42),
.B1(n_46),
.B2(n_146),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_5),
.A2(n_32),
.B1(n_33),
.B2(n_146),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_6),
.A2(n_26),
.B1(n_27),
.B2(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_6),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_6),
.A2(n_49),
.B1(n_50),
.B2(n_117),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_6),
.A2(n_42),
.B1(n_46),
.B2(n_117),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_L g237 ( 
.A1(n_6),
.A2(n_32),
.B1(n_33),
.B2(n_117),
.Y(n_237)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_7),
.Y(n_64)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx10_ASAP7_75t_L g45 ( 
.A(n_9),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_11),
.A2(n_32),
.B1(n_33),
.B2(n_67),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_11),
.Y(n_67)
);

OAI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_11),
.A2(n_26),
.B1(n_27),
.B2(n_67),
.Y(n_75)
);

OAI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_11),
.A2(n_42),
.B1(n_46),
.B2(n_67),
.Y(n_108)
);

OAI22xp33_ASAP7_75t_L g112 ( 
.A1(n_11),
.A2(n_49),
.B1(n_50),
.B2(n_67),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_13),
.A2(n_26),
.B1(n_27),
.B2(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_13),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_13),
.A2(n_32),
.B1(n_33),
.B2(n_119),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_13),
.A2(n_42),
.B1(n_46),
.B2(n_119),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_13),
.A2(n_49),
.B1(n_50),
.B2(n_119),
.Y(n_221)
);

CKINVDCx14_ASAP7_75t_R g137 ( 
.A(n_14),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_14),
.B(n_42),
.C(n_45),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_14),
.A2(n_49),
.B1(n_50),
.B2(n_137),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_14),
.B(n_104),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_14),
.B(n_40),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_14),
.B(n_33),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_14),
.A2(n_33),
.B(n_215),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_14),
.B(n_88),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_14),
.A2(n_26),
.B(n_252),
.Y(n_251)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_15),
.Y(n_51)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_92),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_90),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_81),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_20),
.B(n_81),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_72),
.C(n_76),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_21),
.A2(n_22),
.B1(n_72),
.B2(n_304),
.Y(n_303)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_38),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_23),
.B(n_39),
.C(n_56),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_31),
.B1(n_34),
.B2(n_36),
.Y(n_23)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_24),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_24),
.A2(n_36),
.B(n_87),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_24),
.A2(n_31),
.B1(n_116),
.B2(n_118),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_24),
.A2(n_31),
.B1(n_116),
.B2(n_145),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_24),
.A2(n_118),
.B(n_161),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_24),
.A2(n_31),
.B1(n_145),
.B2(n_251),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_24),
.A2(n_87),
.B(n_290),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_31),
.Y(n_24)
);

OAI22xp33_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_27),
.B1(n_29),
.B2(n_30),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_27),
.B(n_137),
.Y(n_136)
);

NAND3xp33_ASAP7_75t_L g138 ( 
.A(n_27),
.B(n_30),
.C(n_33),
.Y(n_138)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_29),
.Y(n_30)
);

OA22x2_ASAP7_75t_L g31 ( 
.A1(n_29),
.A2(n_30),
.B1(n_32),
.B2(n_33),
.Y(n_31)
);

A2O1A1Ixp33_ASAP7_75t_L g135 ( 
.A1(n_29),
.A2(n_32),
.B(n_136),
.C(n_138),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g72 ( 
.A1(n_31),
.A2(n_34),
.B(n_73),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_31),
.Y(n_88)
);

CKINVDCx6p67_ASAP7_75t_R g33 ( 
.A(n_32),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_32),
.A2(n_33),
.B1(n_62),
.B2(n_63),
.Y(n_70)
);

OAI32xp33_ASAP7_75t_L g213 ( 
.A1(n_33),
.A2(n_50),
.A3(n_63),
.B1(n_214),
.B2(n_216),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_55),
.B1(n_56),
.B2(n_71),
.Y(n_38)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_39),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_39),
.B(n_72),
.C(n_77),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_39),
.A2(n_71),
.B1(n_77),
.B2(n_309),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_47),
.B(n_52),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_40),
.B(n_112),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_40),
.A2(n_47),
.B1(n_180),
.B2(n_181),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_40),
.A2(n_47),
.B1(n_180),
.B2(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_41),
.B(n_48),
.Y(n_47)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_41),
.A2(n_110),
.B(n_111),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_41),
.A2(n_110),
.B1(n_130),
.B2(n_131),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_41),
.A2(n_130),
.B1(n_220),
.B2(n_221),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_41),
.B(n_53),
.Y(n_231)
);

OA22x2_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_44),
.B1(n_45),
.B2(n_46),
.Y(n_41)
);

INVx4_ASAP7_75t_SL g46 ( 
.A(n_42),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_42),
.B(n_103),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_42),
.B(n_193),
.Y(n_192)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

OAI22xp33_ASAP7_75t_L g48 ( 
.A1(n_44),
.A2(n_45),
.B1(n_49),
.B2(n_50),
.Y(n_48)
);

INVx13_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_47),
.B(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_SL g130 ( 
.A(n_47),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_47),
.A2(n_230),
.B(n_231),
.Y(n_229)
);

OA22x2_ASAP7_75t_SL g61 ( 
.A1(n_49),
.A2(n_50),
.B1(n_62),
.B2(n_63),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_49),
.B(n_62),
.Y(n_216)
);

CKINVDCx6p67_ASAP7_75t_R g49 ( 
.A(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_50),
.B(n_185),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_SL g255 ( 
.A1(n_53),
.A2(n_130),
.B(n_155),
.Y(n_255)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_65),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_57),
.A2(n_69),
.B(n_143),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_58),
.B(n_60),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g58 ( 
.A(n_59),
.Y(n_58)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_59),
.A2(n_61),
.B(n_69),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_59),
.A2(n_69),
.B(n_80),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_60),
.B(n_66),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_60),
.A2(n_68),
.B1(n_235),
.B2(n_236),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_60),
.A2(n_68),
.B1(n_78),
.B2(n_296),
.Y(n_295)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_61),
.B(n_70),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_61),
.A2(n_65),
.B(n_164),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_61),
.B(n_137),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_61),
.A2(n_69),
.B1(n_223),
.B2(n_224),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_61),
.A2(n_69),
.B1(n_143),
.B2(n_237),
.Y(n_254)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_68),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_68),
.A2(n_78),
.B(n_79),
.Y(n_77)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_72),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_72),
.A2(n_304),
.B1(n_307),
.B2(n_308),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_74),
.B(n_75),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_75),
.B(n_88),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_76),
.B(n_303),
.Y(n_302)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_77),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_89),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_84),
.B1(n_85),
.B2(n_86),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_84),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_86),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_88),
.B(n_162),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_SL g92 ( 
.A1(n_93),
.A2(n_300),
.B(n_314),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_SL g93 ( 
.A1(n_94),
.A2(n_280),
.B(n_299),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g94 ( 
.A1(n_95),
.A2(n_168),
.B(n_279),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_147),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_96),
.B(n_147),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_121),
.C(n_132),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_97),
.B(n_121),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_99),
.B1(n_113),
.B2(n_114),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_98),
.B(n_115),
.C(n_120),
.Y(n_148)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_109),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_100),
.B(n_109),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_101),
.A2(n_105),
.B(n_107),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_101),
.A2(n_103),
.B(n_125),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_101),
.A2(n_103),
.B1(n_203),
.B2(n_204),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_101),
.A2(n_107),
.B(n_125),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_102),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_102),
.B(n_108),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_102),
.A2(n_104),
.B1(n_106),
.B2(n_140),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_102),
.A2(n_124),
.B(n_176),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_102),
.A2(n_104),
.B1(n_137),
.B2(n_195),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_102),
.A2(n_104),
.B1(n_195),
.B2(n_198),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_103),
.B(n_125),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_103),
.A2(n_127),
.B(n_141),
.Y(n_242)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_104),
.B(n_108),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVxp33_ASAP7_75t_L g294 ( 
.A(n_111),
.Y(n_294)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_120),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_123),
.B1(n_128),
.B2(n_129),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_122),
.B(n_129),
.Y(n_165)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_124),
.B(n_126),
.Y(n_123)
);

INVxp33_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_130),
.A2(n_131),
.B(n_155),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_132),
.B(n_264),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_142),
.C(n_144),
.Y(n_132)
);

FAx1_ASAP7_75t_SL g267 ( 
.A(n_133),
.B(n_142),
.CI(n_144),
.CON(n_267),
.SN(n_267)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_139),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_134),
.A2(n_135),
.B1(n_139),
.B2(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g252 ( 
.A(n_136),
.Y(n_252)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_139),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_148),
.A2(n_149),
.B1(n_150),
.B2(n_167),
.Y(n_147)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_148),
.Y(n_167)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_SL g150 ( 
.A(n_151),
.B(n_157),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_151),
.B(n_157),
.C(n_167),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_153),
.B1(n_154),
.B2(n_156),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_152),
.A2(n_153),
.B1(n_288),
.B2(n_289),
.Y(n_287)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_153),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_153),
.B(n_154),
.Y(n_291)
);

AOI21xp33_ASAP7_75t_L g310 ( 
.A1(n_153),
.A2(n_288),
.B(n_291),
.Y(n_310)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_154),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_158),
.A2(n_159),
.B1(n_165),
.B2(n_166),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_SL g159 ( 
.A(n_160),
.B(n_163),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_160),
.B(n_163),
.C(n_166),
.Y(n_283)
);

CKINVDCx16_ASAP7_75t_R g290 ( 
.A(n_162),
.Y(n_290)
);

CKINVDCx14_ASAP7_75t_R g296 ( 
.A(n_164),
.Y(n_296)
);

CKINVDCx14_ASAP7_75t_R g166 ( 
.A(n_165),
.Y(n_166)
);

AOI321xp33_ASAP7_75t_SL g168 ( 
.A1(n_169),
.A2(n_262),
.A3(n_271),
.B1(n_277),
.B2(n_278),
.C(n_320),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_170),
.A2(n_245),
.B(n_261),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_171),
.A2(n_226),
.B(n_244),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_172),
.A2(n_208),
.B(n_225),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_173),
.A2(n_189),
.B(n_207),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_174),
.B(n_182),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_174),
.B(n_182),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_177),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_175),
.B(n_179),
.C(n_210),
.Y(n_209)
);

CKINVDCx14_ASAP7_75t_R g204 ( 
.A(n_176),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_179),
.Y(n_177)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_178),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_181),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_186),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_183),
.A2(n_184),
.B1(n_186),
.B2(n_187),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_190),
.A2(n_201),
.B(n_206),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_191),
.A2(n_196),
.B(n_200),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_194),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_197),
.B(n_199),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_197),
.B(n_199),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_198),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_205),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_202),
.B(n_205),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_211),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_209),
.B(n_211),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_218),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_212),
.B(n_219),
.C(n_222),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_217),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_213),
.B(n_217),
.Y(n_232)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_222),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_221),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g235 ( 
.A(n_224),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_227),
.B(n_243),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_227),
.B(n_243),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_233),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_232),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_229),
.B(n_232),
.C(n_233),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_231),
.B(n_294),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_SL g233 ( 
.A(n_234),
.B(n_238),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_234),
.B(n_240),
.C(n_241),
.Y(n_258)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_239),
.A2(n_240),
.B1(n_241),
.B2(n_242),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_247),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_246),
.B(n_247),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_248),
.A2(n_249),
.B1(n_256),
.B2(n_257),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_248),
.B(n_258),
.C(n_259),
.Y(n_272)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_253),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_250),
.B(n_254),
.C(n_255),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_255),
.Y(n_253)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_259),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_263),
.B(n_265),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_263),
.B(n_265),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_268),
.C(n_270),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_266),
.A2(n_267),
.B1(n_274),
.B2(n_275),
.Y(n_273)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

BUFx24_ASAP7_75t_SL g317 ( 
.A(n_267),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_268),
.A2(n_269),
.B1(n_270),
.B2(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_270),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_273),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_272),
.B(n_273),
.Y(n_277)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_281),
.B(n_298),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_281),
.B(n_298),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_282),
.A2(n_283),
.B1(n_284),
.B2(n_285),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_282),
.B(n_286),
.C(n_292),
.Y(n_312)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_292),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_291),
.Y(n_286)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_SL g292 ( 
.A1(n_293),
.A2(n_295),
.B(n_297),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_293),
.B(n_295),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_297),
.B(n_306),
.C(n_310),
.Y(n_305)
);

FAx1_ASAP7_75t_SL g313 ( 
.A(n_297),
.B(n_306),
.CI(n_310),
.CON(n_313),
.SN(n_313)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_301),
.B(n_311),
.Y(n_300)
);

AOI21xp33_ASAP7_75t_L g314 ( 
.A1(n_301),
.A2(n_315),
.B(n_316),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_302),
.B(n_305),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_302),
.B(n_305),
.Y(n_316)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_313),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_312),
.B(n_313),
.Y(n_315)
);

BUFx24_ASAP7_75t_SL g318 ( 
.A(n_313),
.Y(n_318)
);


endmodule