module fake_netlist_6_305_n_1005 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_235, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_209, n_98, n_113, n_39, n_63, n_223, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_226, n_228, n_166, n_28, n_184, n_212, n_50, n_158, n_49, n_7, n_210, n_216, n_83, n_206, n_217, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_215, n_178, n_247, n_225, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_227, n_132, n_188, n_102, n_186, n_204, n_245, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_213, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_207, n_2, n_242, n_180, n_19, n_47, n_62, n_29, n_155, n_219, n_75, n_109, n_150, n_233, n_122, n_45, n_205, n_34, n_140, n_218, n_70, n_120, n_234, n_251, n_214, n_37, n_15, n_67, n_33, n_82, n_27, n_236, n_246, n_38, n_110, n_151, n_61, n_112, n_172, n_237, n_81, n_59, n_244, n_181, n_76, n_36, n_182, n_26, n_124, n_238, n_239, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_211, n_64, n_220, n_117, n_118, n_175, n_224, n_48, n_231, n_65, n_230, n_25, n_40, n_93, n_80, n_141, n_240, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_222, n_95, n_179, n_243, n_9, n_248, n_107, n_10, n_71, n_74, n_229, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_249, n_173, n_201, n_250, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_232, n_115, n_12, n_69, n_128, n_241, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_221, n_1005);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_235;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_113;
input n_39;
input n_63;
input n_223;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_226;
input n_228;
input n_166;
input n_28;
input n_184;
input n_212;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_216;
input n_83;
input n_206;
input n_217;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_215;
input n_178;
input n_247;
input n_225;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_227;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_245;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_213;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_242;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_219;
input n_75;
input n_109;
input n_150;
input n_233;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_218;
input n_70;
input n_120;
input n_234;
input n_251;
input n_214;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_236;
input n_246;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_237;
input n_81;
input n_59;
input n_244;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_238;
input n_239;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_211;
input n_64;
input n_220;
input n_117;
input n_118;
input n_175;
input n_224;
input n_48;
input n_231;
input n_65;
input n_230;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_240;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_95;
input n_179;
input n_243;
input n_9;
input n_248;
input n_107;
input n_10;
input n_71;
input n_74;
input n_229;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_249;
input n_173;
input n_201;
input n_250;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_232;
input n_115;
input n_12;
input n_69;
input n_128;
input n_241;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;
input n_221;

output n_1005;

wire n_992;
wire n_591;
wire n_435;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_968;
wire n_909;
wire n_580;
wire n_762;
wire n_881;
wire n_875;
wire n_465;
wire n_680;
wire n_367;
wire n_741;
wire n_760;
wire n_590;
wire n_625;
wire n_661;
wire n_278;
wire n_341;
wire n_362;
wire n_828;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_316;
wire n_419;
wire n_304;
wire n_700;
wire n_694;
wire n_933;
wire n_740;
wire n_578;
wire n_703;
wire n_1003;
wire n_365;
wire n_978;
wire n_384;
wire n_595;
wire n_297;
wire n_627;
wire n_524;
wire n_342;
wire n_820;
wire n_951;
wire n_783;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_310;
wire n_509;
wire n_575;
wire n_368;
wire n_994;
wire n_677;
wire n_969;
wire n_988;
wire n_805;
wire n_396;
wire n_495;
wire n_815;
wire n_350;
wire n_585;
wire n_732;
wire n_974;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_874;
wire n_724;
wire n_673;
wire n_382;
wire n_628;
wire n_883;
wire n_557;
wire n_823;
wire n_349;
wire n_643;
wire n_898;
wire n_617;
wire n_698;
wire n_845;
wire n_255;
wire n_807;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_955;
wire n_865;
wire n_893;
wire n_925;
wire n_485;
wire n_443;
wire n_892;
wire n_768;
wire n_471;
wire n_289;
wire n_935;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_573;
wire n_769;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_963;
wire n_727;
wire n_894;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_832;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_605;
wire n_461;
wire n_873;
wire n_383;
wire n_826;
wire n_669;
wire n_447;
wire n_872;
wire n_300;
wire n_718;
wire n_517;
wire n_747;
wire n_852;
wire n_667;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_621;
wire n_305;
wire n_721;
wire n_996;
wire n_750;
wire n_532;
wire n_742;
wire n_535;
wire n_691;
wire n_544;
wire n_372;
wire n_468;
wire n_901;
wire n_923;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_510;
wire n_837;
wire n_836;
wire n_863;
wire n_601;
wire n_375;
wire n_338;
wire n_522;
wire n_948;
wire n_466;
wire n_704;
wire n_918;
wire n_748;
wire n_506;
wire n_763;
wire n_360;
wire n_945;
wire n_977;
wire n_603;
wire n_991;
wire n_957;
wire n_536;
wire n_895;
wire n_866;
wire n_622;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_658;
wire n_616;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_581;
wire n_428;
wire n_761;
wire n_785;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_987;
wire n_641;
wire n_822;
wire n_693;
wire n_631;
wire n_516;
wire n_720;
wire n_758;
wire n_525;
wire n_842;
wire n_611;
wire n_943;
wire n_491;
wire n_878;
wire n_656;
wire n_772;
wire n_843;
wire n_989;
wire n_797;
wire n_666;
wire n_371;
wire n_795;
wire n_770;
wire n_940;
wire n_567;
wire n_899;
wire n_738;
wire n_405;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_343;
wire n_844;
wire n_448;
wire n_886;
wire n_953;
wire n_1004;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_930;
wire n_888;
wire n_454;
wire n_638;
wire n_910;
wire n_486;
wire n_911;
wire n_381;
wire n_947;
wire n_653;
wire n_887;
wire n_752;
wire n_908;
wire n_944;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_782;
wire n_976;
wire n_490;
wire n_803;
wire n_290;
wire n_809;
wire n_926;
wire n_927;
wire n_839;
wire n_986;
wire n_734;
wire n_708;
wire n_919;
wire n_402;
wire n_352;
wire n_917;
wire n_668;
wire n_478;
wire n_626;
wire n_990;
wire n_574;
wire n_800;
wire n_779;
wire n_929;
wire n_460;
wire n_907;
wire n_854;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_870;
wire n_366;
wire n_904;
wire n_777;
wire n_407;
wire n_913;
wire n_450;
wire n_808;
wire n_867;
wire n_272;
wire n_526;
wire n_921;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_937;
wire n_390;
wire n_473;
wire n_293;
wire n_559;
wire n_334;
wire n_370;
wire n_458;
wire n_650;
wire n_998;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_492;
wire n_972;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_265;
wire n_260;
wire n_313;
wire n_451;
wire n_624;
wire n_824;
wire n_962;
wire n_1000;
wire n_279;
wire n_686;
wire n_796;
wire n_252;
wire n_757;
wire n_594;
wire n_565;
wire n_719;
wire n_356;
wire n_577;
wire n_936;
wire n_552;
wire n_619;
wire n_885;
wire n_455;
wire n_896;
wire n_521;
wire n_363;
wire n_572;
wire n_912;
wire n_395;
wire n_813;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_606;
wire n_393;
wire n_818;
wire n_984;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_884;
wire n_599;
wire n_513;
wire n_855;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_916;
wire n_868;
wire n_570;
wire n_731;
wire n_859;
wire n_406;
wire n_483;
wire n_735;
wire n_934;
wire n_482;
wire n_755;
wire n_931;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_683;
wire n_420;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_958;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_942;
wire n_792;
wire n_880;
wire n_476;
wire n_981;
wire n_714;
wire n_291;
wire n_543;
wire n_889;
wire n_357;
wire n_264;
wire n_263;
wire n_985;
wire n_589;
wire n_860;
wire n_481;
wire n_788;
wire n_819;
wire n_939;
wire n_997;
wire n_821;
wire n_325;
wire n_938;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_831;
wire n_802;
wire n_964;
wire n_982;
wire n_561;
wire n_477;
wire n_549;
wire n_980;
wire n_533;
wire n_954;
wire n_408;
wire n_932;
wire n_806;
wire n_864;
wire n_879;
wire n_959;
wire n_584;
wire n_399;
wire n_979;
wire n_548;
wire n_905;
wire n_282;
wire n_436;
wire n_833;
wire n_523;
wire n_322;
wire n_707;
wire n_993;
wire n_345;
wire n_689;
wire n_409;
wire n_354;
wire n_799;
wire n_505;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_635;
wire n_787;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_966;
wire n_546;
wire n_562;
wire n_386;
wire n_764;
wire n_556;
wire n_692;
wire n_733;
wire n_754;
wire n_941;
wire n_975;
wire n_550;
wire n_487;
wire n_275;
wire n_553;
wire n_652;
wire n_849;
wire n_970;
wire n_560;
wire n_753;
wire n_642;
wire n_995;
wire n_276;
wire n_569;
wire n_441;
wire n_811;
wire n_882;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_269;
wire n_359;
wire n_973;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_790;
wire n_582;
wire n_266;
wire n_296;
wire n_861;
wire n_674;
wire n_857;
wire n_871;
wire n_967;
wire n_775;
wire n_922;
wire n_571;
wire n_268;
wire n_404;
wire n_271;
wire n_651;
wire n_439;
wire n_299;
wire n_518;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_902;
wire n_333;
wire n_588;
wire n_308;
wire n_309;
wire n_914;
wire n_759;
wire n_355;
wire n_426;
wire n_317;
wire n_915;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_285;
wire n_497;
wire n_780;
wire n_773;
wire n_675;
wire n_903;
wire n_257;
wire n_920;
wire n_730;
wire n_655;
wire n_706;
wire n_786;
wire n_670;
wire n_286;
wire n_254;
wire n_834;
wire n_835;
wire n_928;
wire n_850;
wire n_690;
wire n_401;
wire n_324;
wire n_743;
wire n_816;
wire n_766;
wire n_335;
wire n_430;
wire n_1002;
wire n_463;
wire n_545;
wire n_489;
wire n_877;
wire n_604;
wire n_848;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_729;
wire n_876;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_965;
wire n_267;
wire n_438;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_983;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_906;
wire n_688;
wire n_722;
wire n_961;
wire n_862;
wire n_351;
wire n_869;
wire n_437;
wire n_259;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_457;
wire n_391;
wire n_697;
wire n_687;
wire n_364;
wire n_890;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_817;
wire n_950;
wire n_629;
wire n_388;
wire n_858;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_897;
wire n_900;
wire n_846;
wire n_501;
wire n_841;
wire n_956;
wire n_960;
wire n_531;
wire n_827;
wire n_1001;
wire n_663;
wire n_361;
wire n_508;
wire n_856;
wire n_379;
wire n_778;
wire n_332;
wire n_891;
wire n_336;
wire n_410;
wire n_398;
wire n_566;
wire n_554;
wire n_602;
wire n_664;
wire n_949;
wire n_678;
wire n_649;
wire n_283;

BUFx10_ASAP7_75t_L g252 ( 
.A(n_167),
.Y(n_252)
);

CKINVDCx14_ASAP7_75t_R g253 ( 
.A(n_206),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_33),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_187),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_188),
.Y(n_256)
);

OR2x2_ASAP7_75t_L g257 ( 
.A(n_73),
.B(n_10),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_142),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_200),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_239),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_244),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_108),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_109),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_40),
.Y(n_264)
);

BUFx10_ASAP7_75t_L g265 ( 
.A(n_165),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_174),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_28),
.Y(n_267)
);

INVx1_ASAP7_75t_SL g268 ( 
.A(n_193),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_81),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_7),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_145),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_42),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_117),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_100),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_118),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_148),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_154),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_133),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_157),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_13),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_36),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_78),
.Y(n_282)
);

BUFx2_ASAP7_75t_L g283 ( 
.A(n_151),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_197),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_76),
.Y(n_285)
);

BUFx6f_ASAP7_75t_L g286 ( 
.A(n_202),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_162),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_124),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_181),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_236),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_57),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_159),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_177),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_86),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_67),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_144),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_83),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_59),
.Y(n_298)
);

HB1xp67_ASAP7_75t_L g299 ( 
.A(n_210),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_211),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_169),
.Y(n_301)
);

BUFx2_ASAP7_75t_L g302 ( 
.A(n_55),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_96),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_127),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_228),
.Y(n_305)
);

INVx1_ASAP7_75t_SL g306 ( 
.A(n_223),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_64),
.Y(n_307)
);

BUFx3_ASAP7_75t_L g308 ( 
.A(n_47),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_158),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_184),
.Y(n_310)
);

INVx2_ASAP7_75t_SL g311 ( 
.A(n_209),
.Y(n_311)
);

BUFx10_ASAP7_75t_L g312 ( 
.A(n_249),
.Y(n_312)
);

BUFx10_ASAP7_75t_L g313 ( 
.A(n_136),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_237),
.Y(n_314)
);

HB1xp67_ASAP7_75t_L g315 ( 
.A(n_126),
.Y(n_315)
);

BUFx10_ASAP7_75t_L g316 ( 
.A(n_72),
.Y(n_316)
);

NOR2xp67_ASAP7_75t_L g317 ( 
.A(n_134),
.B(n_163),
.Y(n_317)
);

BUFx2_ASAP7_75t_L g318 ( 
.A(n_247),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_14),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_87),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_214),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_125),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_156),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_175),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_178),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_112),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_179),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_213),
.Y(n_328)
);

INVx1_ASAP7_75t_SL g329 ( 
.A(n_131),
.Y(n_329)
);

INVx1_ASAP7_75t_SL g330 ( 
.A(n_150),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_172),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_90),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_106),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_240),
.Y(n_334)
);

INVx1_ASAP7_75t_SL g335 ( 
.A(n_243),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_146),
.Y(n_336)
);

BUFx10_ASAP7_75t_L g337 ( 
.A(n_235),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_121),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_230),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_45),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_170),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_74),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_217),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_189),
.Y(n_344)
);

BUFx10_ASAP7_75t_L g345 ( 
.A(n_245),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_220),
.Y(n_346)
);

BUFx6f_ASAP7_75t_L g347 ( 
.A(n_22),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_171),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_18),
.Y(n_349)
);

NOR2xp67_ASAP7_75t_L g350 ( 
.A(n_82),
.B(n_140),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_98),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_190),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_101),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_104),
.Y(n_354)
);

HB1xp67_ASAP7_75t_L g355 ( 
.A(n_113),
.Y(n_355)
);

HB1xp67_ASAP7_75t_L g356 ( 
.A(n_173),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_122),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_35),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_102),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_238),
.Y(n_360)
);

BUFx6f_ASAP7_75t_L g361 ( 
.A(n_97),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_215),
.Y(n_362)
);

OR2x2_ASAP7_75t_L g363 ( 
.A(n_218),
.B(n_128),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_79),
.Y(n_364)
);

INVx1_ASAP7_75t_SL g365 ( 
.A(n_65),
.Y(n_365)
);

CKINVDCx14_ASAP7_75t_R g366 ( 
.A(n_54),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_48),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_225),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_196),
.Y(n_369)
);

CKINVDCx16_ASAP7_75t_R g370 ( 
.A(n_3),
.Y(n_370)
);

BUFx6f_ASAP7_75t_L g371 ( 
.A(n_242),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_70),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_212),
.Y(n_373)
);

BUFx5_ASAP7_75t_L g374 ( 
.A(n_180),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_186),
.Y(n_375)
);

INVx2_ASAP7_75t_SL g376 ( 
.A(n_95),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_51),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_143),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_119),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_116),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_203),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_89),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_66),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_14),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_205),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_221),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_62),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_246),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_19),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_30),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_75),
.Y(n_391)
);

INVxp33_ASAP7_75t_SL g392 ( 
.A(n_137),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_176),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_24),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_38),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_201),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_71),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_164),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_123),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_229),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_192),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_138),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_198),
.Y(n_403)
);

INVx3_ASAP7_75t_L g404 ( 
.A(n_115),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_20),
.Y(n_405)
);

BUFx2_ASAP7_75t_L g406 ( 
.A(n_3),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_248),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_208),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_135),
.Y(n_409)
);

BUFx2_ASAP7_75t_SL g410 ( 
.A(n_226),
.Y(n_410)
);

NOR2xp67_ASAP7_75t_L g411 ( 
.A(n_88),
.B(n_130),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_149),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_52),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_92),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_94),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_251),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_227),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_141),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_99),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_234),
.Y(n_420)
);

BUFx3_ASAP7_75t_L g421 ( 
.A(n_195),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_182),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_16),
.Y(n_423)
);

BUFx5_ASAP7_75t_L g424 ( 
.A(n_155),
.Y(n_424)
);

BUFx6f_ASAP7_75t_L g425 ( 
.A(n_241),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_168),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_61),
.Y(n_427)
);

NOR2x1_ASAP7_75t_L g428 ( 
.A(n_404),
.B(n_23),
.Y(n_428)
);

BUFx12f_ASAP7_75t_L g429 ( 
.A(n_252),
.Y(n_429)
);

BUFx6f_ASAP7_75t_L g430 ( 
.A(n_270),
.Y(n_430)
);

HB1xp67_ASAP7_75t_L g431 ( 
.A(n_370),
.Y(n_431)
);

AND2x4_ASAP7_75t_L g432 ( 
.A(n_283),
.B(n_0),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_256),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_404),
.B(n_1),
.Y(n_434)
);

CKINVDCx11_ASAP7_75t_R g435 ( 
.A(n_252),
.Y(n_435)
);

AND2x4_ASAP7_75t_L g436 ( 
.A(n_302),
.B(n_2),
.Y(n_436)
);

BUFx2_ASAP7_75t_L g437 ( 
.A(n_406),
.Y(n_437)
);

OA21x2_ASAP7_75t_L g438 ( 
.A1(n_254),
.A2(n_4),
.B(n_5),
.Y(n_438)
);

BUFx6f_ASAP7_75t_L g439 ( 
.A(n_270),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_270),
.Y(n_440)
);

BUFx6f_ASAP7_75t_L g441 ( 
.A(n_347),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_347),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_347),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_318),
.B(n_5),
.Y(n_444)
);

BUFx6f_ASAP7_75t_L g445 ( 
.A(n_286),
.Y(n_445)
);

BUFx6f_ASAP7_75t_L g446 ( 
.A(n_286),
.Y(n_446)
);

HB1xp67_ASAP7_75t_L g447 ( 
.A(n_280),
.Y(n_447)
);

AND2x2_ASAP7_75t_L g448 ( 
.A(n_253),
.B(n_6),
.Y(n_448)
);

BUFx12f_ASAP7_75t_L g449 ( 
.A(n_265),
.Y(n_449)
);

AND2x6_ASAP7_75t_L g450 ( 
.A(n_286),
.B(n_25),
.Y(n_450)
);

INVx3_ASAP7_75t_L g451 ( 
.A(n_312),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_319),
.Y(n_452)
);

BUFx6f_ASAP7_75t_L g453 ( 
.A(n_361),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_389),
.Y(n_454)
);

BUFx12f_ASAP7_75t_L g455 ( 
.A(n_312),
.Y(n_455)
);

OAI22x1_ASAP7_75t_L g456 ( 
.A1(n_423),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_259),
.Y(n_457)
);

BUFx3_ASAP7_75t_L g458 ( 
.A(n_313),
.Y(n_458)
);

INVx2_ASAP7_75t_SL g459 ( 
.A(n_313),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_374),
.Y(n_460)
);

BUFx6f_ASAP7_75t_L g461 ( 
.A(n_361),
.Y(n_461)
);

INVx5_ASAP7_75t_L g462 ( 
.A(n_361),
.Y(n_462)
);

AND2x4_ASAP7_75t_L g463 ( 
.A(n_308),
.B(n_8),
.Y(n_463)
);

BUFx6f_ASAP7_75t_L g464 ( 
.A(n_371),
.Y(n_464)
);

BUFx3_ASAP7_75t_L g465 ( 
.A(n_316),
.Y(n_465)
);

BUFx12f_ASAP7_75t_L g466 ( 
.A(n_316),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_255),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_SL g468 ( 
.A(n_257),
.B(n_9),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_258),
.Y(n_469)
);

AND2x2_ASAP7_75t_L g470 ( 
.A(n_366),
.B(n_10),
.Y(n_470)
);

AOI22xp33_ASAP7_75t_SL g471 ( 
.A1(n_349),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_471)
);

BUFx2_ASAP7_75t_L g472 ( 
.A(n_384),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_260),
.Y(n_473)
);

BUFx6f_ASAP7_75t_L g474 ( 
.A(n_371),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_261),
.Y(n_475)
);

BUFx6f_ASAP7_75t_L g476 ( 
.A(n_371),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_374),
.Y(n_477)
);

AND2x6_ASAP7_75t_L g478 ( 
.A(n_425),
.B(n_26),
.Y(n_478)
);

BUFx2_ASAP7_75t_L g479 ( 
.A(n_405),
.Y(n_479)
);

CKINVDCx16_ASAP7_75t_R g480 ( 
.A(n_277),
.Y(n_480)
);

OR2x2_ASAP7_75t_L g481 ( 
.A(n_299),
.B(n_11),
.Y(n_481)
);

BUFx6f_ASAP7_75t_L g482 ( 
.A(n_425),
.Y(n_482)
);

BUFx6f_ASAP7_75t_L g483 ( 
.A(n_425),
.Y(n_483)
);

INVx3_ASAP7_75t_L g484 ( 
.A(n_337),
.Y(n_484)
);

AND2x4_ASAP7_75t_L g485 ( 
.A(n_421),
.B(n_15),
.Y(n_485)
);

AND2x4_ASAP7_75t_L g486 ( 
.A(n_315),
.B(n_15),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_374),
.Y(n_487)
);

BUFx6f_ASAP7_75t_L g488 ( 
.A(n_337),
.Y(n_488)
);

AND2x4_ASAP7_75t_L g489 ( 
.A(n_355),
.B(n_17),
.Y(n_489)
);

INVx6_ASAP7_75t_L g490 ( 
.A(n_345),
.Y(n_490)
);

BUFx12f_ASAP7_75t_L g491 ( 
.A(n_264),
.Y(n_491)
);

AOI22x1_ASAP7_75t_SL g492 ( 
.A1(n_314),
.A2(n_17),
.B1(n_18),
.B2(n_21),
.Y(n_492)
);

INVxp67_ASAP7_75t_SL g493 ( 
.A(n_356),
.Y(n_493)
);

BUFx6f_ASAP7_75t_L g494 ( 
.A(n_303),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_374),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_262),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_311),
.B(n_21),
.Y(n_497)
);

INVx3_ASAP7_75t_L g498 ( 
.A(n_263),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_267),
.Y(n_499)
);

INVx5_ASAP7_75t_L g500 ( 
.A(n_376),
.Y(n_500)
);

INVx5_ASAP7_75t_L g501 ( 
.A(n_344),
.Y(n_501)
);

AND2x2_ASAP7_75t_L g502 ( 
.A(n_358),
.B(n_22),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_374),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_424),
.Y(n_504)
);

OA21x2_ASAP7_75t_L g505 ( 
.A1(n_271),
.A2(n_27),
.B(n_29),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_281),
.Y(n_506)
);

INVxp67_ASAP7_75t_L g507 ( 
.A(n_284),
.Y(n_507)
);

OAI21x1_ASAP7_75t_L g508 ( 
.A1(n_416),
.A2(n_31),
.B(n_32),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_419),
.B(n_34),
.Y(n_509)
);

AND2x2_ASAP7_75t_SL g510 ( 
.A(n_363),
.B(n_37),
.Y(n_510)
);

BUFx12f_ASAP7_75t_L g511 ( 
.A(n_266),
.Y(n_511)
);

BUFx6f_ASAP7_75t_L g512 ( 
.A(n_285),
.Y(n_512)
);

AND2x4_ASAP7_75t_L g513 ( 
.A(n_288),
.B(n_39),
.Y(n_513)
);

AND2x4_ASAP7_75t_L g514 ( 
.A(n_290),
.B(n_41),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_424),
.Y(n_515)
);

INVx6_ASAP7_75t_L g516 ( 
.A(n_424),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_392),
.B(n_43),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_424),
.Y(n_518)
);

BUFx8_ASAP7_75t_L g519 ( 
.A(n_424),
.Y(n_519)
);

AOI22xp5_ASAP7_75t_L g520 ( 
.A1(n_268),
.A2(n_44),
.B1(n_46),
.B2(n_49),
.Y(n_520)
);

BUFx6f_ASAP7_75t_L g521 ( 
.A(n_292),
.Y(n_521)
);

AND2x2_ASAP7_75t_L g522 ( 
.A(n_306),
.B(n_50),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_445),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_440),
.Y(n_524)
);

BUFx10_ASAP7_75t_L g525 ( 
.A(n_490),
.Y(n_525)
);

INVx3_ASAP7_75t_L g526 ( 
.A(n_430),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_433),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_442),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_457),
.Y(n_529)
);

BUFx3_ASAP7_75t_L g530 ( 
.A(n_491),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_445),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_511),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_435),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_R g534 ( 
.A(n_480),
.B(n_269),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_429),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_449),
.Y(n_536)
);

NAND2xp33_ASAP7_75t_R g537 ( 
.A(n_472),
.B(n_272),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_446),
.Y(n_538)
);

CKINVDCx20_ASAP7_75t_R g539 ( 
.A(n_431),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_430),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_R g541 ( 
.A(n_510),
.B(n_273),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_455),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_446),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_466),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_488),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_439),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_453),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_488),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_472),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_439),
.Y(n_550)
);

HB1xp67_ASAP7_75t_L g551 ( 
.A(n_458),
.Y(n_551)
);

BUFx3_ASAP7_75t_L g552 ( 
.A(n_519),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_479),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_479),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_453),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_461),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_465),
.Y(n_557)
);

INVxp67_ASAP7_75t_L g558 ( 
.A(n_447),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_461),
.Y(n_559)
);

BUFx10_ASAP7_75t_L g560 ( 
.A(n_490),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_451),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_484),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_459),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_441),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_437),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_441),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_493),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_464),
.Y(n_568)
);

BUFx6f_ASAP7_75t_L g569 ( 
.A(n_464),
.Y(n_569)
);

BUFx3_ASAP7_75t_L g570 ( 
.A(n_494),
.Y(n_570)
);

BUFx2_ASAP7_75t_L g571 ( 
.A(n_512),
.Y(n_571)
);

BUFx6f_ASAP7_75t_L g572 ( 
.A(n_474),
.Y(n_572)
);

INVx3_ASAP7_75t_L g573 ( 
.A(n_474),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_500),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_476),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_R g576 ( 
.A(n_468),
.B(n_274),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_476),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_482),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_500),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_494),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_512),
.Y(n_581)
);

AND2x2_ASAP7_75t_L g582 ( 
.A(n_448),
.B(n_329),
.Y(n_582)
);

HB1xp67_ASAP7_75t_L g583 ( 
.A(n_521),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_482),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_521),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_467),
.B(n_469),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_483),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_432),
.Y(n_588)
);

CKINVDCx20_ASAP7_75t_R g589 ( 
.A(n_517),
.Y(n_589)
);

NOR2xp67_ASAP7_75t_L g590 ( 
.A(n_462),
.B(n_293),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_436),
.Y(n_591)
);

BUFx6f_ASAP7_75t_L g592 ( 
.A(n_462),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_507),
.Y(n_593)
);

BUFx3_ASAP7_75t_L g594 ( 
.A(n_473),
.Y(n_594)
);

NOR2xp33_ASAP7_75t_L g595 ( 
.A(n_444),
.B(n_522),
.Y(n_595)
);

BUFx6f_ASAP7_75t_L g596 ( 
.A(n_569),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_583),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_587),
.Y(n_598)
);

INVxp33_ASAP7_75t_L g599 ( 
.A(n_551),
.Y(n_599)
);

NOR2xp67_ASAP7_75t_SL g600 ( 
.A(n_552),
.B(n_438),
.Y(n_600)
);

AO221x1_ASAP7_75t_L g601 ( 
.A1(n_558),
.A2(n_456),
.B1(n_418),
.B2(n_417),
.C(n_295),
.Y(n_601)
);

NOR2xp33_ASAP7_75t_L g602 ( 
.A(n_595),
.B(n_448),
.Y(n_602)
);

AOI22xp33_ASAP7_75t_L g603 ( 
.A1(n_582),
.A2(n_470),
.B1(n_502),
.B2(n_489),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_593),
.B(n_522),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_567),
.B(n_470),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_581),
.B(n_462),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_585),
.B(n_513),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_580),
.B(n_514),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_594),
.Y(n_609)
);

BUFx6f_ASAP7_75t_L g610 ( 
.A(n_569),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_524),
.B(n_501),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g612 ( 
.A(n_558),
.B(n_481),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_528),
.B(n_501),
.Y(n_613)
);

BUFx6f_ASAP7_75t_SL g614 ( 
.A(n_530),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_L g615 ( 
.A(n_561),
.B(n_486),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_592),
.B(n_501),
.Y(n_616)
);

INVxp33_ASAP7_75t_SL g617 ( 
.A(n_545),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_592),
.B(n_502),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_571),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_592),
.B(n_475),
.Y(n_620)
);

NAND2xp33_ASAP7_75t_L g621 ( 
.A(n_541),
.B(n_450),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_SL g622 ( 
.A(n_548),
.B(n_463),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_SL g623 ( 
.A(n_576),
.B(n_485),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_SL g624 ( 
.A(n_562),
.B(n_434),
.Y(n_624)
);

INVx2_ASAP7_75t_SL g625 ( 
.A(n_525),
.Y(n_625)
);

NOR2xp67_ASAP7_75t_L g626 ( 
.A(n_527),
.B(n_498),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_570),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_590),
.B(n_496),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_588),
.B(n_499),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_591),
.B(n_506),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_573),
.Y(n_631)
);

INVxp67_ASAP7_75t_SL g632 ( 
.A(n_573),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_523),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_531),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_572),
.Y(n_635)
);

NOR3xp33_ASAP7_75t_L g636 ( 
.A(n_565),
.B(n_471),
.C(n_497),
.Y(n_636)
);

INVx2_ASAP7_75t_SL g637 ( 
.A(n_525),
.Y(n_637)
);

INVxp67_ASAP7_75t_SL g638 ( 
.A(n_572),
.Y(n_638)
);

INVx2_ASAP7_75t_SL g639 ( 
.A(n_560),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_L g640 ( 
.A(n_563),
.B(n_443),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_538),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_586),
.B(n_516),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_SL g643 ( 
.A(n_529),
.B(n_275),
.Y(n_643)
);

NOR2x1p5_ASAP7_75t_L g644 ( 
.A(n_557),
.B(n_452),
.Y(n_644)
);

INVx2_ASAP7_75t_SL g645 ( 
.A(n_560),
.Y(n_645)
);

NOR2xp33_ASAP7_75t_L g646 ( 
.A(n_589),
.B(n_509),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_SL g647 ( 
.A(n_534),
.B(n_276),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_572),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_540),
.Y(n_649)
);

NOR2xp33_ASAP7_75t_L g650 ( 
.A(n_549),
.B(n_330),
.Y(n_650)
);

INVxp67_ASAP7_75t_L g651 ( 
.A(n_537),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_546),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_586),
.B(n_516),
.Y(n_653)
);

INVx2_ASAP7_75t_SL g654 ( 
.A(n_553),
.Y(n_654)
);

NOR3xp33_ASAP7_75t_L g655 ( 
.A(n_554),
.B(n_365),
.C(n_335),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_543),
.B(n_450),
.Y(n_656)
);

NOR2xp33_ASAP7_75t_L g657 ( 
.A(n_574),
.B(n_454),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_547),
.B(n_555),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_SL g659 ( 
.A(n_579),
.B(n_278),
.Y(n_659)
);

NOR2xp67_ASAP7_75t_L g660 ( 
.A(n_532),
.B(n_520),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_556),
.Y(n_661)
);

HB1xp67_ASAP7_75t_L g662 ( 
.A(n_539),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_559),
.B(n_518),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_568),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_575),
.B(n_460),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_577),
.B(n_515),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_SL g667 ( 
.A(n_535),
.B(n_279),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_578),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_SL g669 ( 
.A(n_536),
.B(n_282),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_550),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_584),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_564),
.Y(n_672)
);

AND2x2_ASAP7_75t_L g673 ( 
.A(n_526),
.B(n_477),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_566),
.Y(n_674)
);

INVxp33_ASAP7_75t_SL g675 ( 
.A(n_533),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_526),
.B(n_487),
.Y(n_676)
);

BUFx2_ASAP7_75t_L g677 ( 
.A(n_662),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_676),
.Y(n_678)
);

INVx5_ASAP7_75t_L g679 ( 
.A(n_596),
.Y(n_679)
);

AOI22xp33_ASAP7_75t_L g680 ( 
.A1(n_602),
.A2(n_438),
.B1(n_478),
.B2(n_450),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_676),
.Y(n_681)
);

BUFx6f_ASAP7_75t_L g682 ( 
.A(n_596),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_673),
.Y(n_683)
);

AOI22xp5_ASAP7_75t_L g684 ( 
.A1(n_646),
.A2(n_289),
.B1(n_291),
.B2(n_287),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_617),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_675),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_SL g687 ( 
.A(n_604),
.B(n_542),
.Y(n_687)
);

OAI22xp33_ASAP7_75t_L g688 ( 
.A1(n_651),
.A2(n_296),
.B1(n_298),
.B2(n_294),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_663),
.Y(n_689)
);

INVx4_ASAP7_75t_L g690 ( 
.A(n_596),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_598),
.Y(n_691)
);

AOI22xp33_ASAP7_75t_L g692 ( 
.A1(n_636),
.A2(n_478),
.B1(n_505),
.B2(n_428),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_663),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_665),
.Y(n_694)
);

AND2x6_ASAP7_75t_SL g695 ( 
.A(n_650),
.B(n_612),
.Y(n_695)
);

AND2x4_ASAP7_75t_L g696 ( 
.A(n_609),
.B(n_632),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_665),
.Y(n_697)
);

AOI22xp33_ASAP7_75t_L g698 ( 
.A1(n_603),
.A2(n_478),
.B1(n_505),
.B2(n_410),
.Y(n_698)
);

AOI22xp5_ASAP7_75t_L g699 ( 
.A1(n_621),
.A2(n_297),
.B1(n_304),
.B2(n_320),
.Y(n_699)
);

AOI21xp5_ASAP7_75t_L g700 ( 
.A1(n_618),
.A2(n_503),
.B(n_495),
.Y(n_700)
);

NOR2xp33_ASAP7_75t_L g701 ( 
.A(n_605),
.B(n_544),
.Y(n_701)
);

BUFx4f_ASAP7_75t_L g702 ( 
.A(n_625),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_642),
.B(n_301),
.Y(n_703)
);

INVx2_ASAP7_75t_SL g704 ( 
.A(n_619),
.Y(n_704)
);

INVx1_ASAP7_75t_SL g705 ( 
.A(n_654),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_SL g706 ( 
.A(n_626),
.B(n_300),
.Y(n_706)
);

HB1xp67_ASAP7_75t_L g707 ( 
.A(n_597),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_SL g708 ( 
.A(n_623),
.B(n_322),
.Y(n_708)
);

AOI211xp5_ASAP7_75t_L g709 ( 
.A1(n_655),
.A2(n_305),
.B(n_307),
.C(n_309),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_649),
.Y(n_710)
);

AOI22xp5_ASAP7_75t_L g711 ( 
.A1(n_615),
.A2(n_377),
.B1(n_323),
.B2(n_325),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_653),
.B(n_600),
.Y(n_712)
);

INVx4_ASAP7_75t_L g713 ( 
.A(n_610),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_652),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_666),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_666),
.Y(n_716)
);

HB1xp67_ASAP7_75t_L g717 ( 
.A(n_629),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_631),
.Y(n_718)
);

NAND2x1p5_ASAP7_75t_L g719 ( 
.A(n_644),
.B(n_508),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_607),
.B(n_608),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_630),
.B(n_310),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_658),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_670),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_624),
.B(n_321),
.Y(n_724)
);

AND2x4_ASAP7_75t_L g725 ( 
.A(n_627),
.B(n_324),
.Y(n_725)
);

NOR2xp67_ASAP7_75t_L g726 ( 
.A(n_637),
.B(n_326),
.Y(n_726)
);

HB1xp67_ASAP7_75t_L g727 ( 
.A(n_599),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_640),
.B(n_327),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_SL g729 ( 
.A(n_660),
.B(n_328),
.Y(n_729)
);

INVx2_ASAP7_75t_SL g730 ( 
.A(n_635),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_SL g731 ( 
.A(n_639),
.B(n_331),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_672),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_674),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_633),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_634),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_638),
.B(n_334),
.Y(n_736)
);

INVxp67_ASAP7_75t_SL g737 ( 
.A(n_610),
.Y(n_737)
);

NOR2x2_ASAP7_75t_L g738 ( 
.A(n_648),
.B(n_492),
.Y(n_738)
);

AND2x4_ASAP7_75t_L g739 ( 
.A(n_641),
.B(n_661),
.Y(n_739)
);

BUFx4f_ASAP7_75t_L g740 ( 
.A(n_645),
.Y(n_740)
);

OR2x6_ASAP7_75t_L g741 ( 
.A(n_622),
.B(n_317),
.Y(n_741)
);

INVx2_ASAP7_75t_SL g742 ( 
.A(n_664),
.Y(n_742)
);

AOI22xp5_ASAP7_75t_L g743 ( 
.A1(n_601),
.A2(n_382),
.B1(n_333),
.B2(n_426),
.Y(n_743)
);

INVx3_ASAP7_75t_L g744 ( 
.A(n_668),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_671),
.Y(n_745)
);

INVx5_ASAP7_75t_L g746 ( 
.A(n_656),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_620),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_606),
.B(n_346),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_611),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_689),
.B(n_647),
.Y(n_750)
);

O2A1O1Ixp5_ASAP7_75t_L g751 ( 
.A1(n_712),
.A2(n_643),
.B(n_659),
.C(n_657),
.Y(n_751)
);

INVx1_ASAP7_75t_SL g752 ( 
.A(n_727),
.Y(n_752)
);

OAI22xp5_ASAP7_75t_L g753 ( 
.A1(n_698),
.A2(n_350),
.B1(n_411),
.B2(n_360),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_683),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_SL g755 ( 
.A(n_720),
.B(n_628),
.Y(n_755)
);

OAI22xp5_ASAP7_75t_L g756 ( 
.A1(n_692),
.A2(n_359),
.B1(n_368),
.B2(n_369),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_691),
.Y(n_757)
);

HB1xp67_ASAP7_75t_L g758 ( 
.A(n_707),
.Y(n_758)
);

BUFx6f_ASAP7_75t_L g759 ( 
.A(n_682),
.Y(n_759)
);

AOI22xp33_ASAP7_75t_L g760 ( 
.A1(n_693),
.A2(n_372),
.B1(n_379),
.B2(n_383),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_710),
.Y(n_761)
);

BUFx6f_ASAP7_75t_L g762 ( 
.A(n_682),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_734),
.Y(n_763)
);

AND2x4_ASAP7_75t_L g764 ( 
.A(n_704),
.B(n_667),
.Y(n_764)
);

AOI21xp5_ASAP7_75t_L g765 ( 
.A1(n_680),
.A2(n_613),
.B(n_616),
.Y(n_765)
);

O2A1O1Ixp33_ASAP7_75t_L g766 ( 
.A1(n_688),
.A2(n_398),
.B(n_408),
.C(n_427),
.Y(n_766)
);

A2O1A1Ixp33_ASAP7_75t_L g767 ( 
.A1(n_694),
.A2(n_397),
.B(n_412),
.C(n_391),
.Y(n_767)
);

OAI22xp5_ASAP7_75t_L g768 ( 
.A1(n_678),
.A2(n_394),
.B1(n_403),
.B2(n_409),
.Y(n_768)
);

BUFx3_ASAP7_75t_L g769 ( 
.A(n_677),
.Y(n_769)
);

NOR2xp67_ASAP7_75t_L g770 ( 
.A(n_686),
.B(n_669),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_SL g771 ( 
.A(n_717),
.B(n_332),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_SL g772 ( 
.A(n_705),
.B(n_336),
.Y(n_772)
);

AOI22xp5_ASAP7_75t_L g773 ( 
.A1(n_697),
.A2(n_413),
.B1(n_338),
.B2(n_422),
.Y(n_773)
);

OAI22xp5_ASAP7_75t_L g774 ( 
.A1(n_681),
.A2(n_715),
.B1(n_716),
.B2(n_722),
.Y(n_774)
);

NOR2x1_ASAP7_75t_R g775 ( 
.A(n_685),
.B(n_339),
.Y(n_775)
);

AOI22xp5_ASAP7_75t_L g776 ( 
.A1(n_749),
.A2(n_385),
.B1(n_341),
.B2(n_420),
.Y(n_776)
);

CKINVDCx11_ASAP7_75t_R g777 ( 
.A(n_695),
.Y(n_777)
);

OAI22xp5_ASAP7_75t_L g778 ( 
.A1(n_747),
.A2(n_381),
.B1(n_342),
.B2(n_415),
.Y(n_778)
);

AOI21xp5_ASAP7_75t_L g779 ( 
.A1(n_703),
.A2(n_380),
.B(n_414),
.Y(n_779)
);

BUFx6f_ASAP7_75t_L g780 ( 
.A(n_682),
.Y(n_780)
);

OAI22xp5_ASAP7_75t_L g781 ( 
.A1(n_724),
.A2(n_386),
.B1(n_343),
.B2(n_407),
.Y(n_781)
);

O2A1O1Ixp5_ASAP7_75t_L g782 ( 
.A1(n_748),
.A2(n_504),
.B(n_402),
.C(n_401),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_721),
.B(n_340),
.Y(n_783)
);

O2A1O1Ixp33_ASAP7_75t_L g784 ( 
.A1(n_728),
.A2(n_400),
.B(n_399),
.C(n_396),
.Y(n_784)
);

INVx4_ASAP7_75t_SL g785 ( 
.A(n_741),
.Y(n_785)
);

AOI21xp5_ASAP7_75t_L g786 ( 
.A1(n_737),
.A2(n_395),
.B(n_393),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_735),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_732),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_714),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_SL g790 ( 
.A(n_696),
.B(n_744),
.Y(n_790)
);

O2A1O1Ixp5_ASAP7_75t_L g791 ( 
.A1(n_708),
.A2(n_390),
.B(n_388),
.C(n_387),
.Y(n_791)
);

O2A1O1Ixp33_ASAP7_75t_L g792 ( 
.A1(n_729),
.A2(n_378),
.B(n_375),
.C(n_373),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_SL g793 ( 
.A(n_701),
.B(n_348),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_746),
.B(n_351),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_SL g795 ( 
.A(n_742),
.B(n_352),
.Y(n_795)
);

AOI21xp5_ASAP7_75t_L g796 ( 
.A1(n_736),
.A2(n_367),
.B(n_364),
.Y(n_796)
);

HB1xp67_ASAP7_75t_L g797 ( 
.A(n_725),
.Y(n_797)
);

AND2x2_ASAP7_75t_L g798 ( 
.A(n_702),
.B(n_353),
.Y(n_798)
);

NOR2x1_ASAP7_75t_L g799 ( 
.A(n_687),
.B(n_614),
.Y(n_799)
);

BUFx6f_ASAP7_75t_L g800 ( 
.A(n_762),
.Y(n_800)
);

BUFx3_ASAP7_75t_L g801 ( 
.A(n_769),
.Y(n_801)
);

AO21x2_ASAP7_75t_L g802 ( 
.A1(n_765),
.A2(n_700),
.B(n_743),
.Y(n_802)
);

BUFx12f_ASAP7_75t_L g803 ( 
.A(n_777),
.Y(n_803)
);

BUFx10_ASAP7_75t_L g804 ( 
.A(n_764),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_763),
.Y(n_805)
);

INVx8_ASAP7_75t_L g806 ( 
.A(n_762),
.Y(n_806)
);

AO21x1_ASAP7_75t_L g807 ( 
.A1(n_753),
.A2(n_719),
.B(n_709),
.Y(n_807)
);

AO21x2_ASAP7_75t_L g808 ( 
.A1(n_756),
.A2(n_706),
.B(n_733),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_774),
.B(n_755),
.Y(n_809)
);

BUFx12f_ASAP7_75t_L g810 ( 
.A(n_759),
.Y(n_810)
);

BUFx3_ASAP7_75t_L g811 ( 
.A(n_759),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_757),
.Y(n_812)
);

BUFx3_ASAP7_75t_L g813 ( 
.A(n_780),
.Y(n_813)
);

OAI21x1_ASAP7_75t_L g814 ( 
.A1(n_782),
.A2(n_718),
.B(n_745),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_761),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_750),
.B(n_746),
.Y(n_816)
);

INVx4_ASAP7_75t_L g817 ( 
.A(n_762),
.Y(n_817)
);

OAI21x1_ASAP7_75t_L g818 ( 
.A1(n_791),
.A2(n_723),
.B(n_699),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_787),
.Y(n_819)
);

BUFx3_ASAP7_75t_L g820 ( 
.A(n_780),
.Y(n_820)
);

BUFx3_ASAP7_75t_L g821 ( 
.A(n_752),
.Y(n_821)
);

OA21x2_ASAP7_75t_L g822 ( 
.A1(n_767),
.A2(n_725),
.B(n_739),
.Y(n_822)
);

AOI21x1_ASAP7_75t_L g823 ( 
.A1(n_794),
.A2(n_739),
.B(n_730),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_789),
.Y(n_824)
);

HB1xp67_ASAP7_75t_L g825 ( 
.A(n_758),
.Y(n_825)
);

INVx3_ASAP7_75t_L g826 ( 
.A(n_754),
.Y(n_826)
);

OAI21x1_ASAP7_75t_L g827 ( 
.A1(n_751),
.A2(n_731),
.B(n_711),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_788),
.Y(n_828)
);

OAI21xp5_ASAP7_75t_L g829 ( 
.A1(n_773),
.A2(n_684),
.B(n_746),
.Y(n_829)
);

BUFx3_ASAP7_75t_L g830 ( 
.A(n_797),
.Y(n_830)
);

BUFx6f_ASAP7_75t_L g831 ( 
.A(n_790),
.Y(n_831)
);

BUFx2_ASAP7_75t_L g832 ( 
.A(n_821),
.Y(n_832)
);

AO21x1_ASAP7_75t_L g833 ( 
.A1(n_809),
.A2(n_784),
.B(n_793),
.Y(n_833)
);

BUFx6f_ASAP7_75t_L g834 ( 
.A(n_800),
.Y(n_834)
);

INVx8_ASAP7_75t_L g835 ( 
.A(n_806),
.Y(n_835)
);

BUFx12f_ASAP7_75t_L g836 ( 
.A(n_810),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_805),
.B(n_783),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_819),
.Y(n_838)
);

AOI21x1_ASAP7_75t_L g839 ( 
.A1(n_823),
.A2(n_768),
.B(n_795),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_828),
.Y(n_840)
);

AND2x2_ASAP7_75t_L g841 ( 
.A(n_821),
.B(n_798),
.Y(n_841)
);

INVx3_ASAP7_75t_L g842 ( 
.A(n_817),
.Y(n_842)
);

AOI22xp33_ASAP7_75t_SL g843 ( 
.A1(n_829),
.A2(n_741),
.B1(n_614),
.B2(n_740),
.Y(n_843)
);

OAI22xp33_ASAP7_75t_L g844 ( 
.A1(n_831),
.A2(n_770),
.B1(n_799),
.B2(n_771),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_812),
.Y(n_845)
);

INVx2_ASAP7_75t_L g846 ( 
.A(n_812),
.Y(n_846)
);

INVx1_ASAP7_75t_SL g847 ( 
.A(n_801),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_815),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_826),
.B(n_815),
.Y(n_849)
);

CKINVDCx11_ASAP7_75t_R g850 ( 
.A(n_803),
.Y(n_850)
);

AOI22xp33_ASAP7_75t_L g851 ( 
.A1(n_807),
.A2(n_760),
.B1(n_781),
.B2(n_772),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_824),
.Y(n_852)
);

AND2x4_ASAP7_75t_L g853 ( 
.A(n_830),
.B(n_785),
.Y(n_853)
);

AND2x2_ASAP7_75t_L g854 ( 
.A(n_830),
.B(n_726),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_825),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_831),
.Y(n_856)
);

AOI22xp33_ASAP7_75t_L g857 ( 
.A1(n_807),
.A2(n_776),
.B1(n_778),
.B2(n_362),
.Y(n_857)
);

INVx1_ASAP7_75t_SL g858 ( 
.A(n_832),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_838),
.Y(n_859)
);

OR2x6_ASAP7_75t_L g860 ( 
.A(n_835),
.B(n_801),
.Y(n_860)
);

AND2x4_ASAP7_75t_L g861 ( 
.A(n_853),
.B(n_811),
.Y(n_861)
);

OR2x2_ASAP7_75t_L g862 ( 
.A(n_855),
.B(n_816),
.Y(n_862)
);

INVx3_ASAP7_75t_L g863 ( 
.A(n_835),
.Y(n_863)
);

CKINVDCx16_ASAP7_75t_R g864 ( 
.A(n_836),
.Y(n_864)
);

INVxp33_ASAP7_75t_SL g865 ( 
.A(n_841),
.Y(n_865)
);

NOR3xp33_ASAP7_75t_SL g866 ( 
.A(n_844),
.B(n_766),
.C(n_357),
.Y(n_866)
);

OR2x2_ASAP7_75t_SL g867 ( 
.A(n_837),
.B(n_831),
.Y(n_867)
);

NAND2xp33_ASAP7_75t_R g868 ( 
.A(n_853),
.B(n_822),
.Y(n_868)
);

OR2x6_ASAP7_75t_L g869 ( 
.A(n_854),
.B(n_806),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_849),
.Y(n_870)
);

NAND2xp33_ASAP7_75t_R g871 ( 
.A(n_856),
.B(n_822),
.Y(n_871)
);

NAND3xp33_ASAP7_75t_SL g872 ( 
.A(n_843),
.B(n_792),
.C(n_779),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_849),
.Y(n_873)
);

AND2x2_ASAP7_75t_L g874 ( 
.A(n_840),
.B(n_804),
.Y(n_874)
);

AND2x4_ASAP7_75t_L g875 ( 
.A(n_847),
.B(n_811),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_846),
.Y(n_876)
);

BUFx2_ASAP7_75t_L g877 ( 
.A(n_834),
.Y(n_877)
);

NOR3xp33_ASAP7_75t_SL g878 ( 
.A(n_844),
.B(n_354),
.C(n_775),
.Y(n_878)
);

OR2x2_ASAP7_75t_L g879 ( 
.A(n_845),
.B(n_813),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_848),
.Y(n_880)
);

OR2x2_ASAP7_75t_L g881 ( 
.A(n_852),
.B(n_813),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_843),
.B(n_804),
.Y(n_882)
);

NAND2xp33_ASAP7_75t_R g883 ( 
.A(n_842),
.B(n_822),
.Y(n_883)
);

AOI21xp5_ASAP7_75t_L g884 ( 
.A1(n_833),
.A2(n_802),
.B(n_827),
.Y(n_884)
);

BUFx3_ASAP7_75t_L g885 ( 
.A(n_875),
.Y(n_885)
);

AOI22xp33_ASAP7_75t_L g886 ( 
.A1(n_865),
.A2(n_857),
.B1(n_851),
.B2(n_808),
.Y(n_886)
);

INVx2_ASAP7_75t_SL g887 ( 
.A(n_860),
.Y(n_887)
);

AND2x2_ASAP7_75t_L g888 ( 
.A(n_874),
.B(n_834),
.Y(n_888)
);

CKINVDCx5p33_ASAP7_75t_R g889 ( 
.A(n_864),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_880),
.Y(n_890)
);

AND2x2_ASAP7_75t_L g891 ( 
.A(n_859),
.B(n_827),
.Y(n_891)
);

AOI22xp33_ASAP7_75t_L g892 ( 
.A1(n_882),
.A2(n_803),
.B1(n_850),
.B2(n_802),
.Y(n_892)
);

AND2x2_ASAP7_75t_L g893 ( 
.A(n_862),
.B(n_820),
.Y(n_893)
);

AND2x2_ASAP7_75t_L g894 ( 
.A(n_879),
.B(n_814),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_858),
.B(n_814),
.Y(n_895)
);

AND2x2_ASAP7_75t_L g896 ( 
.A(n_870),
.B(n_839),
.Y(n_896)
);

AND2x2_ASAP7_75t_L g897 ( 
.A(n_870),
.B(n_818),
.Y(n_897)
);

OR2x2_ASAP7_75t_L g898 ( 
.A(n_867),
.B(n_818),
.Y(n_898)
);

NAND2x1p5_ASAP7_75t_L g899 ( 
.A(n_863),
.B(n_817),
.Y(n_899)
);

AO21x2_ASAP7_75t_L g900 ( 
.A1(n_884),
.A2(n_786),
.B(n_796),
.Y(n_900)
);

AND2x2_ASAP7_75t_L g901 ( 
.A(n_881),
.B(n_800),
.Y(n_901)
);

INVx2_ASAP7_75t_SL g902 ( 
.A(n_860),
.Y(n_902)
);

AND2x4_ASAP7_75t_L g903 ( 
.A(n_873),
.B(n_817),
.Y(n_903)
);

BUFx3_ASAP7_75t_L g904 ( 
.A(n_875),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_876),
.Y(n_905)
);

AOI22xp5_ASAP7_75t_L g906 ( 
.A1(n_878),
.A2(n_850),
.B1(n_713),
.B2(n_806),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_877),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_869),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_871),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_883),
.Y(n_910)
);

HB1xp67_ASAP7_75t_L g911 ( 
.A(n_868),
.Y(n_911)
);

INVx2_ASAP7_75t_L g912 ( 
.A(n_861),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_890),
.Y(n_913)
);

AND2x2_ASAP7_75t_L g914 ( 
.A(n_888),
.B(n_866),
.Y(n_914)
);

OAI22xp5_ASAP7_75t_L g915 ( 
.A1(n_886),
.A2(n_690),
.B1(n_872),
.B2(n_679),
.Y(n_915)
);

INVxp67_ASAP7_75t_L g916 ( 
.A(n_911),
.Y(n_916)
);

INVx3_ASAP7_75t_L g917 ( 
.A(n_898),
.Y(n_917)
);

AND2x2_ASAP7_75t_L g918 ( 
.A(n_907),
.B(n_53),
.Y(n_918)
);

AND2x2_ASAP7_75t_L g919 ( 
.A(n_907),
.B(n_56),
.Y(n_919)
);

AND2x2_ASAP7_75t_L g920 ( 
.A(n_885),
.B(n_58),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_895),
.Y(n_921)
);

OR2x2_ASAP7_75t_L g922 ( 
.A(n_911),
.B(n_60),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_891),
.Y(n_923)
);

AND2x2_ASAP7_75t_L g924 ( 
.A(n_885),
.B(n_63),
.Y(n_924)
);

BUFx2_ASAP7_75t_L g925 ( 
.A(n_904),
.Y(n_925)
);

NOR2xp33_ASAP7_75t_L g926 ( 
.A(n_909),
.B(n_68),
.Y(n_926)
);

NOR3xp33_ASAP7_75t_L g927 ( 
.A(n_908),
.B(n_738),
.C(n_77),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_905),
.Y(n_928)
);

AND2x4_ASAP7_75t_SL g929 ( 
.A(n_903),
.B(n_69),
.Y(n_929)
);

AND2x2_ASAP7_75t_L g930 ( 
.A(n_904),
.B(n_80),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_905),
.Y(n_931)
);

OR2x2_ASAP7_75t_L g932 ( 
.A(n_909),
.B(n_84),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_894),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_897),
.Y(n_934)
);

INVxp67_ASAP7_75t_SL g935 ( 
.A(n_897),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_913),
.Y(n_936)
);

OR2x2_ASAP7_75t_L g937 ( 
.A(n_916),
.B(n_910),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_928),
.Y(n_938)
);

NOR2xp33_ASAP7_75t_L g939 ( 
.A(n_914),
.B(n_887),
.Y(n_939)
);

NAND2x1p5_ASAP7_75t_L g940 ( 
.A(n_925),
.B(n_896),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_SL g941 ( 
.A(n_932),
.B(n_892),
.Y(n_941)
);

AND2x2_ASAP7_75t_L g942 ( 
.A(n_933),
.B(n_887),
.Y(n_942)
);

INVx2_ASAP7_75t_L g943 ( 
.A(n_934),
.Y(n_943)
);

INVx3_ASAP7_75t_L g944 ( 
.A(n_917),
.Y(n_944)
);

AOI22xp33_ASAP7_75t_L g945 ( 
.A1(n_927),
.A2(n_893),
.B1(n_912),
.B2(n_889),
.Y(n_945)
);

INVxp67_ASAP7_75t_SL g946 ( 
.A(n_921),
.Y(n_946)
);

AND2x2_ASAP7_75t_L g947 ( 
.A(n_917),
.B(n_923),
.Y(n_947)
);

AND2x2_ASAP7_75t_L g948 ( 
.A(n_917),
.B(n_902),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_931),
.Y(n_949)
);

OR2x2_ASAP7_75t_L g950 ( 
.A(n_934),
.B(n_912),
.Y(n_950)
);

AND2x2_ASAP7_75t_L g951 ( 
.A(n_935),
.B(n_901),
.Y(n_951)
);

INVx1_ASAP7_75t_SL g952 ( 
.A(n_937),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_936),
.Y(n_953)
);

OAI322xp33_ASAP7_75t_L g954 ( 
.A1(n_941),
.A2(n_946),
.A3(n_926),
.B1(n_922),
.B2(n_939),
.C1(n_949),
.C2(n_938),
.Y(n_954)
);

AOI32xp33_ASAP7_75t_L g955 ( 
.A1(n_945),
.A2(n_915),
.A3(n_929),
.B1(n_930),
.B2(n_924),
.Y(n_955)
);

INVx2_ASAP7_75t_SL g956 ( 
.A(n_942),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_943),
.Y(n_957)
);

NAND4xp75_ASAP7_75t_L g958 ( 
.A(n_941),
.B(n_906),
.C(n_920),
.D(n_919),
.Y(n_958)
);

INVx2_ASAP7_75t_L g959 ( 
.A(n_943),
.Y(n_959)
);

AND2x2_ASAP7_75t_L g960 ( 
.A(n_948),
.B(n_918),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_947),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_951),
.Y(n_962)
);

INVx2_ASAP7_75t_SL g963 ( 
.A(n_956),
.Y(n_963)
);

AOI211xp5_ASAP7_75t_SL g964 ( 
.A1(n_954),
.A2(n_944),
.B(n_950),
.C(n_899),
.Y(n_964)
);

OAI21xp5_ASAP7_75t_L g965 ( 
.A1(n_958),
.A2(n_940),
.B(n_944),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_952),
.B(n_900),
.Y(n_966)
);

AND2x2_ASAP7_75t_L g967 ( 
.A(n_952),
.B(n_85),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_953),
.Y(n_968)
);

INVxp67_ASAP7_75t_L g969 ( 
.A(n_961),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_957),
.Y(n_970)
);

OAI22xp5_ASAP7_75t_L g971 ( 
.A1(n_955),
.A2(n_679),
.B1(n_91),
.B2(n_93),
.Y(n_971)
);

AOI22xp33_ASAP7_75t_L g972 ( 
.A1(n_960),
.A2(n_103),
.B1(n_105),
.B2(n_107),
.Y(n_972)
);

OA22x2_ASAP7_75t_L g973 ( 
.A1(n_962),
.A2(n_959),
.B1(n_110),
.B2(n_111),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_953),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_968),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_974),
.Y(n_976)
);

AND2x2_ASAP7_75t_L g977 ( 
.A(n_963),
.B(n_114),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_970),
.Y(n_978)
);

OR2x2_ASAP7_75t_L g979 ( 
.A(n_969),
.B(n_120),
.Y(n_979)
);

OR2x2_ASAP7_75t_L g980 ( 
.A(n_966),
.B(n_129),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_967),
.Y(n_981)
);

NAND2xp33_ASAP7_75t_SL g982 ( 
.A(n_965),
.B(n_132),
.Y(n_982)
);

NAND2xp33_ASAP7_75t_SL g983 ( 
.A(n_971),
.B(n_964),
.Y(n_983)
);

INVx1_ASAP7_75t_SL g984 ( 
.A(n_973),
.Y(n_984)
);

INVx1_ASAP7_75t_SL g985 ( 
.A(n_972),
.Y(n_985)
);

AOI211xp5_ASAP7_75t_L g986 ( 
.A1(n_983),
.A2(n_139),
.B(n_147),
.C(n_152),
.Y(n_986)
);

NOR2xp33_ASAP7_75t_L g987 ( 
.A(n_984),
.B(n_153),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_975),
.Y(n_988)
);

INVxp67_ASAP7_75t_L g989 ( 
.A(n_987),
.Y(n_989)
);

NOR2xp33_ASAP7_75t_L g990 ( 
.A(n_988),
.B(n_981),
.Y(n_990)
);

NOR3xp33_ASAP7_75t_L g991 ( 
.A(n_986),
.B(n_985),
.C(n_982),
.Y(n_991)
);

AOI211xp5_ASAP7_75t_L g992 ( 
.A1(n_991),
.A2(n_979),
.B(n_980),
.C(n_977),
.Y(n_992)
);

OAI21xp5_ASAP7_75t_SL g993 ( 
.A1(n_989),
.A2(n_976),
.B(n_978),
.Y(n_993)
);

AND2x2_ASAP7_75t_L g994 ( 
.A(n_992),
.B(n_990),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_993),
.Y(n_995)
);

OR2x2_ASAP7_75t_L g996 ( 
.A(n_995),
.B(n_250),
.Y(n_996)
);

CKINVDCx5p33_ASAP7_75t_R g997 ( 
.A(n_996),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_997),
.Y(n_998)
);

CKINVDCx20_ASAP7_75t_R g999 ( 
.A(n_998),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_999),
.B(n_994),
.Y(n_1000)
);

AOI21xp33_ASAP7_75t_SL g1001 ( 
.A1(n_1000),
.A2(n_160),
.B(n_161),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_1001),
.B(n_166),
.Y(n_1002)
);

AOI322xp5_ASAP7_75t_SL g1003 ( 
.A1(n_1002),
.A2(n_183),
.A3(n_185),
.B1(n_191),
.B2(n_194),
.C1(n_199),
.C2(n_204),
.Y(n_1003)
);

AOI222xp33_ASAP7_75t_L g1004 ( 
.A1(n_1003),
.A2(n_207),
.B1(n_216),
.B2(n_219),
.C1(n_222),
.C2(n_224),
.Y(n_1004)
);

AOI22xp5_ASAP7_75t_L g1005 ( 
.A1(n_1004),
.A2(n_231),
.B1(n_232),
.B2(n_233),
.Y(n_1005)
);


endmodule