module real_jpeg_26174_n_18 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_364, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;
input n_364;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_356;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp33_ASAP7_75t_L g34 ( 
.A1(n_0),
.A2(n_35),
.B1(n_36),
.B2(n_38),
.Y(n_34)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

AOI21xp5_ASAP7_75t_L g53 ( 
.A1(n_0),
.A2(n_42),
.B(n_47),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_0),
.B(n_58),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_0),
.A2(n_68),
.B1(n_93),
.B2(n_98),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_0),
.A2(n_110),
.B(n_114),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_0),
.B(n_148),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_1),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_2),
.A2(n_35),
.B1(n_36),
.B2(n_51),
.Y(n_50)
);

CKINVDCx14_ASAP7_75t_R g51 ( 
.A(n_2),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_2),
.A2(n_46),
.B1(n_47),
.B2(n_51),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_2),
.A2(n_51),
.B1(n_110),
.B2(n_111),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_2),
.A2(n_51),
.B1(n_206),
.B2(n_207),
.Y(n_209)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_3),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_L g18 ( 
.A1(n_4),
.A2(n_5),
.B1(n_19),
.B2(n_20),
.Y(n_18)
);

CKINVDCx12_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_6),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_7),
.A2(n_35),
.B1(n_36),
.B2(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_7),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_7),
.A2(n_46),
.B1(n_47),
.B2(n_65),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_7),
.A2(n_65),
.B1(n_110),
.B2(n_111),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_7),
.A2(n_65),
.B1(n_203),
.B2(n_206),
.Y(n_223)
);

INVx8_ASAP7_75t_SL g152 ( 
.A(n_8),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_9),
.A2(n_46),
.B1(n_47),
.B2(n_76),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_9),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_9),
.A2(n_35),
.B1(n_36),
.B2(n_76),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_9),
.A2(n_76),
.B1(n_110),
.B2(n_111),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_9),
.A2(n_76),
.B1(n_175),
.B2(n_263),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_10),
.A2(n_46),
.B1(n_47),
.B2(n_133),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_10),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_10),
.A2(n_35),
.B1(n_36),
.B2(n_133),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_10),
.A2(n_110),
.B1(n_111),
.B2(n_133),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_10),
.A2(n_133),
.B1(n_206),
.B2(n_292),
.Y(n_291)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_11),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_12),
.A2(n_46),
.B1(n_47),
.B2(n_186),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_12),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_12),
.A2(n_35),
.B1(n_36),
.B2(n_186),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_12),
.A2(n_110),
.B1(n_111),
.B2(n_186),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g328 ( 
.A1(n_12),
.A2(n_186),
.B1(n_207),
.B2(n_263),
.Y(n_328)
);

INVx13_ASAP7_75t_L g177 ( 
.A(n_13),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_13),
.B(n_38),
.Y(n_178)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_L g156 ( 
.A1(n_15),
.A2(n_46),
.B1(n_47),
.B2(n_157),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_15),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_15),
.A2(n_35),
.B1(n_36),
.B2(n_157),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g265 ( 
.A1(n_15),
.A2(n_110),
.B1(n_111),
.B2(n_157),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_SL g312 ( 
.A1(n_15),
.A2(n_157),
.B1(n_175),
.B2(n_176),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_16),
.A2(n_46),
.B1(n_47),
.B2(n_73),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_16),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_16),
.A2(n_35),
.B1(n_36),
.B2(n_73),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_16),
.A2(n_73),
.B1(n_110),
.B2(n_111),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_16),
.A2(n_73),
.B1(n_177),
.B2(n_206),
.Y(n_238)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_17),
.Y(n_71)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_17),
.Y(n_78)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_17),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_360),
.C(n_361),
.Y(n_20)
);

OAI21xp5_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_356),
.B(n_359),
.Y(n_21)
);

AOI21xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_342),
.B(n_355),
.Y(n_22)
);

OAI321xp33_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_307),
.A3(n_335),
.B1(n_340),
.B2(n_341),
.C(n_364),
.Y(n_23)
);

AOI311xp33_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_253),
.A3(n_297),
.B(n_301),
.C(n_302),
.Y(n_24)
);

NOR3xp33_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_211),
.C(n_248),
.Y(n_25)
);

AOI21xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_169),
.B(n_210),
.Y(n_26)
);

OAI21xp5_ASAP7_75t_SL g27 ( 
.A1(n_28),
.A2(n_137),
.B(n_168),
.Y(n_27)
);

AOI21xp5_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_104),
.B(n_136),
.Y(n_28)
);

OAI21xp5_ASAP7_75t_SL g29 ( 
.A1(n_30),
.A2(n_79),
.B(n_103),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_54),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_31),
.B(n_54),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_32),
.B(n_52),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_32),
.A2(n_33),
.B1(n_52),
.B2(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_34),
.A2(n_39),
.B1(n_45),
.B2(n_49),
.Y(n_33)
);

OAI22xp33_ASAP7_75t_L g41 ( 
.A1(n_35),
.A2(n_36),
.B1(n_42),
.B2(n_44),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_35),
.A2(n_36),
.B1(n_60),
.B2(n_61),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_35),
.B(n_61),
.Y(n_126)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

A2O1A1Ixp33_ASAP7_75t_SL g52 ( 
.A1(n_36),
.A2(n_38),
.B(n_44),
.C(n_53),
.Y(n_52)
);

OAI32xp33_ASAP7_75t_L g125 ( 
.A1(n_36),
.A2(n_60),
.A3(n_110),
.B1(n_115),
.B2(n_126),
.Y(n_125)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_38),
.B(n_45),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_38),
.B(n_71),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_38),
.B(n_111),
.Y(n_115)
);

OAI21xp33_ASAP7_75t_L g205 ( 
.A1(n_38),
.A2(n_178),
.B(n_206),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_39),
.A2(n_163),
.B(n_164),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_39),
.A2(n_45),
.B1(n_229),
.B2(n_246),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_39),
.A2(n_246),
.B(n_272),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_40),
.A2(n_50),
.B1(n_63),
.B2(n_64),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_40),
.A2(n_63),
.B1(n_64),
.B2(n_121),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_40),
.A2(n_165),
.B(n_197),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_40),
.B(n_231),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_40),
.A2(n_63),
.B(n_165),
.Y(n_316)
);

AND2x2_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_45),
.Y(n_40)
);

INVx13_ASAP7_75t_L g44 ( 
.A(n_42),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_42),
.A2(n_44),
.B1(n_46),
.B2(n_47),
.Y(n_45)
);

BUFx24_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_45),
.B(n_198),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_45),
.A2(n_229),
.B(n_230),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_46),
.B(n_70),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_46),
.B(n_100),
.Y(n_99)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

CKINVDCx16_ASAP7_75t_R g49 ( 
.A(n_50),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_52),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_67),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_56),
.A2(n_57),
.B1(n_62),
.B2(n_66),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_56),
.B(n_66),
.C(n_67),
.Y(n_105)
);

CKINVDCx14_ASAP7_75t_R g56 ( 
.A(n_57),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_58),
.A2(n_117),
.B1(n_143),
.B2(n_144),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_58),
.A2(n_117),
.B1(n_144),
.B2(n_195),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_58),
.B(n_241),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_58),
.A2(n_117),
.B1(n_279),
.B2(n_280),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_L g351 ( 
.A1(n_58),
.A2(n_117),
.B(n_352),
.Y(n_351)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_59),
.A2(n_109),
.B1(n_116),
.B2(n_119),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_59),
.B(n_118),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_59),
.B(n_220),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g264 ( 
.A1(n_59),
.A2(n_265),
.B(n_266),
.Y(n_264)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_60),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_60),
.A2(n_61),
.B1(n_110),
.B2(n_111),
.Y(n_118)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_62),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_63),
.B(n_165),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g67 ( 
.A1(n_68),
.A2(n_72),
.B(n_74),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_68),
.A2(n_83),
.B1(n_93),
.B2(n_94),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_68),
.A2(n_128),
.B(n_129),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_68),
.A2(n_129),
.B(n_227),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_68),
.A2(n_128),
.B(n_155),
.Y(n_269)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_69),
.A2(n_82),
.B1(n_84),
.B2(n_85),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_69),
.B(n_132),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_69),
.A2(n_181),
.B1(n_182),
.B2(n_185),
.Y(n_180)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_70),
.Y(n_155)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx8_ASAP7_75t_L g184 ( 
.A(n_71),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_72),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_74),
.B(n_158),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_75),
.B(n_77),
.Y(n_74)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_75),
.Y(n_128)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

BUFx2_ASAP7_75t_L g131 ( 
.A(n_78),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_89),
.B(n_102),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_87),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_81),
.B(n_87),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_83),
.Y(n_82)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_85),
.Y(n_98)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_86),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g89 ( 
.A1(n_90),
.A2(n_96),
.B(n_101),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_92),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_91),
.B(n_92),
.Y(n_101)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_97),
.B(n_99),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_106),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_105),
.B(n_106),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_107),
.A2(n_124),
.B1(n_134),
.B2(n_135),
.Y(n_106)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_107),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_120),
.B1(n_122),
.B2(n_123),
.Y(n_107)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_108),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_110),
.A2(n_111),
.B1(n_150),
.B2(n_151),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_110),
.B(n_151),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_111),
.Y(n_110)
);

OAI32xp33_ASAP7_75t_L g174 ( 
.A1(n_111),
.A2(n_150),
.A3(n_175),
.B1(n_178),
.B2(n_179),
.Y(n_174)
);

BUFx12f_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

BUFx12f_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_115),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_116),
.A2(n_220),
.B(n_240),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_117),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_117),
.A2(n_195),
.B(n_219),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_117),
.B(n_241),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g317 ( 
.A1(n_117),
.A2(n_280),
.B(n_318),
.Y(n_317)
);

CKINVDCx14_ASAP7_75t_R g143 ( 
.A(n_119),
.Y(n_143)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_120),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_120),
.B(n_123),
.C(n_134),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_121),
.Y(n_163)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_124),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_127),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_125),
.B(n_127),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_132),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_131),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_139),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_138),
.B(n_139),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_140),
.A2(n_141),
.B1(n_159),
.B2(n_160),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_140),
.B(n_162),
.C(n_166),
.Y(n_170)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_SL g141 ( 
.A(n_142),
.B(n_145),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_142),
.B(n_147),
.C(n_153),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_146),
.A2(n_147),
.B1(n_153),
.B2(n_154),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_147),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_148),
.A2(n_200),
.B1(n_205),
.B2(n_209),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_148),
.A2(n_200),
.B1(n_209),
.B2(n_222),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_148),
.B(n_262),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_148),
.B(n_291),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_148),
.A2(n_200),
.B1(n_327),
.B2(n_328),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_SL g360 ( 
.A1(n_148),
.A2(n_200),
.B(n_262),
.Y(n_360)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_149),
.B(n_202),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_149),
.A2(n_201),
.B1(n_223),
.B2(n_238),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_149),
.A2(n_312),
.B(n_313),
.Y(n_311)
);

OAI22xp33_ASAP7_75t_L g202 ( 
.A1(n_150),
.A2(n_151),
.B1(n_203),
.B2(n_204),
.Y(n_202)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_154),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_156),
.B(n_158),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_156),
.Y(n_181)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_161),
.A2(n_162),
.B1(n_166),
.B2(n_167),
.Y(n_160)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_161),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_162),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g281 ( 
.A(n_164),
.B(n_230),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_171),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_170),
.B(n_171),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_192),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_173),
.A2(n_189),
.B1(n_190),
.B2(n_191),
.Y(n_172)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_173),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_173),
.B(n_191),
.C(n_192),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_174),
.A2(n_180),
.B1(n_187),
.B2(n_188),
.Y(n_173)
);

CKINVDCx14_ASAP7_75t_R g188 ( 
.A(n_174),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_174),
.B(n_187),
.Y(n_216)
);

INVx8_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx11_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx8_ASAP7_75t_L g204 ( 
.A(n_177),
.Y(n_204)
);

INVx6_ASAP7_75t_L g208 ( 
.A(n_177),
.Y(n_208)
);

INVx8_ASAP7_75t_L g263 ( 
.A(n_177),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_180),
.Y(n_187)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx5_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_185),
.Y(n_227)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_189),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_199),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_196),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_194),
.B(n_196),
.C(n_199),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_197),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_198),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_200),
.B(n_291),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g348 ( 
.A1(n_200),
.A2(n_328),
.B(n_349),
.Y(n_348)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_201),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_201),
.A2(n_238),
.B(n_261),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_201),
.A2(n_289),
.B(n_290),
.Y(n_288)
);

INVx4_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx8_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx8_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

AOI21xp33_ASAP7_75t_L g303 ( 
.A1(n_212),
.A2(n_304),
.B(n_305),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_232),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g305 ( 
.A(n_213),
.B(n_232),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_224),
.C(n_225),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_214),
.A2(n_215),
.B1(n_251),
.B2(n_252),
.Y(n_250)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_217),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_216),
.B(n_218),
.C(n_221),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_221),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_219),
.Y(n_332)
);

CKINVDCx16_ASAP7_75t_R g352 ( 
.A(n_220),
.Y(n_352)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_SL g252 ( 
.A(n_224),
.B(n_225),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_228),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_226),
.B(n_228),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_232),
.Y(n_299)
);

FAx1_ASAP7_75t_SL g232 ( 
.A(n_233),
.B(n_243),
.CI(n_247),
.CON(n_232),
.SN(n_232)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_234),
.A2(n_235),
.B1(n_236),
.B2(n_242),
.Y(n_233)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_234),
.Y(n_242)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_SL g236 ( 
.A(n_237),
.B(n_239),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_237),
.B(n_239),
.C(n_242),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_240),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_245),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_244),
.B(n_245),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_250),
.Y(n_248)
);

AND2x2_ASAP7_75t_L g304 ( 
.A(n_249),
.B(n_250),
.Y(n_304)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

O2A1O1Ixp33_ASAP7_75t_SL g302 ( 
.A1(n_254),
.A2(n_298),
.B(n_303),
.C(n_306),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_275),
.Y(n_254)
);

AND2x2_ASAP7_75t_L g301 ( 
.A(n_255),
.B(n_275),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_268),
.C(n_274),
.Y(n_255)
);

FAx1_ASAP7_75t_L g300 ( 
.A(n_256),
.B(n_268),
.CI(n_274),
.CON(n_300),
.SN(n_300)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_257),
.A2(n_258),
.B1(n_259),
.B2(n_267),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_257),
.B(n_260),
.C(n_264),
.Y(n_296)
);

CKINVDCx14_ASAP7_75t_R g257 ( 
.A(n_258),
.Y(n_257)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_259),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_SL g259 ( 
.A(n_260),
.B(n_264),
.Y(n_259)
);

AND2x2_ASAP7_75t_L g357 ( 
.A(n_261),
.B(n_313),
.Y(n_357)
);

CKINVDCx16_ASAP7_75t_R g289 ( 
.A(n_262),
.Y(n_289)
);

INVx11_ASAP7_75t_L g292 ( 
.A(n_263),
.Y(n_292)
);

CKINVDCx14_ASAP7_75t_R g279 ( 
.A(n_265),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_266),
.B(n_332),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_269),
.A2(n_270),
.B1(n_271),
.B2(n_273),
.Y(n_268)
);

CKINVDCx16_ASAP7_75t_R g273 ( 
.A(n_269),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_269),
.B(n_271),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_269),
.A2(n_273),
.B1(n_287),
.B2(n_288),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_L g322 ( 
.A1(n_273),
.A2(n_284),
.B(n_288),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_296),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_277),
.A2(n_283),
.B1(n_294),
.B2(n_295),
.Y(n_276)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_277),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_L g277 ( 
.A1(n_278),
.A2(n_281),
.B(n_282),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_278),
.B(n_281),
.Y(n_282)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_282),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_282),
.A2(n_309),
.B1(n_321),
.B2(n_339),
.Y(n_338)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_283),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_283),
.B(n_294),
.C(n_296),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_284),
.A2(n_285),
.B1(n_286),
.B2(n_293),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_286),
.Y(n_293)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_290),
.Y(n_349)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_300),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_299),
.B(n_300),
.Y(n_306)
);

BUFx24_ASAP7_75t_SL g362 ( 
.A(n_300),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_323),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_308),
.B(n_323),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_321),
.C(n_322),
.Y(n_308)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_309),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_310),
.A2(n_311),
.B1(n_314),
.B2(n_320),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_310),
.A2(n_311),
.B1(n_325),
.B2(n_333),
.Y(n_324)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_311),
.B(n_316),
.C(n_317),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_311),
.B(n_333),
.C(n_334),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_312),
.Y(n_327)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_314),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_315),
.A2(n_316),
.B1(n_317),
.B2(n_319),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_315),
.A2(n_316),
.B1(n_330),
.B2(n_331),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_315),
.B(n_326),
.C(n_330),
.Y(n_345)
);

CKINVDCx16_ASAP7_75t_R g315 ( 
.A(n_316),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_317),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_322),
.B(n_338),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_334),
.Y(n_323)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_325),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_SL g325 ( 
.A(n_326),
.B(n_329),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_331),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_336),
.B(n_337),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_336),
.B(n_337),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_343),
.B(n_354),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_SL g355 ( 
.A(n_343),
.B(n_354),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_344),
.A2(n_345),
.B1(n_346),
.B2(n_353),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_344),
.B(n_348),
.C(n_350),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_345),
.Y(n_344)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_346),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_L g346 ( 
.A1(n_347),
.A2(n_348),
.B1(n_350),
.B2(n_351),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_348),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_351),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_357),
.B(n_358),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_SL g359 ( 
.A(n_357),
.B(n_358),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_357),
.Y(n_361)
);


endmodule