module fake_jpeg_26688_n_295 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_295);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_295;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_122;
wire n_75;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_7),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_8),
.B(n_4),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx16f_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_2),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_13),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

INVx1_ASAP7_75t_SL g62 ( 
.A(n_35),
.Y(n_62)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

INVx6_ASAP7_75t_SL g40 ( 
.A(n_29),
.Y(n_40)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_16),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_41),
.B(n_42),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_16),
.Y(n_42)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_44),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_41),
.B(n_42),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_45),
.B(n_50),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_36),
.A2(n_18),
.B1(n_25),
.B2(n_33),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_49),
.A2(n_38),
.B1(n_35),
.B2(n_18),
.Y(n_67)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_51),
.Y(n_85)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_52),
.Y(n_75)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

BUFx2_ASAP7_75t_L g71 ( 
.A(n_53),
.Y(n_71)
);

BUFx2_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

HB1xp67_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

OR2x2_ASAP7_75t_L g55 ( 
.A(n_42),
.B(n_27),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_55),
.B(n_59),
.Y(n_83)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_57),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_36),
.B(n_27),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_36),
.B(n_28),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_60),
.B(n_61),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_38),
.B(n_28),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_35),
.A2(n_18),
.B1(n_25),
.B2(n_32),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_65),
.A2(n_40),
.B1(n_33),
.B2(n_22),
.Y(n_87)
);

O2A1O1Ixp33_ASAP7_75t_L g66 ( 
.A1(n_63),
.A2(n_35),
.B(n_38),
.C(n_25),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_66),
.A2(n_74),
.B(n_86),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_67),
.B(n_87),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_59),
.A2(n_17),
.B1(n_30),
.B2(n_20),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_70),
.A2(n_23),
.B1(n_21),
.B2(n_31),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_63),
.B(n_20),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_73),
.B(n_82),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_49),
.B(n_39),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_54),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_76),
.B(n_80),
.Y(n_106)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_54),
.Y(n_78)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_78),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_56),
.Y(n_80)
);

A2O1A1Ixp33_ASAP7_75t_L g82 ( 
.A1(n_55),
.A2(n_32),
.B(n_21),
.C(n_22),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_50),
.A2(n_33),
.B1(n_22),
.B2(n_21),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_84),
.A2(n_55),
.B1(n_31),
.B2(n_23),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_58),
.B(n_39),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_58),
.B(n_39),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_88),
.B(n_57),
.C(n_52),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_43),
.Y(n_89)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_89),
.Y(n_108)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_62),
.Y(n_90)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_90),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_78),
.A2(n_46),
.B1(n_56),
.B2(n_53),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_92),
.A2(n_46),
.B1(n_47),
.B2(n_48),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_72),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_93),
.B(n_97),
.Y(n_140)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_86),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_94),
.B(n_95),
.Y(n_121)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_86),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_83),
.B(n_84),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_96),
.B(n_102),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_88),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_99),
.A2(n_103),
.B1(n_111),
.B2(n_44),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_67),
.B(n_64),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_100),
.A2(n_37),
.B(n_80),
.Y(n_131)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_88),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_101),
.B(n_104),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_77),
.B(n_74),
.Y(n_102)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_71),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_74),
.B(n_64),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_105),
.B(n_107),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_66),
.B(n_62),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_69),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_110),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_68),
.A2(n_47),
.B1(n_48),
.B2(n_51),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_82),
.B(n_23),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_113),
.B(n_116),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_114),
.B(n_109),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_76),
.B(n_26),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_102),
.B(n_90),
.C(n_68),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_117),
.B(n_142),
.C(n_114),
.Y(n_147)
);

BUFx24_ASAP7_75t_SL g118 ( 
.A(n_112),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_118),
.B(n_130),
.Y(n_171)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_105),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_119),
.B(n_128),
.Y(n_146)
);

OA21x2_ASAP7_75t_L g120 ( 
.A1(n_107),
.A2(n_71),
.B(n_37),
.Y(n_120)
);

AO22x1_ASAP7_75t_L g167 ( 
.A1(n_120),
.A2(n_37),
.B1(n_79),
.B2(n_81),
.Y(n_167)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_108),
.Y(n_122)
);

INVx2_ASAP7_75t_SL g168 ( 
.A(n_122),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_106),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_124),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_106),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_126),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_112),
.B(n_17),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_116),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_131),
.A2(n_132),
.B(n_134),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_109),
.A2(n_0),
.B(n_1),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_111),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_133),
.B(n_137),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_135),
.A2(n_98),
.B1(n_103),
.B2(n_99),
.Y(n_153)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_108),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_136),
.A2(n_79),
.B1(n_30),
.B2(n_17),
.Y(n_170)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_100),
.Y(n_137)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_100),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_139),
.B(n_100),
.Y(n_150)
);

BUFx3_ASAP7_75t_L g141 ( 
.A(n_91),
.Y(n_141)
);

INVx3_ASAP7_75t_SL g165 ( 
.A(n_141),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_94),
.B(n_101),
.C(n_95),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_143),
.A2(n_98),
.B1(n_92),
.B2(n_104),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_138),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_144),
.B(n_127),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_SL g145 ( 
.A(n_135),
.B(n_127),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_145),
.B(n_147),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_133),
.A2(n_139),
.B1(n_137),
.B2(n_119),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_148),
.A2(n_156),
.B1(n_162),
.B2(n_141),
.Y(n_192)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_150),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_129),
.B(n_96),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_151),
.B(n_155),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_142),
.B(n_113),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_152),
.B(n_29),
.C(n_24),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_153),
.Y(n_175)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_138),
.Y(n_155)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_120),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_158),
.B(n_166),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_132),
.A2(n_98),
.B(n_115),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_159),
.A2(n_140),
.B(n_123),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_135),
.A2(n_98),
.B1(n_75),
.B2(n_91),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_161),
.A2(n_163),
.B1(n_172),
.B2(n_121),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_143),
.A2(n_75),
.B1(n_115),
.B2(n_85),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_125),
.A2(n_85),
.B1(n_81),
.B2(n_89),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_124),
.A2(n_24),
.B1(n_30),
.B2(n_17),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_164),
.Y(n_182)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_120),
.Y(n_166)
);

AOI22x1_ASAP7_75t_L g178 ( 
.A1(n_167),
.A2(n_120),
.B1(n_134),
.B2(n_131),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_126),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_169),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_170),
.A2(n_122),
.B1(n_136),
.B2(n_130),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_125),
.A2(n_30),
.B1(n_29),
.B2(n_24),
.Y(n_172)
);

BUFx3_ASAP7_75t_L g173 ( 
.A(n_145),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_173),
.B(n_177),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_174),
.A2(n_181),
.B1(n_188),
.B2(n_162),
.Y(n_210)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_149),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_178),
.A2(n_192),
.B1(n_198),
.B2(n_164),
.Y(n_211)
);

INVx2_ASAP7_75t_SL g179 ( 
.A(n_168),
.Y(n_179)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_179),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_160),
.B(n_128),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_180),
.B(n_183),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_160),
.B(n_154),
.Y(n_184)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_184),
.Y(n_212)
);

BUFx24_ASAP7_75t_SL g185 ( 
.A(n_171),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_185),
.B(n_189),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_158),
.A2(n_117),
.B1(n_129),
.B2(n_121),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_149),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_163),
.Y(n_190)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_190),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_191),
.A2(n_167),
.B(n_172),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_193),
.B(n_168),
.C(n_165),
.Y(n_221)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_146),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_194),
.B(n_146),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_148),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g199 ( 
.A(n_195),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_166),
.A2(n_29),
.B1(n_26),
.B2(n_8),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_SL g201 ( 
.A(n_187),
.B(n_147),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_201),
.B(n_204),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_187),
.B(n_152),
.C(n_161),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_202),
.B(n_216),
.C(n_26),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_SL g203 ( 
.A(n_173),
.B(n_159),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_SL g234 ( 
.A(n_203),
.B(n_29),
.C(n_165),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_188),
.B(n_157),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_191),
.B(n_157),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_205),
.B(n_209),
.Y(n_236)
);

BUFx2_ASAP7_75t_L g207 ( 
.A(n_178),
.Y(n_207)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_207),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_208),
.B(n_220),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_193),
.B(n_151),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_210),
.B(n_182),
.Y(n_231)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_211),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_196),
.B(n_153),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_214),
.B(n_221),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_176),
.B(n_155),
.C(n_150),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_197),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_217),
.B(n_15),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_218),
.A2(n_0),
.B(n_1),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_175),
.A2(n_167),
.B1(n_165),
.B2(n_168),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_221),
.A2(n_175),
.B(n_186),
.Y(n_223)
);

AOI21xp33_ASAP7_75t_L g245 ( 
.A1(n_223),
.A2(n_215),
.B(n_214),
.Y(n_245)
);

AO22x2_ASAP7_75t_L g224 ( 
.A1(n_207),
.A2(n_178),
.B1(n_197),
.B2(n_203),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_224),
.A2(n_233),
.B1(n_213),
.B2(n_199),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_201),
.B(n_181),
.C(n_192),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_225),
.B(n_228),
.Y(n_244)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_219),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_227),
.B(n_10),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_202),
.B(n_196),
.C(n_176),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_231),
.A2(n_6),
.B1(n_14),
.B2(n_12),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_212),
.B(n_179),
.Y(n_232)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_232),
.Y(n_243)
);

A2O1A1Ixp33_ASAP7_75t_SL g233 ( 
.A1(n_218),
.A2(n_182),
.B(n_198),
.C(n_179),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_SL g241 ( 
.A(n_234),
.B(n_205),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_235),
.B(n_0),
.Y(n_253)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_237),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_209),
.B(n_7),
.C(n_14),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_239),
.B(n_206),
.C(n_9),
.Y(n_247)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_240),
.Y(n_252)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_241),
.Y(n_264)
);

OR2x2_ASAP7_75t_L g260 ( 
.A(n_242),
.B(n_249),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_245),
.A2(n_238),
.B(n_229),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_222),
.A2(n_204),
.B1(n_200),
.B2(n_216),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_246),
.A2(n_224),
.B1(n_226),
.B2(n_233),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_247),
.B(n_253),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_235),
.B(n_6),
.C(n_14),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_250),
.B(n_239),
.C(n_233),
.Y(n_255)
);

OAI221xp5_ASAP7_75t_SL g251 ( 
.A1(n_224),
.A2(n_5),
.B1(n_12),
.B2(n_10),
.C(n_9),
.Y(n_251)
);

NOR3xp33_ASAP7_75t_L g261 ( 
.A(n_251),
.B(n_224),
.C(n_233),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_254),
.B(n_10),
.Y(n_257)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_255),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_246),
.B(n_230),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_256),
.B(n_258),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_257),
.B(n_259),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_241),
.B(n_230),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_247),
.B(n_242),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_261),
.B(n_265),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_263),
.A2(n_248),
.B1(n_250),
.B2(n_252),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_244),
.B(n_236),
.C(n_243),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_266),
.B(n_253),
.C(n_236),
.Y(n_272)
);

NOR2xp67_ASAP7_75t_L g269 ( 
.A(n_266),
.B(n_248),
.Y(n_269)
);

NOR2xp67_ASAP7_75t_R g281 ( 
.A(n_269),
.B(n_0),
.Y(n_281)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_260),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_270),
.B(n_271),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_272),
.B(n_275),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_262),
.B(n_255),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_256),
.B(n_12),
.C(n_15),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_276),
.B(n_274),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_268),
.A2(n_260),
.B1(n_264),
.B2(n_258),
.Y(n_277)
);

OR2x2_ASAP7_75t_L g284 ( 
.A(n_277),
.B(n_280),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_273),
.A2(n_15),
.B1(n_2),
.B2(n_3),
.Y(n_280)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_281),
.Y(n_288)
);

AND2x2_ASAP7_75t_L g287 ( 
.A(n_282),
.B(n_283),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_267),
.B(n_2),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_279),
.B(n_270),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_285),
.B(n_286),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_278),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_284),
.B(n_282),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_290),
.A2(n_287),
.B(n_289),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_291),
.A2(n_272),
.B1(n_276),
.B2(n_288),
.Y(n_292)
);

OAI321xp33_ASAP7_75t_L g293 ( 
.A1(n_292),
.A2(n_3),
.A3(n_4),
.B1(n_283),
.B2(n_278),
.C(n_285),
.Y(n_293)
);

BUFx24_ASAP7_75t_SL g294 ( 
.A(n_293),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_294),
.A2(n_3),
.B(n_4),
.Y(n_295)
);


endmodule