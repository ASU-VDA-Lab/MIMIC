module real_aes_659_n_78 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_77, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_78);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_78;
wire n_480;
wire n_113;
wire n_476;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_522;
wire n_485;
wire n_222;
wire n_287;
wire n_357;
wire n_503;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_341;
wire n_232;
wire n_460;
wire n_401;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_320;
wire n_260;
wire n_97;
wire n_186;
wire n_138;
wire n_379;
wire n_453;
wire n_374;
wire n_235;
wire n_399;
wire n_378;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_145;
wire n_415;
wire n_227;
wire n_92;
wire n_519;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_292;
wire n_400;
wire n_116;
wire n_94;
wire n_289;
wire n_462;
wire n_280;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_408;
wire n_184;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_530;
wire n_104;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_506;
wire n_513;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_164;
wire n_231;
wire n_102;
wire n_454;
wire n_122;
wire n_443;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_204;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_331;
wire n_93;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_323;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_368;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_250;
wire n_85;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_402;
wire n_87;
wire n_171;
wire n_531;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_488;
wire n_501;
wire n_251;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_158;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_109;
wire n_203;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_526;
wire n_155;
wire n_243;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_249;
wire n_446;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_180;
wire n_212;
wire n_210;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_103;
wire n_166;
wire n_224;
wire n_151;
wire n_130;
wire n_253;
wire n_459;
wire n_99;
wire n_440;
wire n_525;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_305;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_473;
wire n_465;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_340;
wire n_483;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_206;
wire n_307;
wire n_500;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_264;
wire n_237;
wire n_91;
NAND2xp5_ASAP7_75t_L g314 ( .A(n_0), .B(n_224), .Y(n_314) );
AOI22xp5_ASAP7_75t_L g514 ( .A1(n_0), .A2(n_81), .B1(n_165), .B2(n_515), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_0), .Y(n_515) );
AO22x2_ASAP7_75t_L g102 ( .A1(n_1), .A2(n_55), .B1(n_92), .B2(n_103), .Y(n_102) );
INVx1_ASAP7_75t_L g192 ( .A(n_2), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_3), .B(n_213), .Y(n_267) );
NAND2xp33_ASAP7_75t_SL g260 ( .A(n_4), .B(n_219), .Y(n_260) );
AOI22xp5_ASAP7_75t_L g171 ( .A1(n_5), .A2(n_172), .B1(n_173), .B2(n_179), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_5), .Y(n_172) );
AO22x2_ASAP7_75t_L g99 ( .A1(n_6), .A2(n_18), .B1(n_92), .B2(n_100), .Y(n_99) );
AND2x2_ASAP7_75t_L g265 ( .A(n_7), .B(n_204), .Y(n_265) );
INVx2_ASAP7_75t_L g205 ( .A(n_8), .Y(n_205) );
AOI22xp33_ASAP7_75t_L g151 ( .A1(n_9), .A2(n_57), .B1(n_152), .B2(n_155), .Y(n_151) );
AOI22xp33_ASAP7_75t_L g105 ( .A1(n_10), .A2(n_59), .B1(n_106), .B2(n_111), .Y(n_105) );
AOI221x1_ASAP7_75t_L g254 ( .A1(n_11), .A2(n_208), .B1(n_255), .B2(n_257), .C(n_259), .Y(n_254) );
NAND2xp5_ASAP7_75t_SL g230 ( .A(n_12), .B(n_213), .Y(n_230) );
AOI22xp33_ASAP7_75t_L g117 ( .A1(n_13), .A2(n_46), .B1(n_118), .B2(n_120), .Y(n_117) );
AOI221xp5_ASAP7_75t_SL g207 ( .A1(n_14), .A2(n_31), .B1(n_208), .B2(n_213), .C(n_220), .Y(n_207) );
AOI21xp5_ASAP7_75t_L g268 ( .A1(n_15), .A2(n_208), .B(n_269), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_16), .B(n_224), .Y(n_270) );
AOI22xp33_ASAP7_75t_L g135 ( .A1(n_17), .A2(n_54), .B1(n_136), .B2(n_138), .Y(n_135) );
OAI221xp5_ASAP7_75t_L g184 ( .A1(n_18), .A2(n_55), .B1(n_58), .B2(n_185), .C(n_187), .Y(n_184) );
OR2x2_ASAP7_75t_L g206 ( .A(n_19), .B(n_71), .Y(n_206) );
OA21x2_ASAP7_75t_L g236 ( .A1(n_19), .A2(n_71), .B(n_205), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_20), .B(n_222), .Y(n_234) );
INVxp67_ASAP7_75t_L g253 ( .A(n_21), .Y(n_253) );
AOI22xp33_ASAP7_75t_L g158 ( .A1(n_22), .A2(n_61), .B1(n_159), .B2(n_161), .Y(n_158) );
AND2x2_ASAP7_75t_L g303 ( .A(n_23), .B(n_203), .Y(n_303) );
INVx3_ASAP7_75t_L g92 ( .A(n_24), .Y(n_92) );
AOI21xp5_ASAP7_75t_L g312 ( .A1(n_25), .A2(n_208), .B(n_313), .Y(n_312) );
AOI22xp33_ASAP7_75t_L g124 ( .A1(n_26), .A2(n_60), .B1(n_125), .B2(n_130), .Y(n_124) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_27), .B(n_222), .Y(n_221) );
AOI22xp33_ASAP7_75t_R g80 ( .A1(n_28), .A2(n_81), .B1(n_164), .B2(n_165), .Y(n_80) );
INVx1_ASAP7_75t_L g164 ( .A(n_28), .Y(n_164) );
INVx1_ASAP7_75t_SL g93 ( .A(n_29), .Y(n_93) );
INVx1_ASAP7_75t_L g194 ( .A(n_30), .Y(n_194) );
AND2x2_ASAP7_75t_L g209 ( .A(n_30), .B(n_210), .Y(n_209) );
AND2x2_ASAP7_75t_L g219 ( .A(n_30), .B(n_192), .Y(n_219) );
AOI22xp5_ASAP7_75t_L g287 ( .A1(n_32), .A2(n_64), .B1(n_208), .B2(n_248), .Y(n_287) );
AOI22xp5_ASAP7_75t_L g168 ( .A1(n_33), .A2(n_35), .B1(n_169), .B2(n_170), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_33), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_34), .B(n_224), .Y(n_301) );
INVx1_ASAP7_75t_L g170 ( .A(n_35), .Y(n_170) );
AOI22xp5_ASAP7_75t_L g175 ( .A1(n_36), .A2(n_42), .B1(n_176), .B2(n_177), .Y(n_175) );
INVx1_ASAP7_75t_L g177 ( .A(n_36), .Y(n_177) );
AO22x2_ASAP7_75t_L g95 ( .A1(n_37), .A2(n_58), .B1(n_92), .B2(n_96), .Y(n_95) );
OAI22xp5_ASAP7_75t_L g523 ( .A1(n_38), .A2(n_81), .B1(n_165), .B2(n_524), .Y(n_523) );
CKINVDCx20_ASAP7_75t_R g524 ( .A(n_38), .Y(n_524) );
AND2x2_ASAP7_75t_L g317 ( .A(n_39), .B(n_203), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_40), .B(n_203), .Y(n_226) );
AOI22xp5_ASAP7_75t_L g142 ( .A1(n_41), .A2(n_69), .B1(n_143), .B2(n_147), .Y(n_142) );
INVx1_ASAP7_75t_L g176 ( .A(n_42), .Y(n_176) );
INVx1_ASAP7_75t_L g212 ( .A(n_43), .Y(n_212) );
INVx1_ASAP7_75t_L g216 ( .A(n_43), .Y(n_216) );
INVx1_ASAP7_75t_L g94 ( .A(n_44), .Y(n_94) );
NAND2xp5_ASAP7_75t_SL g302 ( .A(n_45), .B(n_213), .Y(n_302) );
AND2x2_ASAP7_75t_L g281 ( .A(n_47), .B(n_203), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_48), .B(n_222), .Y(n_315) );
AND2x2_ASAP7_75t_SL g237 ( .A(n_49), .B(n_204), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_50), .B(n_224), .Y(n_278) );
AOI21xp5_ASAP7_75t_L g298 ( .A1(n_51), .A2(n_208), .B(n_299), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_52), .B(n_222), .Y(n_271) );
AND2x2_ASAP7_75t_SL g288 ( .A(n_53), .B(n_235), .Y(n_288) );
INVxp33_ASAP7_75t_L g189 ( .A(n_55), .Y(n_189) );
INVx1_ASAP7_75t_L g210 ( .A(n_56), .Y(n_210) );
INVx1_ASAP7_75t_L g218 ( .A(n_56), .Y(n_218) );
INVxp67_ASAP7_75t_L g188 ( .A(n_58), .Y(n_188) );
AOI22xp5_ASAP7_75t_L g173 ( .A1(n_62), .A2(n_174), .B1(n_175), .B2(n_178), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_62), .Y(n_174) );
AOI22xp5_ASAP7_75t_L g286 ( .A1(n_62), .A2(n_65), .B1(n_213), .B2(n_244), .Y(n_286) );
NAND2xp5_ASAP7_75t_SL g279 ( .A(n_63), .B(n_213), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_66), .B(n_224), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_67), .B(n_224), .Y(n_223) );
CKINVDCx20_ASAP7_75t_R g104 ( .A(n_68), .Y(n_104) );
AOI21xp5_ASAP7_75t_L g275 ( .A1(n_70), .A2(n_208), .B(n_276), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_72), .B(n_222), .Y(n_277) );
INVxp67_ASAP7_75t_L g256 ( .A(n_73), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_74), .B(n_213), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_75), .B(n_222), .Y(n_300) );
AOI21xp5_ASAP7_75t_L g231 ( .A1(n_76), .A2(n_208), .B(n_232), .Y(n_231) );
BUFx2_ASAP7_75t_SL g186 ( .A(n_77), .Y(n_186) );
AOI221xp5_ASAP7_75t_L g78 ( .A1(n_79), .A2(n_181), .B1(n_195), .B2(n_510), .C(n_513), .Y(n_78) );
XOR2xp5_ASAP7_75t_L g79 ( .A(n_80), .B(n_166), .Y(n_79) );
HB1xp67_ASAP7_75t_L g81 ( .A(n_82), .Y(n_81) );
INVx2_ASAP7_75t_SL g165 ( .A(n_82), .Y(n_165) );
AND2x2_ASAP7_75t_L g82 ( .A(n_83), .B(n_133), .Y(n_82) );
NOR2xp33_ASAP7_75t_L g83 ( .A(n_84), .B(n_116), .Y(n_83) );
OAI21xp33_ASAP7_75t_SL g84 ( .A1(n_85), .A2(n_104), .B(n_105), .Y(n_84) );
INVx2_ASAP7_75t_L g85 ( .A(n_86), .Y(n_85) );
INVx3_ASAP7_75t_SL g86 ( .A(n_87), .Y(n_86) );
INVx6_ASAP7_75t_L g87 ( .A(n_88), .Y(n_87) );
AND2x2_ASAP7_75t_L g88 ( .A(n_89), .B(n_97), .Y(n_88) );
AND2x4_ASAP7_75t_L g140 ( .A(n_89), .B(n_141), .Y(n_140) );
AND2x4_ASAP7_75t_L g144 ( .A(n_89), .B(n_145), .Y(n_144) );
AND2x2_ASAP7_75t_L g89 ( .A(n_90), .B(n_95), .Y(n_89) );
AND2x2_ASAP7_75t_L g109 ( .A(n_90), .B(n_110), .Y(n_109) );
HB1xp67_ASAP7_75t_L g115 ( .A(n_90), .Y(n_115) );
INVx2_ASAP7_75t_L g123 ( .A(n_90), .Y(n_123) );
OAI22x1_ASAP7_75t_L g90 ( .A1(n_91), .A2(n_92), .B1(n_93), .B2(n_94), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_92), .Y(n_91) );
INVx1_ASAP7_75t_L g96 ( .A(n_92), .Y(n_96) );
INVx2_ASAP7_75t_L g100 ( .A(n_92), .Y(n_100) );
INVx1_ASAP7_75t_L g103 ( .A(n_92), .Y(n_103) );
INVx2_ASAP7_75t_L g110 ( .A(n_95), .Y(n_110) );
AND2x2_ASAP7_75t_L g129 ( .A(n_95), .B(n_123), .Y(n_129) );
BUFx2_ASAP7_75t_L g132 ( .A(n_95), .Y(n_132) );
AND2x4_ASAP7_75t_L g119 ( .A(n_97), .B(n_109), .Y(n_119) );
AND2x4_ASAP7_75t_L g154 ( .A(n_97), .B(n_122), .Y(n_154) );
AND2x2_ASAP7_75t_L g160 ( .A(n_97), .B(n_129), .Y(n_160) );
AND2x4_ASAP7_75t_L g97 ( .A(n_98), .B(n_101), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_99), .Y(n_98) );
AND2x4_ASAP7_75t_L g108 ( .A(n_99), .B(n_101), .Y(n_108) );
AND2x2_ASAP7_75t_L g114 ( .A(n_99), .B(n_102), .Y(n_114) );
INVx1_ASAP7_75t_L g128 ( .A(n_99), .Y(n_128) );
INVxp67_ASAP7_75t_L g141 ( .A(n_101), .Y(n_141) );
INVx2_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
AND2x2_ASAP7_75t_L g127 ( .A(n_102), .B(n_128), .Y(n_127) );
BUFx3_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
AND2x2_ASAP7_75t_L g107 ( .A(n_108), .B(n_109), .Y(n_107) );
AND2x4_ASAP7_75t_L g121 ( .A(n_108), .B(n_122), .Y(n_121) );
AND2x4_ASAP7_75t_L g137 ( .A(n_108), .B(n_129), .Y(n_137) );
AND2x2_ASAP7_75t_L g149 ( .A(n_109), .B(n_127), .Y(n_149) );
AND2x4_ASAP7_75t_L g122 ( .A(n_110), .B(n_123), .Y(n_122) );
INVx2_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
INVx3_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
AND2x2_ASAP7_75t_L g113 ( .A(n_114), .B(n_115), .Y(n_113) );
AND2x4_ASAP7_75t_L g131 ( .A(n_114), .B(n_132), .Y(n_131) );
AND2x4_ASAP7_75t_L g157 ( .A(n_114), .B(n_122), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g116 ( .A(n_117), .B(n_124), .Y(n_116) );
BUFx3_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
BUFx3_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
AND2x4_ASAP7_75t_L g163 ( .A(n_122), .B(n_127), .Y(n_163) );
BUFx6f_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
AND2x2_ASAP7_75t_L g126 ( .A(n_127), .B(n_129), .Y(n_126) );
HB1xp67_ASAP7_75t_L g146 ( .A(n_128), .Y(n_146) );
BUFx2_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
NOR2xp33_ASAP7_75t_L g133 ( .A(n_134), .B(n_150), .Y(n_133) );
NAND2xp5_ASAP7_75t_L g134 ( .A(n_135), .B(n_142), .Y(n_134) );
BUFx3_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
INVx2_ASAP7_75t_SL g138 ( .A(n_139), .Y(n_138) );
INVx6_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
BUFx6f_ASAP7_75t_SL g143 ( .A(n_144), .Y(n_143) );
INVx1_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx2_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx3_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_151), .B(n_158), .Y(n_150) );
INVx2_ASAP7_75t_SL g152 ( .A(n_153), .Y(n_152) );
INVx8_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx2_ASAP7_75t_SL g155 ( .A(n_156), .Y(n_155) );
INVx2_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
BUFx2_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
INVx2_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
INVx8_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
AOI22xp5_ASAP7_75t_L g166 ( .A1(n_167), .A2(n_168), .B1(n_171), .B2(n_180), .Y(n_166) );
CKINVDCx20_ASAP7_75t_R g167 ( .A(n_168), .Y(n_167) );
CKINVDCx20_ASAP7_75t_R g180 ( .A(n_171), .Y(n_180) );
NOR2xp33_ASAP7_75t_L g242 ( .A(n_172), .B(n_243), .Y(n_242) );
CKINVDCx16_ASAP7_75t_R g179 ( .A(n_173), .Y(n_179) );
INVx1_ASAP7_75t_L g178 ( .A(n_175), .Y(n_178) );
CKINVDCx14_ASAP7_75t_R g181 ( .A(n_182), .Y(n_181) );
CKINVDCx20_ASAP7_75t_R g182 ( .A(n_183), .Y(n_182) );
AND3x1_ASAP7_75t_SL g183 ( .A(n_184), .B(n_190), .C(n_193), .Y(n_183) );
INVxp67_ASAP7_75t_L g521 ( .A(n_184), .Y(n_521) );
CKINVDCx8_ASAP7_75t_R g185 ( .A(n_186), .Y(n_185) );
NOR2xp33_ASAP7_75t_L g187 ( .A(n_188), .B(n_189), .Y(n_187) );
CKINVDCx16_ASAP7_75t_R g519 ( .A(n_190), .Y(n_519) );
AOI21xp33_ASAP7_75t_L g529 ( .A1(n_190), .A2(n_530), .B(n_531), .Y(n_529) );
INVx1_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
AND2x2_ASAP7_75t_L g245 ( .A(n_191), .B(n_246), .Y(n_245) );
OR2x2_ASAP7_75t_SL g527 ( .A(n_191), .B(n_193), .Y(n_527) );
HB1xp67_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
AND2x2_ASAP7_75t_L g211 ( .A(n_192), .B(n_212), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_193), .B(n_521), .Y(n_520) );
INVx1_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
NOR2x1p5_ASAP7_75t_L g249 ( .A(n_194), .B(n_250), .Y(n_249) );
INVx1_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
INVx1_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
OR2x6_ASAP7_75t_L g197 ( .A(n_198), .B(n_423), .Y(n_197) );
NAND3xp33_ASAP7_75t_SL g198 ( .A(n_199), .B(n_333), .C(n_373), .Y(n_198) );
O2A1O1Ixp33_ASAP7_75t_L g199 ( .A1(n_200), .A2(n_238), .B(n_262), .C(n_289), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_200), .B(n_338), .Y(n_372) );
NOR2x1p5_ASAP7_75t_L g200 ( .A(n_201), .B(n_227), .Y(n_200) );
BUFx3_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
INVx2_ASAP7_75t_L g308 ( .A(n_202), .Y(n_308) );
INVx2_ASAP7_75t_L g324 ( .A(n_202), .Y(n_324) );
OR2x2_ASAP7_75t_L g336 ( .A(n_202), .B(n_228), .Y(n_336) );
AND2x2_ASAP7_75t_L g350 ( .A(n_202), .B(n_309), .Y(n_350) );
INVx1_ASAP7_75t_L g378 ( .A(n_202), .Y(n_378) );
HB1xp67_ASAP7_75t_L g439 ( .A(n_202), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_202), .B(n_228), .Y(n_484) );
OA21x2_ASAP7_75t_L g202 ( .A1(n_203), .A2(n_207), .B(n_226), .Y(n_202) );
CKINVDCx5p33_ASAP7_75t_R g280 ( .A(n_203), .Y(n_280) );
BUFx6f_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
AND2x2_ASAP7_75t_SL g204 ( .A(n_205), .B(n_206), .Y(n_204) );
AND2x4_ASAP7_75t_L g243 ( .A(n_205), .B(n_206), .Y(n_243) );
AND2x6_ASAP7_75t_L g208 ( .A(n_209), .B(n_211), .Y(n_208) );
BUFx3_ASAP7_75t_L g247 ( .A(n_209), .Y(n_247) );
AND2x6_ASAP7_75t_L g224 ( .A(n_210), .B(n_215), .Y(n_224) );
INVx2_ASAP7_75t_L g251 ( .A(n_210), .Y(n_251) );
AND2x4_ASAP7_75t_L g248 ( .A(n_211), .B(n_249), .Y(n_248) );
AND2x4_ASAP7_75t_L g222 ( .A(n_212), .B(n_217), .Y(n_222) );
INVx2_ASAP7_75t_L g246 ( .A(n_212), .Y(n_246) );
AND2x4_ASAP7_75t_L g213 ( .A(n_214), .B(n_219), .Y(n_213) );
INVx1_ASAP7_75t_L g261 ( .A(n_214), .Y(n_261) );
AND2x4_ASAP7_75t_L g214 ( .A(n_215), .B(n_217), .Y(n_214) );
INVx2_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
INVx2_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
INVx5_ASAP7_75t_L g225 ( .A(n_219), .Y(n_225) );
AOI21xp5_ASAP7_75t_L g220 ( .A1(n_221), .A2(n_223), .B(n_225), .Y(n_220) );
AOI21xp5_ASAP7_75t_L g232 ( .A1(n_225), .A2(n_233), .B(n_234), .Y(n_232) );
AOI21xp5_ASAP7_75t_L g269 ( .A1(n_225), .A2(n_270), .B(n_271), .Y(n_269) );
AOI21xp5_ASAP7_75t_L g276 ( .A1(n_225), .A2(n_277), .B(n_278), .Y(n_276) );
AOI21xp5_ASAP7_75t_L g299 ( .A1(n_225), .A2(n_300), .B(n_301), .Y(n_299) );
AOI21xp5_ASAP7_75t_L g313 ( .A1(n_225), .A2(n_314), .B(n_315), .Y(n_313) );
OR2x2_ASAP7_75t_L g305 ( .A(n_227), .B(n_306), .Y(n_305) );
HB1xp67_ASAP7_75t_L g440 ( .A(n_227), .Y(n_440) );
AND2x2_ASAP7_75t_L g445 ( .A(n_227), .B(n_307), .Y(n_445) );
INVx2_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
AND2x4_ASAP7_75t_L g238 ( .A(n_228), .B(n_239), .Y(n_238) );
OR2x2_ASAP7_75t_L g304 ( .A(n_228), .B(n_240), .Y(n_304) );
OR2x2_ASAP7_75t_L g323 ( .A(n_228), .B(n_324), .Y(n_323) );
INVx2_ASAP7_75t_L g352 ( .A(n_228), .Y(n_352) );
AND2x4_ASAP7_75t_SL g391 ( .A(n_228), .B(n_240), .Y(n_391) );
HB1xp67_ASAP7_75t_L g395 ( .A(n_228), .Y(n_395) );
OR2x2_ASAP7_75t_L g412 ( .A(n_228), .B(n_413), .Y(n_412) );
AND2x2_ASAP7_75t_L g422 ( .A(n_228), .B(n_329), .Y(n_422) );
INVx1_ASAP7_75t_L g451 ( .A(n_228), .Y(n_451) );
OR2x6_ASAP7_75t_L g228 ( .A(n_229), .B(n_237), .Y(n_228) );
AOI21xp5_ASAP7_75t_L g229 ( .A1(n_230), .A2(n_231), .B(n_235), .Y(n_229) );
INVx2_ASAP7_75t_SL g284 ( .A(n_235), .Y(n_284) );
BUFx4f_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
INVx3_ASAP7_75t_L g258 ( .A(n_236), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_238), .B(n_380), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_239), .B(n_309), .Y(n_326) );
AND2x2_ASAP7_75t_L g338 ( .A(n_239), .B(n_339), .Y(n_338) );
OR2x2_ASAP7_75t_L g356 ( .A(n_239), .B(n_323), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_239), .B(n_377), .Y(n_376) );
INVx3_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
AND2x4_ASAP7_75t_L g329 ( .A(n_240), .B(n_330), .Y(n_329) );
AND2x2_ASAP7_75t_L g351 ( .A(n_240), .B(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g386 ( .A(n_240), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_240), .B(n_309), .Y(n_410) );
AND2x4_ASAP7_75t_L g240 ( .A(n_241), .B(n_254), .Y(n_240) );
AOI22xp5_ASAP7_75t_L g241 ( .A1(n_242), .A2(n_244), .B1(n_248), .B2(n_252), .Y(n_241) );
NOR2xp33_ASAP7_75t_L g252 ( .A(n_243), .B(n_253), .Y(n_252) );
NOR2xp33_ASAP7_75t_L g255 ( .A(n_243), .B(n_256), .Y(n_255) );
NOR3xp33_ASAP7_75t_L g259 ( .A(n_243), .B(n_260), .C(n_261), .Y(n_259) );
AOI21xp5_ASAP7_75t_L g266 ( .A1(n_243), .A2(n_267), .B(n_268), .Y(n_266) );
INVx1_ASAP7_75t_L g512 ( .A(n_244), .Y(n_512) );
AND2x4_ASAP7_75t_L g244 ( .A(n_245), .B(n_247), .Y(n_244) );
HB1xp67_ASAP7_75t_L g530 ( .A(n_246), .Y(n_530) );
INVx1_ASAP7_75t_L g532 ( .A(n_247), .Y(n_532) );
INVx3_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
INVx4_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
AOI21x1_ASAP7_75t_L g310 ( .A1(n_258), .A2(n_311), .B(n_317), .Y(n_310) );
AND2x2_ASAP7_75t_L g262 ( .A(n_263), .B(n_272), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_263), .B(n_342), .Y(n_341) );
AND2x4_ASAP7_75t_L g359 ( .A(n_263), .B(n_360), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_263), .B(n_273), .Y(n_364) );
NAND3xp33_ASAP7_75t_L g379 ( .A(n_263), .B(n_380), .C(n_381), .Y(n_379) );
AND2x2_ASAP7_75t_L g427 ( .A(n_263), .B(n_332), .Y(n_427) );
INVx5_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
AND2x2_ASAP7_75t_L g294 ( .A(n_264), .B(n_295), .Y(n_294) );
AND2x4_ASAP7_75t_SL g331 ( .A(n_264), .B(n_332), .Y(n_331) );
INVx2_ASAP7_75t_L g347 ( .A(n_264), .Y(n_347) );
OR2x2_ASAP7_75t_L g370 ( .A(n_264), .B(n_360), .Y(n_370) );
HB1xp67_ASAP7_75t_L g387 ( .A(n_264), .Y(n_387) );
AND2x2_ASAP7_75t_SL g405 ( .A(n_264), .B(n_293), .Y(n_405) );
AND2x4_ASAP7_75t_L g420 ( .A(n_264), .B(n_296), .Y(n_420) );
AND2x2_ASAP7_75t_L g434 ( .A(n_264), .B(n_273), .Y(n_434) );
OR2x2_ASAP7_75t_L g455 ( .A(n_264), .B(n_282), .Y(n_455) );
OR2x6_ASAP7_75t_L g264 ( .A(n_265), .B(n_266), .Y(n_264) );
AND2x2_ASAP7_75t_L g509 ( .A(n_272), .B(n_387), .Y(n_509) );
AND2x2_ASAP7_75t_L g272 ( .A(n_273), .B(n_282), .Y(n_272) );
AND2x4_ASAP7_75t_L g332 ( .A(n_273), .B(n_295), .Y(n_332) );
INVx2_ASAP7_75t_L g343 ( .A(n_273), .Y(n_343) );
AND2x2_ASAP7_75t_L g348 ( .A(n_273), .B(n_293), .Y(n_348) );
HB1xp67_ASAP7_75t_L g381 ( .A(n_273), .Y(n_381) );
OR2x2_ASAP7_75t_L g404 ( .A(n_273), .B(n_296), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_273), .B(n_296), .Y(n_407) );
INVx1_ASAP7_75t_L g416 ( .A(n_273), .Y(n_416) );
AO21x2_ASAP7_75t_L g273 ( .A1(n_274), .A2(n_280), .B(n_281), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_275), .B(n_279), .Y(n_274) );
AO21x2_ASAP7_75t_L g296 ( .A1(n_280), .A2(n_297), .B(n_303), .Y(n_296) );
AO21x2_ASAP7_75t_L g360 ( .A1(n_280), .A2(n_297), .B(n_303), .Y(n_360) );
AND2x2_ASAP7_75t_L g319 ( .A(n_282), .B(n_296), .Y(n_319) );
BUFx2_ASAP7_75t_L g368 ( .A(n_282), .Y(n_368) );
AND2x2_ASAP7_75t_L g463 ( .A(n_282), .B(n_343), .Y(n_463) );
INVx2_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
BUFx6f_ASAP7_75t_L g293 ( .A(n_283), .Y(n_293) );
AOI21x1_ASAP7_75t_L g283 ( .A1(n_284), .A2(n_285), .B(n_288), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_286), .B(n_287), .Y(n_285) );
OAI221xp5_ASAP7_75t_L g289 ( .A1(n_290), .A2(n_304), .B1(n_305), .B2(n_318), .C(n_320), .Y(n_289) );
INVx1_ASAP7_75t_SL g290 ( .A(n_291), .Y(n_290) );
AND2x2_ASAP7_75t_L g291 ( .A(n_292), .B(n_294), .Y(n_291) );
NOR2x1_ASAP7_75t_L g365 ( .A(n_292), .B(n_366), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_292), .B(n_359), .Y(n_399) );
OR2x2_ASAP7_75t_L g411 ( .A(n_292), .B(n_407), .Y(n_411) );
OR2x2_ASAP7_75t_L g414 ( .A(n_292), .B(n_415), .Y(n_414) );
OR2x2_ASAP7_75t_L g503 ( .A(n_292), .B(n_504), .Y(n_503) );
INVx2_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
AND2x4_ASAP7_75t_L g342 ( .A(n_293), .B(n_343), .Y(n_342) );
OA33x2_ASAP7_75t_L g375 ( .A1(n_293), .A2(n_336), .A3(n_376), .B1(n_379), .B2(n_382), .B3(n_385), .Y(n_375) );
OR2x2_ASAP7_75t_L g406 ( .A(n_293), .B(n_407), .Y(n_406) );
OR2x2_ASAP7_75t_L g430 ( .A(n_293), .B(n_431), .Y(n_430) );
OR2x2_ASAP7_75t_L g438 ( .A(n_293), .B(n_439), .Y(n_438) );
AND2x2_ASAP7_75t_L g458 ( .A(n_293), .B(n_332), .Y(n_458) );
NOR2xp33_ASAP7_75t_L g496 ( .A(n_293), .B(n_347), .Y(n_496) );
INVx2_ASAP7_75t_L g366 ( .A(n_294), .Y(n_366) );
AOI322xp5_ASAP7_75t_L g436 ( .A1(n_294), .A2(n_349), .A3(n_437), .B1(n_440), .B2(n_441), .C1(n_443), .C2(n_445), .Y(n_436) );
INVx2_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
HB1xp67_ASAP7_75t_L g465 ( .A(n_296), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_298), .B(n_302), .Y(n_297) );
OR2x2_ASAP7_75t_L g418 ( .A(n_304), .B(n_397), .Y(n_418) );
NOR2xp33_ASAP7_75t_L g470 ( .A(n_304), .B(n_471), .Y(n_470) );
INVx1_ASAP7_75t_SL g491 ( .A(n_304), .Y(n_491) );
INVx1_ASAP7_75t_SL g357 ( .A(n_305), .Y(n_357) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
AND2x2_ASAP7_75t_L g390 ( .A(n_307), .B(n_391), .Y(n_390) );
AND2x2_ASAP7_75t_L g307 ( .A(n_308), .B(n_309), .Y(n_307) );
INVx2_ASAP7_75t_L g330 ( .A(n_309), .Y(n_330) );
INVx1_ASAP7_75t_L g339 ( .A(n_309), .Y(n_339) );
INVx1_ASAP7_75t_L g380 ( .A(n_309), .Y(n_380) );
OR2x2_ASAP7_75t_L g397 ( .A(n_309), .B(n_324), .Y(n_397) );
HB1xp67_ASAP7_75t_L g472 ( .A(n_309), .Y(n_472) );
INVx3_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_312), .B(n_316), .Y(n_311) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
AND2x2_ASAP7_75t_SL g441 ( .A(n_319), .B(n_442), .Y(n_441) );
OAI21xp5_ASAP7_75t_SL g320 ( .A1(n_321), .A2(n_327), .B(n_331), .Y(n_320) );
A2O1A1Ixp33_ASAP7_75t_L g394 ( .A1(n_321), .A2(n_395), .B(n_396), .C(n_398), .Y(n_394) );
AND2x4_ASAP7_75t_L g321 ( .A(n_322), .B(n_325), .Y(n_321) );
INVx2_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
OR2x2_ASAP7_75t_L g459 ( .A(n_323), .B(n_460), .Y(n_459) );
HB1xp67_ASAP7_75t_L g328 ( .A(n_324), .Y(n_328) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
OR2x2_ASAP7_75t_L g483 ( .A(n_326), .B(n_484), .Y(n_483) );
AND2x2_ASAP7_75t_L g327 ( .A(n_328), .B(n_329), .Y(n_327) );
AND2x2_ASAP7_75t_SL g452 ( .A(n_329), .B(n_453), .Y(n_452) );
INVx1_ASAP7_75t_L g460 ( .A(n_329), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_329), .B(n_451), .Y(n_468) );
INVx3_ASAP7_75t_SL g393 ( .A(n_332), .Y(n_393) );
AOI221xp5_ASAP7_75t_L g333 ( .A1(n_334), .A2(n_340), .B1(n_344), .B2(n_349), .C(n_353), .Y(n_333) );
INVx1_ASAP7_75t_SL g334 ( .A(n_335), .Y(n_334) );
OR2x2_ASAP7_75t_L g335 ( .A(n_336), .B(n_337), .Y(n_335) );
INVx1_ASAP7_75t_SL g337 ( .A(n_338), .Y(n_337) );
HB1xp67_ASAP7_75t_L g384 ( .A(n_339), .Y(n_384) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
AOI21xp5_ASAP7_75t_L g447 ( .A1(n_342), .A2(n_369), .B(n_441), .Y(n_447) );
AND2x2_ASAP7_75t_L g473 ( .A(n_342), .B(n_420), .Y(n_473) );
HB1xp67_ASAP7_75t_L g361 ( .A(n_343), .Y(n_361) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_346), .B(n_348), .Y(n_345) );
INVx2_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_347), .B(n_463), .Y(n_462) );
OR2x2_ASAP7_75t_L g482 ( .A(n_347), .B(n_404), .Y(n_482) );
AND2x2_ASAP7_75t_L g349 ( .A(n_350), .B(n_351), .Y(n_349) );
INVx2_ASAP7_75t_L g431 ( .A(n_350), .Y(n_431) );
OAI21xp33_ASAP7_75t_L g353 ( .A1(n_354), .A2(n_358), .B(n_362), .Y(n_353) );
NOR2xp33_ASAP7_75t_L g354 ( .A(n_355), .B(n_357), .Y(n_354) );
INVx1_ASAP7_75t_SL g355 ( .A(n_356), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_359), .B(n_361), .Y(n_358) );
INVx2_ASAP7_75t_L g504 ( .A(n_359), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_360), .B(n_416), .Y(n_415) );
AND2x2_ASAP7_75t_L g433 ( .A(n_360), .B(n_434), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_361), .B(n_383), .Y(n_382) );
OAI31xp33_ASAP7_75t_SL g362 ( .A1(n_363), .A2(n_365), .A3(n_367), .B(n_371), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_366), .B(n_393), .Y(n_392) );
AND2x2_ASAP7_75t_L g367 ( .A(n_368), .B(n_369), .Y(n_367) );
OR2x2_ASAP7_75t_L g444 ( .A(n_368), .B(n_370), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_368), .B(n_420), .Y(n_499) );
INVx1_ASAP7_75t_SL g369 ( .A(n_370), .Y(n_369) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
NOR5xp2_ASAP7_75t_L g373 ( .A(n_374), .B(n_388), .C(n_400), .D(n_409), .E(n_417), .Y(n_373) );
INVxp67_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
HB1xp67_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_378), .B(n_380), .Y(n_413) );
INVx1_ASAP7_75t_L g453 ( .A(n_378), .Y(n_453) );
INVxp67_ASAP7_75t_SL g490 ( .A(n_378), .Y(n_490) );
INVx1_ASAP7_75t_L g442 ( .A(n_381), .Y(n_442) );
INVxp67_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
NAND2xp33_ASAP7_75t_SL g385 ( .A(n_386), .B(n_387), .Y(n_385) );
OAI321xp33_ASAP7_75t_L g425 ( .A1(n_386), .A2(n_426), .A3(n_428), .B1(n_432), .B2(n_435), .C(n_436), .Y(n_425) );
INVx1_ASAP7_75t_L g479 ( .A(n_387), .Y(n_479) );
OAI21xp33_ASAP7_75t_L g388 ( .A1(n_389), .A2(n_392), .B(n_394), .Y(n_388) );
INVx1_ASAP7_75t_SL g389 ( .A(n_390), .Y(n_389) );
AOI22xp33_ASAP7_75t_L g469 ( .A1(n_390), .A2(n_463), .B1(n_470), .B2(n_473), .Y(n_469) );
AND2x2_ASAP7_75t_L g498 ( .A(n_391), .B(n_472), .Y(n_498) );
INVx1_ASAP7_75t_L g408 ( .A(n_396), .Y(n_408) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
AOI21xp5_ASAP7_75t_L g400 ( .A1(n_401), .A2(n_406), .B(n_408), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
AND2x2_ASAP7_75t_L g402 ( .A(n_403), .B(n_405), .Y(n_402) );
INVx2_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
OAI22xp5_ASAP7_75t_L g417 ( .A1(n_407), .A2(n_418), .B1(n_419), .B2(n_421), .Y(n_417) );
INVx1_ASAP7_75t_L g480 ( .A(n_407), .Y(n_480) );
OAI22xp5_ASAP7_75t_L g409 ( .A1(n_410), .A2(n_411), .B1(n_412), .B2(n_414), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_416), .B(n_420), .Y(n_419) );
OAI221xp5_ASAP7_75t_L g494 ( .A1(n_418), .A2(n_495), .B1(n_497), .B2(n_499), .C(n_500), .Y(n_494) );
INVx1_ASAP7_75t_L g501 ( .A(n_418), .Y(n_501) );
OAI221xp5_ASAP7_75t_L g475 ( .A1(n_419), .A2(n_476), .B1(n_483), .B2(n_485), .C(n_486), .Y(n_475) );
OAI21xp5_ASAP7_75t_L g446 ( .A1(n_421), .A2(n_447), .B(n_448), .Y(n_446) );
INVx2_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_424), .B(n_474), .Y(n_423) );
NOR3xp33_ASAP7_75t_L g424 ( .A(n_425), .B(n_446), .C(n_464), .Y(n_424) );
INVx2_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
HB1xp67_ASAP7_75t_L g493 ( .A(n_427), .Y(n_493) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx3_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g492 ( .A(n_435), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_437), .B(n_467), .Y(n_466) );
INVx1_ASAP7_75t_SL g437 ( .A(n_438), .Y(n_437) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx1_ASAP7_75t_L g485 ( .A(n_445), .Y(n_485) );
AOI21xp5_ASAP7_75t_L g448 ( .A1(n_449), .A2(n_454), .B(n_456), .Y(n_448) );
INVxp67_ASAP7_75t_L g506 ( .A(n_449), .Y(n_506) );
AND2x2_ASAP7_75t_L g449 ( .A(n_450), .B(n_452), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx2_ASAP7_75t_SL g461 ( .A(n_452), .Y(n_461) );
INVx1_ASAP7_75t_SL g454 ( .A(n_455), .Y(n_454) );
OAI22xp33_ASAP7_75t_L g456 ( .A1(n_457), .A2(n_459), .B1(n_461), .B2(n_462), .Y(n_456) );
INVx2_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
OAI21xp33_ASAP7_75t_L g464 ( .A1(n_465), .A2(n_466), .B(n_469), .Y(n_464) );
INVx1_ASAP7_75t_SL g467 ( .A(n_468), .Y(n_467) );
INVx1_ASAP7_75t_L g507 ( .A(n_470), .Y(n_507) );
INVx1_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
NOR3xp33_ASAP7_75t_L g474 ( .A(n_475), .B(n_494), .C(n_505), .Y(n_474) );
NOR2xp33_ASAP7_75t_L g476 ( .A(n_477), .B(n_481), .Y(n_476) );
INVx2_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
NAND2xp5_ASAP7_75t_SL g478 ( .A(n_479), .B(n_480), .Y(n_478) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
OAI21xp5_ASAP7_75t_SL g486 ( .A1(n_487), .A2(n_492), .B(n_493), .Y(n_486) );
INVx1_ASAP7_75t_SL g487 ( .A(n_488), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_489), .B(n_491), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
INVx1_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
INVxp67_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
OAI21xp5_ASAP7_75t_L g500 ( .A1(n_498), .A2(n_501), .B(n_502), .Y(n_500) );
INVx1_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
AOI21xp33_ASAP7_75t_L g505 ( .A1(n_506), .A2(n_507), .B(n_508), .Y(n_505) );
INVx1_ASAP7_75t_SL g508 ( .A(n_509), .Y(n_508) );
CKINVDCx20_ASAP7_75t_R g510 ( .A(n_511), .Y(n_510) );
HB1xp67_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
OAI222xp33_ASAP7_75t_L g513 ( .A1(n_514), .A2(n_515), .B1(n_516), .B2(n_522), .C1(n_525), .C2(n_528), .Y(n_513) );
CKINVDCx20_ASAP7_75t_R g516 ( .A(n_517), .Y(n_516) );
CKINVDCx20_ASAP7_75t_R g517 ( .A(n_518), .Y(n_517) );
OR2x2_ASAP7_75t_L g518 ( .A(n_519), .B(n_520), .Y(n_518) );
CKINVDCx20_ASAP7_75t_R g522 ( .A(n_523), .Y(n_522) );
CKINVDCx20_ASAP7_75t_R g525 ( .A(n_526), .Y(n_525) );
INVx2_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
INVx1_ASAP7_75t_SL g528 ( .A(n_529), .Y(n_528) );
INVxp67_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
endmodule