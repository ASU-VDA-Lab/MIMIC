module fake_jpeg_10247_n_109 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_109);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_109;

wire n_10;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_106;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx12f_ASAP7_75t_L g10 ( 
.A(n_3),
.Y(n_10)
);

BUFx3_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_7),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_1),
.Y(n_13)
);

BUFx16f_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_7),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx1_ASAP7_75t_SL g20 ( 
.A(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_21),
.B(n_22),
.Y(n_28)
);

OR2x2_ASAP7_75t_L g22 ( 
.A(n_13),
.B(n_0),
.Y(n_22)
);

AND2x2_ASAP7_75t_L g23 ( 
.A(n_14),
.B(n_0),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g34 ( 
.A(n_23),
.B(n_20),
.C(n_19),
.Y(n_34)
);

OR2x2_ASAP7_75t_L g24 ( 
.A(n_13),
.B(n_1),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_24),
.B(n_26),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_25),
.Y(n_30)
);

INVx13_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_27),
.A2(n_20),
.B1(n_18),
.B2(n_19),
.Y(n_33)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_29),
.B(n_32),
.Y(n_39)
);

AO22x1_ASAP7_75t_SL g31 ( 
.A1(n_23),
.A2(n_14),
.B1(n_17),
.B2(n_18),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_31),
.A2(n_20),
.B1(n_23),
.B2(n_26),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_33),
.A2(n_31),
.B1(n_27),
.B2(n_16),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_34),
.B(n_22),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_36),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_37),
.B(n_40),
.Y(n_48)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_28),
.B(n_22),
.Y(n_41)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_42),
.B(n_24),
.Y(n_54)
);

OAI22xp33_ASAP7_75t_L g43 ( 
.A1(n_31),
.A2(n_27),
.B1(n_23),
.B2(n_18),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_43),
.A2(n_45),
.B1(n_21),
.B2(n_30),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_24),
.Y(n_44)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_29),
.B(n_22),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_46),
.B(n_47),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_35),
.B(n_34),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_45),
.A2(n_31),
.B1(n_30),
.B2(n_21),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_49),
.A2(n_51),
.B1(n_37),
.B2(n_42),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g50 ( 
.A(n_39),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_50),
.B(n_57),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_54),
.B(n_56),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_38),
.B(n_10),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_L g58 ( 
.A1(n_44),
.A2(n_24),
.B(n_36),
.Y(n_58)
);

AOI21xp5_ASAP7_75t_L g67 ( 
.A1(n_58),
.A2(n_16),
.B(n_15),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_59),
.A2(n_69),
.B1(n_55),
.B2(n_53),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_60),
.B(n_65),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_55),
.A2(n_40),
.B1(n_37),
.B2(n_47),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_61),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_52),
.B(n_46),
.C(n_41),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_62),
.B(n_66),
.C(n_12),
.Y(n_76)
);

NOR2x1_ASAP7_75t_L g64 ( 
.A(n_58),
.B(n_32),
.Y(n_64)
);

NAND3xp33_ASAP7_75t_L g75 ( 
.A(n_64),
.B(n_53),
.C(n_2),
.Y(n_75)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_57),
.B(n_38),
.C(n_32),
.Y(n_66)
);

XNOR2xp5_ASAP7_75t_L g70 ( 
.A(n_67),
.B(n_48),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_51),
.A2(n_30),
.B1(n_15),
.B2(n_12),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_70),
.B(n_71),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_68),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_63),
.Y(n_72)
);

AO221x1_ASAP7_75t_L g85 ( 
.A1(n_72),
.A2(n_11),
.B1(n_10),
.B2(n_32),
.C(n_4),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_73),
.A2(n_60),
.B1(n_69),
.B2(n_59),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_65),
.B(n_50),
.Y(n_74)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_74),
.Y(n_80)
);

OAI322xp33_ASAP7_75t_L g87 ( 
.A1(n_75),
.A2(n_77),
.A3(n_9),
.B1(n_2),
.B2(n_3),
.C1(n_4),
.C2(n_5),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_76),
.B(n_67),
.C(n_62),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_61),
.B(n_17),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_81),
.A2(n_84),
.B1(n_78),
.B2(n_11),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g90 ( 
.A1(n_82),
.A2(n_78),
.B(n_73),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_79),
.A2(n_64),
.B1(n_66),
.B2(n_17),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_85),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_76),
.B(n_32),
.C(n_25),
.Y(n_86)
);

XOR2xp5_ASAP7_75t_L g89 ( 
.A(n_86),
.B(n_77),
.Y(n_89)
);

NAND3xp33_ASAP7_75t_L g93 ( 
.A(n_87),
.B(n_9),
.C(n_3),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g88 ( 
.A(n_82),
.B(n_70),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_88),
.B(n_89),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_90),
.A2(n_83),
.B(n_80),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_80),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_91),
.B(n_94),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_93),
.A2(n_8),
.B1(n_5),
.B2(n_6),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_97),
.B(n_98),
.Y(n_102)
);

AOI322xp5_ASAP7_75t_L g98 ( 
.A1(n_91),
.A2(n_84),
.A3(n_86),
.B1(n_11),
.B2(n_17),
.C1(n_25),
.C2(n_10),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_99),
.B(n_93),
.Y(n_100)
);

A2O1A1Ixp33_ASAP7_75t_L g104 ( 
.A1(n_100),
.A2(n_103),
.B(n_96),
.C(n_10),
.Y(n_104)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_95),
.Y(n_101)
);

AOI322xp5_ASAP7_75t_L g105 ( 
.A1(n_101),
.A2(n_1),
.A3(n_6),
.B1(n_7),
.B2(n_9),
.C1(n_25),
.C2(n_102),
.Y(n_105)
);

OR2x2_ASAP7_75t_L g103 ( 
.A(n_98),
.B(n_92),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_104),
.B(n_105),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_103),
.B(n_6),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_106),
.B(n_101),
.C(n_1),
.Y(n_107)
);

OR2x2_ASAP7_75t_L g109 ( 
.A(n_107),
.B(n_108),
.Y(n_109)
);


endmodule