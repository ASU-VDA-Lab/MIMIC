module fake_jpeg_26219_n_253 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_253);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_253;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_15),
.Y(n_17)
);

BUFx2_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx10_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_35),
.B(n_38),
.Y(n_45)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_31),
.B(n_0),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_31),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

BUFx24_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_43),
.B(n_27),
.Y(n_48)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_36),
.A2(n_28),
.B1(n_26),
.B2(n_42),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_46),
.A2(n_63),
.B1(n_44),
.B2(n_38),
.Y(n_77)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_39),
.B(n_30),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_50),
.B(n_52),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_30),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_53),
.B(n_62),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_38),
.B(n_33),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_55),
.B(n_56),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_36),
.A2(n_26),
.B1(n_31),
.B2(n_18),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_57),
.A2(n_59),
.B1(n_27),
.B2(n_21),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_41),
.B(n_25),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_58),
.B(n_65),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_36),
.A2(n_20),
.B1(n_21),
.B2(n_19),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_40),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_60),
.B(n_40),
.Y(n_69)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_44),
.A2(n_25),
.B1(n_33),
.B2(n_32),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_41),
.B(n_17),
.Y(n_65)
);

OAI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_64),
.A2(n_43),
.B1(n_37),
.B2(n_35),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_66),
.A2(n_74),
.B1(n_64),
.B2(n_59),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_68),
.B(n_73),
.Y(n_120)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_69),
.Y(n_114)
);

BUFx10_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_71),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_56),
.A2(n_43),
.B1(n_37),
.B2(n_35),
.Y(n_74)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_75),
.Y(n_101)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_61),
.Y(n_76)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_76),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_SL g107 ( 
.A(n_77),
.B(n_87),
.C(n_88),
.Y(n_107)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_78),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_56),
.B(n_50),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_81),
.B(n_92),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_60),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_82),
.B(n_89),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_48),
.B(n_44),
.C(n_40),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_83),
.B(n_62),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_54),
.A2(n_35),
.B1(n_17),
.B2(n_22),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_84),
.Y(n_103)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_55),
.Y(n_85)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_85),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_63),
.A2(n_32),
.B1(n_22),
.B2(n_23),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_86),
.A2(n_90),
.B(n_85),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_54),
.A2(n_23),
.B1(n_34),
.B2(n_31),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_64),
.A2(n_34),
.B1(n_24),
.B2(n_27),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_47),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_65),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_90),
.B(n_96),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_91),
.B(n_96),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_52),
.B(n_27),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_58),
.B(n_29),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_93),
.B(n_95),
.Y(n_115)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_51),
.Y(n_94)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_94),
.Y(n_121)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_57),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_57),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_98),
.A2(n_118),
.B1(n_93),
.B2(n_71),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_100),
.B(n_116),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_70),
.B(n_47),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_102),
.A2(n_105),
.B(n_110),
.Y(n_137)
);

OR2x2_ASAP7_75t_L g104 ( 
.A(n_72),
.B(n_41),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_104),
.A2(n_106),
.B(n_109),
.Y(n_148)
);

A2O1A1Ixp33_ASAP7_75t_L g106 ( 
.A1(n_81),
.A2(n_46),
.B(n_49),
.C(n_53),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_68),
.A2(n_73),
.B(n_67),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_95),
.A2(n_49),
.B(n_61),
.Y(n_110)
);

INVx1_ASAP7_75t_SL g111 ( 
.A(n_86),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_111),
.B(n_82),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_67),
.A2(n_61),
.B(n_1),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_113),
.A2(n_0),
.B(n_2),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_70),
.B(n_47),
.Y(n_116)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_119),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_123),
.B(n_124),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_110),
.Y(n_124)
);

OR2x2_ASAP7_75t_L g150 ( 
.A(n_125),
.B(n_104),
.Y(n_150)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_108),
.Y(n_126)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_126),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_111),
.A2(n_91),
.B1(n_83),
.B2(n_79),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_127),
.A2(n_129),
.B1(n_140),
.B2(n_121),
.Y(n_163)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_99),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_128),
.B(n_131),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_122),
.A2(n_79),
.B1(n_92),
.B2(n_94),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_114),
.B(n_80),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_130),
.B(n_132),
.Y(n_159)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_99),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_113),
.B(n_80),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_L g133 ( 
.A1(n_107),
.A2(n_78),
.B1(n_89),
.B2(n_75),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_133),
.A2(n_139),
.B1(n_103),
.B2(n_115),
.Y(n_160)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_106),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_134),
.B(n_135),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_97),
.B(n_72),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_107),
.A2(n_78),
.B1(n_76),
.B2(n_71),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_138),
.A2(n_101),
.B1(n_112),
.B2(n_19),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_98),
.A2(n_71),
.B1(n_41),
.B2(n_21),
.Y(n_140)
);

O2A1O1Ixp33_ASAP7_75t_L g141 ( 
.A1(n_103),
.A2(n_24),
.B(n_41),
.C(n_21),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_141),
.B(n_145),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_120),
.Y(n_142)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_142),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_117),
.B(n_20),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_143),
.B(n_146),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_L g165 ( 
.A1(n_144),
.A2(n_112),
.B1(n_101),
.B2(n_108),
.Y(n_165)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_98),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_117),
.B(n_20),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_115),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_147),
.B(n_149),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_97),
.B(n_20),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_150),
.A2(n_160),
.B(n_165),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_126),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_156),
.B(n_174),
.Y(n_189)
);

AOI322xp5_ASAP7_75t_L g161 ( 
.A1(n_148),
.A2(n_105),
.A3(n_109),
.B1(n_102),
.B2(n_100),
.C1(n_116),
.C2(n_118),
.Y(n_161)
);

AO21x1_ASAP7_75t_L g176 ( 
.A1(n_161),
.A2(n_170),
.B(n_134),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_136),
.B(n_102),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_SL g183 ( 
.A(n_162),
.B(n_169),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_163),
.B(n_164),
.Y(n_187)
);

NOR2x1_ASAP7_75t_L g164 ( 
.A(n_139),
.B(n_121),
.Y(n_164)
);

OR2x2_ASAP7_75t_L g166 ( 
.A(n_129),
.B(n_24),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_166),
.A2(n_172),
.B(n_0),
.Y(n_186)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_149),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_168),
.B(n_173),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_SL g169 ( 
.A(n_148),
.B(n_29),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_124),
.A2(n_19),
.B1(n_29),
.B2(n_4),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_171),
.A2(n_141),
.B1(n_142),
.B2(n_123),
.Y(n_177)
);

OR2x2_ASAP7_75t_L g172 ( 
.A(n_140),
.B(n_29),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_137),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_137),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_162),
.B(n_136),
.C(n_147),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_175),
.B(n_181),
.C(n_188),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_176),
.B(n_184),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_177),
.A2(n_186),
.B1(n_193),
.B2(n_153),
.Y(n_201)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_152),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_178),
.A2(n_179),
.B(n_192),
.Y(n_205)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_152),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_173),
.B(n_174),
.C(n_163),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_164),
.A2(n_145),
.B1(n_127),
.B2(n_135),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_182),
.A2(n_185),
.B1(n_166),
.B2(n_157),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_168),
.A2(n_144),
.B1(n_131),
.B2(n_128),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_153),
.B(n_3),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_151),
.B(n_16),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_190),
.Y(n_196)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_151),
.Y(n_191)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_191),
.Y(n_198)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_167),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_160),
.A2(n_14),
.B1(n_15),
.B2(n_5),
.Y(n_193)
);

OA21x2_ASAP7_75t_L g194 ( 
.A1(n_155),
.A2(n_3),
.B(n_4),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_194),
.A2(n_150),
.B(n_6),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_189),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_197),
.B(n_200),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_199),
.B(n_202),
.Y(n_215)
);

INVx13_ASAP7_75t_L g200 ( 
.A(n_180),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_201),
.A2(n_203),
.B1(n_206),
.B2(n_208),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_185),
.A2(n_169),
.B1(n_171),
.B2(n_157),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_193),
.A2(n_158),
.B1(n_159),
.B2(n_155),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_204),
.B(n_207),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_187),
.A2(n_167),
.B1(n_156),
.B2(n_172),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_182),
.A2(n_154),
.B1(n_6),
.B2(n_7),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_177),
.A2(n_154),
.B1(n_6),
.B2(n_8),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_209),
.A2(n_3),
.B1(n_9),
.B2(n_10),
.Y(n_220)
);

BUFx24_ASAP7_75t_SL g210 ( 
.A(n_188),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_210),
.A2(n_175),
.B(n_186),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_211),
.B(n_216),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_195),
.B(n_181),
.C(n_178),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_212),
.B(n_217),
.C(n_221),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_195),
.B(n_176),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_205),
.B(n_179),
.C(n_180),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_197),
.A2(n_184),
.B(n_194),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_218),
.B(n_208),
.C(n_204),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_205),
.A2(n_192),
.B(n_194),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_219),
.A2(n_207),
.B(n_198),
.Y(n_228)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_220),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_199),
.B(n_183),
.C(n_10),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_214),
.B(n_196),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_223),
.B(n_224),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_219),
.B(n_200),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_225),
.B(n_216),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_222),
.A2(n_198),
.B1(n_202),
.B2(n_206),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_226),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_228),
.A2(n_213),
.B(n_215),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_212),
.B(n_183),
.C(n_10),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_230),
.B(n_13),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_217),
.B(n_9),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_231),
.B(n_9),
.Y(n_236)
);

NAND3xp33_ASAP7_75t_SL g242 ( 
.A(n_234),
.B(n_232),
.C(n_227),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_235),
.B(n_239),
.Y(n_243)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_236),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_224),
.A2(n_221),
.B(n_215),
.Y(n_238)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_238),
.Y(n_244)
);

AND2x4_ASAP7_75t_SL g240 ( 
.A(n_237),
.B(n_232),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_240),
.B(n_242),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_244),
.A2(n_233),
.B(n_236),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_245),
.B(n_246),
.C(n_12),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_243),
.B(n_229),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_241),
.B(n_11),
.Y(n_248)
);

OR2x2_ASAP7_75t_L g249 ( 
.A(n_248),
.B(n_12),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_249),
.A2(n_250),
.B(n_247),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_251),
.B(n_246),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_252),
.B(n_12),
.Y(n_253)
);


endmodule