module fake_jpeg_11266_n_551 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_551);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_551;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_17),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_2),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

INVx2_ASAP7_75t_SL g38 ( 
.A(n_4),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_1),
.Y(n_40)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_4),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_0),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

CKINVDCx14_ASAP7_75t_R g46 ( 
.A(n_7),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_12),
.Y(n_47)
);

INVx1_ASAP7_75t_SL g48 ( 
.A(n_2),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_5),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_0),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_8),
.Y(n_51)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_15),
.Y(n_52)
);

INVx4_ASAP7_75t_SL g53 ( 
.A(n_24),
.Y(n_53)
);

INVx2_ASAP7_75t_SL g150 ( 
.A(n_53),
.Y(n_150)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_29),
.Y(n_54)
);

BUFx2_ASAP7_75t_L g146 ( 
.A(n_54),
.Y(n_146)
);

INVx13_ASAP7_75t_L g55 ( 
.A(n_52),
.Y(n_55)
);

INVx1_ASAP7_75t_SL g144 ( 
.A(n_55),
.Y(n_144)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_31),
.Y(n_56)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_56),
.Y(n_107)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_31),
.Y(n_57)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_57),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_24),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_58),
.Y(n_116)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_31),
.Y(n_59)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_59),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_24),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_60),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_24),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_61),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_25),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_62),
.Y(n_167)
);

OR2x2_ASAP7_75t_L g63 ( 
.A(n_39),
.B(n_10),
.Y(n_63)
);

NAND2xp33_ASAP7_75t_SL g125 ( 
.A(n_63),
.B(n_68),
.Y(n_125)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_64),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_25),
.Y(n_65)
);

INVx6_ASAP7_75t_L g137 ( 
.A(n_65),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_25),
.Y(n_66)
);

INVx6_ASAP7_75t_L g154 ( 
.A(n_66),
.Y(n_154)
);

INVx2_ASAP7_75t_SL g67 ( 
.A(n_36),
.Y(n_67)
);

HB1xp67_ASAP7_75t_L g147 ( 
.A(n_67),
.Y(n_147)
);

OR2x2_ASAP7_75t_L g68 ( 
.A(n_39),
.B(n_10),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_51),
.Y(n_69)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_69),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_25),
.Y(n_70)
);

INVx8_ASAP7_75t_L g121 ( 
.A(n_70),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_20),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g134 ( 
.A(n_71),
.Y(n_134)
);

HAxp5_ASAP7_75t_SL g72 ( 
.A(n_46),
.B(n_0),
.CON(n_72),
.SN(n_72)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_72),
.B(n_100),
.Y(n_132)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_29),
.Y(n_73)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_73),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_32),
.Y(n_74)
);

INVx8_ASAP7_75t_L g122 ( 
.A(n_74),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_32),
.Y(n_75)
);

INVx3_ASAP7_75t_SL g164 ( 
.A(n_75),
.Y(n_164)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_20),
.Y(n_76)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_76),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_32),
.Y(n_77)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_77),
.Y(n_139)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_20),
.Y(n_78)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_78),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_32),
.Y(n_79)
);

INVx5_ASAP7_75t_L g170 ( 
.A(n_79),
.Y(n_170)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_29),
.Y(n_80)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_80),
.Y(n_142)
);

BUFx24_ASAP7_75t_L g81 ( 
.A(n_52),
.Y(n_81)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_81),
.Y(n_126)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_35),
.Y(n_82)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_82),
.Y(n_143)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_51),
.Y(n_83)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_83),
.Y(n_138)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_35),
.Y(n_84)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_84),
.Y(n_145)
);

BUFx12_ASAP7_75t_L g85 ( 
.A(n_26),
.Y(n_85)
);

INVx6_ASAP7_75t_SL g160 ( 
.A(n_85),
.Y(n_160)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_36),
.Y(n_86)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_86),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_37),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g172 ( 
.A(n_87),
.Y(n_172)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_27),
.Y(n_88)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_88),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_37),
.Y(n_89)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_89),
.Y(n_109)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_36),
.Y(n_90)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_90),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_37),
.Y(n_91)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_91),
.Y(n_111)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_27),
.Y(n_92)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_92),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_41),
.Y(n_93)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_93),
.Y(n_112)
);

INVx13_ASAP7_75t_L g94 ( 
.A(n_46),
.Y(n_94)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_94),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_41),
.Y(n_95)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_95),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_19),
.B(n_10),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_96),
.B(n_16),
.Y(n_141)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_35),
.Y(n_97)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_97),
.Y(n_157)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_26),
.Y(n_98)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_98),
.Y(n_171)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_26),
.Y(n_99)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_99),
.Y(n_163)
);

BUFx12f_ASAP7_75t_L g100 ( 
.A(n_30),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_27),
.Y(n_101)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_101),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_30),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_102),
.B(n_105),
.Y(n_161)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_41),
.Y(n_103)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_103),
.Y(n_120)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_22),
.Y(n_104)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_104),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_30),
.Y(n_105)
);

NAND2x1_ASAP7_75t_L g106 ( 
.A(n_22),
.B(n_10),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_106),
.B(n_48),
.Y(n_113)
);

NAND3xp33_ASAP7_75t_L g178 ( 
.A(n_113),
.B(n_117),
.C(n_94),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_81),
.A2(n_48),
.B1(n_34),
.B2(n_22),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_115),
.B(n_7),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_63),
.B(n_19),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_67),
.A2(n_48),
.B1(n_38),
.B2(n_72),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_123),
.A2(n_127),
.B1(n_131),
.B2(n_153),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_68),
.A2(n_34),
.B1(n_49),
.B2(n_47),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_124),
.A2(n_136),
.B1(n_149),
.B2(n_152),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_58),
.A2(n_34),
.B1(n_49),
.B2(n_47),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_85),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_130),
.B(n_166),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_86),
.A2(n_38),
.B1(n_43),
.B2(n_42),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_60),
.A2(n_21),
.B1(n_28),
.B2(n_38),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_141),
.B(n_156),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_61),
.A2(n_77),
.B1(n_79),
.B2(n_62),
.Y(n_149)
);

OAI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_65),
.A2(n_50),
.B1(n_45),
.B2(n_44),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_90),
.A2(n_38),
.B1(n_43),
.B2(n_42),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_106),
.B(n_21),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_103),
.A2(n_42),
.B1(n_43),
.B2(n_23),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_165),
.A2(n_169),
.B1(n_33),
.B2(n_44),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_100),
.B(n_28),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_87),
.A2(n_40),
.B1(n_23),
.B2(n_50),
.Y(n_169)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_120),
.Y(n_173)
);

INVx1_ASAP7_75t_SL g260 ( 
.A(n_173),
.Y(n_260)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_172),
.Y(n_174)
);

INVx4_ASAP7_75t_L g246 ( 
.A(n_174),
.Y(n_246)
);

BUFx3_ASAP7_75t_L g175 ( 
.A(n_160),
.Y(n_175)
);

INVx5_ASAP7_75t_L g288 ( 
.A(n_175),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_147),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_177),
.B(n_178),
.Y(n_248)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_135),
.Y(n_179)
);

HB1xp67_ASAP7_75t_L g250 ( 
.A(n_179),
.Y(n_250)
);

OAI22xp33_ASAP7_75t_L g180 ( 
.A1(n_169),
.A2(n_89),
.B1(n_95),
.B2(n_93),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_180),
.A2(n_198),
.B1(n_212),
.B2(n_225),
.Y(n_258)
);

BUFx3_ASAP7_75t_L g181 ( 
.A(n_134),
.Y(n_181)
);

INVx3_ASAP7_75t_L g237 ( 
.A(n_181),
.Y(n_237)
);

HB1xp67_ASAP7_75t_L g182 ( 
.A(n_163),
.Y(n_182)
);

HB1xp67_ASAP7_75t_L g280 ( 
.A(n_182),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_161),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_183),
.B(n_194),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_108),
.B(n_40),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_184),
.B(n_229),
.Y(n_252)
);

INVx4_ASAP7_75t_L g186 ( 
.A(n_171),
.Y(n_186)
);

INVx3_ASAP7_75t_L g272 ( 
.A(n_186),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_116),
.Y(n_187)
);

INVx8_ASAP7_75t_L g249 ( 
.A(n_187),
.Y(n_249)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_114),
.Y(n_188)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_188),
.Y(n_236)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_148),
.Y(n_189)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_189),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_116),
.Y(n_190)
);

INVx3_ASAP7_75t_L g277 ( 
.A(n_190),
.Y(n_277)
);

INVx6_ASAP7_75t_L g191 ( 
.A(n_151),
.Y(n_191)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_191),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_125),
.B(n_100),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_192),
.B(n_193),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_132),
.B(n_53),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_148),
.Y(n_194)
);

INVx8_ASAP7_75t_L g195 ( 
.A(n_151),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_195),
.Y(n_275)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_159),
.Y(n_196)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_196),
.Y(n_243)
);

O2A1O1Ixp33_ASAP7_75t_L g197 ( 
.A1(n_123),
.A2(n_55),
.B(n_33),
.C(n_50),
.Y(n_197)
);

OA22x2_ASAP7_75t_L g273 ( 
.A1(n_197),
.A2(n_223),
.B1(n_168),
.B2(n_11),
.Y(n_273)
);

HB1xp67_ASAP7_75t_L g199 ( 
.A(n_150),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g235 ( 
.A(n_199),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_144),
.A2(n_91),
.B1(n_33),
.B2(n_45),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_200),
.Y(n_276)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_107),
.Y(n_201)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_201),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_146),
.Y(n_202)
);

CKINVDCx14_ASAP7_75t_R g278 ( 
.A(n_202),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_129),
.B(n_44),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_203),
.B(n_215),
.Y(n_268)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_118),
.Y(n_204)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_204),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_144),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_205),
.B(n_213),
.Y(n_262)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_119),
.Y(n_207)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_207),
.Y(n_259)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_162),
.Y(n_208)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_208),
.Y(n_279)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_158),
.Y(n_209)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_209),
.Y(n_282)
);

HB1xp67_ASAP7_75t_L g210 ( 
.A(n_150),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g256 ( 
.A(n_210),
.Y(n_256)
);

BUFx3_ASAP7_75t_L g211 ( 
.A(n_134),
.Y(n_211)
);

CKINVDCx14_ASAP7_75t_R g289 ( 
.A(n_211),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_165),
.A2(n_75),
.B1(n_74),
.B2(n_70),
.Y(n_212)
);

INVx5_ASAP7_75t_L g213 ( 
.A(n_109),
.Y(n_213)
);

BUFx2_ASAP7_75t_L g214 ( 
.A(n_171),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_214),
.B(n_216),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_140),
.B(n_45),
.Y(n_215)
);

CKINVDCx14_ASAP7_75t_R g216 ( 
.A(n_126),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_133),
.Y(n_217)
);

NAND2xp33_ASAP7_75t_SL g245 ( 
.A(n_217),
.B(n_224),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_158),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_SL g253 ( 
.A1(n_218),
.A2(n_220),
.B1(n_231),
.B2(n_234),
.Y(n_253)
);

INVx8_ASAP7_75t_L g220 ( 
.A(n_167),
.Y(n_220)
);

HB1xp67_ASAP7_75t_L g221 ( 
.A(n_157),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_221),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_152),
.A2(n_66),
.B1(n_2),
.B2(n_3),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_222),
.A2(n_230),
.B1(n_167),
.B2(n_154),
.Y(n_251)
);

OA22x2_ASAP7_75t_L g223 ( 
.A1(n_109),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_138),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_131),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_225)
);

INVx13_ASAP7_75t_L g226 ( 
.A(n_146),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_226),
.Y(n_266)
);

BUFx8_ASAP7_75t_L g227 ( 
.A(n_164),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_227),
.Y(n_267)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_164),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_228),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_121),
.B(n_6),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_137),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_230)
);

BUFx3_ASAP7_75t_L g231 ( 
.A(n_172),
.Y(n_231)
);

OAI22xp33_ASAP7_75t_SL g232 ( 
.A1(n_153),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_232),
.A2(n_225),
.B1(n_180),
.B2(n_197),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_128),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_233),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_219),
.B(n_143),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_239),
.B(n_265),
.C(n_274),
.Y(n_330)
);

OAI22xp33_ASAP7_75t_L g241 ( 
.A1(n_222),
.A2(n_112),
.B1(n_111),
.B2(n_155),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_241),
.A2(n_251),
.B1(n_284),
.B2(n_287),
.Y(n_299)
);

OAI22xp33_ASAP7_75t_SL g242 ( 
.A1(n_206),
.A2(n_111),
.B1(n_155),
.B2(n_112),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_242),
.A2(n_228),
.B1(n_213),
.B2(n_173),
.Y(n_295)
);

AOI22xp33_ASAP7_75t_L g247 ( 
.A1(n_206),
.A2(n_121),
.B1(n_122),
.B2(n_110),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_247),
.A2(n_283),
.B1(n_281),
.B2(n_290),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_184),
.B(n_157),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_257),
.B(n_263),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_229),
.B(n_122),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_176),
.B(n_145),
.C(n_142),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_201),
.B(n_154),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_270),
.B(n_218),
.Y(n_300)
);

AND2x2_ASAP7_75t_L g316 ( 
.A(n_273),
.B(n_281),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_234),
.B(n_137),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_233),
.A2(n_170),
.B1(n_139),
.B2(n_12),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_230),
.A2(n_170),
.B1(n_139),
.B2(n_13),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_179),
.B(n_9),
.C(n_11),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_285),
.B(n_202),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_223),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_226),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_290),
.B(n_266),
.Y(n_338)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_270),
.Y(n_292)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_292),
.Y(n_341)
);

OAI21xp5_ASAP7_75t_L g293 ( 
.A1(n_264),
.A2(n_185),
.B(n_175),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_L g366 ( 
.A1(n_293),
.A2(n_296),
.B(n_306),
.Y(n_366)
);

XOR2xp5_ASAP7_75t_L g354 ( 
.A(n_294),
.B(n_325),
.Y(n_354)
);

AOI22xp33_ASAP7_75t_L g343 ( 
.A1(n_295),
.A2(n_335),
.B1(n_266),
.B2(n_256),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_276),
.A2(n_223),
.B(n_207),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_258),
.A2(n_223),
.B1(n_204),
.B2(n_191),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_297),
.A2(n_321),
.B1(n_324),
.B2(n_326),
.Y(n_344)
);

OAI32xp33_ASAP7_75t_L g298 ( 
.A1(n_252),
.A2(n_214),
.A3(n_186),
.B1(n_220),
.B2(n_195),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_298),
.B(n_300),
.Y(n_361)
);

OAI32xp33_ASAP7_75t_L g301 ( 
.A1(n_252),
.A2(n_209),
.A3(n_190),
.B1(n_187),
.B2(n_227),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_301),
.B(n_302),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_263),
.B(n_174),
.Y(n_302)
);

CKINVDCx14_ASAP7_75t_R g303 ( 
.A(n_262),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_303),
.B(n_311),
.Y(n_340)
);

INVx3_ASAP7_75t_L g304 ( 
.A(n_249),
.Y(n_304)
);

BUFx2_ASAP7_75t_L g359 ( 
.A(n_304),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_274),
.B(n_211),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g374 ( 
.A(n_305),
.B(n_308),
.Y(n_374)
);

OAI21xp5_ASAP7_75t_L g306 ( 
.A1(n_276),
.A2(n_181),
.B(n_231),
.Y(n_306)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_240),
.Y(n_307)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_307),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_257),
.B(n_13),
.Y(n_308)
);

O2A1O1Ixp33_ASAP7_75t_L g309 ( 
.A1(n_286),
.A2(n_227),
.B(n_14),
.C(n_15),
.Y(n_309)
);

AND2x2_ASAP7_75t_L g371 ( 
.A(n_309),
.B(n_328),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_265),
.A2(n_13),
.B1(n_14),
.B2(n_16),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_L g348 ( 
.A1(n_310),
.A2(n_332),
.B1(n_235),
.B2(n_249),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_261),
.B(n_14),
.Y(n_311)
);

INVxp67_ASAP7_75t_L g312 ( 
.A(n_269),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_312),
.B(n_313),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_239),
.B(n_16),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_243),
.Y(n_314)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_314),
.Y(n_353)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_243),
.Y(n_315)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_315),
.Y(n_377)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_279),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_317),
.B(n_318),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_250),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_286),
.B(n_18),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_319),
.B(n_320),
.Y(n_362)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_279),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_258),
.A2(n_18),
.B1(n_16),
.B2(n_17),
.Y(n_321)
);

AOI22xp33_ASAP7_75t_SL g322 ( 
.A1(n_251),
.A2(n_18),
.B1(n_267),
.B2(n_288),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g363 ( 
.A(n_322),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_268),
.B(n_18),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_323),
.B(n_327),
.Y(n_364)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_253),
.B(n_245),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_273),
.A2(n_241),
.B1(n_283),
.B2(n_248),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_280),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_244),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_L g329 ( 
.A1(n_273),
.A2(n_284),
.B1(n_287),
.B2(n_240),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_329),
.A2(n_334),
.B1(n_336),
.B2(n_272),
.Y(n_352)
);

AND2x2_ASAP7_75t_SL g331 ( 
.A(n_273),
.B(n_236),
.Y(n_331)
);

INVxp67_ASAP7_75t_L g376 ( 
.A(n_331),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_236),
.A2(n_271),
.B1(n_255),
.B2(n_254),
.Y(n_332)
);

CKINVDCx14_ASAP7_75t_R g333 ( 
.A(n_278),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_SL g356 ( 
.A1(n_333),
.A2(n_335),
.B(n_312),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_282),
.A2(n_271),
.B1(n_285),
.B2(n_260),
.Y(n_334)
);

CKINVDCx16_ASAP7_75t_R g335 ( 
.A(n_267),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_L g336 ( 
.A1(n_282),
.A2(n_255),
.B1(n_275),
.B2(n_277),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_L g337 ( 
.A1(n_289),
.A2(n_238),
.B(n_260),
.Y(n_337)
);

AOI21xp5_ASAP7_75t_SL g347 ( 
.A1(n_337),
.A2(n_275),
.B(n_288),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_338),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_244),
.B(n_259),
.Y(n_339)
);

MAJx2_ASAP7_75t_L g365 ( 
.A(n_339),
.B(n_237),
.C(n_330),
.Y(n_365)
);

INVxp67_ASAP7_75t_L g388 ( 
.A(n_343),
.Y(n_388)
);

AO22x1_ASAP7_75t_L g345 ( 
.A1(n_331),
.A2(n_238),
.B1(n_254),
.B2(n_259),
.Y(n_345)
);

A2O1A1Ixp33_ASAP7_75t_SL g390 ( 
.A1(n_345),
.A2(n_370),
.B(n_320),
.C(n_328),
.Y(n_390)
);

OAI21xp5_ASAP7_75t_SL g411 ( 
.A1(n_347),
.A2(n_345),
.B(n_371),
.Y(n_411)
);

AOI22xp5_ASAP7_75t_L g403 ( 
.A1(n_348),
.A2(n_358),
.B1(n_372),
.B2(n_373),
.Y(n_403)
);

BUFx3_ASAP7_75t_L g350 ( 
.A(n_304),
.Y(n_350)
);

INVx1_ASAP7_75t_SL g407 ( 
.A(n_350),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_339),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_351),
.B(n_357),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_L g412 ( 
.A1(n_352),
.A2(n_355),
.B1(n_378),
.B2(n_381),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_316),
.A2(n_277),
.B1(n_246),
.B2(n_272),
.Y(n_355)
);

INVxp67_ASAP7_75t_L g417 ( 
.A(n_356),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_332),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_L g358 ( 
.A1(n_299),
.A2(n_237),
.B1(n_246),
.B2(n_292),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_365),
.B(n_374),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_336),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_367),
.Y(n_400)
);

INVx13_ASAP7_75t_L g369 ( 
.A(n_309),
.Y(n_369)
);

CKINVDCx14_ASAP7_75t_R g391 ( 
.A(n_369),
.Y(n_391)
);

OAI21xp33_ASAP7_75t_SL g370 ( 
.A1(n_331),
.A2(n_296),
.B(n_319),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_L g372 ( 
.A1(n_299),
.A2(n_291),
.B1(n_316),
.B2(n_331),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_L g373 ( 
.A1(n_291),
.A2(n_316),
.B1(n_302),
.B2(n_329),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_330),
.A2(n_297),
.B1(n_324),
.B2(n_305),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_375),
.A2(n_379),
.B1(n_380),
.B2(n_373),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_326),
.A2(n_325),
.B1(n_321),
.B2(n_334),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_SL g379 ( 
.A1(n_300),
.A2(n_295),
.B1(n_308),
.B2(n_301),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_SL g380 ( 
.A1(n_298),
.A2(n_310),
.B1(n_313),
.B2(n_306),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_294),
.A2(n_327),
.B1(n_337),
.B2(n_293),
.Y(n_381)
);

AOI21xp5_ASAP7_75t_L g382 ( 
.A1(n_366),
.A2(n_318),
.B(n_314),
.Y(n_382)
);

A2O1A1Ixp33_ASAP7_75t_SL g425 ( 
.A1(n_382),
.A2(n_390),
.B(n_394),
.C(n_347),
.Y(n_425)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_360),
.Y(n_383)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_383),
.Y(n_423)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_360),
.Y(n_384)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_384),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_354),
.B(n_315),
.C(n_317),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_385),
.B(n_393),
.C(n_397),
.Y(n_432)
);

CKINVDCx16_ASAP7_75t_R g386 ( 
.A(n_340),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g424 ( 
.A(n_386),
.B(n_387),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_340),
.Y(n_387)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_353),
.Y(n_389)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_389),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_SL g392 ( 
.A(n_349),
.B(n_323),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_SL g443 ( 
.A(n_392),
.B(n_416),
.Y(n_443)
);

XOR2xp5_ASAP7_75t_L g393 ( 
.A(n_354),
.B(n_307),
.Y(n_393)
);

AOI21xp5_ASAP7_75t_L g394 ( 
.A1(n_366),
.A2(n_376),
.B(n_356),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_353),
.Y(n_395)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_395),
.Y(n_446)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_377),
.Y(n_396)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_396),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_365),
.B(n_381),
.C(n_375),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_344),
.A2(n_378),
.B1(n_368),
.B2(n_361),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_399),
.B(n_404),
.Y(n_419)
);

XNOR2x1_ASAP7_75t_L g418 ( 
.A(n_401),
.B(n_358),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_SL g402 ( 
.A1(n_380),
.A2(n_379),
.B1(n_372),
.B2(n_363),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_L g426 ( 
.A1(n_402),
.A2(n_409),
.B1(n_403),
.B2(n_398),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_SL g404 ( 
.A1(n_344),
.A2(n_368),
.B1(n_361),
.B2(n_352),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_377),
.Y(n_405)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_405),
.Y(n_427)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_346),
.Y(n_406)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_406),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_365),
.B(n_374),
.Y(n_408)
);

XOR2xp5_ASAP7_75t_L g421 ( 
.A(n_408),
.B(n_362),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_357),
.A2(n_367),
.B1(n_351),
.B2(n_341),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_410),
.B(n_371),
.Y(n_436)
);

AOI21xp5_ASAP7_75t_L g428 ( 
.A1(n_411),
.A2(n_371),
.B(n_347),
.Y(n_428)
);

A2O1A1O1Ixp25_ASAP7_75t_L g413 ( 
.A1(n_341),
.A2(n_349),
.B(n_370),
.C(n_362),
.D(n_364),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_413),
.B(n_414),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_342),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_346),
.Y(n_415)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_415),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_342),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_SL g473 ( 
.A(n_418),
.B(n_421),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_L g422 ( 
.A(n_393),
.B(n_345),
.Y(n_422)
);

XOR2xp5_ASAP7_75t_L g451 ( 
.A(n_422),
.B(n_429),
.Y(n_451)
);

INVxp67_ASAP7_75t_L g460 ( 
.A(n_425),
.Y(n_460)
);

INVxp67_ASAP7_75t_L g469 ( 
.A(n_426),
.Y(n_469)
);

AOI21xp5_ASAP7_75t_L g470 ( 
.A1(n_428),
.A2(n_442),
.B(n_447),
.Y(n_470)
);

XNOR2xp5_ASAP7_75t_SL g429 ( 
.A(n_401),
.B(n_408),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_L g431 ( 
.A1(n_402),
.A2(n_355),
.B1(n_364),
.B2(n_369),
.Y(n_431)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_431),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_L g434 ( 
.A(n_385),
.B(n_348),
.Y(n_434)
);

XOR2xp5_ASAP7_75t_L g454 ( 
.A(n_434),
.B(n_439),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_436),
.B(n_438),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_403),
.A2(n_369),
.B1(n_371),
.B2(n_359),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_L g439 ( 
.A(n_397),
.B(n_350),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_410),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_SL g461 ( 
.A(n_440),
.B(n_389),
.Y(n_461)
);

AOI22xp33_ASAP7_75t_SL g442 ( 
.A1(n_417),
.A2(n_350),
.B1(n_359),
.B2(n_388),
.Y(n_442)
);

AND2x2_ASAP7_75t_L g444 ( 
.A(n_400),
.B(n_359),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_444),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_400),
.B(n_383),
.Y(n_445)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_445),
.Y(n_462)
);

OAI21xp5_ASAP7_75t_L g447 ( 
.A1(n_394),
.A2(n_417),
.B(n_411),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_SL g448 ( 
.A1(n_409),
.A2(n_404),
.B1(n_399),
.B2(n_382),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_448),
.B(n_388),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_432),
.B(n_412),
.C(n_384),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_L g480 ( 
.A(n_449),
.B(n_456),
.Y(n_480)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_445),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_SL g483 ( 
.A(n_453),
.B(n_465),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_L g456 ( 
.A(n_432),
.B(n_413),
.Y(n_456)
);

XNOR2xp5_ASAP7_75t_L g457 ( 
.A(n_434),
.B(n_421),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_L g493 ( 
.A(n_457),
.B(n_464),
.Y(n_493)
);

OAI22xp5_ASAP7_75t_SL g494 ( 
.A1(n_458),
.A2(n_455),
.B1(n_428),
.B2(n_470),
.Y(n_494)
);

BUFx6f_ASAP7_75t_L g459 ( 
.A(n_423),
.Y(n_459)
);

INVx6_ASAP7_75t_L g481 ( 
.A(n_459),
.Y(n_481)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_461),
.Y(n_479)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_430),
.Y(n_463)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_463),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_429),
.B(n_390),
.Y(n_464)
);

CKINVDCx20_ASAP7_75t_R g465 ( 
.A(n_444),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_439),
.B(n_390),
.C(n_415),
.Y(n_466)
);

XOR2xp5_ASAP7_75t_L g484 ( 
.A(n_466),
.B(n_468),
.Y(n_484)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_424),
.Y(n_467)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_467),
.Y(n_490)
);

XOR2xp5_ASAP7_75t_L g468 ( 
.A(n_422),
.B(n_418),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_L g471 ( 
.A(n_448),
.B(n_390),
.Y(n_471)
);

XOR2xp5_ASAP7_75t_L g488 ( 
.A(n_471),
.B(n_472),
.Y(n_488)
);

XOR2xp5_ASAP7_75t_L g472 ( 
.A(n_419),
.B(n_390),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_444),
.B(n_406),
.Y(n_474)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_474),
.Y(n_491)
);

XOR2x2_ASAP7_75t_L g475 ( 
.A(n_464),
.B(n_473),
.Y(n_475)
);

AOI21xp5_ASAP7_75t_L g510 ( 
.A1(n_475),
.A2(n_489),
.B(n_427),
.Y(n_510)
);

OAI22xp5_ASAP7_75t_L g476 ( 
.A1(n_469),
.A2(n_443),
.B1(n_450),
.B2(n_433),
.Y(n_476)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_476),
.Y(n_502)
);

CKINVDCx16_ASAP7_75t_R g477 ( 
.A(n_474),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g504 ( 
.A(n_477),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_452),
.B(n_435),
.Y(n_478)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_478),
.Y(n_509)
);

AOI22xp5_ASAP7_75t_L g485 ( 
.A1(n_469),
.A2(n_438),
.B1(n_419),
.B2(n_436),
.Y(n_485)
);

OAI22xp5_ASAP7_75t_SL g496 ( 
.A1(n_485),
.A2(n_470),
.B1(n_460),
.B2(n_449),
.Y(n_496)
);

XNOR2x1_ASAP7_75t_L g486 ( 
.A(n_466),
.B(n_425),
.Y(n_486)
);

XOR2xp5_ASAP7_75t_L g500 ( 
.A(n_486),
.B(n_492),
.Y(n_500)
);

CKINVDCx16_ASAP7_75t_R g487 ( 
.A(n_455),
.Y(n_487)
);

HB1xp67_ASAP7_75t_L g498 ( 
.A(n_487),
.Y(n_498)
);

XOR2x2_ASAP7_75t_L g489 ( 
.A(n_473),
.B(n_447),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_462),
.B(n_441),
.Y(n_492)
);

AOI22xp5_ASAP7_75t_L g511 ( 
.A1(n_494),
.A2(n_495),
.B1(n_446),
.B2(n_396),
.Y(n_511)
);

OAI22xp5_ASAP7_75t_L g495 ( 
.A1(n_458),
.A2(n_391),
.B1(n_441),
.B2(n_435),
.Y(n_495)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_496),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_480),
.B(n_454),
.C(n_457),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_SL g521 ( 
.A(n_497),
.B(n_506),
.Y(n_521)
);

OAI22xp5_ASAP7_75t_SL g499 ( 
.A1(n_485),
.A2(n_460),
.B1(n_471),
.B2(n_472),
.Y(n_499)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_499),
.Y(n_513)
);

AOI22xp5_ASAP7_75t_SL g501 ( 
.A1(n_494),
.A2(n_425),
.B1(n_468),
.B2(n_456),
.Y(n_501)
);

OAI22xp5_ASAP7_75t_SL g514 ( 
.A1(n_501),
.A2(n_507),
.B1(n_511),
.B2(n_486),
.Y(n_514)
);

OAI21xp5_ASAP7_75t_L g503 ( 
.A1(n_491),
.A2(n_425),
.B(n_459),
.Y(n_503)
);

OAI21xp5_ASAP7_75t_L g519 ( 
.A1(n_503),
.A2(n_510),
.B(n_488),
.Y(n_519)
);

OAI22xp5_ASAP7_75t_SL g505 ( 
.A1(n_483),
.A2(n_427),
.B1(n_420),
.B2(n_437),
.Y(n_505)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_505),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_480),
.B(n_454),
.C(n_451),
.Y(n_506)
);

AOI22xp5_ASAP7_75t_SL g507 ( 
.A1(n_491),
.A2(n_489),
.B1(n_478),
.B2(n_479),
.Y(n_507)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_484),
.B(n_451),
.C(n_420),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_508),
.B(n_493),
.C(n_407),
.Y(n_523)
);

OAI22xp5_ASAP7_75t_SL g512 ( 
.A1(n_492),
.A2(n_395),
.B1(n_405),
.B2(n_407),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_512),
.B(n_488),
.Y(n_516)
);

XOR2xp5_ASAP7_75t_L g529 ( 
.A(n_514),
.B(n_519),
.Y(n_529)
);

CKINVDCx14_ASAP7_75t_R g515 ( 
.A(n_498),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_515),
.B(n_516),
.Y(n_535)
);

OAI22xp5_ASAP7_75t_L g520 ( 
.A1(n_502),
.A2(n_490),
.B1(n_482),
.B2(n_481),
.Y(n_520)
);

XNOR2xp5_ASAP7_75t_L g534 ( 
.A(n_520),
.B(n_522),
.Y(n_534)
);

AOI21xp5_ASAP7_75t_L g522 ( 
.A1(n_507),
.A2(n_475),
.B(n_484),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_523),
.B(n_525),
.Y(n_527)
);

OAI21xp5_ASAP7_75t_L g524 ( 
.A1(n_503),
.A2(n_493),
.B(n_481),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_SL g532 ( 
.A(n_524),
.B(n_526),
.Y(n_532)
);

NOR2xp67_ASAP7_75t_L g525 ( 
.A(n_508),
.B(n_497),
.Y(n_525)
);

OAI21xp5_ASAP7_75t_L g526 ( 
.A1(n_510),
.A2(n_499),
.B(n_509),
.Y(n_526)
);

MAJIxp5_ASAP7_75t_L g528 ( 
.A(n_518),
.B(n_506),
.C(n_511),
.Y(n_528)
);

AOI21xp5_ASAP7_75t_L g536 ( 
.A1(n_528),
.A2(n_531),
.B(n_524),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_521),
.B(n_504),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_530),
.B(n_533),
.Y(n_538)
);

MAJIxp5_ASAP7_75t_L g531 ( 
.A(n_518),
.B(n_496),
.C(n_500),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_513),
.B(n_509),
.Y(n_533)
);

AND2x2_ASAP7_75t_L g543 ( 
.A(n_536),
.B(n_540),
.Y(n_543)
);

AOI21xp5_ASAP7_75t_L g537 ( 
.A1(n_527),
.A2(n_526),
.B(n_519),
.Y(n_537)
);

OAI21xp5_ASAP7_75t_SL g544 ( 
.A1(n_537),
.A2(n_522),
.B(n_531),
.Y(n_544)
);

INVx11_ASAP7_75t_L g539 ( 
.A(n_535),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_539),
.B(n_541),
.Y(n_542)
);

AO21x1_ASAP7_75t_L g540 ( 
.A1(n_532),
.A2(n_517),
.B(n_514),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_528),
.B(n_523),
.Y(n_541)
);

MAJIxp5_ASAP7_75t_L g546 ( 
.A(n_544),
.B(n_538),
.C(n_534),
.Y(n_546)
);

NAND4xp25_ASAP7_75t_L g545 ( 
.A(n_542),
.B(n_538),
.C(n_543),
.D(n_529),
.Y(n_545)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_545),
.Y(n_547)
);

MAJIxp5_ASAP7_75t_L g548 ( 
.A(n_547),
.B(n_546),
.C(n_529),
.Y(n_548)
);

NOR3xp33_ASAP7_75t_L g549 ( 
.A(n_548),
.B(n_500),
.C(n_512),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_549),
.B(n_505),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_L g551 ( 
.A(n_550),
.B(n_501),
.Y(n_551)
);


endmodule