module fake_jpeg_1986_n_260 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_260);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_260;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

BUFx2_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx5_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx8_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_5),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_16),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_4),
.Y(n_32)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_0),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_0),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_37),
.Y(n_40)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_40),
.Y(n_80)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_43),
.Y(n_81)
);

INVx3_ASAP7_75t_SL g44 ( 
.A(n_25),
.Y(n_44)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_44),
.Y(n_84)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_25),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_46),
.Y(n_97)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_26),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_26),
.Y(n_48)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_48),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_21),
.Y(n_49)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_29),
.B(n_17),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_50),
.B(n_54),
.Y(n_64)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_24),
.Y(n_51)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_51),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_31),
.B(n_1),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_52),
.B(n_34),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_18),
.B(n_1),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_53),
.B(n_58),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_29),
.B(n_17),
.Y(n_54)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_26),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_55),
.B(n_56),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_21),
.Y(n_56)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_24),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_57),
.B(n_59),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_18),
.B(n_1),
.Y(n_58)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_24),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_19),
.B(n_16),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_60),
.B(n_62),
.Y(n_83)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_20),
.Y(n_61)
);

HAxp5_ASAP7_75t_SL g76 ( 
.A(n_61),
.B(n_33),
.CON(n_76),
.SN(n_76)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_22),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_18),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_63),
.B(n_27),
.Y(n_73)
);

NAND2x1_ASAP7_75t_L g67 ( 
.A(n_53),
.B(n_24),
.Y(n_67)
);

A2O1A1Ixp33_ASAP7_75t_L g129 ( 
.A1(n_67),
.A2(n_93),
.B(n_15),
.C(n_11),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_42),
.A2(n_20),
.B1(n_22),
.B2(n_27),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_71),
.A2(n_87),
.B1(n_92),
.B2(n_45),
.Y(n_103)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_73),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_58),
.A2(n_21),
.B1(n_30),
.B2(n_23),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_74),
.A2(n_79),
.B1(n_56),
.B2(n_46),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_40),
.A2(n_23),
.B1(n_30),
.B2(n_39),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g128 ( 
.A1(n_75),
.A2(n_77),
.B1(n_86),
.B2(n_9),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_76),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_49),
.A2(n_23),
.B1(n_30),
.B2(n_39),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_63),
.B(n_38),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_78),
.B(n_85),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_49),
.A2(n_55),
.B1(n_47),
.B2(n_27),
.Y(n_79)
);

OAI21xp33_ASAP7_75t_L g85 ( 
.A1(n_44),
.A2(n_36),
.B(n_35),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_44),
.A2(n_34),
.B1(n_32),
.B2(n_28),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_42),
.A2(n_36),
.B1(n_35),
.B2(n_31),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_56),
.B(n_38),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_88),
.B(n_89),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_62),
.B(n_32),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_90),
.B(n_95),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_42),
.A2(n_28),
.B1(n_3),
.B2(n_5),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_56),
.B(n_2),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_51),
.B(n_2),
.Y(n_95)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_80),
.Y(n_98)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_98),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_64),
.B(n_59),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_102),
.B(n_108),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_103),
.Y(n_141)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_80),
.Y(n_104)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_104),
.Y(n_151)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_84),
.Y(n_105)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_105),
.Y(n_132)
);

AO22x1_ASAP7_75t_L g106 ( 
.A1(n_79),
.A2(n_74),
.B1(n_94),
.B2(n_84),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_106),
.B(n_122),
.Y(n_142)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_94),
.Y(n_107)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_107),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_90),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_89),
.B(n_57),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_109),
.B(n_112),
.Y(n_154)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_94),
.Y(n_110)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_110),
.Y(n_144)
);

INVx8_ASAP7_75t_L g111 ( 
.A(n_96),
.Y(n_111)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_111),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_70),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_78),
.Y(n_113)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_113),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_97),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_114),
.Y(n_150)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_88),
.Y(n_115)
);

INVx1_ASAP7_75t_SL g134 ( 
.A(n_115),
.Y(n_134)
);

O2A1O1Ixp33_ASAP7_75t_L g116 ( 
.A1(n_67),
.A2(n_43),
.B(n_61),
.C(n_41),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_116),
.B(n_126),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_118),
.A2(n_69),
.B1(n_66),
.B2(n_82),
.Y(n_147)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_68),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_119),
.Y(n_146)
);

OA22x2_ASAP7_75t_SL g121 ( 
.A1(n_67),
.A2(n_48),
.B1(n_3),
.B2(n_6),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_121),
.Y(n_139)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_65),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_91),
.A2(n_48),
.B1(n_6),
.B2(n_7),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_123),
.Y(n_140)
);

BUFx12f_ASAP7_75t_L g124 ( 
.A(n_82),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_124),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_91),
.A2(n_48),
.B1(n_7),
.B2(n_8),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_125),
.A2(n_127),
.B1(n_93),
.B2(n_65),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_83),
.B(n_2),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_73),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_L g131 ( 
.A1(n_128),
.A2(n_81),
.B1(n_68),
.B2(n_69),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_129),
.B(n_10),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_130),
.A2(n_136),
.B1(n_145),
.B2(n_147),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_131),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_99),
.B(n_97),
.C(n_72),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_133),
.B(n_124),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_113),
.A2(n_66),
.B1(n_72),
.B2(n_81),
.Y(n_136)
);

NAND2xp33_ASAP7_75t_L g159 ( 
.A(n_143),
.B(n_125),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_99),
.A2(n_118),
.B1(n_115),
.B2(n_101),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_106),
.A2(n_66),
.B1(n_76),
.B2(n_96),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_149),
.A2(n_107),
.B1(n_123),
.B2(n_127),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_154),
.A2(n_112),
.B(n_117),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_156),
.A2(n_160),
.B(n_179),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_138),
.B(n_108),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_157),
.Y(n_190)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_132),
.Y(n_158)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_158),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_159),
.B(n_168),
.Y(n_181)
);

A2O1A1O1Ixp25_ASAP7_75t_L g160 ( 
.A1(n_139),
.A2(n_129),
.B(n_120),
.C(n_116),
.D(n_121),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_145),
.A2(n_106),
.B1(n_121),
.B2(n_110),
.Y(n_162)
);

OAI21xp33_ASAP7_75t_SL g192 ( 
.A1(n_162),
.A2(n_167),
.B(n_149),
.Y(n_192)
);

BUFx2_ASAP7_75t_L g163 ( 
.A(n_155),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_163),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_165),
.B(n_169),
.Y(n_186)
);

HB1xp67_ASAP7_75t_L g166 ( 
.A(n_146),
.Y(n_166)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_166),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_142),
.A2(n_100),
.B1(n_122),
.B2(n_98),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_134),
.B(n_105),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_153),
.B(n_104),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_142),
.A2(n_111),
.B1(n_114),
.B2(n_119),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_170),
.B(n_171),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_142),
.A2(n_124),
.B1(n_13),
.B2(n_14),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_132),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_172),
.B(n_173),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_150),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_174),
.B(n_176),
.Y(n_193)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_148),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_175),
.B(n_178),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_134),
.B(n_11),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_150),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_177),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_153),
.A2(n_124),
.B1(n_13),
.B2(n_15),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_146),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_173),
.A2(n_141),
.B(n_135),
.Y(n_182)
);

AOI22x1_ASAP7_75t_L g210 ( 
.A1(n_182),
.A2(n_183),
.B1(n_136),
.B2(n_178),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_173),
.A2(n_141),
.B(n_162),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_156),
.A2(n_135),
.B(n_143),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_185),
.A2(n_191),
.B(n_194),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_169),
.B(n_133),
.C(n_144),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_187),
.B(n_137),
.C(n_172),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_160),
.A2(n_174),
.B(n_170),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_192),
.A2(n_161),
.B1(n_165),
.B2(n_164),
.Y(n_202)
);

NAND2x1_ASAP7_75t_L g194 ( 
.A(n_167),
.B(n_144),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_161),
.A2(n_147),
.B(n_152),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_197),
.B(n_171),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_187),
.B(n_198),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_200),
.B(n_207),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_190),
.B(n_177),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_201),
.B(n_209),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_202),
.A2(n_208),
.B1(n_188),
.B2(n_181),
.Y(n_222)
);

BUFx24_ASAP7_75t_SL g203 ( 
.A(n_185),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_203),
.B(n_214),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_204),
.B(n_211),
.C(n_180),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_186),
.A2(n_191),
.B1(n_197),
.B2(n_183),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_205),
.A2(n_183),
.B1(n_186),
.B2(n_182),
.Y(n_217)
);

AND2x4_ASAP7_75t_L g225 ( 
.A(n_206),
.B(n_210),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_SL g207 ( 
.A(n_198),
.B(n_137),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_192),
.A2(n_140),
.B1(n_164),
.B2(n_130),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_193),
.B(n_148),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_187),
.B(n_158),
.C(n_175),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_180),
.Y(n_212)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_212),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_193),
.B(n_151),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_189),
.B(n_179),
.Y(n_215)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_215),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_217),
.A2(n_208),
.B1(n_210),
.B2(n_207),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_218),
.B(n_220),
.C(n_226),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_211),
.B(n_184),
.C(n_182),
.Y(n_220)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_222),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_202),
.A2(n_185),
.B1(n_181),
.B2(n_188),
.Y(n_224)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_224),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_204),
.B(n_184),
.C(n_194),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_227),
.A2(n_213),
.B(n_205),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_229),
.B(n_232),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_231),
.A2(n_225),
.B1(n_196),
.B2(n_194),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_225),
.A2(n_210),
.B(n_200),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_218),
.B(n_189),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_233),
.B(n_235),
.Y(n_243)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_223),
.Y(n_235)
);

CKINVDCx16_ASAP7_75t_R g236 ( 
.A(n_221),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_236),
.A2(n_219),
.B1(n_226),
.B2(n_195),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_237),
.B(n_238),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_230),
.B(n_220),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_230),
.B(n_216),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_SL g244 ( 
.A(n_239),
.B(n_231),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_240),
.B(n_242),
.Y(n_245)
);

NOR2xp67_ASAP7_75t_L g242 ( 
.A(n_234),
.B(n_216),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_244),
.B(n_239),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_241),
.A2(n_225),
.B1(n_228),
.B2(n_229),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_246),
.A2(n_247),
.B(n_232),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_243),
.B(n_228),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_249),
.B(n_250),
.C(n_251),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_245),
.A2(n_225),
.B1(n_238),
.B2(n_237),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_246),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_252),
.B(n_248),
.C(n_194),
.Y(n_254)
);

AOI21x1_ASAP7_75t_L g256 ( 
.A1(n_254),
.A2(n_196),
.B(n_163),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_SL g255 ( 
.A1(n_250),
.A2(n_195),
.B(n_199),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_255),
.B(n_155),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_256),
.B(n_257),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_SL g259 ( 
.A1(n_258),
.A2(n_253),
.B(n_151),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_259),
.B(n_15),
.Y(n_260)
);


endmodule