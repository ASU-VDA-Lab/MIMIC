module fake_jpeg_15472_n_81 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_81);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_81;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_80;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

NAND2xp5_ASAP7_75t_L g10 ( 
.A(n_8),
.B(n_9),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_3),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_8),
.Y(n_12)
);

INVx4_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_6),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

AND2x2_ASAP7_75t_SL g22 ( 
.A(n_10),
.B(n_0),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_22),
.B(n_24),
.Y(n_31)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

HB1xp67_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_13),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_25)
);

OR2x2_ASAP7_75t_L g34 ( 
.A(n_25),
.B(n_29),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_10),
.B(n_2),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_26),
.B(n_28),
.Y(n_36)
);

OAI22xp33_ASAP7_75t_SL g27 ( 
.A1(n_13),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_27),
.B(n_4),
.Y(n_35)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_22),
.B(n_17),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_30),
.B(n_12),
.Y(n_50)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_28),
.Y(n_32)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

NOR2x1_ASAP7_75t_L g33 ( 
.A(n_22),
.B(n_21),
.Y(n_33)
);

NOR3xp33_ASAP7_75t_L g46 ( 
.A(n_33),
.B(n_35),
.C(n_11),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_22),
.B(n_16),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_38),
.B(n_18),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_L g39 ( 
.A1(n_31),
.A2(n_25),
.B(n_26),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_49),
.C(n_36),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_34),
.A2(n_29),
.B1(n_23),
.B2(n_20),
.Y(n_40)
);

NOR3xp33_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_43),
.C(n_46),
.Y(n_55)
);

O2A1O1Ixp33_ASAP7_75t_L g41 ( 
.A1(n_33),
.A2(n_21),
.B(n_11),
.C(n_18),
.Y(n_41)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

OAI21xp33_ASAP7_75t_L g57 ( 
.A1(n_42),
.A2(n_47),
.B(n_48),
.Y(n_57)
);

OR2x2_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_24),
.Y(n_43)
);

BUFx12_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

OAI21xp33_ASAP7_75t_L g47 ( 
.A1(n_31),
.A2(n_14),
.B(n_20),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_34),
.A2(n_12),
.B1(n_17),
.B2(n_15),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_38),
.B(n_19),
.C(n_15),
.Y(n_49)
);

HAxp5_ASAP7_75t_SL g53 ( 
.A(n_50),
.B(n_35),
.CON(n_53),
.SN(n_53)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_53),
.B(n_54),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_43),
.B(n_36),
.Y(n_54)
);

XOR2xp5_ASAP7_75t_L g63 ( 
.A(n_56),
.B(n_37),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_42),
.B(n_34),
.Y(n_58)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_58),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g59 ( 
.A(n_52),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_59),
.B(n_60),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_SL g60 ( 
.A1(n_51),
.A2(n_39),
.B(n_41),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_SL g62 ( 
.A1(n_54),
.A2(n_40),
.B(n_49),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_62),
.B(n_63),
.C(n_45),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_51),
.A2(n_58),
.B1(n_56),
.B2(n_55),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_65),
.A2(n_37),
.B1(n_52),
.B2(n_19),
.Y(n_69)
);

XOR2xp5_ASAP7_75t_L g66 ( 
.A(n_63),
.B(n_57),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_68),
.A2(n_69),
.B1(n_67),
.B2(n_61),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_64),
.B(n_44),
.C(n_7),
.Y(n_70)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_70),
.Y(n_73)
);

AO221x1_ASAP7_75t_L g72 ( 
.A1(n_69),
.A2(n_59),
.B1(n_44),
.B2(n_4),
.C(n_60),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_72),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_SL g75 ( 
.A1(n_71),
.A2(n_66),
.B(n_4),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_75),
.B(n_73),
.Y(n_77)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_74),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_76),
.Y(n_78)
);

INVxp67_ASAP7_75t_SL g79 ( 
.A(n_77),
.Y(n_79)
);

BUFx24_ASAP7_75t_SL g80 ( 
.A(n_79),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_80),
.B(n_78),
.Y(n_81)
);


endmodule