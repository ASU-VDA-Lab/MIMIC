module real_aes_268_n_98 (n_17, n_28, n_76, n_56, n_34, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_98);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_98;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_357;
wire n_287;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_421;
wire n_319;
wire n_555;
wire n_766;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_786;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_791;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_808;
wire n_770;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_417;
wire n_363;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_527;
wire n_769;
wire n_434;
wire n_502;
wire n_505;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_768;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_749;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_789;
wire n_268;
wire n_544;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_639;
wire n_587;
wire n_546;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
NAND2xp5_ASAP7_75t_SL g190 ( .A(n_0), .B(n_123), .Y(n_190) );
AOI21xp5_ASAP7_75t_L g153 ( .A1(n_1), .A2(n_132), .B(n_154), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g781 ( .A(n_2), .B(n_782), .Y(n_781) );
NAND2xp5_ASAP7_75t_SL g202 ( .A(n_3), .B(n_139), .Y(n_202) );
INVx1_ASAP7_75t_L g130 ( .A(n_4), .Y(n_130) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_5), .B(n_139), .Y(n_177) );
NAND2xp5_ASAP7_75t_SL g462 ( .A(n_6), .B(n_143), .Y(n_462) );
INVx1_ASAP7_75t_L g496 ( .A(n_7), .Y(n_496) );
CKINVDCx16_ASAP7_75t_R g782 ( .A(n_8), .Y(n_782) );
CKINVDCx5p33_ASAP7_75t_R g534 ( .A(n_9), .Y(n_534) );
NAND2xp33_ASAP7_75t_L g140 ( .A(n_10), .B(n_141), .Y(n_140) );
INVx2_ASAP7_75t_L g120 ( .A(n_11), .Y(n_120) );
AOI221x1_ASAP7_75t_L g218 ( .A1(n_12), .A2(n_24), .B1(n_123), .B2(n_132), .C(n_219), .Y(n_218) );
CKINVDCx16_ASAP7_75t_R g105 ( .A(n_13), .Y(n_105) );
NAND2xp5_ASAP7_75t_SL g122 ( .A(n_14), .B(n_123), .Y(n_122) );
AO21x2_ASAP7_75t_L g117 ( .A1(n_15), .A2(n_118), .B(n_121), .Y(n_117) );
INVx1_ASAP7_75t_L g471 ( .A(n_16), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_17), .B(n_157), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_18), .B(n_139), .Y(n_166) );
AO21x1_ASAP7_75t_L g197 ( .A1(n_19), .A2(n_123), .B(n_198), .Y(n_197) );
INVx1_ASAP7_75t_L g108 ( .A(n_20), .Y(n_108) );
INVx1_ASAP7_75t_L g469 ( .A(n_21), .Y(n_469) );
INVx1_ASAP7_75t_SL g479 ( .A(n_22), .Y(n_479) );
NAND2xp5_ASAP7_75t_SL g562 ( .A(n_23), .B(n_124), .Y(n_562) );
NAND2x1_ASAP7_75t_L g188 ( .A(n_25), .B(n_139), .Y(n_188) );
AOI33xp33_ASAP7_75t_L g508 ( .A1(n_26), .A2(n_51), .A3(n_446), .B1(n_451), .B2(n_509), .B3(n_510), .Y(n_508) );
NAND2x1_ASAP7_75t_L g176 ( .A(n_27), .B(n_141), .Y(n_176) );
INVx1_ASAP7_75t_L g528 ( .A(n_28), .Y(n_528) );
OA21x2_ASAP7_75t_L g119 ( .A1(n_29), .A2(n_84), .B(n_120), .Y(n_119) );
OR2x2_ASAP7_75t_L g144 ( .A(n_29), .B(n_84), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_30), .B(n_454), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_31), .B(n_141), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g138 ( .A(n_32), .B(n_139), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_33), .B(n_141), .Y(n_201) );
AOI21xp5_ASAP7_75t_L g207 ( .A1(n_34), .A2(n_132), .B(n_208), .Y(n_207) );
AND2x2_ASAP7_75t_L g129 ( .A(n_35), .B(n_130), .Y(n_129) );
AND2x2_ASAP7_75t_L g133 ( .A(n_35), .B(n_134), .Y(n_133) );
INVx1_ASAP7_75t_L g445 ( .A(n_35), .Y(n_445) );
OR2x6_ASAP7_75t_L g106 ( .A(n_36), .B(n_107), .Y(n_106) );
CKINVDCx20_ASAP7_75t_R g530 ( .A(n_37), .Y(n_530) );
NAND2xp5_ASAP7_75t_SL g211 ( .A(n_38), .B(n_123), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_39), .B(n_454), .Y(n_516) );
AOI22xp5_ASAP7_75t_L g555 ( .A1(n_40), .A2(n_143), .B1(n_150), .B2(n_556), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_41), .B(n_564), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_42), .B(n_124), .Y(n_480) );
CKINVDCx20_ASAP7_75t_R g170 ( .A(n_43), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_44), .B(n_141), .Y(n_209) );
CKINVDCx20_ASAP7_75t_R g801 ( .A(n_45), .Y(n_801) );
NAND2xp5_ASAP7_75t_SL g498 ( .A(n_46), .B(n_118), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_47), .B(n_124), .Y(n_497) );
AOI21xp5_ASAP7_75t_L g174 ( .A1(n_48), .A2(n_132), .B(n_175), .Y(n_174) );
CKINVDCx5p33_ASAP7_75t_R g559 ( .A(n_49), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_50), .B(n_141), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_52), .B(n_124), .Y(n_520) );
INVx1_ASAP7_75t_L g126 ( .A(n_53), .Y(n_126) );
INVx1_ASAP7_75t_L g136 ( .A(n_53), .Y(n_136) );
AND2x2_ASAP7_75t_L g521 ( .A(n_54), .B(n_157), .Y(n_521) );
AOI221xp5_ASAP7_75t_L g494 ( .A1(n_55), .A2(n_72), .B1(n_443), .B2(n_454), .C(n_495), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_56), .B(n_454), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_57), .B(n_139), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_58), .B(n_150), .Y(n_536) );
AOI21xp5_ASAP7_75t_SL g442 ( .A1(n_59), .A2(n_443), .B(n_448), .Y(n_442) );
AOI21xp5_ASAP7_75t_L g186 ( .A1(n_60), .A2(n_132), .B(n_187), .Y(n_186) );
INVx1_ASAP7_75t_L g465 ( .A(n_61), .Y(n_465) );
AO21x1_ASAP7_75t_L g199 ( .A1(n_62), .A2(n_132), .B(n_200), .Y(n_199) );
NAND2xp5_ASAP7_75t_SL g152 ( .A(n_63), .B(n_123), .Y(n_152) );
INVx1_ASAP7_75t_L g519 ( .A(n_64), .Y(n_519) );
NAND2xp5_ASAP7_75t_SL g178 ( .A(n_65), .B(n_123), .Y(n_178) );
AOI21xp5_ASAP7_75t_L g517 ( .A1(n_66), .A2(n_443), .B(n_518), .Y(n_517) );
AND2x2_ASAP7_75t_L g212 ( .A(n_67), .B(n_158), .Y(n_212) );
INVx1_ASAP7_75t_L g128 ( .A(n_68), .Y(n_128) );
INVx1_ASAP7_75t_L g134 ( .A(n_68), .Y(n_134) );
AND2x2_ASAP7_75t_L g180 ( .A(n_69), .B(n_149), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_70), .B(n_454), .Y(n_511) );
AOI22xp33_ASAP7_75t_L g768 ( .A1(n_71), .A2(n_100), .B1(n_769), .B2(n_773), .Y(n_768) );
AND2x2_ASAP7_75t_L g481 ( .A(n_73), .B(n_149), .Y(n_481) );
INVx1_ASAP7_75t_L g466 ( .A(n_74), .Y(n_466) );
AOI21xp5_ASAP7_75t_L g477 ( .A1(n_75), .A2(n_443), .B(n_478), .Y(n_477) );
A2O1A1Ixp33_ASAP7_75t_L g560 ( .A1(n_76), .A2(n_443), .B(n_503), .C(n_561), .Y(n_560) );
INVx1_ASAP7_75t_L g109 ( .A(n_77), .Y(n_109) );
AND2x2_ASAP7_75t_L g148 ( .A(n_78), .B(n_149), .Y(n_148) );
NAND2xp5_ASAP7_75t_SL g168 ( .A(n_79), .B(n_123), .Y(n_168) );
AND2x2_ASAP7_75t_SL g440 ( .A(n_80), .B(n_149), .Y(n_440) );
AOI22xp5_ASAP7_75t_L g505 ( .A1(n_81), .A2(n_443), .B1(n_506), .B2(n_507), .Y(n_505) );
AOI222xp33_ASAP7_75t_L g98 ( .A1(n_82), .A2(n_99), .B1(n_775), .B2(n_786), .C1(n_802), .C2(n_806), .Y(n_98) );
OAI22xp5_ASAP7_75t_SL g788 ( .A1(n_82), .A2(n_789), .B1(n_790), .B2(n_791), .Y(n_788) );
INVx1_ASAP7_75t_L g790 ( .A(n_82), .Y(n_790) );
AND2x2_ASAP7_75t_L g198 ( .A(n_83), .B(n_143), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_85), .B(n_141), .Y(n_167) );
AND2x2_ASAP7_75t_L g192 ( .A(n_86), .B(n_149), .Y(n_192) );
INVx1_ASAP7_75t_L g449 ( .A(n_87), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_88), .B(n_139), .Y(n_210) );
AOI21xp5_ASAP7_75t_L g164 ( .A1(n_89), .A2(n_132), .B(n_165), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_90), .B(n_141), .Y(n_220) );
CKINVDCx20_ASAP7_75t_R g100 ( .A(n_91), .Y(n_100) );
AND2x2_ASAP7_75t_L g512 ( .A(n_92), .B(n_149), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_93), .B(n_139), .Y(n_155) );
A2O1A1Ixp33_ASAP7_75t_L g525 ( .A1(n_94), .A2(n_526), .B(n_527), .C(n_529), .Y(n_525) );
BUFx2_ASAP7_75t_L g783 ( .A(n_95), .Y(n_783) );
BUFx2_ASAP7_75t_SL g810 ( .A(n_95), .Y(n_810) );
AOI21xp5_ASAP7_75t_L g131 ( .A1(n_96), .A2(n_132), .B(n_137), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_97), .B(n_124), .Y(n_452) );
OAI21xp5_ASAP7_75t_L g99 ( .A1(n_100), .A2(n_101), .B(n_768), .Y(n_99) );
INVx1_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
OAI22xp5_ASAP7_75t_L g102 ( .A1(n_103), .A2(n_110), .B1(n_433), .B2(n_766), .Y(n_102) );
INVx3_ASAP7_75t_SL g771 ( .A(n_103), .Y(n_771) );
CKINVDCx5p33_ASAP7_75t_R g103 ( .A(n_104), .Y(n_103) );
AND2x6_ASAP7_75t_SL g104 ( .A(n_105), .B(n_106), .Y(n_104) );
OR2x6_ASAP7_75t_SL g766 ( .A(n_105), .B(n_767), .Y(n_766) );
OR2x2_ASAP7_75t_L g774 ( .A(n_105), .B(n_106), .Y(n_774) );
NAND2xp5_ASAP7_75t_L g785 ( .A(n_105), .B(n_767), .Y(n_785) );
CKINVDCx5p33_ASAP7_75t_R g767 ( .A(n_106), .Y(n_767) );
NAND2xp5_ASAP7_75t_L g107 ( .A(n_108), .B(n_109), .Y(n_107) );
INVx2_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
OAI22xp5_ASAP7_75t_SL g769 ( .A1(n_111), .A2(n_766), .B1(n_770), .B2(n_772), .Y(n_769) );
INVx1_ASAP7_75t_L g789 ( .A(n_111), .Y(n_789) );
INVx2_ASAP7_75t_L g792 ( .A(n_111), .Y(n_792) );
AND2x4_ASAP7_75t_L g111 ( .A(n_112), .B(n_354), .Y(n_111) );
NOR3xp33_ASAP7_75t_SL g112 ( .A(n_113), .B(n_266), .C(n_306), .Y(n_112) );
OAI221xp5_ASAP7_75t_L g113 ( .A1(n_114), .A2(n_181), .B1(n_230), .B2(n_245), .C(n_248), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
AND2x2_ASAP7_75t_L g115 ( .A(n_116), .B(n_145), .Y(n_115) );
INVx2_ASAP7_75t_L g263 ( .A(n_116), .Y(n_263) );
AND2x2_ASAP7_75t_L g293 ( .A(n_116), .B(n_294), .Y(n_293) );
BUFx3_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
AND2x2_ASAP7_75t_L g231 ( .A(n_117), .B(n_232), .Y(n_231) );
OR2x2_ASAP7_75t_L g238 ( .A(n_117), .B(n_171), .Y(n_238) );
INVx2_ASAP7_75t_L g244 ( .A(n_117), .Y(n_244) );
AND2x2_ASAP7_75t_L g253 ( .A(n_117), .B(n_147), .Y(n_253) );
INVx1_ASAP7_75t_L g269 ( .A(n_117), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_117), .B(n_315), .Y(n_314) );
OA21x2_ASAP7_75t_L g493 ( .A1(n_118), .A2(n_494), .B(n_498), .Y(n_493) );
INVx2_ASAP7_75t_SL g503 ( .A(n_118), .Y(n_503) );
BUFx4f_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVx3_ASAP7_75t_L g150 ( .A(n_119), .Y(n_150) );
AND2x4_ASAP7_75t_L g143 ( .A(n_120), .B(n_144), .Y(n_143) );
AND2x2_ASAP7_75t_SL g158 ( .A(n_120), .B(n_144), .Y(n_158) );
AOI21xp5_ASAP7_75t_L g121 ( .A1(n_122), .A2(n_131), .B(n_143), .Y(n_121) );
AND2x4_ASAP7_75t_L g123 ( .A(n_124), .B(n_129), .Y(n_123) );
INVx1_ASAP7_75t_L g467 ( .A(n_124), .Y(n_467) );
AND2x4_ASAP7_75t_L g124 ( .A(n_125), .B(n_127), .Y(n_124) );
AND2x6_ASAP7_75t_L g141 ( .A(n_125), .B(n_134), .Y(n_141) );
INVx2_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
AND2x4_ASAP7_75t_L g139 ( .A(n_127), .B(n_136), .Y(n_139) );
INVx2_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
INVx5_ASAP7_75t_L g142 ( .A(n_129), .Y(n_142) );
HB1xp67_ASAP7_75t_L g529 ( .A(n_129), .Y(n_529) );
AND2x2_ASAP7_75t_L g135 ( .A(n_130), .B(n_136), .Y(n_135) );
HB1xp67_ASAP7_75t_L g456 ( .A(n_130), .Y(n_456) );
AND2x6_ASAP7_75t_L g132 ( .A(n_133), .B(n_135), .Y(n_132) );
BUFx3_ASAP7_75t_L g457 ( .A(n_133), .Y(n_457) );
INVx2_ASAP7_75t_L g447 ( .A(n_134), .Y(n_447) );
AND2x4_ASAP7_75t_L g443 ( .A(n_135), .B(n_444), .Y(n_443) );
INVx2_ASAP7_75t_L g451 ( .A(n_136), .Y(n_451) );
AOI21xp5_ASAP7_75t_L g137 ( .A1(n_138), .A2(n_140), .B(n_142), .Y(n_137) );
INVxp67_ASAP7_75t_L g472 ( .A(n_139), .Y(n_472) );
INVxp67_ASAP7_75t_L g470 ( .A(n_141), .Y(n_470) );
AOI21xp5_ASAP7_75t_L g154 ( .A1(n_142), .A2(n_155), .B(n_156), .Y(n_154) );
AOI21xp5_ASAP7_75t_L g165 ( .A1(n_142), .A2(n_166), .B(n_167), .Y(n_165) );
AOI21xp5_ASAP7_75t_L g175 ( .A1(n_142), .A2(n_176), .B(n_177), .Y(n_175) );
AOI21xp5_ASAP7_75t_L g187 ( .A1(n_142), .A2(n_188), .B(n_189), .Y(n_187) );
AOI21xp5_ASAP7_75t_L g200 ( .A1(n_142), .A2(n_201), .B(n_202), .Y(n_200) );
AOI21xp5_ASAP7_75t_L g208 ( .A1(n_142), .A2(n_209), .B(n_210), .Y(n_208) );
AOI21xp5_ASAP7_75t_L g219 ( .A1(n_142), .A2(n_220), .B(n_221), .Y(n_219) );
O2A1O1Ixp33_ASAP7_75t_L g448 ( .A1(n_142), .A2(n_449), .B(n_450), .C(n_452), .Y(n_448) );
NOR2xp33_ASAP7_75t_L g473 ( .A(n_142), .B(n_143), .Y(n_473) );
O2A1O1Ixp33_ASAP7_75t_SL g478 ( .A1(n_142), .A2(n_450), .B(n_479), .C(n_480), .Y(n_478) );
O2A1O1Ixp33_ASAP7_75t_SL g495 ( .A1(n_142), .A2(n_450), .B(n_496), .C(n_497), .Y(n_495) );
INVx1_ASAP7_75t_L g506 ( .A(n_142), .Y(n_506) );
O2A1O1Ixp33_ASAP7_75t_L g518 ( .A1(n_142), .A2(n_450), .B(n_519), .C(n_520), .Y(n_518) );
AOI21xp5_ASAP7_75t_L g561 ( .A1(n_142), .A2(n_562), .B(n_563), .Y(n_561) );
INVx1_ASAP7_75t_SL g162 ( .A(n_143), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_143), .B(n_204), .Y(n_203) );
AOI21xp5_ASAP7_75t_L g441 ( .A1(n_143), .A2(n_442), .B(n_453), .Y(n_441) );
AND2x2_ASAP7_75t_SL g145 ( .A(n_146), .B(n_159), .Y(n_145) );
INVx4_ASAP7_75t_L g234 ( .A(n_146), .Y(n_234) );
AND2x2_ASAP7_75t_L g265 ( .A(n_146), .B(n_172), .Y(n_265) );
AND2x2_ASAP7_75t_L g341 ( .A(n_146), .B(n_315), .Y(n_341) );
NAND2x1p5_ASAP7_75t_L g383 ( .A(n_146), .B(n_171), .Y(n_383) );
INVx5_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_147), .B(n_171), .Y(n_270) );
AND2x2_ASAP7_75t_L g294 ( .A(n_147), .B(n_172), .Y(n_294) );
BUFx2_ASAP7_75t_L g310 ( .A(n_147), .Y(n_310) );
NOR2x1_ASAP7_75t_SL g413 ( .A(n_147), .B(n_315), .Y(n_413) );
OR2x6_ASAP7_75t_L g147 ( .A(n_148), .B(n_151), .Y(n_147) );
INVx3_ASAP7_75t_L g191 ( .A(n_149), .Y(n_191) );
OAI22xp5_ASAP7_75t_L g524 ( .A1(n_149), .A2(n_191), .B1(n_525), .B2(n_530), .Y(n_524) );
INVx4_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_150), .B(n_533), .Y(n_532) );
AOI21xp5_ASAP7_75t_L g151 ( .A1(n_152), .A2(n_153), .B(n_157), .Y(n_151) );
CKINVDCx5p33_ASAP7_75t_R g179 ( .A(n_157), .Y(n_179) );
OA21x2_ASAP7_75t_L g217 ( .A1(n_157), .A2(n_218), .B(n_222), .Y(n_217) );
OA21x2_ASAP7_75t_L g280 ( .A1(n_157), .A2(n_218), .B(n_222), .Y(n_280) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx2_ASAP7_75t_L g290 ( .A(n_159), .Y(n_290) );
AOI221xp5_ASAP7_75t_L g356 ( .A1(n_159), .A2(n_357), .B1(n_359), .B2(n_361), .C(n_366), .Y(n_356) );
AND2x2_ASAP7_75t_L g376 ( .A(n_159), .B(n_269), .Y(n_376) );
AND2x4_ASAP7_75t_L g159 ( .A(n_160), .B(n_171), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx2_ASAP7_75t_L g232 ( .A(n_161), .Y(n_232) );
INVx1_ASAP7_75t_L g285 ( .A(n_161), .Y(n_285) );
AO21x2_ASAP7_75t_L g161 ( .A1(n_162), .A2(n_163), .B(n_169), .Y(n_161) );
NOR2xp33_ASAP7_75t_L g169 ( .A(n_162), .B(n_170), .Y(n_169) );
AO21x2_ASAP7_75t_L g315 ( .A1(n_162), .A2(n_163), .B(n_169), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_164), .B(n_168), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_171), .B(n_242), .Y(n_241) );
AND2x2_ASAP7_75t_L g254 ( .A(n_171), .B(n_242), .Y(n_254) );
INVx2_ASAP7_75t_L g296 ( .A(n_171), .Y(n_296) );
AND2x2_ASAP7_75t_L g429 ( .A(n_171), .B(n_244), .Y(n_429) );
INVx4_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
HB1xp67_ASAP7_75t_L g286 ( .A(n_172), .Y(n_286) );
AO21x2_ASAP7_75t_L g172 ( .A1(n_173), .A2(n_179), .B(n_180), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_174), .B(n_178), .Y(n_173) );
AO21x2_ASAP7_75t_L g474 ( .A1(n_179), .A2(n_475), .B(n_481), .Y(n_474) );
NOR3xp33_ASAP7_75t_L g181 ( .A(n_182), .B(n_213), .C(n_228), .Y(n_181) );
AND2x2_ASAP7_75t_L g182 ( .A(n_183), .B(n_193), .Y(n_182) );
INVx2_ASAP7_75t_L g343 ( .A(n_183), .Y(n_343) );
AND2x2_ASAP7_75t_L g388 ( .A(n_183), .B(n_265), .Y(n_388) );
BUFx2_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
INVx1_ASAP7_75t_L g333 ( .A(n_184), .Y(n_333) );
AND2x4_ASAP7_75t_SL g348 ( .A(n_184), .B(n_260), .Y(n_348) );
AO21x2_ASAP7_75t_L g184 ( .A1(n_185), .A2(n_191), .B(n_192), .Y(n_184) );
AO21x2_ASAP7_75t_L g227 ( .A1(n_185), .A2(n_191), .B(n_192), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_186), .B(n_190), .Y(n_185) );
AO21x2_ASAP7_75t_L g205 ( .A1(n_191), .A2(n_206), .B(n_212), .Y(n_205) );
AO21x2_ASAP7_75t_L g225 ( .A1(n_191), .A2(n_206), .B(n_212), .Y(n_225) );
AO21x2_ASAP7_75t_L g514 ( .A1(n_191), .A2(n_515), .B(n_521), .Y(n_514) );
AO21x2_ASAP7_75t_L g544 ( .A1(n_191), .A2(n_515), .B(n_521), .Y(n_544) );
INVx2_ASAP7_75t_L g302 ( .A(n_193), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_193), .B(n_332), .Y(n_358) );
AND2x4_ASAP7_75t_L g391 ( .A(n_193), .B(n_338), .Y(n_391) );
AND2x4_ASAP7_75t_L g193 ( .A(n_194), .B(n_205), .Y(n_193) );
AND2x2_ASAP7_75t_L g229 ( .A(n_194), .B(n_224), .Y(n_229) );
OR2x2_ASAP7_75t_L g259 ( .A(n_194), .B(n_260), .Y(n_259) );
AND2x2_ASAP7_75t_SL g328 ( .A(n_194), .B(n_280), .Y(n_328) );
INVx2_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
BUFx2_ASAP7_75t_L g273 ( .A(n_195), .Y(n_273) );
INVx2_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
INVx2_ASAP7_75t_L g247 ( .A(n_196), .Y(n_247) );
OAI21x1_ASAP7_75t_SL g196 ( .A1(n_197), .A2(n_199), .B(n_203), .Y(n_196) );
INVx1_ASAP7_75t_L g204 ( .A(n_198), .Y(n_204) );
INVx2_ASAP7_75t_L g260 ( .A(n_205), .Y(n_260) );
NAND2xp5_ASAP7_75t_SL g206 ( .A(n_207), .B(n_211), .Y(n_206) );
NOR2xp33_ASAP7_75t_L g422 ( .A(n_213), .B(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_215), .B(n_223), .Y(n_214) );
AND2x2_ASAP7_75t_L g228 ( .A(n_215), .B(n_229), .Y(n_228) );
OR2x2_ASAP7_75t_L g301 ( .A(n_215), .B(n_302), .Y(n_301) );
INVx1_ASAP7_75t_L g386 ( .A(n_215), .Y(n_386) );
BUFx2_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
AND2x4_ASAP7_75t_L g246 ( .A(n_216), .B(n_247), .Y(n_246) );
AND2x2_ASAP7_75t_L g365 ( .A(n_216), .B(n_225), .Y(n_365) );
AND2x2_ASAP7_75t_L g369 ( .A(n_216), .B(n_235), .Y(n_369) );
INVx2_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
INVx2_ASAP7_75t_L g338 ( .A(n_217), .Y(n_338) );
HB1xp67_ASAP7_75t_L g406 ( .A(n_217), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_223), .B(n_246), .Y(n_322) );
AND2x2_ASAP7_75t_L g223 ( .A(n_224), .B(n_226), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_224), .B(n_247), .Y(n_432) );
INVx2_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
AND2x2_ASAP7_75t_L g236 ( .A(n_225), .B(n_227), .Y(n_236) );
AND2x2_ASAP7_75t_L g318 ( .A(n_225), .B(n_280), .Y(n_318) );
AND2x2_ASAP7_75t_L g337 ( .A(n_225), .B(n_226), .Y(n_337) );
BUFx2_ASAP7_75t_L g258 ( .A(n_226), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_226), .B(n_318), .Y(n_317) );
INVx2_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
BUFx3_ASAP7_75t_L g235 ( .A(n_227), .Y(n_235) );
INVxp67_ASAP7_75t_L g278 ( .A(n_227), .Y(n_278) );
INVx1_ASAP7_75t_L g251 ( .A(n_229), .Y(n_251) );
AND2x2_ASAP7_75t_L g287 ( .A(n_229), .B(n_258), .Y(n_287) );
NAND2xp33_ASAP7_75t_L g368 ( .A(n_229), .B(n_369), .Y(n_368) );
AND2x2_ASAP7_75t_L g405 ( .A(n_229), .B(n_406), .Y(n_405) );
AOI221xp5_ASAP7_75t_L g230 ( .A1(n_231), .A2(n_233), .B1(n_236), .B2(n_237), .C(n_239), .Y(n_230) );
AND2x2_ASAP7_75t_L g334 ( .A(n_231), .B(n_234), .Y(n_334) );
AND2x2_ASAP7_75t_SL g353 ( .A(n_231), .B(n_294), .Y(n_353) );
AND2x2_ASAP7_75t_L g371 ( .A(n_231), .B(n_296), .Y(n_371) );
AND2x2_ASAP7_75t_L g426 ( .A(n_231), .B(n_265), .Y(n_426) );
INVx1_ASAP7_75t_L g242 ( .A(n_232), .Y(n_242) );
HB1xp67_ASAP7_75t_L g298 ( .A(n_232), .Y(n_298) );
CKINVDCx16_ASAP7_75t_R g378 ( .A(n_233), .Y(n_378) );
AND2x4_ASAP7_75t_L g233 ( .A(n_234), .B(n_235), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_234), .B(n_244), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_234), .B(n_285), .Y(n_360) );
AND2x2_ASAP7_75t_L g327 ( .A(n_235), .B(n_328), .Y(n_327) );
INVx1_ASAP7_75t_SL g363 ( .A(n_235), .Y(n_363) );
AND2x2_ASAP7_75t_L g272 ( .A(n_236), .B(n_273), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_236), .B(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g414 ( .A(n_236), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_236), .B(n_338), .Y(n_424) );
AND2x4_ASAP7_75t_L g340 ( .A(n_237), .B(n_341), .Y(n_340) );
INVx2_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
OR2x2_ASAP7_75t_L g411 ( .A(n_238), .B(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
OR2x2_ASAP7_75t_L g240 ( .A(n_241), .B(n_243), .Y(n_240) );
OR2x2_ASAP7_75t_L g282 ( .A(n_243), .B(n_283), .Y(n_282) );
OR2x2_ASAP7_75t_L g289 ( .A(n_244), .B(n_290), .Y(n_289) );
AND2x2_ASAP7_75t_L g320 ( .A(n_244), .B(n_294), .Y(n_320) );
AND2x2_ASAP7_75t_L g394 ( .A(n_244), .B(n_315), .Y(n_394) );
INVx1_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
AND2x2_ASAP7_75t_L g342 ( .A(n_246), .B(n_343), .Y(n_342) );
OAI32xp33_ASAP7_75t_L g407 ( .A1(n_246), .A2(n_408), .A3(n_410), .B1(n_411), .B2(n_414), .Y(n_407) );
AND2x4_ASAP7_75t_L g279 ( .A(n_247), .B(n_280), .Y(n_279) );
OR2x2_ASAP7_75t_L g377 ( .A(n_247), .B(n_280), .Y(n_377) );
AOI22xp5_ASAP7_75t_L g248 ( .A1(n_249), .A2(n_252), .B1(n_255), .B2(n_261), .Y(n_248) );
INVxp67_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
O2A1O1Ixp33_ASAP7_75t_SL g366 ( .A1(n_250), .A2(n_264), .B(n_367), .C(n_368), .Y(n_366) );
HB1xp67_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
OR2x2_ASAP7_75t_L g350 ( .A(n_251), .B(n_278), .Y(n_350) );
INVx1_ASAP7_75t_SL g421 ( .A(n_252), .Y(n_421) );
AND2x4_ASAP7_75t_L g252 ( .A(n_253), .B(n_254), .Y(n_252) );
AND2x4_ASAP7_75t_L g324 ( .A(n_254), .B(n_263), .Y(n_324) );
AOI221xp5_ASAP7_75t_L g402 ( .A1(n_254), .A2(n_403), .B1(n_404), .B2(n_405), .C(n_407), .Y(n_402) );
INVx1_ASAP7_75t_SL g255 ( .A(n_256), .Y(n_255) );
OR2x2_ASAP7_75t_L g256 ( .A(n_257), .B(n_259), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
NOR2xp33_ASAP7_75t_L g330 ( .A(n_259), .B(n_331), .Y(n_330) );
INVx1_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
OAI22xp33_ASAP7_75t_L g344 ( .A1(n_262), .A2(n_292), .B1(n_345), .B2(n_346), .Y(n_344) );
OR2x2_ASAP7_75t_L g262 ( .A(n_263), .B(n_264), .Y(n_262) );
OAI211xp5_ASAP7_75t_SL g380 ( .A1(n_263), .A2(n_381), .B(n_389), .C(n_402), .Y(n_380) );
INVx2_ASAP7_75t_SL g264 ( .A(n_265), .Y(n_264) );
AND2x2_ASAP7_75t_L g300 ( .A(n_265), .B(n_269), .Y(n_300) );
OAI211xp5_ASAP7_75t_SL g266 ( .A1(n_267), .A2(n_271), .B(n_274), .C(n_303), .Y(n_266) );
OR2x2_ASAP7_75t_L g267 ( .A(n_268), .B(n_270), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
AND2x2_ASAP7_75t_L g297 ( .A(n_269), .B(n_298), .Y(n_297) );
AND2x2_ASAP7_75t_L g417 ( .A(n_269), .B(n_413), .Y(n_417) );
OAI32xp33_ASAP7_75t_L g374 ( .A1(n_270), .A2(n_375), .A3(n_377), .B1(n_378), .B2(n_379), .Y(n_374) );
INVx1_ASAP7_75t_SL g271 ( .A(n_272), .Y(n_271) );
AND2x2_ASAP7_75t_SL g364 ( .A(n_273), .B(n_365), .Y(n_364) );
AOI221xp5_ASAP7_75t_L g274 ( .A1(n_275), .A2(n_281), .B1(n_287), .B2(n_288), .C(n_291), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
NAND2xp5_ASAP7_75t_SL g276 ( .A(n_277), .B(n_279), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
OR2x2_ASAP7_75t_L g431 ( .A(n_278), .B(n_432), .Y(n_431) );
NAND2xp5_ASAP7_75t_SL g345 ( .A(n_279), .B(n_343), .Y(n_345) );
A2O1A1O1Ixp25_ASAP7_75t_L g416 ( .A1(n_279), .A2(n_348), .B(n_364), .C(n_410), .D(n_417), .Y(n_416) );
AOI31xp33_ASAP7_75t_L g418 ( .A1(n_279), .A2(n_300), .A3(n_410), .B(n_417), .Y(n_418) );
AND2x2_ASAP7_75t_L g332 ( .A(n_280), .B(n_333), .Y(n_332) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
NAND2xp5_ASAP7_75t_SL g420 ( .A(n_282), .B(n_421), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_284), .B(n_286), .Y(n_283) );
INVx2_ASAP7_75t_L g409 ( .A(n_284), .Y(n_409) );
INVx2_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
AND2x2_ASAP7_75t_L g404 ( .A(n_285), .B(n_296), .Y(n_404) );
INVx1_ASAP7_75t_L g319 ( .A(n_287), .Y(n_319) );
AND2x2_ASAP7_75t_L g304 ( .A(n_288), .B(n_305), .Y(n_304) );
INVx2_ASAP7_75t_SL g288 ( .A(n_289), .Y(n_288) );
AOI31xp33_ASAP7_75t_L g291 ( .A1(n_292), .A2(n_295), .A3(n_299), .B(n_301), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_294), .B(n_409), .Y(n_408) );
AND2x2_ASAP7_75t_L g427 ( .A(n_294), .B(n_373), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_296), .B(n_297), .Y(n_295) );
AND2x2_ASAP7_75t_L g372 ( .A(n_296), .B(n_373), .Y(n_372) );
INVx1_ASAP7_75t_L g398 ( .A(n_296), .Y(n_398) );
INVxp67_ASAP7_75t_L g367 ( .A(n_297), .Y(n_367) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
INVx2_ASAP7_75t_L g305 ( .A(n_301), .Y(n_305) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
NAND3xp33_ASAP7_75t_SL g306 ( .A(n_307), .B(n_323), .C(n_339), .Y(n_306) );
AOI22xp5_ASAP7_75t_L g307 ( .A1(n_308), .A2(n_316), .B1(n_320), .B2(n_321), .Y(n_307) );
INVxp67_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_310), .B(n_311), .Y(n_309) );
INVx2_ASAP7_75t_L g393 ( .A(n_310), .Y(n_393) );
INVx1_ASAP7_75t_SL g311 ( .A(n_312), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
INVxp67_ASAP7_75t_SL g373 ( .A(n_314), .Y(n_373) );
INVxp67_ASAP7_75t_SL g399 ( .A(n_314), .Y(n_399) );
OR2x2_ASAP7_75t_L g400 ( .A(n_314), .B(n_383), .Y(n_400) );
NAND2xp33_ASAP7_75t_L g316 ( .A(n_317), .B(n_319), .Y(n_316) );
INVx1_ASAP7_75t_L g351 ( .A(n_318), .Y(n_351) );
INVx1_ASAP7_75t_SL g321 ( .A(n_322), .Y(n_321) );
AOI22xp33_ASAP7_75t_L g323 ( .A1(n_324), .A2(n_325), .B1(n_334), .B2(n_335), .Y(n_323) );
NAND2xp5_ASAP7_75t_SL g325 ( .A(n_326), .B(n_329), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
INVx1_ASAP7_75t_SL g331 ( .A(n_332), .Y(n_331) );
AOI221xp5_ASAP7_75t_L g370 ( .A1(n_332), .A2(n_337), .B1(n_371), .B2(n_372), .C(n_374), .Y(n_370) );
INVx2_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
NAND2x1_ASAP7_75t_L g336 ( .A(n_337), .B(n_338), .Y(n_336) );
INVx1_ASAP7_75t_L g410 ( .A(n_337), .Y(n_410) );
AND2x2_ASAP7_75t_L g347 ( .A(n_338), .B(n_348), .Y(n_347) );
O2A1O1Ixp33_ASAP7_75t_SL g395 ( .A1(n_338), .A2(n_396), .B(n_400), .C(n_401), .Y(n_395) );
AOI211xp5_ASAP7_75t_L g339 ( .A1(n_340), .A2(n_342), .B(n_344), .C(n_349), .Y(n_339) );
AND2x2_ASAP7_75t_L g390 ( .A(n_343), .B(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
INVx1_ASAP7_75t_L g401 ( .A(n_348), .Y(n_401) );
AOI21xp33_ASAP7_75t_SL g349 ( .A1(n_350), .A2(n_351), .B(n_352), .Y(n_349) );
INVx2_ASAP7_75t_SL g352 ( .A(n_353), .Y(n_352) );
NOR3xp33_ASAP7_75t_L g354 ( .A(n_355), .B(n_380), .C(n_415), .Y(n_354) );
NAND2xp5_ASAP7_75t_SL g355 ( .A(n_356), .B(n_370), .Y(n_355) );
INVx1_ASAP7_75t_SL g357 ( .A(n_358), .Y(n_357) );
INVxp67_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
NAND2xp5_ASAP7_75t_SL g362 ( .A(n_363), .B(n_364), .Y(n_362) );
INVx1_ASAP7_75t_L g379 ( .A(n_364), .Y(n_379) );
INVxp67_ASAP7_75t_L g403 ( .A(n_368), .Y(n_403) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx1_ASAP7_75t_SL g387 ( .A(n_377), .Y(n_387) );
AOI22xp5_ASAP7_75t_L g381 ( .A1(n_382), .A2(n_384), .B1(n_387), .B2(n_388), .Y(n_381) );
INVx2_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
AOI21xp5_ASAP7_75t_L g389 ( .A1(n_390), .A2(n_392), .B(n_395), .Y(n_389) );
AND2x2_ASAP7_75t_L g392 ( .A(n_393), .B(n_394), .Y(n_392) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
AND2x2_ASAP7_75t_L g397 ( .A(n_398), .B(n_399), .Y(n_397) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
AND2x2_ASAP7_75t_L g428 ( .A(n_413), .B(n_429), .Y(n_428) );
OAI221xp5_ASAP7_75t_L g415 ( .A1(n_416), .A2(n_418), .B1(n_419), .B2(n_422), .C(n_425), .Y(n_415) );
INVxp67_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
OAI31xp33_ASAP7_75t_SL g425 ( .A1(n_426), .A2(n_427), .A3(n_428), .B(n_430), .Y(n_425) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g772 ( .A(n_433), .Y(n_772) );
NAND3x1_ASAP7_75t_L g433 ( .A(n_434), .B(n_653), .C(n_730), .Y(n_433) );
AND2x2_ASAP7_75t_L g434 ( .A(n_435), .B(n_605), .Y(n_434) );
NOR2xp67_ASAP7_75t_L g435 ( .A(n_436), .B(n_545), .Y(n_435) );
AOI22xp33_ASAP7_75t_L g436 ( .A1(n_437), .A2(n_482), .B1(n_489), .B2(n_538), .Y(n_436) );
OR2x2_ASAP7_75t_L g437 ( .A(n_438), .B(n_458), .Y(n_437) );
NOR2xp67_ASAP7_75t_SL g588 ( .A(n_438), .B(n_589), .Y(n_588) );
AND2x4_ASAP7_75t_L g603 ( .A(n_438), .B(n_604), .Y(n_603) );
NOR2x1_ASAP7_75t_L g620 ( .A(n_438), .B(n_621), .Y(n_620) );
AND2x4_ASAP7_75t_SL g660 ( .A(n_438), .B(n_661), .Y(n_660) );
INVx4_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
NAND2xp5_ASAP7_75t_SL g487 ( .A(n_439), .B(n_488), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_439), .B(n_566), .Y(n_565) );
INVx2_ASAP7_75t_L g595 ( .A(n_439), .Y(n_595) );
BUFx6f_ASAP7_75t_L g600 ( .A(n_439), .Y(n_600) );
AND2x2_ASAP7_75t_L g629 ( .A(n_439), .B(n_569), .Y(n_629) );
OR2x2_ASAP7_75t_L g633 ( .A(n_439), .B(n_474), .Y(n_633) );
AND2x4_ASAP7_75t_L g646 ( .A(n_439), .B(n_604), .Y(n_646) );
NOR2x1_ASAP7_75t_SL g648 ( .A(n_439), .B(n_461), .Y(n_648) );
AND2x2_ASAP7_75t_L g676 ( .A(n_439), .B(n_554), .Y(n_676) );
OR2x6_ASAP7_75t_L g439 ( .A(n_440), .B(n_441), .Y(n_439) );
INVxp67_ASAP7_75t_L g535 ( .A(n_443), .Y(n_535) );
NOR2x1p5_ASAP7_75t_L g444 ( .A(n_445), .B(n_446), .Y(n_444) );
INVx1_ASAP7_75t_L g510 ( .A(n_446), .Y(n_510) );
INVx3_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
OR2x6_ASAP7_75t_L g450 ( .A(n_447), .B(n_451), .Y(n_450) );
OAI22xp5_ASAP7_75t_L g464 ( .A1(n_450), .A2(n_465), .B1(n_466), .B2(n_467), .Y(n_464) );
INVxp67_ASAP7_75t_L g526 ( .A(n_450), .Y(n_526) );
INVx2_ASAP7_75t_L g564 ( .A(n_450), .Y(n_564) );
AND2x2_ASAP7_75t_L g455 ( .A(n_451), .B(n_456), .Y(n_455) );
INVxp33_ASAP7_75t_L g509 ( .A(n_451), .Y(n_509) );
INVx1_ASAP7_75t_L g537 ( .A(n_454), .Y(n_537) );
AND2x4_ASAP7_75t_L g454 ( .A(n_455), .B(n_457), .Y(n_454) );
INVx1_ASAP7_75t_L g557 ( .A(n_455), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_457), .Y(n_558) );
NOR2xp33_ASAP7_75t_L g643 ( .A(n_458), .B(n_644), .Y(n_643) );
INVx1_ASAP7_75t_SL g458 ( .A(n_459), .Y(n_458) );
AOI22xp5_ASAP7_75t_L g733 ( .A1(n_459), .A2(n_734), .B1(n_736), .B2(n_739), .Y(n_733) );
AND2x2_ASAP7_75t_L g459 ( .A(n_460), .B(n_474), .Y(n_459) );
INVx1_ASAP7_75t_L g488 ( .A(n_460), .Y(n_488) );
AND2x2_ASAP7_75t_L g591 ( .A(n_460), .B(n_592), .Y(n_591) );
AND2x4_ASAP7_75t_L g596 ( .A(n_460), .B(n_554), .Y(n_596) );
INVx3_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
AND2x2_ASAP7_75t_L g553 ( .A(n_461), .B(n_554), .Y(n_553) );
INVx2_ASAP7_75t_L g569 ( .A(n_461), .Y(n_569) );
AND2x2_ASAP7_75t_L g602 ( .A(n_461), .B(n_474), .Y(n_602) );
AND2x4_ASAP7_75t_L g461 ( .A(n_462), .B(n_463), .Y(n_461) );
OAI21xp5_ASAP7_75t_L g463 ( .A1(n_464), .A2(n_468), .B(n_473), .Y(n_463) );
NOR2xp33_ASAP7_75t_L g527 ( .A(n_467), .B(n_528), .Y(n_527) );
OAI22xp5_ASAP7_75t_L g468 ( .A1(n_469), .A2(n_470), .B1(n_471), .B2(n_472), .Y(n_468) );
INVx2_ASAP7_75t_L g486 ( .A(n_474), .Y(n_486) );
HB1xp67_ASAP7_75t_L g571 ( .A(n_474), .Y(n_571) );
INVx1_ASAP7_75t_L g590 ( .A(n_474), .Y(n_590) );
HB1xp67_ASAP7_75t_L g659 ( .A(n_474), .Y(n_659) );
INVx1_ASAP7_75t_L g671 ( .A(n_474), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_476), .B(n_477), .Y(n_475) );
INVx1_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
OAI31xp33_ASAP7_75t_SL g725 ( .A1(n_483), .A2(n_726), .A3(n_727), .B(n_728), .Y(n_725) );
NOR2x1_ASAP7_75t_L g483 ( .A(n_484), .B(n_487), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
OR2x2_ASAP7_75t_L g650 ( .A(n_485), .B(n_552), .Y(n_650) );
HB1xp67_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
INVx2_ASAP7_75t_L g566 ( .A(n_486), .Y(n_566) );
AND2x4_ASAP7_75t_SL g686 ( .A(n_488), .B(n_590), .Y(n_686) );
OAI21xp5_ASAP7_75t_L g606 ( .A1(n_489), .A2(n_607), .B(n_610), .Y(n_606) );
OR2x2_ASAP7_75t_L g489 ( .A(n_490), .B(n_499), .Y(n_489) );
INVx2_ASAP7_75t_L g579 ( .A(n_490), .Y(n_579) );
INVx3_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
NAND2x1p5_ASAP7_75t_L g706 ( .A(n_491), .B(n_614), .Y(n_706) );
BUFx3_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
AND2x2_ASAP7_75t_L g616 ( .A(n_492), .B(n_522), .Y(n_616) );
INVx1_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
INVxp67_ASAP7_75t_L g541 ( .A(n_493), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_493), .B(n_502), .Y(n_576) );
AND2x4_ASAP7_75t_L g586 ( .A(n_493), .B(n_587), .Y(n_586) );
AND2x2_ASAP7_75t_L g631 ( .A(n_493), .B(n_523), .Y(n_631) );
INVx2_ASAP7_75t_L g639 ( .A(n_493), .Y(n_639) );
INVx1_ASAP7_75t_L g738 ( .A(n_493), .Y(n_738) );
HB1xp67_ASAP7_75t_L g747 ( .A(n_493), .Y(n_747) );
INVx1_ASAP7_75t_L g684 ( .A(n_499), .Y(n_684) );
NAND2x1p5_ASAP7_75t_L g499 ( .A(n_500), .B(n_513), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
AND2x2_ASAP7_75t_L g540 ( .A(n_501), .B(n_541), .Y(n_540) );
AND2x4_ASAP7_75t_L g679 ( .A(n_501), .B(n_614), .Y(n_679) );
AND2x2_ASAP7_75t_L g696 ( .A(n_501), .B(n_514), .Y(n_696) );
INVx2_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_502), .B(n_544), .Y(n_719) );
AO21x2_ASAP7_75t_L g502 ( .A1(n_503), .A2(n_504), .B(n_512), .Y(n_502) );
AO21x2_ASAP7_75t_L g549 ( .A1(n_503), .A2(n_504), .B(n_512), .Y(n_549) );
NAND2xp5_ASAP7_75t_SL g504 ( .A(n_505), .B(n_511), .Y(n_504) );
INVx1_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
AND2x2_ASAP7_75t_L g642 ( .A(n_513), .B(n_540), .Y(n_642) );
AND2x2_ASAP7_75t_L g513 ( .A(n_514), .B(n_522), .Y(n_513) );
INVx2_ASAP7_75t_L g548 ( .A(n_514), .Y(n_548) );
NOR2xp67_ASAP7_75t_L g729 ( .A(n_514), .B(n_522), .Y(n_729) );
NOR2x1_ASAP7_75t_L g737 ( .A(n_514), .B(n_738), .Y(n_737) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_516), .B(n_517), .Y(n_515) );
AND2x2_ASAP7_75t_L g645 ( .A(n_522), .B(n_549), .Y(n_645) );
INVx2_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_523), .B(n_544), .Y(n_543) );
INVx1_ASAP7_75t_L g574 ( .A(n_523), .Y(n_574) );
AND2x4_ASAP7_75t_L g638 ( .A(n_523), .B(n_639), .Y(n_638) );
INVx1_ASAP7_75t_L g668 ( .A(n_523), .Y(n_668) );
OR2x2_ASAP7_75t_L g523 ( .A(n_524), .B(n_531), .Y(n_523) );
OAI22xp5_ASAP7_75t_L g531 ( .A1(n_532), .A2(n_535), .B1(n_536), .B2(n_537), .Y(n_531) );
INVx1_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
HB1xp67_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
OAI221xp5_ASAP7_75t_L g689 ( .A1(n_539), .A2(n_552), .B1(n_690), .B2(n_691), .C(n_692), .Y(n_689) );
NAND2x1p5_ASAP7_75t_L g539 ( .A(n_540), .B(n_542), .Y(n_539) );
AND2x2_ASAP7_75t_L g666 ( .A(n_540), .B(n_667), .Y(n_666) );
BUFx2_ASAP7_75t_L g709 ( .A(n_540), .Y(n_709) );
INVx2_ASAP7_75t_SL g542 ( .A(n_543), .Y(n_542) );
OR2x2_ASAP7_75t_L g652 ( .A(n_543), .B(n_576), .Y(n_652) );
INVx3_ASAP7_75t_L g614 ( .A(n_544), .Y(n_614) );
AND2x2_ASAP7_75t_L g746 ( .A(n_544), .B(n_747), .Y(n_746) );
NAND3xp33_ASAP7_75t_SL g545 ( .A(n_546), .B(n_577), .C(n_593), .Y(n_545) );
AOI22xp5_ASAP7_75t_L g546 ( .A1(n_547), .A2(n_550), .B1(n_567), .B2(n_572), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_547), .B(n_582), .Y(n_581) );
AND2x2_ASAP7_75t_L g677 ( .A(n_547), .B(n_678), .Y(n_677) );
AND2x2_ASAP7_75t_L g688 ( .A(n_547), .B(n_583), .Y(n_688) );
AND2x2_ASAP7_75t_L g758 ( .A(n_547), .B(n_631), .Y(n_758) );
AND2x4_ASAP7_75t_L g547 ( .A(n_548), .B(n_549), .Y(n_547) );
INVx2_ASAP7_75t_L g587 ( .A(n_549), .Y(n_587) );
INVx1_ASAP7_75t_L g636 ( .A(n_549), .Y(n_636) );
INVxp67_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
OAI222xp33_ASAP7_75t_L g703 ( .A1(n_551), .A2(n_704), .B1(n_705), .B2(n_707), .C1(n_708), .C2(n_710), .Y(n_703) );
OR2x2_ASAP7_75t_L g551 ( .A(n_552), .B(n_565), .Y(n_551) );
NOR2xp33_ASAP7_75t_L g578 ( .A(n_552), .B(n_579), .Y(n_578) );
NOR2x1_ASAP7_75t_L g711 ( .A(n_552), .B(n_712), .Y(n_711) );
INVx2_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
AND2x2_ASAP7_75t_L g670 ( .A(n_553), .B(n_671), .Y(n_670) );
AND2x2_ASAP7_75t_L g726 ( .A(n_553), .B(n_600), .Y(n_726) );
INVx2_ASAP7_75t_L g592 ( .A(n_554), .Y(n_592) );
INVx1_ASAP7_75t_L g604 ( .A(n_554), .Y(n_604) );
HB1xp67_ASAP7_75t_L g661 ( .A(n_554), .Y(n_661) );
AND2x2_ASAP7_75t_L g554 ( .A(n_555), .B(n_560), .Y(n_554) );
NOR3xp33_ASAP7_75t_L g556 ( .A(n_557), .B(n_558), .C(n_559), .Y(n_556) );
HB1xp67_ASAP7_75t_L g609 ( .A(n_566), .Y(n_609) );
INVx3_ASAP7_75t_L g628 ( .A(n_566), .Y(n_628) );
INVx1_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
INVx2_ASAP7_75t_L g694 ( .A(n_568), .Y(n_694) );
NAND2x1_ASAP7_75t_L g568 ( .A(n_569), .B(n_570), .Y(n_568) );
INVx1_ASAP7_75t_L g681 ( .A(n_570), .Y(n_681) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
AND2x2_ASAP7_75t_L g572 ( .A(n_573), .B(n_575), .Y(n_572) );
INVx1_ASAP7_75t_L g682 ( .A(n_573), .Y(n_682) );
INVx1_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
INVx2_ASAP7_75t_L g583 ( .A(n_574), .Y(n_583) );
AND2x2_ASAP7_75t_L g701 ( .A(n_574), .B(n_586), .Y(n_701) );
AND2x2_ASAP7_75t_L g764 ( .A(n_574), .B(n_696), .Y(n_764) );
AND2x2_ASAP7_75t_L g693 ( .A(n_575), .B(n_613), .Y(n_693) );
INVx1_ASAP7_75t_L g704 ( .A(n_575), .Y(n_704) );
AND2x2_ASAP7_75t_L g721 ( .A(n_575), .B(n_668), .Y(n_721) );
INVx2_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
AOI22xp5_ASAP7_75t_L g577 ( .A1(n_578), .A2(n_580), .B1(n_584), .B2(n_588), .Y(n_577) );
OAI21xp5_ASAP7_75t_L g593 ( .A1(n_580), .A2(n_594), .B(n_597), .Y(n_593) );
INVx1_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
AND2x2_ASAP7_75t_L g625 ( .A(n_583), .B(n_586), .Y(n_625) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
AND2x4_ASAP7_75t_L g728 ( .A(n_586), .B(n_729), .Y(n_728) );
BUFx2_ASAP7_75t_L g691 ( .A(n_589), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_590), .B(n_591), .Y(n_589) );
HB1xp67_ASAP7_75t_L g619 ( .A(n_590), .Y(n_619) );
AND2x2_ASAP7_75t_SL g599 ( .A(n_591), .B(n_600), .Y(n_599) );
INVx2_ASAP7_75t_L g664 ( .A(n_591), .Y(n_664) );
AND2x2_ASAP7_75t_L g762 ( .A(n_591), .B(n_659), .Y(n_762) );
INVx1_ASAP7_75t_L g717 ( .A(n_592), .Y(n_717) );
INVx1_ASAP7_75t_L g623 ( .A(n_594), .Y(n_623) );
AND2x2_ASAP7_75t_L g594 ( .A(n_595), .B(n_596), .Y(n_594) );
INVx1_ASAP7_75t_L g712 ( .A(n_595), .Y(n_712) );
INVx4_ASAP7_75t_L g621 ( .A(n_596), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_598), .B(n_601), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
AOI32xp33_ASAP7_75t_L g692 ( .A1(n_599), .A2(n_693), .A3(n_694), .B1(n_695), .B2(n_696), .Y(n_692) );
AND2x2_ASAP7_75t_L g687 ( .A(n_600), .B(n_602), .Y(n_687) );
O2A1O1Ixp33_ASAP7_75t_SL g750 ( .A1(n_600), .A2(n_751), .B(n_752), .C(n_754), .Y(n_750) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_602), .B(n_603), .Y(n_601) );
AND2x2_ASAP7_75t_SL g715 ( .A(n_602), .B(n_716), .Y(n_715) );
INVx1_ASAP7_75t_L g754 ( .A(n_602), .Y(n_754) );
AND2x2_ASAP7_75t_L g608 ( .A(n_603), .B(n_609), .Y(n_608) );
INVx1_ASAP7_75t_L g735 ( .A(n_603), .Y(n_735) );
AND2x2_ASAP7_75t_L g741 ( .A(n_603), .B(n_628), .Y(n_741) );
NOR3x1_ASAP7_75t_L g605 ( .A(n_606), .B(n_622), .C(n_640), .Y(n_605) );
INVx1_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_611), .B(n_617), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
OR2x2_ASAP7_75t_L g612 ( .A(n_613), .B(n_615), .Y(n_612) );
AND2x2_ASAP7_75t_L g630 ( .A(n_613), .B(n_631), .Y(n_630) );
AND2x2_ASAP7_75t_L g673 ( .A(n_613), .B(n_638), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_613), .B(n_659), .Y(n_700) );
INVx3_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
INVx2_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_619), .B(n_620), .Y(n_618) );
NOR2xp33_ASAP7_75t_L g727 ( .A(n_621), .B(n_628), .Y(n_727) );
INVx2_ASAP7_75t_L g749 ( .A(n_621), .Y(n_749) );
OAI21xp5_ASAP7_75t_L g622 ( .A1(n_623), .A2(n_624), .B(n_626), .Y(n_622) );
OAI221xp5_ASAP7_75t_L g713 ( .A1(n_623), .A2(n_714), .B1(n_718), .B2(n_720), .C(n_725), .Y(n_713) );
OAI22xp5_ASAP7_75t_L g743 ( .A1(n_624), .A2(n_744), .B1(n_745), .B2(n_748), .Y(n_743) );
INVx3_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
AOI22xp5_ASAP7_75t_L g626 ( .A1(n_627), .A2(n_630), .B1(n_632), .B2(n_634), .Y(n_626) );
AND2x2_ASAP7_75t_L g627 ( .A(n_628), .B(n_629), .Y(n_627) );
AND2x2_ASAP7_75t_L g672 ( .A(n_628), .B(n_648), .Y(n_672) );
INVx1_ASAP7_75t_L g678 ( .A(n_628), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_628), .B(n_646), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g765 ( .A(n_631), .B(n_699), .Y(n_765) );
NAND2x1_ASAP7_75t_L g748 ( .A(n_632), .B(n_749), .Y(n_748) );
INVx2_ASAP7_75t_SL g632 ( .A(n_633), .Y(n_632) );
NOR2x1_ASAP7_75t_L g663 ( .A(n_633), .B(n_664), .Y(n_663) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
OR2x2_ASAP7_75t_L g635 ( .A(n_636), .B(n_637), .Y(n_635) );
NAND2x1_ASAP7_75t_SL g751 ( .A(n_636), .B(n_638), .Y(n_751) );
NAND2xp5_ASAP7_75t_L g757 ( .A(n_636), .B(n_736), .Y(n_757) );
OR2x2_ASAP7_75t_L g718 ( .A(n_637), .B(n_719), .Y(n_718) );
INVx3_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
AND2x2_ASAP7_75t_L g753 ( .A(n_638), .B(n_679), .Y(n_753) );
NAND2xp5_ASAP7_75t_SL g640 ( .A(n_641), .B(n_647), .Y(n_640) );
OAI21xp33_ASAP7_75t_SL g641 ( .A1(n_642), .A2(n_643), .B(n_646), .Y(n_641) );
OR2x2_ASAP7_75t_L g705 ( .A(n_644), .B(n_706), .Y(n_705) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
AND2x2_ASAP7_75t_L g739 ( .A(n_645), .B(n_737), .Y(n_739) );
AND2x2_ASAP7_75t_SL g685 ( .A(n_646), .B(n_686), .Y(n_685) );
INVx2_ASAP7_75t_L g695 ( .A(n_646), .Y(n_695) );
OAI21xp33_ASAP7_75t_L g647 ( .A1(n_648), .A2(n_649), .B(n_651), .Y(n_647) );
AND2x2_ASAP7_75t_L g680 ( .A(n_648), .B(n_681), .Y(n_680) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
INVx1_ASAP7_75t_SL g651 ( .A(n_652), .Y(n_651) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_655), .B(n_697), .Y(n_654) );
NOR3xp33_ASAP7_75t_SL g655 ( .A(n_656), .B(n_674), .C(n_689), .Y(n_655) );
A2O1A1Ixp33_ASAP7_75t_L g656 ( .A1(n_657), .A2(n_662), .B(n_665), .C(n_669), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_658), .B(n_660), .Y(n_657) );
BUFx2_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
BUFx2_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
INVx1_ASAP7_75t_SL g723 ( .A(n_668), .Y(n_723) );
AND2x2_ASAP7_75t_L g736 ( .A(n_668), .B(n_737), .Y(n_736) );
OAI21xp5_ASAP7_75t_L g669 ( .A1(n_670), .A2(n_672), .B(n_673), .Y(n_669) );
INVx1_ASAP7_75t_L g744 ( .A(n_670), .Y(n_744) );
OAI21xp5_ASAP7_75t_SL g674 ( .A1(n_675), .A2(n_682), .B(n_683), .Y(n_674) );
AOI22xp5_ASAP7_75t_L g675 ( .A1(n_676), .A2(n_677), .B1(n_679), .B2(n_680), .Y(n_675) );
HB1xp67_ASAP7_75t_L g702 ( .A(n_676), .Y(n_702) );
AOI22xp5_ASAP7_75t_L g683 ( .A1(n_684), .A2(n_685), .B1(n_687), .B2(n_688), .Y(n_683) );
INVx1_ASAP7_75t_SL g690 ( .A(n_688), .Y(n_690) );
NOR2xp33_ASAP7_75t_L g734 ( .A(n_694), .B(n_735), .Y(n_734) );
OAI22xp33_ASAP7_75t_SL g760 ( .A1(n_695), .A2(n_761), .B1(n_763), .B2(n_765), .Y(n_760) );
AOI211x1_ASAP7_75t_L g697 ( .A1(n_698), .A2(n_702), .B(n_703), .C(n_713), .Y(n_697) );
AND2x2_ASAP7_75t_L g698 ( .A(n_699), .B(n_701), .Y(n_698) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
INVx1_ASAP7_75t_SL g714 ( .A(n_715), .Y(n_714) );
OAI21xp5_ASAP7_75t_L g755 ( .A1(n_715), .A2(n_756), .B(n_758), .Y(n_755) );
INVx2_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
INVx1_ASAP7_75t_L g724 ( .A(n_719), .Y(n_724) );
NOR2xp67_ASAP7_75t_L g720 ( .A(n_721), .B(n_722), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g740 ( .A(n_722), .B(n_741), .Y(n_740) );
AND2x2_ASAP7_75t_L g722 ( .A(n_723), .B(n_724), .Y(n_722) );
INVx1_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
NAND4xp25_ASAP7_75t_L g731 ( .A(n_732), .B(n_742), .C(n_755), .D(n_759), .Y(n_731) );
AND2x2_ASAP7_75t_L g732 ( .A(n_733), .B(n_740), .Y(n_732) );
NOR2xp33_ASAP7_75t_L g742 ( .A(n_743), .B(n_750), .Y(n_742) );
INVxp67_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
INVx2_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
INVx1_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
INVx1_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
INVx2_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
INVx1_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
INVx4_ASAP7_75t_SL g770 ( .A(n_771), .Y(n_770) );
INVx3_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
INVx1_ASAP7_75t_SL g775 ( .A(n_776), .Y(n_775) );
INVx1_ASAP7_75t_L g776 ( .A(n_777), .Y(n_776) );
AND2x2_ASAP7_75t_L g777 ( .A(n_778), .B(n_784), .Y(n_777) );
INVxp67_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
NAND2xp5_ASAP7_75t_SL g779 ( .A(n_780), .B(n_783), .Y(n_779) );
INVx2_ASAP7_75t_L g780 ( .A(n_781), .Y(n_780) );
OR2x2_ASAP7_75t_SL g805 ( .A(n_781), .B(n_783), .Y(n_805) );
AOI21xp5_ASAP7_75t_L g807 ( .A1(n_781), .A2(n_808), .B(n_811), .Y(n_807) );
BUFx2_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
BUFx2_ASAP7_75t_R g795 ( .A(n_785), .Y(n_795) );
BUFx3_ASAP7_75t_L g800 ( .A(n_785), .Y(n_800) );
BUFx2_ASAP7_75t_L g812 ( .A(n_785), .Y(n_812) );
INVxp67_ASAP7_75t_L g786 ( .A(n_787), .Y(n_786) );
AOI21xp5_ASAP7_75t_L g787 ( .A1(n_788), .A2(n_793), .B(n_796), .Y(n_787) );
INVx1_ASAP7_75t_L g791 ( .A(n_792), .Y(n_791) );
INVx1_ASAP7_75t_SL g793 ( .A(n_794), .Y(n_793) );
INVx1_ASAP7_75t_SL g794 ( .A(n_795), .Y(n_794) );
NOR2xp33_ASAP7_75t_SL g796 ( .A(n_797), .B(n_801), .Y(n_796) );
INVx1_ASAP7_75t_SL g797 ( .A(n_798), .Y(n_797) );
BUFx2_ASAP7_75t_L g798 ( .A(n_799), .Y(n_798) );
CKINVDCx20_ASAP7_75t_R g799 ( .A(n_800), .Y(n_799) );
CKINVDCx9p33_ASAP7_75t_R g802 ( .A(n_803), .Y(n_802) );
INVx2_ASAP7_75t_L g803 ( .A(n_804), .Y(n_803) );
INVx1_ASAP7_75t_L g804 ( .A(n_805), .Y(n_804) );
INVx1_ASAP7_75t_SL g806 ( .A(n_807), .Y(n_806) );
CKINVDCx11_ASAP7_75t_R g808 ( .A(n_809), .Y(n_808) );
CKINVDCx8_ASAP7_75t_R g809 ( .A(n_810), .Y(n_809) );
INVx2_ASAP7_75t_L g811 ( .A(n_812), .Y(n_811) );
endmodule