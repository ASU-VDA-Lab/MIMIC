module fake_aes_1900_n_600 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_17, n_63, n_14, n_10, n_15, n_56, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_51, n_29, n_43, n_7, n_40, n_27, n_39, n_600);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_51;
input n_29;
input n_43;
input n_7;
input n_40;
input n_27;
input n_39;
output n_600;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_590;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_73;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_593;
wire n_554;
wire n_447;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_72;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_69;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_446;
wire n_342;
wire n_423;
wire n_370;
wire n_589;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_70;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_75;
wire n_376;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_583;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_74;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_71;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_68;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVxp33_ASAP7_75t_SL g68 ( .A(n_38), .Y(n_68) );
INVxp67_ASAP7_75t_SL g69 ( .A(n_35), .Y(n_69) );
INVxp33_ASAP7_75t_L g70 ( .A(n_12), .Y(n_70) );
INVxp67_ASAP7_75t_SL g71 ( .A(n_11), .Y(n_71) );
INVx1_ASAP7_75t_L g72 ( .A(n_43), .Y(n_72) );
INVx2_ASAP7_75t_SL g73 ( .A(n_58), .Y(n_73) );
INVx2_ASAP7_75t_L g74 ( .A(n_37), .Y(n_74) );
INVx1_ASAP7_75t_L g75 ( .A(n_11), .Y(n_75) );
CKINVDCx20_ASAP7_75t_R g76 ( .A(n_30), .Y(n_76) );
CKINVDCx20_ASAP7_75t_R g77 ( .A(n_52), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_14), .Y(n_78) );
INVxp33_ASAP7_75t_L g79 ( .A(n_59), .Y(n_79) );
INVxp67_ASAP7_75t_SL g80 ( .A(n_9), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_21), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_10), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_25), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_24), .Y(n_84) );
CKINVDCx16_ASAP7_75t_R g85 ( .A(n_6), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_42), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_3), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_64), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_63), .Y(n_89) );
INVxp67_ASAP7_75t_SL g90 ( .A(n_36), .Y(n_90) );
CKINVDCx5p33_ASAP7_75t_R g91 ( .A(n_53), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_20), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_46), .Y(n_93) );
INVxp67_ASAP7_75t_L g94 ( .A(n_19), .Y(n_94) );
INVxp33_ASAP7_75t_SL g95 ( .A(n_34), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_6), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_62), .Y(n_97) );
CKINVDCx5p33_ASAP7_75t_R g98 ( .A(n_18), .Y(n_98) );
INVx2_ASAP7_75t_L g99 ( .A(n_49), .Y(n_99) );
INVxp67_ASAP7_75t_SL g100 ( .A(n_27), .Y(n_100) );
INVxp33_ASAP7_75t_SL g101 ( .A(n_48), .Y(n_101) );
INVx2_ASAP7_75t_SL g102 ( .A(n_47), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_15), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_26), .Y(n_104) );
CKINVDCx20_ASAP7_75t_R g105 ( .A(n_51), .Y(n_105) );
CKINVDCx20_ASAP7_75t_R g106 ( .A(n_17), .Y(n_106) );
NOR2xp67_ASAP7_75t_L g107 ( .A(n_65), .B(n_56), .Y(n_107) );
CKINVDCx20_ASAP7_75t_R g108 ( .A(n_2), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_1), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_10), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_61), .Y(n_111) );
INVxp67_ASAP7_75t_SL g112 ( .A(n_33), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_7), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_66), .Y(n_114) );
NOR2xp67_ASAP7_75t_L g115 ( .A(n_40), .B(n_29), .Y(n_115) );
INVx2_ASAP7_75t_L g116 ( .A(n_74), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_81), .Y(n_117) );
NOR2xp33_ASAP7_75t_L g118 ( .A(n_73), .B(n_0), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_81), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_83), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_83), .Y(n_121) );
CKINVDCx5p33_ASAP7_75t_R g122 ( .A(n_76), .Y(n_122) );
INVx3_ASAP7_75t_L g123 ( .A(n_84), .Y(n_123) );
NAND2xp5_ASAP7_75t_L g124 ( .A(n_73), .B(n_0), .Y(n_124) );
CKINVDCx5p33_ASAP7_75t_R g125 ( .A(n_77), .Y(n_125) );
NOR2xp33_ASAP7_75t_L g126 ( .A(n_102), .B(n_1), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_84), .Y(n_127) );
CKINVDCx5p33_ASAP7_75t_R g128 ( .A(n_105), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_86), .Y(n_129) );
NOR2xp33_ASAP7_75t_R g130 ( .A(n_91), .B(n_32), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_86), .Y(n_131) );
CKINVDCx5p33_ASAP7_75t_R g132 ( .A(n_91), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_92), .Y(n_133) );
CKINVDCx5p33_ASAP7_75t_R g134 ( .A(n_68), .Y(n_134) );
BUFx6f_ASAP7_75t_L g135 ( .A(n_74), .Y(n_135) );
BUFx2_ASAP7_75t_L g136 ( .A(n_98), .Y(n_136) );
BUFx2_ASAP7_75t_L g137 ( .A(n_98), .Y(n_137) );
NAND2xp5_ASAP7_75t_SL g138 ( .A(n_102), .B(n_2), .Y(n_138) );
INVx4_ASAP7_75t_L g139 ( .A(n_99), .Y(n_139) );
AND2x2_ASAP7_75t_L g140 ( .A(n_70), .B(n_3), .Y(n_140) );
INVx2_ASAP7_75t_L g141 ( .A(n_99), .Y(n_141) );
INVx2_ASAP7_75t_L g142 ( .A(n_92), .Y(n_142) );
CKINVDCx5p33_ASAP7_75t_R g143 ( .A(n_68), .Y(n_143) );
AND2x2_ASAP7_75t_L g144 ( .A(n_85), .B(n_4), .Y(n_144) );
HB1xp67_ASAP7_75t_L g145 ( .A(n_94), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_111), .Y(n_146) );
AND2x2_ASAP7_75t_L g147 ( .A(n_79), .B(n_4), .Y(n_147) );
AND2x4_ASAP7_75t_L g148 ( .A(n_75), .B(n_5), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_111), .Y(n_149) );
INVx2_ASAP7_75t_L g150 ( .A(n_114), .Y(n_150) );
CKINVDCx5p33_ASAP7_75t_R g151 ( .A(n_95), .Y(n_151) );
INVx6_ASAP7_75t_L g152 ( .A(n_95), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_114), .Y(n_153) );
AOI22xp5_ASAP7_75t_L g154 ( .A1(n_106), .A2(n_5), .B1(n_7), .B2(n_8), .Y(n_154) );
AND2x2_ASAP7_75t_L g155 ( .A(n_75), .B(n_82), .Y(n_155) );
BUFx6f_ASAP7_75t_L g156 ( .A(n_72), .Y(n_156) );
CKINVDCx5p33_ASAP7_75t_R g157 ( .A(n_101), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_88), .Y(n_158) );
BUFx3_ASAP7_75t_L g159 ( .A(n_156), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_148), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_148), .Y(n_161) );
NOR2xp33_ASAP7_75t_L g162 ( .A(n_152), .B(n_97), .Y(n_162) );
AND3x1_ASAP7_75t_L g163 ( .A(n_154), .B(n_82), .C(n_110), .Y(n_163) );
INVx2_ASAP7_75t_L g164 ( .A(n_135), .Y(n_164) );
AND2x2_ASAP7_75t_L g165 ( .A(n_136), .B(n_110), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_148), .Y(n_166) );
INVx2_ASAP7_75t_L g167 ( .A(n_135), .Y(n_167) );
AND2x4_ASAP7_75t_L g168 ( .A(n_155), .B(n_78), .Y(n_168) );
BUFx6f_ASAP7_75t_L g169 ( .A(n_135), .Y(n_169) );
INVx8_ASAP7_75t_L g170 ( .A(n_148), .Y(n_170) );
INVxp67_ASAP7_75t_L g171 ( .A(n_136), .Y(n_171) );
INVxp67_ASAP7_75t_L g172 ( .A(n_137), .Y(n_172) );
INVx1_ASAP7_75t_SL g173 ( .A(n_137), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_155), .Y(n_174) );
OAI22xp33_ASAP7_75t_L g175 ( .A1(n_154), .A2(n_78), .B1(n_113), .B2(n_71), .Y(n_175) );
AND2x2_ASAP7_75t_L g176 ( .A(n_145), .B(n_113), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_124), .Y(n_177) );
OR2x4_ASAP7_75t_L g178 ( .A(n_158), .B(n_96), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_124), .Y(n_179) );
BUFx2_ASAP7_75t_L g180 ( .A(n_132), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_123), .Y(n_181) );
OR2x2_ASAP7_75t_L g182 ( .A(n_140), .B(n_80), .Y(n_182) );
AND2x4_ASAP7_75t_L g183 ( .A(n_117), .B(n_87), .Y(n_183) );
INVx2_ASAP7_75t_L g184 ( .A(n_135), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_123), .Y(n_185) );
INVx2_ASAP7_75t_L g186 ( .A(n_135), .Y(n_186) );
INVx2_ASAP7_75t_L g187 ( .A(n_135), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_152), .B(n_101), .Y(n_188) );
INVx2_ASAP7_75t_L g189 ( .A(n_156), .Y(n_189) );
NAND2x1p5_ASAP7_75t_L g190 ( .A(n_147), .B(n_103), .Y(n_190) );
INVx6_ASAP7_75t_L g191 ( .A(n_139), .Y(n_191) );
CKINVDCx5p33_ASAP7_75t_R g192 ( .A(n_122), .Y(n_192) );
BUFx6f_ASAP7_75t_L g193 ( .A(n_156), .Y(n_193) );
CKINVDCx5p33_ASAP7_75t_R g194 ( .A(n_125), .Y(n_194) );
NAND3x1_ASAP7_75t_L g195 ( .A(n_144), .B(n_109), .C(n_108), .Y(n_195) );
INVx1_ASAP7_75t_L g196 ( .A(n_123), .Y(n_196) );
AND2x2_ASAP7_75t_L g197 ( .A(n_147), .B(n_100), .Y(n_197) );
OAI221xp5_ASAP7_75t_L g198 ( .A1(n_117), .A2(n_69), .B1(n_112), .B2(n_90), .C(n_104), .Y(n_198) );
NOR2x1p5_ASAP7_75t_L g199 ( .A(n_128), .B(n_89), .Y(n_199) );
NAND3x1_ASAP7_75t_L g200 ( .A(n_144), .B(n_93), .C(n_9), .Y(n_200) );
INVx2_ASAP7_75t_L g201 ( .A(n_156), .Y(n_201) );
NOR2xp33_ASAP7_75t_L g202 ( .A(n_152), .B(n_115), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_123), .Y(n_203) );
BUFx2_ASAP7_75t_L g204 ( .A(n_134), .Y(n_204) );
NAND2x1p5_ASAP7_75t_L g205 ( .A(n_140), .B(n_107), .Y(n_205) );
AND2x2_ASAP7_75t_L g206 ( .A(n_152), .B(n_8), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_142), .Y(n_207) );
NOR2xp33_ASAP7_75t_L g208 ( .A(n_152), .B(n_39), .Y(n_208) );
AND2x4_ASAP7_75t_L g209 ( .A(n_119), .B(n_12), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_142), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_142), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_158), .B(n_13), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_150), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_150), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_150), .Y(n_215) );
OR2x2_ASAP7_75t_SL g216 ( .A(n_119), .B(n_13), .Y(n_216) );
AOI22xp5_ASAP7_75t_L g217 ( .A1(n_143), .A2(n_14), .B1(n_15), .B2(n_16), .Y(n_217) );
AND2x2_ASAP7_75t_L g218 ( .A(n_120), .B(n_16), .Y(n_218) );
INVx8_ASAP7_75t_L g219 ( .A(n_151), .Y(n_219) );
OR2x2_ASAP7_75t_L g220 ( .A(n_120), .B(n_17), .Y(n_220) );
INVx1_ASAP7_75t_L g221 ( .A(n_181), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_177), .B(n_157), .Y(n_222) );
INVx3_ASAP7_75t_L g223 ( .A(n_170), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_179), .B(n_131), .Y(n_224) );
NOR3xp33_ASAP7_75t_SL g225 ( .A(n_175), .B(n_138), .C(n_118), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_209), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_209), .Y(n_227) );
INVx2_ASAP7_75t_L g228 ( .A(n_189), .Y(n_228) );
CKINVDCx5p33_ASAP7_75t_R g229 ( .A(n_192), .Y(n_229) );
NAND2x1p5_ASAP7_75t_L g230 ( .A(n_209), .B(n_218), .Y(n_230) );
INVx2_ASAP7_75t_L g231 ( .A(n_201), .Y(n_231) );
AND2x4_ASAP7_75t_L g232 ( .A(n_168), .B(n_133), .Y(n_232) );
INVx2_ASAP7_75t_SL g233 ( .A(n_170), .Y(n_233) );
INVx4_ASAP7_75t_L g234 ( .A(n_170), .Y(n_234) );
INVx1_ASAP7_75t_SL g235 ( .A(n_173), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_185), .Y(n_236) );
NAND2xp33_ASAP7_75t_R g237 ( .A(n_192), .B(n_130), .Y(n_237) );
AND2x2_ASAP7_75t_L g238 ( .A(n_197), .B(n_133), .Y(n_238) );
CKINVDCx5p33_ASAP7_75t_R g239 ( .A(n_194), .Y(n_239) );
CKINVDCx5p33_ASAP7_75t_R g240 ( .A(n_194), .Y(n_240) );
NOR2xp33_ASAP7_75t_R g241 ( .A(n_219), .B(n_126), .Y(n_241) );
BUFx3_ASAP7_75t_L g242 ( .A(n_170), .Y(n_242) );
AND2x2_ASAP7_75t_L g243 ( .A(n_197), .B(n_121), .Y(n_243) );
NAND3xp33_ASAP7_75t_L g244 ( .A(n_171), .B(n_121), .C(n_153), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_174), .Y(n_245) );
BUFx6f_ASAP7_75t_L g246 ( .A(n_193), .Y(n_246) );
BUFx2_ASAP7_75t_L g247 ( .A(n_172), .Y(n_247) );
INVx4_ASAP7_75t_L g248 ( .A(n_191), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_218), .Y(n_249) );
NAND2xp5_ASAP7_75t_SL g250 ( .A(n_188), .B(n_153), .Y(n_250) );
NOR3xp33_ASAP7_75t_SL g251 ( .A(n_198), .B(n_127), .C(n_129), .Y(n_251) );
INVxp33_ASAP7_75t_L g252 ( .A(n_180), .Y(n_252) );
BUFx2_ASAP7_75t_L g253 ( .A(n_204), .Y(n_253) );
AND3x1_ASAP7_75t_L g254 ( .A(n_217), .B(n_127), .C(n_149), .Y(n_254) );
NOR3xp33_ASAP7_75t_SL g255 ( .A(n_202), .B(n_149), .C(n_146), .Y(n_255) );
CKINVDCx8_ASAP7_75t_R g256 ( .A(n_219), .Y(n_256) );
AND2x2_ASAP7_75t_L g257 ( .A(n_168), .B(n_146), .Y(n_257) );
INVx2_ASAP7_75t_L g258 ( .A(n_201), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_220), .Y(n_259) );
BUFx3_ASAP7_75t_L g260 ( .A(n_191), .Y(n_260) );
NOR3xp33_ASAP7_75t_SL g261 ( .A(n_202), .B(n_131), .C(n_129), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_168), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_196), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_162), .B(n_139), .Y(n_264) );
BUFx2_ASAP7_75t_L g265 ( .A(n_190), .Y(n_265) );
AND2x6_ASAP7_75t_SL g266 ( .A(n_176), .B(n_18), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_162), .B(n_139), .Y(n_267) );
INVx4_ASAP7_75t_L g268 ( .A(n_191), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_183), .B(n_139), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_183), .B(n_141), .Y(n_270) );
NOR3xp33_ASAP7_75t_SL g271 ( .A(n_212), .B(n_19), .C(n_156), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_183), .B(n_141), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_203), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_165), .B(n_141), .Y(n_274) );
BUFx12f_ASAP7_75t_SL g275 ( .A(n_165), .Y(n_275) );
BUFx6f_ASAP7_75t_L g276 ( .A(n_193), .Y(n_276) );
NOR3xp33_ASAP7_75t_SL g277 ( .A(n_163), .B(n_156), .C(n_116), .Y(n_277) );
BUFx3_ASAP7_75t_L g278 ( .A(n_206), .Y(n_278) );
INVxp67_ASAP7_75t_L g279 ( .A(n_176), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_207), .Y(n_280) );
INVx2_ASAP7_75t_L g281 ( .A(n_193), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_210), .Y(n_282) );
NAND2xp5_ASAP7_75t_SL g283 ( .A(n_160), .B(n_116), .Y(n_283) );
INVx1_ASAP7_75t_SL g284 ( .A(n_219), .Y(n_284) );
BUFx6f_ASAP7_75t_L g285 ( .A(n_234), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_221), .Y(n_286) );
INVx3_ASAP7_75t_L g287 ( .A(n_234), .Y(n_287) );
INVx2_ASAP7_75t_L g288 ( .A(n_221), .Y(n_288) );
AND2x2_ASAP7_75t_L g289 ( .A(n_235), .B(n_190), .Y(n_289) );
INVx3_ASAP7_75t_L g290 ( .A(n_234), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_236), .Y(n_291) );
INVx2_ASAP7_75t_L g292 ( .A(n_236), .Y(n_292) );
AOI21xp33_ASAP7_75t_L g293 ( .A1(n_226), .A2(n_208), .B(n_166), .Y(n_293) );
INVx2_ASAP7_75t_L g294 ( .A(n_280), .Y(n_294) );
INVx3_ASAP7_75t_L g295 ( .A(n_223), .Y(n_295) );
BUFx2_ASAP7_75t_L g296 ( .A(n_242), .Y(n_296) );
INVx2_ASAP7_75t_L g297 ( .A(n_280), .Y(n_297) );
CKINVDCx11_ASAP7_75t_R g298 ( .A(n_256), .Y(n_298) );
INVx1_ASAP7_75t_SL g299 ( .A(n_242), .Y(n_299) );
BUFx3_ASAP7_75t_L g300 ( .A(n_223), .Y(n_300) );
INVx3_ASAP7_75t_L g301 ( .A(n_223), .Y(n_301) );
AND2x4_ASAP7_75t_SL g302 ( .A(n_233), .B(n_206), .Y(n_302) );
BUFx12f_ASAP7_75t_L g303 ( .A(n_253), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_224), .B(n_230), .Y(n_304) );
OR2x6_ASAP7_75t_L g305 ( .A(n_230), .B(n_219), .Y(n_305) );
AOI21xp5_ASAP7_75t_L g306 ( .A1(n_250), .A2(n_161), .B(n_208), .Y(n_306) );
AOI21xp5_ASAP7_75t_L g307 ( .A1(n_283), .A2(n_178), .B(n_182), .Y(n_307) );
AND2x4_ASAP7_75t_L g308 ( .A(n_233), .B(n_199), .Y(n_308) );
OR2x2_ASAP7_75t_SL g309 ( .A(n_256), .B(n_182), .Y(n_309) );
NAND2x1p5_ASAP7_75t_L g310 ( .A(n_227), .B(n_215), .Y(n_310) );
INVx3_ASAP7_75t_L g311 ( .A(n_248), .Y(n_311) );
OR2x6_ASAP7_75t_L g312 ( .A(n_230), .B(n_200), .Y(n_312) );
INVx4_ASAP7_75t_L g313 ( .A(n_232), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_282), .Y(n_314) );
AND2x2_ASAP7_75t_L g315 ( .A(n_238), .B(n_214), .Y(n_315) );
INVx2_ASAP7_75t_SL g316 ( .A(n_232), .Y(n_316) );
BUFx3_ASAP7_75t_L g317 ( .A(n_260), .Y(n_317) );
AOI22xp33_ASAP7_75t_L g318 ( .A1(n_278), .A2(n_205), .B1(n_213), .B2(n_211), .Y(n_318) );
OR2x2_ASAP7_75t_L g319 ( .A(n_253), .B(n_216), .Y(n_319) );
INVx2_ASAP7_75t_SL g320 ( .A(n_232), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_282), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_238), .B(n_178), .Y(n_322) );
INVx2_ASAP7_75t_SL g323 ( .A(n_265), .Y(n_323) );
AOI22xp33_ASAP7_75t_L g324 ( .A1(n_278), .A2(n_205), .B1(n_116), .B2(n_159), .Y(n_324) );
AND2x2_ASAP7_75t_L g325 ( .A(n_243), .B(n_195), .Y(n_325) );
BUFx6f_ASAP7_75t_L g326 ( .A(n_246), .Y(n_326) );
OAI22xp33_ASAP7_75t_L g327 ( .A1(n_252), .A2(n_195), .B1(n_200), .B2(n_159), .Y(n_327) );
AND2x2_ASAP7_75t_L g328 ( .A(n_243), .B(n_187), .Y(n_328) );
AND2x4_ASAP7_75t_L g329 ( .A(n_249), .B(n_22), .Y(n_329) );
BUFx2_ASAP7_75t_L g330 ( .A(n_275), .Y(n_330) );
OAI22xp5_ASAP7_75t_L g331 ( .A1(n_259), .A2(n_187), .B1(n_186), .B2(n_184), .Y(n_331) );
AOI22xp33_ASAP7_75t_L g332 ( .A1(n_262), .A2(n_186), .B1(n_184), .B2(n_167), .Y(n_332) );
INVx1_ASAP7_75t_SL g333 ( .A(n_247), .Y(n_333) );
AND2x2_ASAP7_75t_L g334 ( .A(n_257), .B(n_247), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_263), .Y(n_335) );
A2O1A1Ixp33_ASAP7_75t_L g336 ( .A1(n_306), .A2(n_261), .B(n_255), .C(n_225), .Y(n_336) );
CKINVDCx5p33_ASAP7_75t_R g337 ( .A(n_298), .Y(n_337) );
BUFx3_ASAP7_75t_L g338 ( .A(n_285), .Y(n_338) );
INVx6_ASAP7_75t_L g339 ( .A(n_285), .Y(n_339) );
OAI222xp33_ASAP7_75t_L g340 ( .A1(n_312), .A2(n_239), .B1(n_240), .B2(n_229), .C1(n_284), .C2(n_265), .Y(n_340) );
AND2x2_ASAP7_75t_L g341 ( .A(n_315), .B(n_257), .Y(n_341) );
OAI22xp33_ASAP7_75t_L g342 ( .A1(n_333), .A2(n_240), .B1(n_239), .B2(n_229), .Y(n_342) );
AOI22xp33_ASAP7_75t_L g343 ( .A1(n_312), .A2(n_275), .B1(n_222), .B2(n_279), .Y(n_343) );
OR2x2_ASAP7_75t_L g344 ( .A(n_333), .B(n_252), .Y(n_344) );
INVx2_ASAP7_75t_L g345 ( .A(n_288), .Y(n_345) );
AND2x4_ASAP7_75t_L g346 ( .A(n_305), .B(n_245), .Y(n_346) );
INVx6_ASAP7_75t_L g347 ( .A(n_285), .Y(n_347) );
BUFx3_ASAP7_75t_L g348 ( .A(n_285), .Y(n_348) );
OAI22xp33_ASAP7_75t_L g349 ( .A1(n_312), .A2(n_237), .B1(n_244), .B2(n_274), .Y(n_349) );
INVx2_ASAP7_75t_SL g350 ( .A(n_285), .Y(n_350) );
NAND2x1_ASAP7_75t_L g351 ( .A(n_294), .B(n_273), .Y(n_351) );
INVx3_ASAP7_75t_SL g352 ( .A(n_305), .Y(n_352) );
AND2x2_ASAP7_75t_L g353 ( .A(n_315), .B(n_251), .Y(n_353) );
OAI22xp5_ASAP7_75t_L g354 ( .A1(n_304), .A2(n_272), .B1(n_270), .B2(n_269), .Y(n_354) );
AND2x4_ASAP7_75t_L g355 ( .A(n_305), .B(n_277), .Y(n_355) );
BUFx2_ASAP7_75t_L g356 ( .A(n_303), .Y(n_356) );
AO31x2_ASAP7_75t_L g357 ( .A1(n_294), .A2(n_164), .A3(n_167), .B(n_264), .Y(n_357) );
AOI22xp33_ASAP7_75t_L g358 ( .A1(n_312), .A2(n_241), .B1(n_260), .B2(n_267), .Y(n_358) );
NAND3xp33_ASAP7_75t_SL g359 ( .A(n_319), .B(n_271), .C(n_266), .Y(n_359) );
AND2x2_ASAP7_75t_L g360 ( .A(n_334), .B(n_254), .Y(n_360) );
BUFx12f_ASAP7_75t_L g361 ( .A(n_303), .Y(n_361) );
NOR2xp33_ASAP7_75t_L g362 ( .A(n_319), .B(n_248), .Y(n_362) );
BUFx3_ASAP7_75t_L g363 ( .A(n_285), .Y(n_363) );
OAI22xp5_ASAP7_75t_L g364 ( .A1(n_304), .A2(n_248), .B1(n_268), .B2(n_231), .Y(n_364) );
HB1xp67_ASAP7_75t_L g365 ( .A(n_303), .Y(n_365) );
AND2x4_ASAP7_75t_L g366 ( .A(n_305), .B(n_268), .Y(n_366) );
OR2x2_ASAP7_75t_L g367 ( .A(n_334), .B(n_268), .Y(n_367) );
INVx2_ASAP7_75t_L g368 ( .A(n_345), .Y(n_368) );
INVx2_ASAP7_75t_L g369 ( .A(n_345), .Y(n_369) );
AOI221xp5_ASAP7_75t_L g370 ( .A1(n_353), .A2(n_327), .B1(n_325), .B2(n_322), .C(n_307), .Y(n_370) );
AOI22xp33_ASAP7_75t_SL g371 ( .A1(n_356), .A2(n_312), .B1(n_325), .B2(n_305), .Y(n_371) );
OAI211xp5_ASAP7_75t_L g372 ( .A1(n_343), .A2(n_318), .B(n_324), .C(n_322), .Y(n_372) );
OAI22xp33_ASAP7_75t_L g373 ( .A1(n_352), .A2(n_323), .B1(n_316), .B2(n_320), .Y(n_373) );
AOI22xp33_ASAP7_75t_L g374 ( .A1(n_359), .A2(n_289), .B1(n_329), .B2(n_308), .Y(n_374) );
BUFx3_ASAP7_75t_L g375 ( .A(n_352), .Y(n_375) );
AOI222xp33_ASAP7_75t_L g376 ( .A1(n_360), .A2(n_289), .B1(n_308), .B2(n_335), .C1(n_330), .C2(n_314), .Y(n_376) );
HB1xp67_ASAP7_75t_L g377 ( .A(n_344), .Y(n_377) );
AOI22xp33_ASAP7_75t_L g378 ( .A1(n_353), .A2(n_329), .B1(n_308), .B2(n_320), .Y(n_378) );
OAI22xp5_ASAP7_75t_L g379 ( .A1(n_352), .A2(n_309), .B1(n_294), .B2(n_297), .Y(n_379) );
AOI22xp33_ASAP7_75t_SL g380 ( .A1(n_356), .A2(n_329), .B1(n_330), .B2(n_309), .Y(n_380) );
AND2x2_ASAP7_75t_L g381 ( .A(n_341), .B(n_297), .Y(n_381) );
AOI21xp5_ASAP7_75t_L g382 ( .A1(n_336), .A2(n_293), .B(n_326), .Y(n_382) );
CKINVDCx14_ASAP7_75t_R g383 ( .A(n_337), .Y(n_383) );
INVx2_ASAP7_75t_L g384 ( .A(n_351), .Y(n_384) );
INVx1_ASAP7_75t_SL g385 ( .A(n_344), .Y(n_385) );
OAI22xp5_ASAP7_75t_L g386 ( .A1(n_354), .A2(n_297), .B1(n_321), .B2(n_314), .Y(n_386) );
OAI22xp5_ASAP7_75t_L g387 ( .A1(n_346), .A2(n_321), .B1(n_292), .B2(n_288), .Y(n_387) );
AOI22xp33_ASAP7_75t_L g388 ( .A1(n_360), .A2(n_329), .B1(n_308), .B2(n_316), .Y(n_388) );
AND2x4_ASAP7_75t_SL g389 ( .A(n_346), .B(n_313), .Y(n_389) );
AOI22xp33_ASAP7_75t_L g390 ( .A1(n_346), .A2(n_313), .B1(n_335), .B2(n_286), .Y(n_390) );
INVx2_ASAP7_75t_L g391 ( .A(n_351), .Y(n_391) );
BUFx6f_ASAP7_75t_L g392 ( .A(n_363), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_341), .Y(n_393) );
AND2x4_ASAP7_75t_L g394 ( .A(n_346), .B(n_286), .Y(n_394) );
AO21x2_ASAP7_75t_L g395 ( .A1(n_349), .A2(n_293), .B(n_291), .Y(n_395) );
AND2x2_ASAP7_75t_L g396 ( .A(n_381), .B(n_288), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_368), .Y(n_397) );
AND2x4_ASAP7_75t_L g398 ( .A(n_394), .B(n_363), .Y(n_398) );
INVx2_ASAP7_75t_L g399 ( .A(n_368), .Y(n_399) );
INVx2_ASAP7_75t_L g400 ( .A(n_368), .Y(n_400) );
OAI332xp33_ASAP7_75t_L g401 ( .A1(n_393), .A2(n_342), .A3(n_323), .B1(n_362), .B2(n_367), .B3(n_291), .C1(n_340), .C2(n_331), .Y(n_401) );
AOI22xp5_ASAP7_75t_L g402 ( .A1(n_387), .A2(n_355), .B1(n_358), .B2(n_366), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_393), .B(n_367), .Y(n_403) );
AOI221xp5_ASAP7_75t_L g404 ( .A1(n_370), .A2(n_365), .B1(n_331), .B2(n_313), .C(n_355), .Y(n_404) );
OAI211xp5_ASAP7_75t_L g405 ( .A1(n_380), .A2(n_337), .B(n_313), .C(n_296), .Y(n_405) );
BUFx3_ASAP7_75t_L g406 ( .A(n_375), .Y(n_406) );
OAI211xp5_ASAP7_75t_SL g407 ( .A1(n_376), .A2(n_299), .B(n_295), .C(n_301), .Y(n_407) );
OAI221xp5_ASAP7_75t_L g408 ( .A1(n_374), .A2(n_310), .B1(n_299), .B2(n_296), .C(n_295), .Y(n_408) );
NAND4xp25_ASAP7_75t_L g409 ( .A(n_376), .B(n_355), .C(n_328), .D(n_366), .Y(n_409) );
AND2x2_ASAP7_75t_L g410 ( .A(n_381), .B(n_292), .Y(n_410) );
AND2x2_ASAP7_75t_L g411 ( .A(n_394), .B(n_292), .Y(n_411) );
INVx2_ASAP7_75t_L g412 ( .A(n_369), .Y(n_412) );
INVx2_ASAP7_75t_L g413 ( .A(n_369), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_369), .Y(n_414) );
AOI33xp33_ASAP7_75t_L g415 ( .A1(n_385), .A2(n_328), .A3(n_302), .B1(n_164), .B2(n_366), .B3(n_332), .Y(n_415) );
AND2x2_ASAP7_75t_L g416 ( .A(n_394), .B(n_363), .Y(n_416) );
OAI221xp5_ASAP7_75t_L g417 ( .A1(n_378), .A2(n_310), .B1(n_301), .B2(n_295), .C(n_364), .Y(n_417) );
AOI211xp5_ASAP7_75t_SL g418 ( .A1(n_379), .A2(n_366), .B(n_361), .C(n_287), .Y(n_418) );
AOI211xp5_ASAP7_75t_L g419 ( .A1(n_379), .A2(n_350), .B(n_338), .C(n_348), .Y(n_419) );
OAI211xp5_ASAP7_75t_L g420 ( .A1(n_371), .A2(n_370), .B(n_388), .C(n_377), .Y(n_420) );
INVx2_ASAP7_75t_SL g421 ( .A(n_389), .Y(n_421) );
HB1xp67_ASAP7_75t_L g422 ( .A(n_385), .Y(n_422) );
AOI221xp5_ASAP7_75t_SL g423 ( .A1(n_387), .A2(n_295), .B1(n_301), .B2(n_311), .C(n_169), .Y(n_423) );
AOI22xp33_ASAP7_75t_SL g424 ( .A1(n_375), .A2(n_361), .B1(n_339), .B2(n_347), .Y(n_424) );
OR2x2_ASAP7_75t_L g425 ( .A(n_386), .B(n_350), .Y(n_425) );
INVx2_ASAP7_75t_L g426 ( .A(n_384), .Y(n_426) );
INVx2_ASAP7_75t_L g427 ( .A(n_384), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_384), .Y(n_428) );
INVxp67_ASAP7_75t_L g429 ( .A(n_375), .Y(n_429) );
INVx4_ASAP7_75t_L g430 ( .A(n_406), .Y(n_430) );
AOI33xp33_ASAP7_75t_L g431 ( .A1(n_424), .A2(n_390), .A3(n_389), .B1(n_373), .B2(n_391), .B3(n_302), .Y(n_431) );
OR2x2_ASAP7_75t_L g432 ( .A(n_422), .B(n_386), .Y(n_432) );
OR2x2_ASAP7_75t_L g433 ( .A(n_409), .B(n_391), .Y(n_433) );
AND2x2_ASAP7_75t_L g434 ( .A(n_397), .B(n_395), .Y(n_434) );
INVx2_ASAP7_75t_L g435 ( .A(n_426), .Y(n_435) );
AND2x4_ASAP7_75t_L g436 ( .A(n_428), .B(n_392), .Y(n_436) );
INVx2_ASAP7_75t_L g437 ( .A(n_426), .Y(n_437) );
INVxp67_ASAP7_75t_SL g438 ( .A(n_399), .Y(n_438) );
HB1xp67_ASAP7_75t_L g439 ( .A(n_426), .Y(n_439) );
AOI222xp33_ASAP7_75t_L g440 ( .A1(n_407), .A2(n_389), .B1(n_372), .B2(n_302), .C1(n_338), .C2(n_348), .Y(n_440) );
OAI222xp33_ASAP7_75t_L g441 ( .A1(n_402), .A2(n_383), .B1(n_382), .B2(n_310), .C1(n_395), .C2(n_287), .Y(n_441) );
INVx2_ASAP7_75t_L g442 ( .A(n_427), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_427), .Y(n_443) );
BUFx3_ASAP7_75t_L g444 ( .A(n_406), .Y(n_444) );
INVx1_ASAP7_75t_SL g445 ( .A(n_406), .Y(n_445) );
AOI22xp33_ASAP7_75t_L g446 ( .A1(n_409), .A2(n_395), .B1(n_392), .B2(n_347), .Y(n_446) );
AND2x2_ASAP7_75t_L g447 ( .A(n_414), .B(n_392), .Y(n_447) );
AOI31xp33_ASAP7_75t_L g448 ( .A1(n_418), .A2(n_392), .A3(n_347), .B(n_339), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_427), .Y(n_449) );
NOR2xp33_ASAP7_75t_L g450 ( .A(n_401), .B(n_347), .Y(n_450) );
HB1xp67_ASAP7_75t_L g451 ( .A(n_399), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_399), .B(n_392), .Y(n_452) );
AND2x2_ASAP7_75t_L g453 ( .A(n_400), .B(n_392), .Y(n_453) );
BUFx2_ASAP7_75t_L g454 ( .A(n_425), .Y(n_454) );
INVx2_ASAP7_75t_SL g455 ( .A(n_400), .Y(n_455) );
INVxp67_ASAP7_75t_SL g456 ( .A(n_400), .Y(n_456) );
INVx2_ASAP7_75t_L g457 ( .A(n_412), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_425), .Y(n_458) );
O2A1O1Ixp5_ASAP7_75t_SL g459 ( .A1(n_420), .A2(n_311), .B(n_301), .C(n_357), .Y(n_459) );
INVxp67_ASAP7_75t_SL g460 ( .A(n_412), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_413), .B(n_357), .Y(n_461) );
AND2x2_ASAP7_75t_L g462 ( .A(n_413), .B(n_357), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_396), .Y(n_463) );
INVx1_ASAP7_75t_SL g464 ( .A(n_398), .Y(n_464) );
INVx2_ASAP7_75t_L g465 ( .A(n_396), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_410), .Y(n_466) );
NOR2x1_ASAP7_75t_L g467 ( .A(n_405), .B(n_290), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_411), .B(n_339), .Y(n_468) );
NOR3xp33_ASAP7_75t_L g469 ( .A(n_401), .B(n_290), .C(n_287), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_403), .B(n_317), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_416), .B(n_23), .Y(n_471) );
INVx3_ASAP7_75t_L g472 ( .A(n_398), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_402), .B(n_317), .Y(n_473) );
NOR2xp33_ASAP7_75t_L g474 ( .A(n_450), .B(n_429), .Y(n_474) );
INVx4_ASAP7_75t_L g475 ( .A(n_430), .Y(n_475) );
INVx2_ASAP7_75t_L g476 ( .A(n_455), .Y(n_476) );
HB1xp67_ASAP7_75t_L g477 ( .A(n_451), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_463), .B(n_418), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_463), .B(n_415), .Y(n_479) );
AND2x4_ASAP7_75t_SL g480 ( .A(n_430), .B(n_398), .Y(n_480) );
OR2x2_ASAP7_75t_L g481 ( .A(n_465), .B(n_421), .Y(n_481) );
AOI22xp33_ASAP7_75t_L g482 ( .A1(n_469), .A2(n_404), .B1(n_408), .B2(n_421), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_466), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_432), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_432), .Y(n_485) );
OAI221xp5_ASAP7_75t_L g486 ( .A1(n_446), .A2(n_419), .B1(n_423), .B2(n_417), .C(n_287), .Y(n_486) );
NAND2x1p5_ASAP7_75t_L g487 ( .A(n_430), .B(n_290), .Y(n_487) );
INVx3_ASAP7_75t_L g488 ( .A(n_430), .Y(n_488) );
AOI21xp33_ASAP7_75t_L g489 ( .A1(n_440), .A2(n_423), .B(n_317), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_458), .B(n_311), .Y(n_490) );
AND2x2_ASAP7_75t_L g491 ( .A(n_468), .B(n_28), .Y(n_491) );
NOR2xp33_ASAP7_75t_L g492 ( .A(n_433), .B(n_31), .Y(n_492) );
OR2x2_ASAP7_75t_L g493 ( .A(n_464), .B(n_290), .Y(n_493) );
NOR3xp33_ASAP7_75t_L g494 ( .A(n_469), .B(n_300), .C(n_281), .Y(n_494) );
AND2x2_ASAP7_75t_L g495 ( .A(n_444), .B(n_41), .Y(n_495) );
OAI32xp33_ASAP7_75t_L g496 ( .A1(n_433), .A2(n_300), .A3(n_45), .B1(n_50), .B2(n_54), .Y(n_496) );
NOR2xp33_ASAP7_75t_L g497 ( .A(n_441), .B(n_44), .Y(n_497) );
AND2x2_ASAP7_75t_L g498 ( .A(n_444), .B(n_55), .Y(n_498) );
CKINVDCx5p33_ASAP7_75t_R g499 ( .A(n_444), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_462), .B(n_169), .Y(n_500) );
NAND2xp33_ASAP7_75t_SL g501 ( .A(n_431), .B(n_326), .Y(n_501) );
NOR2xp33_ASAP7_75t_L g502 ( .A(n_441), .B(n_57), .Y(n_502) );
NAND4xp25_ASAP7_75t_L g503 ( .A(n_446), .B(n_300), .C(n_228), .D(n_258), .Y(n_503) );
OR2x2_ASAP7_75t_L g504 ( .A(n_455), .B(n_60), .Y(n_504) );
HB1xp67_ASAP7_75t_L g505 ( .A(n_439), .Y(n_505) );
AOI22xp33_ASAP7_75t_L g506 ( .A1(n_440), .A2(n_326), .B1(n_276), .B2(n_246), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_443), .Y(n_507) );
NAND2xp33_ASAP7_75t_SL g508 ( .A(n_454), .B(n_326), .Y(n_508) );
INVx2_ASAP7_75t_L g509 ( .A(n_435), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_443), .Y(n_510) );
INVx1_ASAP7_75t_SL g511 ( .A(n_499), .Y(n_511) );
AOI22xp33_ASAP7_75t_L g512 ( .A1(n_494), .A2(n_473), .B1(n_472), .B2(n_470), .Y(n_512) );
OAI211xp5_ASAP7_75t_SL g513 ( .A1(n_482), .A2(n_467), .B(n_470), .C(n_445), .Y(n_513) );
OAI21xp5_ASAP7_75t_L g514 ( .A1(n_494), .A2(n_467), .B(n_459), .Y(n_514) );
NAND2xp67_ASAP7_75t_L g515 ( .A(n_480), .B(n_471), .Y(n_515) );
XOR2x2_ASAP7_75t_L g516 ( .A(n_475), .B(n_471), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_484), .B(n_434), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_485), .B(n_434), .Y(n_518) );
OAI22xp5_ASAP7_75t_L g519 ( .A1(n_482), .A2(n_448), .B1(n_472), .B2(n_473), .Y(n_519) );
INVx2_ASAP7_75t_L g520 ( .A(n_477), .Y(n_520) );
OAI221xp5_ASAP7_75t_L g521 ( .A1(n_501), .A2(n_448), .B1(n_461), .B2(n_460), .C(n_438), .Y(n_521) );
INVx1_ASAP7_75t_SL g522 ( .A(n_480), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_483), .Y(n_523) );
INVx1_ASAP7_75t_SL g524 ( .A(n_475), .Y(n_524) );
INVx1_ASAP7_75t_SL g525 ( .A(n_488), .Y(n_525) );
AOI21xp33_ASAP7_75t_SL g526 ( .A1(n_497), .A2(n_472), .B(n_461), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_507), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_510), .Y(n_528) );
OAI22xp33_ASAP7_75t_L g529 ( .A1(n_503), .A2(n_472), .B1(n_460), .B2(n_438), .Y(n_529) );
NAND2xp33_ASAP7_75t_L g530 ( .A(n_506), .B(n_457), .Y(n_530) );
OAI22xp5_ASAP7_75t_L g531 ( .A1(n_506), .A2(n_456), .B1(n_449), .B2(n_457), .Y(n_531) );
NOR3xp33_ASAP7_75t_L g532 ( .A(n_497), .B(n_452), .C(n_449), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_479), .B(n_447), .Y(n_533) );
AO21x1_ASAP7_75t_L g534 ( .A1(n_508), .A2(n_436), .B(n_457), .Y(n_534) );
AND2x4_ASAP7_75t_L g535 ( .A(n_488), .B(n_436), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_478), .B(n_447), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_505), .Y(n_537) );
INVx2_ASAP7_75t_L g538 ( .A(n_509), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_481), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_490), .B(n_442), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_509), .Y(n_541) );
OAI22xp5_ASAP7_75t_L g542 ( .A1(n_502), .A2(n_437), .B1(n_442), .B2(n_435), .Y(n_542) );
INVx2_ASAP7_75t_L g543 ( .A(n_476), .Y(n_543) );
AOI221xp5_ASAP7_75t_L g544 ( .A1(n_474), .A2(n_442), .B1(n_437), .B2(n_435), .C(n_453), .Y(n_544) );
INVxp67_ASAP7_75t_L g545 ( .A(n_508), .Y(n_545) );
OAI21xp33_ASAP7_75t_L g546 ( .A1(n_521), .A2(n_502), .B(n_492), .Y(n_546) );
NOR2xp33_ASAP7_75t_L g547 ( .A(n_533), .B(n_492), .Y(n_547) );
O2A1O1Ixp33_ASAP7_75t_L g548 ( .A1(n_513), .A2(n_489), .B(n_486), .C(n_496), .Y(n_548) );
NAND2xp5_ASAP7_75t_SL g549 ( .A(n_529), .B(n_487), .Y(n_549) );
INVx1_ASAP7_75t_SL g550 ( .A(n_511), .Y(n_550) );
AOI221xp5_ASAP7_75t_L g551 ( .A1(n_519), .A2(n_521), .B1(n_526), .B2(n_544), .C(n_513), .Y(n_551) );
XNOR2xp5_ASAP7_75t_L g552 ( .A(n_516), .B(n_515), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_539), .B(n_517), .Y(n_553) );
INVx2_ASAP7_75t_L g554 ( .A(n_520), .Y(n_554) );
NOR2xp33_ASAP7_75t_L g555 ( .A(n_536), .B(n_491), .Y(n_555) );
INVx1_ASAP7_75t_SL g556 ( .A(n_524), .Y(n_556) );
NOR2xp67_ASAP7_75t_SL g557 ( .A(n_514), .B(n_504), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_523), .Y(n_558) );
INVx1_ASAP7_75t_SL g559 ( .A(n_522), .Y(n_559) );
INVxp67_ASAP7_75t_L g560 ( .A(n_525), .Y(n_560) );
AOI21xp5_ASAP7_75t_L g561 ( .A1(n_529), .A2(n_498), .B(n_495), .Y(n_561) );
NOR2xp33_ASAP7_75t_L g562 ( .A(n_518), .B(n_493), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_537), .B(n_500), .Y(n_563) );
INVx1_ASAP7_75t_SL g564 ( .A(n_535), .Y(n_564) );
AO22x2_ASAP7_75t_L g565 ( .A1(n_559), .A2(n_545), .B1(n_528), .B2(n_527), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_558), .Y(n_566) );
AOI22xp33_ASAP7_75t_L g567 ( .A1(n_546), .A2(n_532), .B1(n_530), .B2(n_542), .Y(n_567) );
NAND4xp25_ASAP7_75t_L g568 ( .A(n_551), .B(n_512), .C(n_544), .D(n_531), .Y(n_568) );
INVxp67_ASAP7_75t_L g569 ( .A(n_556), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_553), .Y(n_570) );
AND2x2_ASAP7_75t_L g571 ( .A(n_564), .B(n_543), .Y(n_571) );
NAND2x1_ASAP7_75t_L g572 ( .A(n_561), .B(n_541), .Y(n_572) );
O2A1O1Ixp33_ASAP7_75t_L g573 ( .A1(n_548), .A2(n_534), .B(n_540), .C(n_538), .Y(n_573) );
AOI22xp33_ASAP7_75t_L g574 ( .A1(n_547), .A2(n_552), .B1(n_549), .B2(n_555), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_554), .Y(n_575) );
AOI22xp5_ASAP7_75t_L g576 ( .A1(n_547), .A2(n_326), .B1(n_246), .B2(n_276), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_563), .Y(n_577) );
AND2x2_ASAP7_75t_L g578 ( .A(n_571), .B(n_560), .Y(n_578) );
AOI221xp5_ASAP7_75t_L g579 ( .A1(n_568), .A2(n_573), .B1(n_574), .B2(n_565), .C(n_570), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_566), .Y(n_580) );
OR2x2_ASAP7_75t_L g581 ( .A(n_577), .B(n_562), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_568), .B(n_557), .Y(n_582) );
XOR2xp5_ASAP7_75t_L g583 ( .A(n_567), .B(n_67), .Y(n_583) );
OAI22xp5_ASAP7_75t_SL g584 ( .A1(n_575), .A2(n_276), .B1(n_574), .B2(n_552), .Y(n_584) );
NAND3xp33_ASAP7_75t_SL g585 ( .A(n_576), .B(n_572), .C(n_573), .Y(n_585) );
NOR2xp33_ASAP7_75t_L g586 ( .A(n_569), .B(n_550), .Y(n_586) );
NOR3xp33_ASAP7_75t_L g587 ( .A(n_568), .B(n_573), .C(n_551), .Y(n_587) );
NOR4xp25_ASAP7_75t_L g588 ( .A(n_574), .B(n_550), .C(n_573), .D(n_568), .Y(n_588) );
AND4x1_ASAP7_75t_L g589 ( .A(n_588), .B(n_587), .C(n_579), .D(n_582), .Y(n_589) );
INVx2_ASAP7_75t_L g590 ( .A(n_580), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_581), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_578), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_591), .Y(n_593) );
XNOR2x1_ASAP7_75t_L g594 ( .A(n_589), .B(n_583), .Y(n_594) );
NOR3xp33_ASAP7_75t_SL g595 ( .A(n_591), .B(n_584), .C(n_585), .Y(n_595) );
INVx2_ASAP7_75t_SL g596 ( .A(n_593), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_594), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_597), .B(n_592), .Y(n_598) );
AOI22xp5_ASAP7_75t_SL g599 ( .A1(n_598), .A2(n_596), .B1(n_595), .B2(n_586), .Y(n_599) );
AOI21xp33_ASAP7_75t_L g600 ( .A1(n_599), .A2(n_596), .B(n_590), .Y(n_600) );
endmodule