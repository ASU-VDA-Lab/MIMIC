module fake_netlist_6_2348_n_1196 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1196);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1196;

wire n_992;
wire n_591;
wire n_435;
wire n_1115;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_968;
wire n_909;
wire n_580;
wire n_762;
wire n_1030;
wire n_881;
wire n_875;
wire n_209;
wire n_367;
wire n_465;
wire n_680;
wire n_741;
wire n_760;
wire n_1008;
wire n_1027;
wire n_590;
wire n_625;
wire n_661;
wire n_1189;
wire n_223;
wire n_278;
wire n_1079;
wire n_341;
wire n_362;
wire n_226;
wire n_828;
wire n_208;
wire n_462;
wire n_1033;
wire n_1052;
wire n_607;
wire n_671;
wire n_726;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_1103;
wire n_933;
wire n_740;
wire n_1038;
wire n_578;
wire n_703;
wire n_1003;
wire n_365;
wire n_978;
wire n_1061;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_820;
wire n_1044;
wire n_951;
wire n_783;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_188;
wire n_1164;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_368;
wire n_575;
wire n_994;
wire n_1072;
wire n_677;
wire n_988;
wire n_969;
wire n_805;
wire n_1151;
wire n_396;
wire n_495;
wire n_1065;
wire n_815;
wire n_350;
wire n_1100;
wire n_585;
wire n_732;
wire n_974;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_874;
wire n_480;
wire n_724;
wire n_1128;
wire n_382;
wire n_673;
wire n_1020;
wire n_180;
wire n_1009;
wire n_1042;
wire n_1071;
wire n_628;
wire n_1067;
wire n_1160;
wire n_883;
wire n_557;
wire n_823;
wire n_1132;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_898;
wire n_1074;
wire n_1032;
wire n_845;
wire n_255;
wire n_807;
wire n_1036;
wire n_739;
wire n_400;
wire n_955;
wire n_284;
wire n_337;
wire n_865;
wire n_1138;
wire n_893;
wire n_214;
wire n_925;
wire n_485;
wire n_1099;
wire n_1026;
wire n_443;
wire n_1101;
wire n_246;
wire n_892;
wire n_768;
wire n_1097;
wire n_471;
wire n_289;
wire n_935;
wire n_1192;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_1130;
wire n_181;
wire n_1127;
wire n_182;
wire n_238;
wire n_1095;
wire n_573;
wire n_769;
wire n_202;
wire n_320;
wire n_639;
wire n_963;
wire n_676;
wire n_327;
wire n_794;
wire n_727;
wire n_894;
wire n_369;
wire n_1120;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_832;
wire n_353;
wire n_1187;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_230;
wire n_605;
wire n_461;
wire n_873;
wire n_383;
wire n_826;
wire n_1024;
wire n_669;
wire n_200;
wire n_447;
wire n_872;
wire n_1139;
wire n_198;
wire n_300;
wire n_718;
wire n_179;
wire n_248;
wire n_222;
wire n_517;
wire n_1018;
wire n_1172;
wire n_747;
wire n_852;
wire n_667;
wire n_229;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_1105;
wire n_621;
wire n_305;
wire n_1037;
wire n_721;
wire n_996;
wire n_750;
wire n_532;
wire n_742;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_901;
wire n_504;
wire n_923;
wire n_314;
wire n_1140;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_183;
wire n_510;
wire n_837;
wire n_836;
wire n_1015;
wire n_863;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_948;
wire n_466;
wire n_704;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1057;
wire n_1147;
wire n_360;
wire n_945;
wire n_977;
wire n_603;
wire n_1005;
wire n_991;
wire n_957;
wire n_235;
wire n_1143;
wire n_536;
wire n_895;
wire n_1126;
wire n_866;
wire n_622;
wire n_191;
wire n_340;
wire n_710;
wire n_1108;
wire n_387;
wire n_1182;
wire n_452;
wire n_658;
wire n_616;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_1119;
wire n_581;
wire n_761;
wire n_428;
wire n_785;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_987;
wire n_641;
wire n_822;
wire n_693;
wire n_1056;
wire n_631;
wire n_516;
wire n_720;
wire n_758;
wire n_842;
wire n_525;
wire n_1163;
wire n_1173;
wire n_1180;
wire n_1116;
wire n_611;
wire n_943;
wire n_1168;
wire n_491;
wire n_843;
wire n_772;
wire n_656;
wire n_989;
wire n_1174;
wire n_797;
wire n_666;
wire n_1016;
wire n_371;
wire n_795;
wire n_770;
wire n_940;
wire n_567;
wire n_899;
wire n_189;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_1035;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_197;
wire n_844;
wire n_886;
wire n_343;
wire n_953;
wire n_448;
wire n_1017;
wire n_1004;
wire n_1094;
wire n_1176;
wire n_1190;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_1022;
wire n_1083;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_930;
wire n_888;
wire n_1112;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_1181;
wire n_910;
wire n_486;
wire n_911;
wire n_381;
wire n_947;
wire n_236;
wire n_653;
wire n_887;
wire n_1117;
wire n_1087;
wire n_752;
wire n_908;
wire n_944;
wire n_713;
wire n_648;
wire n_657;
wire n_1049;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_976;
wire n_490;
wire n_803;
wire n_290;
wire n_220;
wire n_809;
wire n_1043;
wire n_1011;
wire n_224;
wire n_926;
wire n_927;
wire n_986;
wire n_839;
wire n_734;
wire n_1088;
wire n_708;
wire n_196;
wire n_919;
wire n_1081;
wire n_402;
wire n_352;
wire n_917;
wire n_668;
wire n_478;
wire n_626;
wire n_990;
wire n_574;
wire n_779;
wire n_800;
wire n_929;
wire n_460;
wire n_1084;
wire n_1171;
wire n_1104;
wire n_907;
wire n_854;
wire n_1058;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_1122;
wire n_374;
wire n_659;
wire n_709;
wire n_870;
wire n_366;
wire n_904;
wire n_777;
wire n_407;
wire n_913;
wire n_450;
wire n_808;
wire n_867;
wire n_272;
wire n_526;
wire n_1109;
wire n_921;
wire n_185;
wire n_712;
wire n_1183;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_937;
wire n_390;
wire n_473;
wire n_1193;
wire n_1148;
wire n_293;
wire n_1054;
wire n_334;
wire n_559;
wire n_370;
wire n_1161;
wire n_458;
wire n_1070;
wire n_1085;
wire n_232;
wire n_650;
wire n_998;
wire n_1046;
wire n_717;
wire n_1145;
wire n_330;
wire n_771;
wire n_1121;
wire n_1152;
wire n_470;
wire n_475;
wire n_924;
wire n_1102;
wire n_298;
wire n_492;
wire n_972;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_1149;
wire n_564;
wire n_1178;
wire n_260;
wire n_265;
wire n_313;
wire n_451;
wire n_624;
wire n_1184;
wire n_824;
wire n_962;
wire n_1073;
wire n_1000;
wire n_279;
wire n_686;
wire n_796;
wire n_1041;
wire n_252;
wire n_757;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_1195;
wire n_356;
wire n_577;
wire n_936;
wire n_184;
wire n_552;
wire n_1186;
wire n_1062;
wire n_619;
wire n_885;
wire n_455;
wire n_216;
wire n_896;
wire n_521;
wire n_363;
wire n_572;
wire n_912;
wire n_395;
wire n_813;
wire n_592;
wire n_1090;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_1156;
wire n_606;
wire n_393;
wire n_818;
wire n_984;
wire n_411;
wire n_1142;
wire n_503;
wire n_716;
wire n_623;
wire n_1048;
wire n_1123;
wire n_884;
wire n_599;
wire n_513;
wire n_855;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_916;
wire n_227;
wire n_1078;
wire n_868;
wire n_570;
wire n_731;
wire n_859;
wire n_406;
wire n_735;
wire n_483;
wire n_204;
wire n_934;
wire n_482;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_474;
wire n_261;
wire n_608;
wire n_620;
wire n_683;
wire n_811;
wire n_630;
wire n_312;
wire n_394;
wire n_878;
wire n_420;
wire n_519;
wire n_541;
wire n_512;
wire n_958;
wire n_292;
wire n_307;
wire n_469;
wire n_1137;
wire n_433;
wire n_500;
wire n_942;
wire n_792;
wire n_880;
wire n_476;
wire n_981;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_1144;
wire n_889;
wire n_357;
wire n_264;
wire n_263;
wire n_985;
wire n_589;
wire n_860;
wire n_481;
wire n_1162;
wire n_788;
wire n_819;
wire n_939;
wire n_997;
wire n_821;
wire n_325;
wire n_938;
wire n_1068;
wire n_767;
wire n_804;
wire n_329;
wire n_600;
wire n_464;
wire n_831;
wire n_802;
wire n_982;
wire n_964;
wire n_561;
wire n_477;
wire n_549;
wire n_980;
wire n_533;
wire n_954;
wire n_1075;
wire n_408;
wire n_932;
wire n_806;
wire n_864;
wire n_879;
wire n_959;
wire n_237;
wire n_584;
wire n_1110;
wire n_244;
wire n_399;
wire n_243;
wire n_979;
wire n_548;
wire n_905;
wire n_282;
wire n_436;
wire n_833;
wire n_211;
wire n_523;
wire n_707;
wire n_322;
wire n_993;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_240;
wire n_1155;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_1133;
wire n_635;
wire n_787;
wire n_1194;
wire n_311;
wire n_1064;
wire n_403;
wire n_1080;
wire n_723;
wire n_253;
wire n_634;
wire n_1051;
wire n_583;
wire n_596;
wire n_1146;
wire n_546;
wire n_562;
wire n_1141;
wire n_966;
wire n_249;
wire n_201;
wire n_386;
wire n_764;
wire n_1039;
wire n_556;
wire n_1034;
wire n_1086;
wire n_1066;
wire n_692;
wire n_733;
wire n_1158;
wire n_754;
wire n_1136;
wire n_941;
wire n_975;
wire n_1031;
wire n_487;
wire n_550;
wire n_241;
wire n_1125;
wire n_275;
wire n_553;
wire n_652;
wire n_849;
wire n_970;
wire n_1107;
wire n_560;
wire n_1014;
wire n_753;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_569;
wire n_1092;
wire n_441;
wire n_221;
wire n_882;
wire n_1060;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_1111;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_269;
wire n_193;
wire n_359;
wire n_973;
wire n_346;
wire n_1053;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_1029;
wire n_418;
wire n_1093;
wire n_618;
wire n_1055;
wire n_790;
wire n_1106;
wire n_582;
wire n_199;
wire n_1167;
wire n_266;
wire n_296;
wire n_861;
wire n_674;
wire n_857;
wire n_871;
wire n_967;
wire n_775;
wire n_922;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_1153;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_1069;
wire n_1185;
wire n_453;
wire n_612;
wire n_633;
wire n_1170;
wire n_665;
wire n_902;
wire n_333;
wire n_588;
wire n_215;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_914;
wire n_759;
wire n_1047;
wire n_1010;
wire n_355;
wire n_1165;
wire n_426;
wire n_317;
wire n_1040;
wire n_915;
wire n_632;
wire n_702;
wire n_1166;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_1131;
wire n_502;
wire n_1175;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_1006;
wire n_373;
wire n_1012;
wire n_195;
wire n_497;
wire n_285;
wire n_780;
wire n_773;
wire n_675;
wire n_920;
wire n_257;
wire n_903;
wire n_730;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_670;
wire n_286;
wire n_203;
wire n_254;
wire n_207;
wire n_834;
wire n_242;
wire n_835;
wire n_928;
wire n_690;
wire n_850;
wire n_1089;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_766;
wire n_743;
wire n_816;
wire n_1157;
wire n_335;
wire n_430;
wire n_1002;
wire n_463;
wire n_1188;
wire n_545;
wire n_489;
wire n_877;
wire n_205;
wire n_604;
wire n_848;
wire n_251;
wire n_1019;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_1096;
wire n_1063;
wire n_729;
wire n_1091;
wire n_876;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_965;
wire n_267;
wire n_438;
wire n_1124;
wire n_339;
wire n_784;
wire n_315;
wire n_515;
wire n_434;
wire n_983;
wire n_288;
wire n_427;
wire n_1059;
wire n_479;
wire n_598;
wire n_496;
wire n_422;
wire n_696;
wire n_906;
wire n_688;
wire n_722;
wire n_1077;
wire n_961;
wire n_862;
wire n_351;
wire n_869;
wire n_437;
wire n_1082;
wire n_259;
wire n_1154;
wire n_1113;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_1098;
wire n_697;
wire n_687;
wire n_364;
wire n_890;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_817;
wire n_950;
wire n_629;
wire n_388;
wire n_190;
wire n_858;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_187;
wire n_900;
wire n_897;
wire n_846;
wire n_501;
wire n_841;
wire n_956;
wire n_960;
wire n_531;
wire n_827;
wire n_1001;
wire n_361;
wire n_508;
wire n_663;
wire n_856;
wire n_1050;
wire n_379;
wire n_778;
wire n_1025;
wire n_1134;
wire n_1177;
wire n_332;
wire n_891;
wire n_336;
wire n_1150;
wire n_398;
wire n_410;
wire n_1129;
wire n_1191;
wire n_566;
wire n_554;
wire n_602;
wire n_1013;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_664;
wire n_949;
wire n_678;
wire n_192;
wire n_1007;
wire n_649;
wire n_283;

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_165),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_51),
.Y(n_180)
);

CKINVDCx14_ASAP7_75t_R g181 ( 
.A(n_67),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_95),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_83),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_152),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_37),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_172),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_92),
.Y(n_187)
);

BUFx2_ASAP7_75t_SL g188 ( 
.A(n_94),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_127),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_3),
.Y(n_190)
);

BUFx3_ASAP7_75t_L g191 ( 
.A(n_99),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_54),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_60),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_70),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_23),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_12),
.Y(n_196)
);

BUFx3_ASAP7_75t_L g197 ( 
.A(n_58),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_12),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_120),
.Y(n_199)
);

INVx1_ASAP7_75t_SL g200 ( 
.A(n_77),
.Y(n_200)
);

HB1xp67_ASAP7_75t_L g201 ( 
.A(n_0),
.Y(n_201)
);

BUFx3_ASAP7_75t_L g202 ( 
.A(n_143),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_114),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_90),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_89),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_65),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_105),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_128),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_39),
.Y(n_209)
);

BUFx10_ASAP7_75t_L g210 ( 
.A(n_170),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_100),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_111),
.Y(n_212)
);

BUFx5_ASAP7_75t_L g213 ( 
.A(n_118),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_55),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_173),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_141),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_3),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_32),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_26),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_168),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_26),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_61),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_43),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_1),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_49),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_101),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_82),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_146),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_79),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_16),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_30),
.Y(n_231)
);

INVx2_ASAP7_75t_SL g232 ( 
.A(n_86),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_102),
.Y(n_233)
);

BUFx3_ASAP7_75t_L g234 ( 
.A(n_27),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_14),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_167),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_234),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_179),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_180),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_201),
.Y(n_240)
);

BUFx3_ASAP7_75t_L g241 ( 
.A(n_191),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_183),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_185),
.Y(n_243)
);

BUFx3_ASAP7_75t_L g244 ( 
.A(n_191),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_186),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_234),
.Y(n_246)
);

HB1xp67_ASAP7_75t_L g247 ( 
.A(n_190),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_189),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_194),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_195),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_224),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_213),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_199),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_204),
.Y(n_254)
);

INVxp67_ASAP7_75t_SL g255 ( 
.A(n_197),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_205),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_207),
.Y(n_257)
);

BUFx6f_ASAP7_75t_L g258 ( 
.A(n_214),
.Y(n_258)
);

BUFx10_ASAP7_75t_L g259 ( 
.A(n_214),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_209),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_230),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_211),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_226),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_228),
.Y(n_264)
);

CKINVDCx14_ASAP7_75t_R g265 ( 
.A(n_181),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_182),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_237),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_258),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_237),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_266),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_258),
.Y(n_271)
);

NOR2xp67_ASAP7_75t_L g272 ( 
.A(n_238),
.B(n_208),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_239),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_246),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_242),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_246),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_250),
.Y(n_277)
);

INVxp33_ASAP7_75t_SL g278 ( 
.A(n_243),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_245),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_248),
.Y(n_280)
);

INVx1_ASAP7_75t_SL g281 ( 
.A(n_249),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_250),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_251),
.Y(n_283)
);

INVx4_ASAP7_75t_R g284 ( 
.A(n_241),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_253),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_254),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_251),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_261),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_261),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_259),
.Y(n_290)
);

HB1xp67_ASAP7_75t_L g291 ( 
.A(n_247),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_259),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_259),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_259),
.Y(n_294)
);

OR2x2_ASAP7_75t_L g295 ( 
.A(n_244),
.B(n_231),
.Y(n_295)
);

BUFx3_ASAP7_75t_L g296 ( 
.A(n_244),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_244),
.Y(n_297)
);

HB1xp67_ASAP7_75t_L g298 ( 
.A(n_256),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_241),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_257),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_260),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_262),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_255),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_258),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_263),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_264),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_265),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_240),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_258),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_258),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_258),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_252),
.Y(n_312)
);

HB1xp67_ASAP7_75t_L g313 ( 
.A(n_252),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_266),
.Y(n_314)
);

BUFx3_ASAP7_75t_L g315 ( 
.A(n_244),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_258),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_266),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_270),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_313),
.Y(n_319)
);

BUFx6f_ASAP7_75t_L g320 ( 
.A(n_271),
.Y(n_320)
);

INVxp67_ASAP7_75t_SL g321 ( 
.A(n_296),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_312),
.Y(n_322)
);

INVxp33_ASAP7_75t_L g323 ( 
.A(n_291),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_267),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_317),
.Y(n_325)
);

INVxp67_ASAP7_75t_SL g326 ( 
.A(n_296),
.Y(n_326)
);

INVxp67_ASAP7_75t_SL g327 ( 
.A(n_315),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_286),
.Y(n_328)
);

INVx1_ASAP7_75t_SL g329 ( 
.A(n_270),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_269),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_274),
.Y(n_331)
);

INVx2_ASAP7_75t_SL g332 ( 
.A(n_315),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_268),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_276),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_277),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_268),
.Y(n_336)
);

INVxp67_ASAP7_75t_SL g337 ( 
.A(n_297),
.Y(n_337)
);

INVxp33_ASAP7_75t_L g338 ( 
.A(n_295),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_301),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_287),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_R g341 ( 
.A(n_307),
.B(n_181),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_288),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_289),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_314),
.Y(n_344)
);

BUFx3_ASAP7_75t_L g345 ( 
.A(n_299),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_282),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_282),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_283),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_283),
.Y(n_349)
);

INVxp67_ASAP7_75t_SL g350 ( 
.A(n_271),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_295),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_304),
.Y(n_352)
);

BUFx6f_ASAP7_75t_L g353 ( 
.A(n_271),
.Y(n_353)
);

NOR2xp67_ASAP7_75t_L g354 ( 
.A(n_273),
.B(n_232),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_314),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_309),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_316),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_316),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_271),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_273),
.Y(n_360)
);

HB1xp67_ASAP7_75t_L g361 ( 
.A(n_308),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_303),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_310),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_307),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_310),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_290),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_325),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_338),
.B(n_278),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_324),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_324),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_330),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_328),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_330),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_339),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_360),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_323),
.B(n_281),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_319),
.B(n_275),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_331),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_355),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_333),
.Y(n_380)
);

BUFx2_ASAP7_75t_L g381 ( 
.A(n_361),
.Y(n_381)
);

NOR2xp67_ASAP7_75t_L g382 ( 
.A(n_364),
.B(n_275),
.Y(n_382)
);

HB1xp67_ASAP7_75t_L g383 ( 
.A(n_351),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_319),
.B(n_279),
.Y(n_384)
);

HB1xp67_ASAP7_75t_L g385 ( 
.A(n_332),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_331),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_343),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_343),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_346),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_318),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_347),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_318),
.Y(n_392)
);

CKINVDCx16_ASAP7_75t_R g393 ( 
.A(n_341),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_348),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_344),
.Y(n_395)
);

BUFx6f_ASAP7_75t_SL g396 ( 
.A(n_366),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_344),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_349),
.Y(n_398)
);

HB1xp67_ASAP7_75t_L g399 ( 
.A(n_332),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_335),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_364),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_329),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_362),
.B(n_279),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_345),
.Y(n_404)
);

INVxp67_ASAP7_75t_L g405 ( 
.A(n_345),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_362),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_321),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_326),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_327),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_340),
.Y(n_410)
);

CKINVDCx16_ASAP7_75t_R g411 ( 
.A(n_342),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_389),
.Y(n_412)
);

AND2x4_ASAP7_75t_L g413 ( 
.A(n_400),
.B(n_337),
.Y(n_413)
);

BUFx6f_ASAP7_75t_L g414 ( 
.A(n_369),
.Y(n_414)
);

BUFx2_ASAP7_75t_L g415 ( 
.A(n_406),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_380),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_380),
.Y(n_417)
);

AND2x4_ASAP7_75t_L g418 ( 
.A(n_391),
.B(n_334),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_370),
.Y(n_419)
);

AND2x4_ASAP7_75t_L g420 ( 
.A(n_394),
.B(n_322),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_398),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_371),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_SL g423 ( 
.A(n_403),
.B(n_363),
.Y(n_423)
);

AND2x2_ASAP7_75t_L g424 ( 
.A(n_373),
.B(n_378),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_386),
.Y(n_425)
);

INVx2_ASAP7_75t_SL g426 ( 
.A(n_385),
.Y(n_426)
);

INVx6_ASAP7_75t_L g427 ( 
.A(n_393),
.Y(n_427)
);

BUFx6f_ASAP7_75t_L g428 ( 
.A(n_387),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_388),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_383),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_399),
.B(n_363),
.Y(n_431)
);

BUFx2_ASAP7_75t_L g432 ( 
.A(n_381),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_405),
.Y(n_433)
);

BUFx3_ASAP7_75t_L g434 ( 
.A(n_404),
.Y(n_434)
);

BUFx2_ASAP7_75t_L g435 ( 
.A(n_381),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_410),
.Y(n_436)
);

INVx3_ASAP7_75t_L g437 ( 
.A(n_410),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_407),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_407),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_408),
.Y(n_440)
);

OAI22x1_ASAP7_75t_L g441 ( 
.A1(n_392),
.A2(n_308),
.B1(n_285),
.B2(n_300),
.Y(n_441)
);

OA21x2_ASAP7_75t_L g442 ( 
.A1(n_377),
.A2(n_356),
.B(n_352),
.Y(n_442)
);

AND2x2_ASAP7_75t_L g443 ( 
.A(n_376),
.B(n_365),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_408),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_409),
.B(n_365),
.Y(n_445)
);

AND2x4_ASAP7_75t_L g446 ( 
.A(n_409),
.B(n_322),
.Y(n_446)
);

AND2x2_ASAP7_75t_L g447 ( 
.A(n_384),
.B(n_298),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_396),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_396),
.Y(n_449)
);

INVx3_ASAP7_75t_L g450 ( 
.A(n_411),
.Y(n_450)
);

INVxp67_ASAP7_75t_L g451 ( 
.A(n_368),
.Y(n_451)
);

AOI22xp5_ASAP7_75t_SL g452 ( 
.A1(n_402),
.A2(n_235),
.B1(n_187),
.B2(n_206),
.Y(n_452)
);

INVxp67_ASAP7_75t_L g453 ( 
.A(n_396),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_382),
.B(n_354),
.Y(n_454)
);

INVx2_ASAP7_75t_SL g455 ( 
.A(n_392),
.Y(n_455)
);

BUFx6f_ASAP7_75t_L g456 ( 
.A(n_401),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_395),
.B(n_272),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_395),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_397),
.B(n_280),
.Y(n_459)
);

OA21x2_ASAP7_75t_L g460 ( 
.A1(n_397),
.A2(n_356),
.B(n_352),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_401),
.B(n_280),
.Y(n_461)
);

AOI22xp5_ASAP7_75t_L g462 ( 
.A1(n_390),
.A2(n_302),
.B1(n_305),
.B2(n_306),
.Y(n_462)
);

INVx3_ASAP7_75t_L g463 ( 
.A(n_367),
.Y(n_463)
);

BUFx6f_ASAP7_75t_L g464 ( 
.A(n_367),
.Y(n_464)
);

INVx4_ASAP7_75t_L g465 ( 
.A(n_374),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_374),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_372),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_375),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_379),
.Y(n_469)
);

AND2x4_ASAP7_75t_L g470 ( 
.A(n_400),
.B(n_359),
.Y(n_470)
);

OAI22xp5_ASAP7_75t_L g471 ( 
.A1(n_403),
.A2(n_182),
.B1(n_233),
.B2(n_220),
.Y(n_471)
);

AND2x4_ASAP7_75t_L g472 ( 
.A(n_400),
.B(n_359),
.Y(n_472)
);

OR2x2_ASAP7_75t_L g473 ( 
.A(n_411),
.B(n_285),
.Y(n_473)
);

CKINVDCx8_ASAP7_75t_R g474 ( 
.A(n_392),
.Y(n_474)
);

BUFx3_ASAP7_75t_L g475 ( 
.A(n_404),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_389),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_389),
.Y(n_477)
);

BUFx6f_ASAP7_75t_L g478 ( 
.A(n_369),
.Y(n_478)
);

BUFx6f_ASAP7_75t_L g479 ( 
.A(n_369),
.Y(n_479)
);

AND2x6_ASAP7_75t_L g480 ( 
.A(n_369),
.B(n_184),
.Y(n_480)
);

OAI21x1_ASAP7_75t_L g481 ( 
.A1(n_380),
.A2(n_358),
.B(n_357),
.Y(n_481)
);

AND2x4_ASAP7_75t_L g482 ( 
.A(n_400),
.B(n_333),
.Y(n_482)
);

AND2x4_ASAP7_75t_L g483 ( 
.A(n_400),
.B(n_336),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_369),
.B(n_300),
.Y(n_484)
);

AND2x4_ASAP7_75t_L g485 ( 
.A(n_400),
.B(n_197),
.Y(n_485)
);

CKINVDCx6p67_ASAP7_75t_R g486 ( 
.A(n_375),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_389),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_369),
.B(n_302),
.Y(n_488)
);

BUFx2_ASAP7_75t_L g489 ( 
.A(n_406),
.Y(n_489)
);

BUFx6f_ASAP7_75t_L g490 ( 
.A(n_369),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_392),
.Y(n_491)
);

HB1xp67_ASAP7_75t_L g492 ( 
.A(n_381),
.Y(n_492)
);

BUFx6f_ASAP7_75t_L g493 ( 
.A(n_369),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_380),
.Y(n_494)
);

OAI22xp5_ASAP7_75t_SL g495 ( 
.A1(n_390),
.A2(n_235),
.B1(n_187),
.B2(n_233),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_389),
.Y(n_496)
);

AND2x2_ASAP7_75t_L g497 ( 
.A(n_403),
.B(n_305),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_389),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_416),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_443),
.B(n_306),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_416),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_443),
.B(n_350),
.Y(n_502)
);

BUFx2_ASAP7_75t_L g503 ( 
.A(n_432),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_424),
.B(n_292),
.Y(n_504)
);

HB1xp67_ASAP7_75t_L g505 ( 
.A(n_432),
.Y(n_505)
);

HB1xp67_ASAP7_75t_L g506 ( 
.A(n_435),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_419),
.B(n_293),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_417),
.Y(n_508)
);

BUFx2_ASAP7_75t_L g509 ( 
.A(n_435),
.Y(n_509)
);

OAI21x1_ASAP7_75t_L g510 ( 
.A1(n_481),
.A2(n_236),
.B(n_184),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_SL g511 ( 
.A(n_414),
.B(n_206),
.Y(n_511)
);

INVx4_ASAP7_75t_L g512 ( 
.A(n_414),
.Y(n_512)
);

AND2x4_ASAP7_75t_L g513 ( 
.A(n_418),
.B(n_36),
.Y(n_513)
);

AND2x4_ASAP7_75t_L g514 ( 
.A(n_418),
.B(n_38),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_494),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_419),
.B(n_422),
.Y(n_516)
);

AND2x2_ASAP7_75t_L g517 ( 
.A(n_422),
.B(n_425),
.Y(n_517)
);

BUFx6f_ASAP7_75t_L g518 ( 
.A(n_414),
.Y(n_518)
);

AND2x2_ASAP7_75t_L g519 ( 
.A(n_425),
.B(n_294),
.Y(n_519)
);

AND2x2_ASAP7_75t_L g520 ( 
.A(n_429),
.B(n_192),
.Y(n_520)
);

INVx3_ASAP7_75t_L g521 ( 
.A(n_414),
.Y(n_521)
);

BUFx2_ASAP7_75t_L g522 ( 
.A(n_492),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_423),
.B(n_428),
.Y(n_523)
);

AND2x2_ASAP7_75t_L g524 ( 
.A(n_447),
.B(n_193),
.Y(n_524)
);

OAI22xp5_ASAP7_75t_SL g525 ( 
.A1(n_495),
.A2(n_220),
.B1(n_196),
.B2(n_198),
.Y(n_525)
);

INVx3_ASAP7_75t_L g526 ( 
.A(n_428),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_SL g527 ( 
.A(n_428),
.B(n_311),
.Y(n_527)
);

CKINVDCx20_ASAP7_75t_R g528 ( 
.A(n_486),
.Y(n_528)
);

INVx3_ASAP7_75t_L g529 ( 
.A(n_478),
.Y(n_529)
);

AND2x2_ASAP7_75t_L g530 ( 
.A(n_447),
.B(n_203),
.Y(n_530)
);

BUFx2_ASAP7_75t_L g531 ( 
.A(n_415),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_SL g532 ( 
.A(n_478),
.B(n_320),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_500),
.B(n_451),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_500),
.B(n_497),
.Y(n_534)
);

AND2x2_ASAP7_75t_L g535 ( 
.A(n_524),
.B(n_436),
.Y(n_535)
);

AND2x2_ASAP7_75t_L g536 ( 
.A(n_524),
.B(n_436),
.Y(n_536)
);

OAI22xp33_ASAP7_75t_SL g537 ( 
.A1(n_511),
.A2(n_471),
.B1(n_423),
.B2(n_437),
.Y(n_537)
);

AO22x2_ASAP7_75t_L g538 ( 
.A1(n_511),
.A2(n_497),
.B1(n_437),
.B2(n_466),
.Y(n_538)
);

AOI22x1_ASAP7_75t_SL g539 ( 
.A1(n_528),
.A2(n_491),
.B1(n_468),
.B2(n_463),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_L g540 ( 
.A(n_505),
.B(n_445),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_517),
.Y(n_541)
);

AND2x2_ASAP7_75t_L g542 ( 
.A(n_524),
.B(n_439),
.Y(n_542)
);

AND2x2_ASAP7_75t_L g543 ( 
.A(n_530),
.B(n_439),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_SL g544 ( 
.A(n_523),
.B(n_478),
.Y(n_544)
);

BUFx10_ASAP7_75t_L g545 ( 
.A(n_513),
.Y(n_545)
);

AO22x2_ASAP7_75t_L g546 ( 
.A1(n_523),
.A2(n_437),
.B1(n_458),
.B2(n_463),
.Y(n_546)
);

INVx3_ASAP7_75t_L g547 ( 
.A(n_512),
.Y(n_547)
);

OAI22xp33_ASAP7_75t_L g548 ( 
.A1(n_504),
.A2(n_431),
.B1(n_502),
.B2(n_458),
.Y(n_548)
);

OAI22xp5_ASAP7_75t_SL g549 ( 
.A1(n_525),
.A2(n_491),
.B1(n_459),
.B2(n_461),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_515),
.Y(n_550)
);

AND2x2_ASAP7_75t_SL g551 ( 
.A(n_513),
.B(n_514),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_516),
.Y(n_552)
);

OAI22xp33_ASAP7_75t_SL g553 ( 
.A1(n_504),
.A2(n_488),
.B1(n_484),
.B2(n_440),
.Y(n_553)
);

INVxp33_ASAP7_75t_L g554 ( 
.A(n_505),
.Y(n_554)
);

AOI22xp5_ASAP7_75t_L g555 ( 
.A1(n_525),
.A2(n_462),
.B1(n_455),
.B2(n_473),
.Y(n_555)
);

OA22x2_ASAP7_75t_L g556 ( 
.A1(n_506),
.A2(n_509),
.B1(n_503),
.B2(n_522),
.Y(n_556)
);

AOI22xp5_ASAP7_75t_L g557 ( 
.A1(n_513),
.A2(n_455),
.B1(n_473),
.B2(n_450),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_516),
.Y(n_558)
);

NOR2xp33_ASAP7_75t_L g559 ( 
.A(n_506),
.B(n_438),
.Y(n_559)
);

AOI22xp5_ASAP7_75t_L g560 ( 
.A1(n_513),
.A2(n_450),
.B1(n_463),
.B2(n_441),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_499),
.Y(n_561)
);

AND2x2_ASAP7_75t_L g562 ( 
.A(n_530),
.B(n_444),
.Y(n_562)
);

AND2x2_ASAP7_75t_L g563 ( 
.A(n_530),
.B(n_446),
.Y(n_563)
);

AOI22xp5_ASAP7_75t_L g564 ( 
.A1(n_513),
.A2(n_450),
.B1(n_441),
.B2(n_467),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_515),
.Y(n_565)
);

AND2x2_ASAP7_75t_L g566 ( 
.A(n_503),
.B(n_446),
.Y(n_566)
);

AOI22xp5_ASAP7_75t_L g567 ( 
.A1(n_514),
.A2(n_467),
.B1(n_457),
.B2(n_469),
.Y(n_567)
);

OAI22xp33_ASAP7_75t_L g568 ( 
.A1(n_502),
.A2(n_456),
.B1(n_421),
.B2(n_412),
.Y(n_568)
);

OAI22xp33_ASAP7_75t_L g569 ( 
.A1(n_507),
.A2(n_456),
.B1(n_477),
.B2(n_476),
.Y(n_569)
);

AOI22xp5_ASAP7_75t_L g570 ( 
.A1(n_514),
.A2(n_469),
.B1(n_446),
.B2(n_465),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_561),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_SL g572 ( 
.A(n_553),
.B(n_479),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_550),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_565),
.Y(n_574)
);

CKINVDCx20_ASAP7_75t_R g575 ( 
.A(n_539),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_534),
.B(n_509),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_541),
.Y(n_577)
);

INVx5_ASAP7_75t_L g578 ( 
.A(n_547),
.Y(n_578)
);

AO21x2_ASAP7_75t_L g579 ( 
.A1(n_548),
.A2(n_510),
.B(n_527),
.Y(n_579)
);

INVx4_ASAP7_75t_L g580 ( 
.A(n_547),
.Y(n_580)
);

CKINVDCx11_ASAP7_75t_R g581 ( 
.A(n_545),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_552),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_SL g583 ( 
.A(n_568),
.B(n_479),
.Y(n_583)
);

INVx6_ASAP7_75t_L g584 ( 
.A(n_545),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_542),
.Y(n_585)
);

INVx2_ASAP7_75t_SL g586 ( 
.A(n_566),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_533),
.B(n_430),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_558),
.Y(n_588)
);

OAI22xp33_ASAP7_75t_L g589 ( 
.A1(n_555),
.A2(n_415),
.B1(n_489),
.B2(n_456),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_543),
.Y(n_590)
);

OR2x6_ASAP7_75t_L g591 ( 
.A(n_556),
.B(n_512),
.Y(n_591)
);

HB1xp67_ASAP7_75t_L g592 ( 
.A(n_563),
.Y(n_592)
);

INVxp33_ASAP7_75t_SL g593 ( 
.A(n_549),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_533),
.B(n_433),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_535),
.Y(n_595)
);

INVx8_ASAP7_75t_L g596 ( 
.A(n_536),
.Y(n_596)
);

INVx2_ASAP7_75t_SL g597 ( 
.A(n_556),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_544),
.Y(n_598)
);

INVx3_ASAP7_75t_L g599 ( 
.A(n_551),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_562),
.B(n_540),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_544),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_546),
.Y(n_602)
);

AOI22xp33_ASAP7_75t_L g603 ( 
.A1(n_537),
.A2(n_531),
.B1(n_520),
.B2(n_519),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_L g604 ( 
.A(n_554),
.B(n_531),
.Y(n_604)
);

BUFx2_ASAP7_75t_L g605 ( 
.A(n_546),
.Y(n_605)
);

NOR2xp33_ASAP7_75t_L g606 ( 
.A(n_554),
.B(n_522),
.Y(n_606)
);

INVx5_ASAP7_75t_L g607 ( 
.A(n_551),
.Y(n_607)
);

NOR2xp33_ASAP7_75t_L g608 ( 
.A(n_540),
.B(n_489),
.Y(n_608)
);

AOI21x1_ASAP7_75t_L g609 ( 
.A1(n_546),
.A2(n_510),
.B(n_442),
.Y(n_609)
);

CKINVDCx20_ASAP7_75t_R g610 ( 
.A(n_560),
.Y(n_610)
);

AO21x2_ASAP7_75t_L g611 ( 
.A1(n_548),
.A2(n_510),
.B(n_527),
.Y(n_611)
);

INVx4_ASAP7_75t_L g612 ( 
.A(n_538),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_559),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_559),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_538),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_538),
.Y(n_616)
);

BUFx3_ASAP7_75t_L g617 ( 
.A(n_557),
.Y(n_617)
);

AND2x2_ASAP7_75t_L g618 ( 
.A(n_567),
.B(n_433),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_570),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_568),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_SL g621 ( 
.A(n_569),
.B(n_479),
.Y(n_621)
);

AOI22xp5_ASAP7_75t_L g622 ( 
.A1(n_564),
.A2(n_468),
.B1(n_465),
.B2(n_456),
.Y(n_622)
);

INVx3_ASAP7_75t_L g623 ( 
.A(n_569),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_561),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_533),
.B(n_519),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_539),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_SL g627 ( 
.A(n_553),
.B(n_479),
.Y(n_627)
);

AOI21x1_ASAP7_75t_L g628 ( 
.A1(n_546),
.A2(n_442),
.B(n_532),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_550),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_SL g630 ( 
.A(n_553),
.B(n_490),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_533),
.B(n_519),
.Y(n_631)
);

NAND3xp33_ASAP7_75t_L g632 ( 
.A(n_567),
.B(n_452),
.C(n_454),
.Y(n_632)
);

BUFx2_ASAP7_75t_L g633 ( 
.A(n_566),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_533),
.B(n_413),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_SL g635 ( 
.A(n_553),
.B(n_490),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_533),
.B(n_413),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_550),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_550),
.Y(n_638)
);

AND3x2_ASAP7_75t_L g639 ( 
.A(n_533),
.B(n_453),
.C(n_449),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_561),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_533),
.B(n_413),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_550),
.Y(n_642)
);

INVxp67_ASAP7_75t_SL g643 ( 
.A(n_540),
.Y(n_643)
);

OAI22xp5_ASAP7_75t_L g644 ( 
.A1(n_567),
.A2(n_474),
.B1(n_465),
.B2(n_427),
.Y(n_644)
);

OAI22xp5_ASAP7_75t_L g645 ( 
.A1(n_567),
.A2(n_474),
.B1(n_427),
.B2(n_426),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_550),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_550),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_539),
.Y(n_648)
);

INVx3_ASAP7_75t_L g649 ( 
.A(n_545),
.Y(n_649)
);

INVx2_ASAP7_75t_SL g650 ( 
.A(n_566),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_571),
.Y(n_651)
);

NOR2xp33_ASAP7_75t_L g652 ( 
.A(n_634),
.B(n_514),
.Y(n_652)
);

AND2x4_ASAP7_75t_L g653 ( 
.A(n_633),
.B(n_514),
.Y(n_653)
);

AOI22xp33_ASAP7_75t_L g654 ( 
.A1(n_593),
.A2(n_520),
.B1(n_210),
.B2(n_202),
.Y(n_654)
);

OR2x6_ASAP7_75t_L g655 ( 
.A(n_591),
.B(n_512),
.Y(n_655)
);

INVx4_ASAP7_75t_SL g656 ( 
.A(n_584),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_582),
.B(n_499),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_624),
.Y(n_658)
);

INVx8_ASAP7_75t_L g659 ( 
.A(n_596),
.Y(n_659)
);

AOI22xp33_ASAP7_75t_L g660 ( 
.A1(n_593),
.A2(n_520),
.B1(n_210),
.B2(n_202),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_582),
.B(n_501),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_574),
.Y(n_662)
);

INVx4_ASAP7_75t_SL g663 ( 
.A(n_584),
.Y(n_663)
);

INVx4_ASAP7_75t_L g664 ( 
.A(n_581),
.Y(n_664)
);

INVx5_ASAP7_75t_L g665 ( 
.A(n_584),
.Y(n_665)
);

AND2x2_ASAP7_75t_L g666 ( 
.A(n_592),
.B(n_460),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_640),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_574),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_588),
.B(n_501),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_626),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_588),
.B(n_643),
.Y(n_671)
);

INVx4_ASAP7_75t_L g672 ( 
.A(n_581),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_629),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_629),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_L g675 ( 
.A(n_636),
.B(n_490),
.Y(n_675)
);

BUFx2_ASAP7_75t_L g676 ( 
.A(n_596),
.Y(n_676)
);

BUFx3_ASAP7_75t_L g677 ( 
.A(n_596),
.Y(n_677)
);

AND2x2_ASAP7_75t_L g678 ( 
.A(n_586),
.B(n_460),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_625),
.B(n_508),
.Y(n_679)
);

OR2x2_ASAP7_75t_L g680 ( 
.A(n_600),
.B(n_434),
.Y(n_680)
);

OR2x2_ASAP7_75t_L g681 ( 
.A(n_631),
.B(n_434),
.Y(n_681)
);

BUFx6f_ASAP7_75t_L g682 ( 
.A(n_650),
.Y(n_682)
);

NAND3x1_ASAP7_75t_L g683 ( 
.A(n_622),
.B(n_448),
.C(n_215),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_598),
.Y(n_684)
);

BUFx6f_ASAP7_75t_L g685 ( 
.A(n_639),
.Y(n_685)
);

BUFx3_ASAP7_75t_L g686 ( 
.A(n_606),
.Y(n_686)
);

AND2x4_ASAP7_75t_L g687 ( 
.A(n_577),
.B(n_529),
.Y(n_687)
);

INVx2_ASAP7_75t_SL g688 ( 
.A(n_585),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_598),
.Y(n_689)
);

BUFx10_ASAP7_75t_L g690 ( 
.A(n_608),
.Y(n_690)
);

AND2x6_ASAP7_75t_L g691 ( 
.A(n_599),
.B(n_518),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_620),
.B(n_508),
.Y(n_692)
);

HAxp5_ASAP7_75t_SL g693 ( 
.A(n_632),
.B(n_486),
.CON(n_693),
.SN(n_693)
);

NAND2xp5_ASAP7_75t_SL g694 ( 
.A(n_607),
.B(n_518),
.Y(n_694)
);

AND2x2_ASAP7_75t_L g695 ( 
.A(n_576),
.B(n_460),
.Y(n_695)
);

OR2x6_ASAP7_75t_L g696 ( 
.A(n_591),
.B(n_512),
.Y(n_696)
);

INVx3_ASAP7_75t_L g697 ( 
.A(n_577),
.Y(n_697)
);

INVx4_ASAP7_75t_L g698 ( 
.A(n_578),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_637),
.Y(n_699)
);

AOI22xp33_ASAP7_75t_L g700 ( 
.A1(n_617),
.A2(n_210),
.B1(n_218),
.B2(n_217),
.Y(n_700)
);

AND2x4_ASAP7_75t_L g701 ( 
.A(n_591),
.B(n_607),
.Y(n_701)
);

AOI21x1_ASAP7_75t_L g702 ( 
.A1(n_609),
.A2(n_442),
.B(n_532),
.Y(n_702)
);

OR2x6_ASAP7_75t_L g703 ( 
.A(n_583),
.B(n_512),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_601),
.Y(n_704)
);

AND2x6_ASAP7_75t_L g705 ( 
.A(n_599),
.B(n_518),
.Y(n_705)
);

BUFx3_ASAP7_75t_L g706 ( 
.A(n_606),
.Y(n_706)
);

INVx6_ASAP7_75t_L g707 ( 
.A(n_578),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_573),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_SL g709 ( 
.A(n_607),
.B(n_623),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_637),
.Y(n_710)
);

NOR2xp33_ASAP7_75t_L g711 ( 
.A(n_641),
.B(n_490),
.Y(n_711)
);

INVx5_ASAP7_75t_L g712 ( 
.A(n_578),
.Y(n_712)
);

AND2x2_ASAP7_75t_L g713 ( 
.A(n_576),
.B(n_485),
.Y(n_713)
);

NOR2xp33_ASAP7_75t_L g714 ( 
.A(n_608),
.B(n_493),
.Y(n_714)
);

NOR2xp33_ASAP7_75t_L g715 ( 
.A(n_617),
.B(n_493),
.Y(n_715)
);

INVx3_ASAP7_75t_L g716 ( 
.A(n_649),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_SL g717 ( 
.A(n_589),
.B(n_464),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_602),
.Y(n_718)
);

AND2x2_ASAP7_75t_L g719 ( 
.A(n_590),
.B(n_485),
.Y(n_719)
);

INVx3_ASAP7_75t_L g720 ( 
.A(n_649),
.Y(n_720)
);

AND2x4_ASAP7_75t_L g721 ( 
.A(n_607),
.B(n_529),
.Y(n_721)
);

INVx4_ASAP7_75t_L g722 ( 
.A(n_578),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_595),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_638),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_597),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_638),
.Y(n_726)
);

AND2x2_ASAP7_75t_L g727 ( 
.A(n_604),
.B(n_485),
.Y(n_727)
);

INVx4_ASAP7_75t_L g728 ( 
.A(n_580),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_642),
.Y(n_729)
);

A2O1A1Ixp33_ASAP7_75t_L g730 ( 
.A1(n_654),
.A2(n_623),
.B(n_603),
.C(n_644),
.Y(n_730)
);

INVx3_ASAP7_75t_L g731 ( 
.A(n_716),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_SL g732 ( 
.A(n_685),
.B(n_618),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_671),
.B(n_605),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_686),
.B(n_604),
.Y(n_734)
);

BUFx6f_ASAP7_75t_SL g735 ( 
.A(n_664),
.Y(n_735)
);

AND2x2_ASAP7_75t_L g736 ( 
.A(n_706),
.B(n_613),
.Y(n_736)
);

NOR2xp67_ASAP7_75t_L g737 ( 
.A(n_665),
.B(n_612),
.Y(n_737)
);

NAND2x1_ASAP7_75t_L g738 ( 
.A(n_707),
.B(n_580),
.Y(n_738)
);

NOR2xp33_ASAP7_75t_L g739 ( 
.A(n_680),
.B(n_475),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_671),
.B(n_594),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_SL g741 ( 
.A(n_685),
.B(n_464),
.Y(n_741)
);

BUFx6f_ASAP7_75t_L g742 ( 
.A(n_682),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_SL g743 ( 
.A(n_685),
.B(n_464),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_695),
.B(n_614),
.Y(n_744)
);

BUFx6f_ASAP7_75t_SL g745 ( 
.A(n_664),
.Y(n_745)
);

INVx8_ASAP7_75t_L g746 ( 
.A(n_659),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_651),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_681),
.B(n_587),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_708),
.B(n_619),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_658),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_675),
.B(n_619),
.Y(n_751)
);

NAND2xp33_ASAP7_75t_L g752 ( 
.A(n_654),
.B(n_464),
.Y(n_752)
);

NOR2xp33_ASAP7_75t_L g753 ( 
.A(n_690),
.B(n_475),
.Y(n_753)
);

HB1xp67_ASAP7_75t_L g754 ( 
.A(n_718),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_675),
.B(n_603),
.Y(n_755)
);

AND2x2_ASAP7_75t_L g756 ( 
.A(n_690),
.B(n_612),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_711),
.B(n_572),
.Y(n_757)
);

NAND2xp33_ASAP7_75t_L g758 ( 
.A(n_660),
.B(n_683),
.Y(n_758)
);

BUFx6f_ASAP7_75t_SL g759 ( 
.A(n_672),
.Y(n_759)
);

AND2x2_ASAP7_75t_L g760 ( 
.A(n_727),
.B(n_612),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_711),
.B(n_572),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_SL g762 ( 
.A(n_715),
.B(n_645),
.Y(n_762)
);

NOR2xp33_ASAP7_75t_L g763 ( 
.A(n_713),
.B(n_427),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_SL g764 ( 
.A(n_715),
.B(n_652),
.Y(n_764)
);

BUFx5_ASAP7_75t_L g765 ( 
.A(n_691),
.Y(n_765)
);

INVx2_ASAP7_75t_SL g766 ( 
.A(n_682),
.Y(n_766)
);

INVxp67_ASAP7_75t_L g767 ( 
.A(n_682),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_684),
.B(n_615),
.Y(n_768)
);

NOR2xp67_ASAP7_75t_L g769 ( 
.A(n_665),
.B(n_627),
.Y(n_769)
);

AND2x2_ASAP7_75t_SL g770 ( 
.A(n_701),
.B(n_616),
.Y(n_770)
);

BUFx6f_ASAP7_75t_L g771 ( 
.A(n_677),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_667),
.Y(n_772)
);

NOR2xp33_ASAP7_75t_L g773 ( 
.A(n_670),
.B(n_427),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_652),
.B(n_627),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_679),
.B(n_630),
.Y(n_775)
);

NOR2xp33_ASAP7_75t_L g776 ( 
.A(n_672),
.B(n_648),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_689),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_679),
.B(n_630),
.Y(n_778)
);

NOR2xp33_ASAP7_75t_L g779 ( 
.A(n_714),
.B(n_575),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_688),
.B(n_635),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_723),
.B(n_635),
.Y(n_781)
);

AND2x2_ASAP7_75t_SL g782 ( 
.A(n_701),
.B(n_616),
.Y(n_782)
);

NOR2xp33_ASAP7_75t_L g783 ( 
.A(n_714),
.B(n_575),
.Y(n_783)
);

NAND2x1_ASAP7_75t_L g784 ( 
.A(n_707),
.B(n_580),
.Y(n_784)
);

INVx4_ASAP7_75t_L g785 ( 
.A(n_665),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_666),
.B(n_610),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_704),
.Y(n_787)
);

NOR2xp33_ASAP7_75t_L g788 ( 
.A(n_676),
.B(n_610),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_726),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_662),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_668),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_SL g792 ( 
.A(n_665),
.B(n_583),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_673),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_SL g794 ( 
.A(n_717),
.B(n_621),
.Y(n_794)
);

INVx3_ASAP7_75t_L g795 ( 
.A(n_716),
.Y(n_795)
);

NOR2xp33_ASAP7_75t_L g796 ( 
.A(n_719),
.B(n_426),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_697),
.B(n_642),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_697),
.Y(n_798)
);

INVxp67_ASAP7_75t_L g799 ( 
.A(n_736),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_754),
.Y(n_800)
);

NOR2xp33_ASAP7_75t_L g801 ( 
.A(n_753),
.B(n_720),
.Y(n_801)
);

NOR2xp33_ASAP7_75t_L g802 ( 
.A(n_748),
.B(n_720),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_SL g803 ( 
.A(n_771),
.B(n_656),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_SL g804 ( 
.A(n_771),
.B(n_656),
.Y(n_804)
);

BUFx3_ASAP7_75t_L g805 ( 
.A(n_742),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_SL g806 ( 
.A(n_771),
.B(n_656),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_740),
.B(n_751),
.Y(n_807)
);

BUFx3_ASAP7_75t_L g808 ( 
.A(n_742),
.Y(n_808)
);

NOR2xp33_ASAP7_75t_L g809 ( 
.A(n_734),
.B(n_725),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_747),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_750),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_SL g812 ( 
.A(n_774),
.B(n_663),
.Y(n_812)
);

AOI22xp33_ASAP7_75t_L g813 ( 
.A1(n_758),
.A2(n_700),
.B1(n_660),
.B2(n_653),
.Y(n_813)
);

NOR3xp33_ASAP7_75t_L g814 ( 
.A(n_752),
.B(n_709),
.C(n_693),
.Y(n_814)
);

OR2x2_ASAP7_75t_L g815 ( 
.A(n_733),
.B(n_655),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_744),
.B(n_709),
.Y(n_816)
);

INVx4_ASAP7_75t_L g817 ( 
.A(n_735),
.Y(n_817)
);

NOR2xp33_ASAP7_75t_L g818 ( 
.A(n_739),
.B(n_653),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_733),
.B(n_678),
.Y(n_819)
);

INVx2_ASAP7_75t_SL g820 ( 
.A(n_742),
.Y(n_820)
);

OR2x6_ASAP7_75t_L g821 ( 
.A(n_746),
.B(n_655),
.Y(n_821)
);

AOI21xp5_ASAP7_75t_L g822 ( 
.A1(n_792),
.A2(n_621),
.B(n_694),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_SL g823 ( 
.A(n_764),
.B(n_796),
.Y(n_823)
);

BUFx4f_ASAP7_75t_L g824 ( 
.A(n_746),
.Y(n_824)
);

BUFx8_ASAP7_75t_L g825 ( 
.A(n_735),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_772),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_757),
.B(n_761),
.Y(n_827)
);

NOR2xp33_ASAP7_75t_L g828 ( 
.A(n_779),
.B(n_659),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_789),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_SL g830 ( 
.A(n_783),
.B(n_663),
.Y(n_830)
);

AND2x4_ASAP7_75t_L g831 ( 
.A(n_737),
.B(n_655),
.Y(n_831)
);

INVx3_ASAP7_75t_L g832 ( 
.A(n_731),
.Y(n_832)
);

INVx3_ASAP7_75t_L g833 ( 
.A(n_731),
.Y(n_833)
);

NAND3xp33_ASAP7_75t_L g834 ( 
.A(n_730),
.B(n_700),
.C(n_216),
.Y(n_834)
);

NAND2xp33_ASAP7_75t_L g835 ( 
.A(n_746),
.B(n_659),
.Y(n_835)
);

NOR2xp33_ASAP7_75t_L g836 ( 
.A(n_788),
.B(n_728),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_777),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_775),
.B(n_674),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_SL g839 ( 
.A(n_732),
.B(n_663),
.Y(n_839)
);

BUFx6f_ASAP7_75t_L g840 ( 
.A(n_766),
.Y(n_840)
);

NOR2xp33_ASAP7_75t_L g841 ( 
.A(n_763),
.B(n_728),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_778),
.B(n_699),
.Y(n_842)
);

NOR2xp33_ASAP7_75t_L g843 ( 
.A(n_767),
.B(n_721),
.Y(n_843)
);

NOR2x1p5_ASAP7_75t_L g844 ( 
.A(n_755),
.B(n_692),
.Y(n_844)
);

NOR3xp33_ASAP7_75t_L g845 ( 
.A(n_741),
.B(n_694),
.C(n_692),
.Y(n_845)
);

AOI22xp5_ASAP7_75t_L g846 ( 
.A1(n_762),
.A2(n_696),
.B1(n_721),
.B2(n_703),
.Y(n_846)
);

INVxp33_ASAP7_75t_L g847 ( 
.A(n_773),
.Y(n_847)
);

AOI22xp5_ASAP7_75t_L g848 ( 
.A1(n_745),
.A2(n_696),
.B1(n_703),
.B2(n_691),
.Y(n_848)
);

INVx2_ASAP7_75t_SL g849 ( 
.A(n_795),
.Y(n_849)
);

OR2x2_ASAP7_75t_L g850 ( 
.A(n_768),
.B(n_696),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_749),
.B(n_710),
.Y(n_851)
);

BUFx3_ASAP7_75t_L g852 ( 
.A(n_776),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_790),
.Y(n_853)
);

AND2x6_ASAP7_75t_SL g854 ( 
.A(n_745),
.B(n_703),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_781),
.B(n_724),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_791),
.Y(n_856)
);

INVx4_ASAP7_75t_L g857 ( 
.A(n_759),
.Y(n_857)
);

AOI22xp5_ASAP7_75t_L g858 ( 
.A1(n_759),
.A2(n_705),
.B1(n_691),
.B2(n_707),
.Y(n_858)
);

AOI22xp5_ASAP7_75t_L g859 ( 
.A1(n_794),
.A2(n_705),
.B1(n_691),
.B2(n_579),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_793),
.B(n_729),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_787),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_786),
.B(n_657),
.Y(n_862)
);

HB1xp67_ASAP7_75t_L g863 ( 
.A(n_780),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_SL g864 ( 
.A(n_756),
.B(n_712),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_760),
.B(n_657),
.Y(n_865)
);

NOR2xp33_ASAP7_75t_SL g866 ( 
.A(n_785),
.B(n_698),
.Y(n_866)
);

BUFx8_ASAP7_75t_L g867 ( 
.A(n_798),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_797),
.B(n_661),
.Y(n_868)
);

INVx8_ASAP7_75t_L g869 ( 
.A(n_795),
.Y(n_869)
);

A2O1A1Ixp33_ASAP7_75t_L g870 ( 
.A1(n_769),
.A2(n_236),
.B(n_212),
.C(n_223),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_768),
.B(n_661),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_770),
.B(n_669),
.Y(n_872)
);

NOR2xp67_ASAP7_75t_L g873 ( 
.A(n_785),
.B(n_712),
.Y(n_873)
);

INVxp67_ASAP7_75t_L g874 ( 
.A(n_863),
.Y(n_874)
);

AO22x2_ASAP7_75t_L g875 ( 
.A1(n_800),
.A2(n_743),
.B1(n_784),
.B2(n_738),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_810),
.Y(n_876)
);

BUFx6f_ASAP7_75t_L g877 ( 
.A(n_824),
.Y(n_877)
);

BUFx6f_ASAP7_75t_SL g878 ( 
.A(n_817),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_811),
.Y(n_879)
);

AND2x2_ASAP7_75t_L g880 ( 
.A(n_799),
.B(n_782),
.Y(n_880)
);

AND2x2_ASAP7_75t_L g881 ( 
.A(n_815),
.B(n_765),
.Y(n_881)
);

OAI221xp5_ASAP7_75t_L g882 ( 
.A1(n_834),
.A2(n_769),
.B1(n_219),
.B2(n_221),
.C(n_737),
.Y(n_882)
);

AND2x2_ASAP7_75t_SL g883 ( 
.A(n_814),
.B(n_698),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_829),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_SL g885 ( 
.A(n_817),
.B(n_765),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_853),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_807),
.B(n_765),
.Y(n_887)
);

NOR2xp33_ASAP7_75t_L g888 ( 
.A(n_847),
.B(n_765),
.Y(n_888)
);

AO22x2_ASAP7_75t_L g889 ( 
.A1(n_837),
.A2(n_722),
.B1(n_687),
.B2(n_669),
.Y(n_889)
);

BUFx8_ASAP7_75t_L g890 ( 
.A(n_852),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_856),
.Y(n_891)
);

OR2x6_ASAP7_75t_L g892 ( 
.A(n_857),
.B(n_722),
.Y(n_892)
);

AO22x2_ASAP7_75t_L g893 ( 
.A1(n_861),
.A2(n_687),
.B1(n_765),
.B2(n_647),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_827),
.B(n_579),
.Y(n_894)
);

NAND2x1p5_ASAP7_75t_L g895 ( 
.A(n_824),
.B(n_712),
.Y(n_895)
);

OAI221xp5_ASAP7_75t_L g896 ( 
.A1(n_813),
.A2(n_229),
.B1(n_222),
.B2(n_227),
.C(n_188),
.Y(n_896)
);

INVxp67_ASAP7_75t_L g897 ( 
.A(n_809),
.Y(n_897)
);

NAND2x1p5_ASAP7_75t_L g898 ( 
.A(n_803),
.B(n_712),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_844),
.B(n_802),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_SL g900 ( 
.A(n_857),
.B(n_646),
.Y(n_900)
);

AND2x4_ASAP7_75t_L g901 ( 
.A(n_831),
.B(n_864),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_826),
.Y(n_902)
);

AND2x4_ASAP7_75t_L g903 ( 
.A(n_831),
.B(n_705),
.Y(n_903)
);

HB1xp67_ASAP7_75t_L g904 ( 
.A(n_850),
.Y(n_904)
);

AO22x2_ASAP7_75t_L g905 ( 
.A1(n_849),
.A2(n_647),
.B1(n_646),
.B2(n_498),
.Y(n_905)
);

AO22x2_ASAP7_75t_L g906 ( 
.A1(n_822),
.A2(n_496),
.B1(n_487),
.B2(n_507),
.Y(n_906)
);

AO22x2_ASAP7_75t_L g907 ( 
.A1(n_839),
.A2(n_529),
.B1(n_521),
.B2(n_526),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_860),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_855),
.Y(n_909)
);

CKINVDCx5p33_ASAP7_75t_R g910 ( 
.A(n_825),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_838),
.Y(n_911)
);

CKINVDCx5p33_ASAP7_75t_R g912 ( 
.A(n_825),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_842),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_851),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_832),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_833),
.Y(n_916)
);

OR2x2_ASAP7_75t_L g917 ( 
.A(n_819),
.B(n_611),
.Y(n_917)
);

AO22x2_ASAP7_75t_L g918 ( 
.A1(n_833),
.A2(n_529),
.B1(n_521),
.B2(n_526),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_871),
.Y(n_919)
);

HB1xp67_ASAP7_75t_L g920 ( 
.A(n_816),
.Y(n_920)
);

AO22x2_ASAP7_75t_L g921 ( 
.A1(n_812),
.A2(n_529),
.B1(n_521),
.B2(n_526),
.Y(n_921)
);

AND2x2_ASAP7_75t_L g922 ( 
.A(n_865),
.B(n_611),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_868),
.Y(n_923)
);

AOI21xp5_ASAP7_75t_L g924 ( 
.A1(n_896),
.A2(n_870),
.B(n_835),
.Y(n_924)
);

INVx1_ASAP7_75t_SL g925 ( 
.A(n_910),
.Y(n_925)
);

INVx2_ASAP7_75t_SL g926 ( 
.A(n_890),
.Y(n_926)
);

A2O1A1Ixp33_ASAP7_75t_L g927 ( 
.A1(n_882),
.A2(n_823),
.B(n_828),
.C(n_836),
.Y(n_927)
);

BUFx6f_ASAP7_75t_L g928 ( 
.A(n_877),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_923),
.B(n_872),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_923),
.B(n_862),
.Y(n_930)
);

INVx5_ASAP7_75t_L g931 ( 
.A(n_877),
.Y(n_931)
);

AOI21xp5_ASAP7_75t_L g932 ( 
.A1(n_906),
.A2(n_806),
.B(n_804),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_919),
.B(n_845),
.Y(n_933)
);

AND2x4_ASAP7_75t_L g934 ( 
.A(n_901),
.B(n_821),
.Y(n_934)
);

AOI22xp5_ASAP7_75t_L g935 ( 
.A1(n_883),
.A2(n_888),
.B1(n_906),
.B2(n_901),
.Y(n_935)
);

INVx2_ASAP7_75t_L g936 ( 
.A(n_876),
.Y(n_936)
);

AOI21xp5_ASAP7_75t_L g937 ( 
.A1(n_885),
.A2(n_830),
.B(n_866),
.Y(n_937)
);

BUFx6f_ASAP7_75t_L g938 ( 
.A(n_877),
.Y(n_938)
);

NOR2x1_ASAP7_75t_R g939 ( 
.A(n_912),
.B(n_805),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_919),
.B(n_801),
.Y(n_940)
);

CKINVDCx5p33_ASAP7_75t_R g941 ( 
.A(n_878),
.Y(n_941)
);

INVx4_ASAP7_75t_L g942 ( 
.A(n_892),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_876),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_920),
.B(n_846),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_911),
.B(n_859),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_915),
.Y(n_946)
);

AOI21xp5_ASAP7_75t_L g947 ( 
.A1(n_900),
.A2(n_821),
.B(n_848),
.Y(n_947)
);

AOI21xp5_ASAP7_75t_L g948 ( 
.A1(n_875),
.A2(n_873),
.B(n_858),
.Y(n_948)
);

NOR2xp33_ASAP7_75t_L g949 ( 
.A(n_897),
.B(n_818),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_913),
.B(n_854),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_SL g951 ( 
.A(n_899),
.B(n_840),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_909),
.B(n_869),
.Y(n_952)
);

A2O1A1Ixp33_ASAP7_75t_L g953 ( 
.A1(n_894),
.A2(n_841),
.B(n_843),
.C(n_873),
.Y(n_953)
);

INVx2_ASAP7_75t_L g954 ( 
.A(n_916),
.Y(n_954)
);

AOI21xp5_ASAP7_75t_L g955 ( 
.A1(n_875),
.A2(n_869),
.B(n_820),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_879),
.Y(n_956)
);

NOR2xp33_ASAP7_75t_L g957 ( 
.A(n_890),
.B(n_867),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_874),
.B(n_840),
.Y(n_958)
);

NOR2xp33_ASAP7_75t_L g959 ( 
.A(n_887),
.B(n_867),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_914),
.B(n_908),
.Y(n_960)
);

AOI21xp5_ASAP7_75t_L g961 ( 
.A1(n_892),
.A2(n_889),
.B(n_907),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_922),
.B(n_904),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_902),
.B(n_840),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_884),
.B(n_808),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_SL g965 ( 
.A(n_898),
.B(n_628),
.Y(n_965)
);

NOR2xp33_ASAP7_75t_SL g966 ( 
.A(n_895),
.B(n_705),
.Y(n_966)
);

AOI21xp5_ASAP7_75t_L g967 ( 
.A1(n_889),
.A2(n_200),
.B(n_418),
.Y(n_967)
);

AOI21xp5_ASAP7_75t_L g968 ( 
.A1(n_907),
.A2(n_225),
.B(n_214),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_SL g969 ( 
.A(n_903),
.B(n_213),
.Y(n_969)
);

AOI21xp5_ASAP7_75t_L g970 ( 
.A1(n_921),
.A2(n_225),
.B(n_214),
.Y(n_970)
);

O2A1O1Ixp33_ASAP7_75t_L g971 ( 
.A1(n_917),
.A2(n_0),
.B(n_1),
.C(n_2),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_886),
.B(n_213),
.Y(n_972)
);

AOI21x1_ASAP7_75t_L g973 ( 
.A1(n_905),
.A2(n_918),
.B(n_893),
.Y(n_973)
);

BUFx6f_ASAP7_75t_L g974 ( 
.A(n_903),
.Y(n_974)
);

AOI21xp5_ASAP7_75t_L g975 ( 
.A1(n_921),
.A2(n_225),
.B(n_420),
.Y(n_975)
);

A2O1A1Ixp33_ASAP7_75t_L g976 ( 
.A1(n_881),
.A2(n_225),
.B(n_4),
.C(n_5),
.Y(n_976)
);

NOR2xp33_ASAP7_75t_L g977 ( 
.A(n_880),
.B(n_2),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_891),
.B(n_213),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_905),
.Y(n_979)
);

HB1xp67_ASAP7_75t_L g980 ( 
.A(n_874),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_876),
.Y(n_981)
);

INVx2_ASAP7_75t_SL g982 ( 
.A(n_890),
.Y(n_982)
);

AND2x4_ASAP7_75t_L g983 ( 
.A(n_979),
.B(n_702),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_943),
.Y(n_984)
);

O2A1O1Ixp33_ASAP7_75t_L g985 ( 
.A1(n_976),
.A2(n_4),
.B(n_5),
.C(n_6),
.Y(n_985)
);

INVx2_ASAP7_75t_L g986 ( 
.A(n_936),
.Y(n_986)
);

INVx2_ASAP7_75t_SL g987 ( 
.A(n_931),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_933),
.B(n_213),
.Y(n_988)
);

BUFx12f_ASAP7_75t_L g989 ( 
.A(n_941),
.Y(n_989)
);

INVxp67_ASAP7_75t_L g990 ( 
.A(n_980),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_945),
.B(n_213),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_930),
.B(n_213),
.Y(n_992)
);

BUFx3_ASAP7_75t_L g993 ( 
.A(n_926),
.Y(n_993)
);

INVx2_ASAP7_75t_L g994 ( 
.A(n_981),
.Y(n_994)
);

AND3x1_ASAP7_75t_SL g995 ( 
.A(n_939),
.B(n_956),
.C(n_935),
.Y(n_995)
);

NOR2xp33_ASAP7_75t_R g996 ( 
.A(n_982),
.B(n_6),
.Y(n_996)
);

O2A1O1Ixp33_ASAP7_75t_L g997 ( 
.A1(n_971),
.A2(n_7),
.B(n_8),
.C(n_9),
.Y(n_997)
);

INVx2_ASAP7_75t_SL g998 ( 
.A(n_931),
.Y(n_998)
);

AND2x6_ASAP7_75t_L g999 ( 
.A(n_928),
.B(n_521),
.Y(n_999)
);

INVx2_ASAP7_75t_L g1000 ( 
.A(n_973),
.Y(n_1000)
);

BUFx3_ASAP7_75t_L g1001 ( 
.A(n_931),
.Y(n_1001)
);

INVx2_ASAP7_75t_L g1002 ( 
.A(n_946),
.Y(n_1002)
);

INVx2_ASAP7_75t_L g1003 ( 
.A(n_954),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_SL g1004 ( 
.A(n_990),
.B(n_942),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_991),
.B(n_950),
.Y(n_1005)
);

NOR2x1_ASAP7_75t_L g1006 ( 
.A(n_1001),
.B(n_957),
.Y(n_1006)
);

AOI21x1_ASAP7_75t_L g1007 ( 
.A1(n_1000),
.A2(n_978),
.B(n_972),
.Y(n_1007)
);

OAI22xp5_ASAP7_75t_L g1008 ( 
.A1(n_993),
.A2(n_967),
.B1(n_953),
.B2(n_944),
.Y(n_1008)
);

OAI21xp33_ASAP7_75t_L g1009 ( 
.A1(n_997),
.A2(n_929),
.B(n_940),
.Y(n_1009)
);

OAI21x1_ASAP7_75t_L g1010 ( 
.A1(n_1000),
.A2(n_948),
.B(n_955),
.Y(n_1010)
);

AOI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_985),
.A2(n_924),
.B(n_927),
.Y(n_1011)
);

AND2x2_ASAP7_75t_L g1012 ( 
.A(n_993),
.B(n_974),
.Y(n_1012)
);

BUFx6f_ASAP7_75t_L g1013 ( 
.A(n_989),
.Y(n_1013)
);

NOR2xp33_ASAP7_75t_L g1014 ( 
.A(n_989),
.B(n_925),
.Y(n_1014)
);

AOI21x1_ASAP7_75t_L g1015 ( 
.A1(n_987),
.A2(n_951),
.B(n_968),
.Y(n_1015)
);

AOI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_988),
.A2(n_969),
.B(n_961),
.Y(n_1016)
);

OAI22x1_ASAP7_75t_L g1017 ( 
.A1(n_987),
.A2(n_977),
.B1(n_949),
.B2(n_959),
.Y(n_1017)
);

A2O1A1Ixp33_ASAP7_75t_L g1018 ( 
.A1(n_995),
.A2(n_932),
.B(n_937),
.C(n_947),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_998),
.B(n_960),
.Y(n_1019)
);

NOR2xp33_ASAP7_75t_L g1020 ( 
.A(n_1001),
.B(n_928),
.Y(n_1020)
);

CKINVDCx6p67_ASAP7_75t_R g1021 ( 
.A(n_996),
.Y(n_1021)
);

NOR2xp33_ASAP7_75t_L g1022 ( 
.A(n_998),
.B(n_928),
.Y(n_1022)
);

O2A1O1Ixp33_ASAP7_75t_SL g1023 ( 
.A1(n_992),
.A2(n_958),
.B(n_952),
.C(n_963),
.Y(n_1023)
);

OAI22xp5_ASAP7_75t_L g1024 ( 
.A1(n_984),
.A2(n_974),
.B1(n_970),
.B2(n_975),
.Y(n_1024)
);

OR2x2_ASAP7_75t_L g1025 ( 
.A(n_1003),
.B(n_962),
.Y(n_1025)
);

INVxp67_ASAP7_75t_L g1026 ( 
.A(n_984),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_994),
.Y(n_1027)
);

OAI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_1002),
.A2(n_965),
.B(n_964),
.Y(n_1028)
);

AO31x2_ASAP7_75t_L g1029 ( 
.A1(n_1018),
.A2(n_994),
.A3(n_986),
.B(n_1002),
.Y(n_1029)
);

AND2x2_ASAP7_75t_L g1030 ( 
.A(n_1006),
.B(n_974),
.Y(n_1030)
);

INVx4_ASAP7_75t_L g1031 ( 
.A(n_1013),
.Y(n_1031)
);

NOR2xp33_ASAP7_75t_SL g1032 ( 
.A(n_1021),
.B(n_938),
.Y(n_1032)
);

INVx3_ASAP7_75t_L g1033 ( 
.A(n_1013),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_SL g1034 ( 
.A(n_1008),
.B(n_934),
.Y(n_1034)
);

NAND2x1p5_ASAP7_75t_L g1035 ( 
.A(n_1012),
.B(n_938),
.Y(n_1035)
);

INVx2_ASAP7_75t_L g1036 ( 
.A(n_1033),
.Y(n_1036)
);

AND2x4_ASAP7_75t_L g1037 ( 
.A(n_1030),
.B(n_1013),
.Y(n_1037)
);

AND2x2_ASAP7_75t_L g1038 ( 
.A(n_1037),
.B(n_1033),
.Y(n_1038)
);

OAI21x1_ASAP7_75t_L g1039 ( 
.A1(n_1036),
.A2(n_1010),
.B(n_1035),
.Y(n_1039)
);

OAI21x1_ASAP7_75t_L g1040 ( 
.A1(n_1037),
.A2(n_1034),
.B(n_1004),
.Y(n_1040)
);

INVx1_ASAP7_75t_SL g1041 ( 
.A(n_1038),
.Y(n_1041)
);

BUFx2_ASAP7_75t_L g1042 ( 
.A(n_1040),
.Y(n_1042)
);

BUFx2_ASAP7_75t_L g1043 ( 
.A(n_1040),
.Y(n_1043)
);

BUFx2_ASAP7_75t_SL g1044 ( 
.A(n_1041),
.Y(n_1044)
);

BUFx8_ASAP7_75t_SL g1045 ( 
.A(n_1042),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_1044),
.Y(n_1046)
);

BUFx2_ASAP7_75t_R g1047 ( 
.A(n_1045),
.Y(n_1047)
);

AND2x2_ASAP7_75t_L g1048 ( 
.A(n_1046),
.B(n_1031),
.Y(n_1048)
);

AOI21x1_ASAP7_75t_SL g1049 ( 
.A1(n_1047),
.A2(n_1031),
.B(n_1005),
.Y(n_1049)
);

BUFx3_ASAP7_75t_L g1050 ( 
.A(n_1048),
.Y(n_1050)
);

OAI21xp5_ASAP7_75t_SL g1051 ( 
.A1(n_1049),
.A2(n_1043),
.B(n_1011),
.Y(n_1051)
);

AO21x2_ASAP7_75t_L g1052 ( 
.A1(n_1051),
.A2(n_1039),
.B(n_1014),
.Y(n_1052)
);

AND2x4_ASAP7_75t_L g1053 ( 
.A(n_1050),
.B(n_1039),
.Y(n_1053)
);

AND2x2_ASAP7_75t_L g1054 ( 
.A(n_1052),
.B(n_1032),
.Y(n_1054)
);

AO32x2_ASAP7_75t_L g1055 ( 
.A1(n_1052),
.A2(n_1029),
.A3(n_1024),
.B1(n_1022),
.B2(n_1020),
.Y(n_1055)
);

AND2x2_ASAP7_75t_L g1056 ( 
.A(n_1054),
.B(n_1053),
.Y(n_1056)
);

AND2x2_ASAP7_75t_L g1057 ( 
.A(n_1055),
.B(n_1029),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_1054),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_1057),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_1056),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_1056),
.Y(n_1061)
);

A2O1A1Ixp33_ASAP7_75t_L g1062 ( 
.A1(n_1060),
.A2(n_1058),
.B(n_1053),
.C(n_1026),
.Y(n_1062)
);

INVx2_ASAP7_75t_L g1063 ( 
.A(n_1061),
.Y(n_1063)
);

AOI22xp33_ASAP7_75t_L g1064 ( 
.A1(n_1063),
.A2(n_1059),
.B1(n_1017),
.B2(n_1027),
.Y(n_1064)
);

INVx2_ASAP7_75t_L g1065 ( 
.A(n_1062),
.Y(n_1065)
);

AOI22xp33_ASAP7_75t_L g1066 ( 
.A1(n_1064),
.A2(n_938),
.B1(n_1016),
.B2(n_1019),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_1065),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_1067),
.B(n_1029),
.Y(n_1068)
);

INVx1_ASAP7_75t_SL g1069 ( 
.A(n_1066),
.Y(n_1069)
);

AND2x2_ASAP7_75t_L g1070 ( 
.A(n_1069),
.B(n_1025),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_1068),
.B(n_1009),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_1070),
.Y(n_1072)
);

OAI33xp33_ASAP7_75t_L g1073 ( 
.A1(n_1071),
.A2(n_7),
.A3(n_8),
.B1(n_9),
.B2(n_10),
.B3(n_11),
.Y(n_1073)
);

OR2x2_ASAP7_75t_L g1074 ( 
.A(n_1072),
.B(n_1028),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_1073),
.Y(n_1075)
);

INVx2_ASAP7_75t_L g1076 ( 
.A(n_1072),
.Y(n_1076)
);

AND2x2_ASAP7_75t_L g1077 ( 
.A(n_1076),
.B(n_1007),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_1074),
.Y(n_1078)
);

INVxp67_ASAP7_75t_SL g1079 ( 
.A(n_1075),
.Y(n_1079)
);

OR2x2_ASAP7_75t_L g1080 ( 
.A(n_1077),
.B(n_10),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_1079),
.Y(n_1081)
);

INVxp67_ASAP7_75t_L g1082 ( 
.A(n_1080),
.Y(n_1082)
);

NOR2xp33_ASAP7_75t_L g1083 ( 
.A(n_1081),
.B(n_1078),
.Y(n_1083)
);

AND2x2_ASAP7_75t_L g1084 ( 
.A(n_1082),
.B(n_1003),
.Y(n_1084)
);

AOI22xp33_ASAP7_75t_L g1085 ( 
.A1(n_1083),
.A2(n_983),
.B1(n_986),
.B2(n_480),
.Y(n_1085)
);

AOI221xp5_ASAP7_75t_L g1086 ( 
.A1(n_1084),
.A2(n_1085),
.B1(n_1023),
.B2(n_284),
.C(n_15),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_1084),
.Y(n_1087)
);

INVx1_ASAP7_75t_SL g1088 ( 
.A(n_1087),
.Y(n_1088)
);

AOI22xp5_ASAP7_75t_L g1089 ( 
.A1(n_1086),
.A2(n_983),
.B1(n_13),
.B2(n_14),
.Y(n_1089)
);

AOI32xp33_ASAP7_75t_L g1090 ( 
.A1(n_1088),
.A2(n_11),
.A3(n_13),
.B1(n_15),
.B2(n_16),
.Y(n_1090)
);

AOI21xp5_ASAP7_75t_L g1091 ( 
.A1(n_1089),
.A2(n_17),
.B(n_18),
.Y(n_1091)
);

O2A1O1Ixp33_ASAP7_75t_L g1092 ( 
.A1(n_1091),
.A2(n_17),
.B(n_18),
.C(n_19),
.Y(n_1092)
);

NAND3xp33_ASAP7_75t_L g1093 ( 
.A(n_1090),
.B(n_19),
.C(n_20),
.Y(n_1093)
);

OAI32xp33_ASAP7_75t_L g1094 ( 
.A1(n_1091),
.A2(n_20),
.A3(n_21),
.B1(n_22),
.B2(n_23),
.Y(n_1094)
);

OR2x2_ASAP7_75t_L g1095 ( 
.A(n_1093),
.B(n_21),
.Y(n_1095)
);

INVx2_ASAP7_75t_L g1096 ( 
.A(n_1094),
.Y(n_1096)
);

INVx2_ASAP7_75t_L g1097 ( 
.A(n_1092),
.Y(n_1097)
);

CKINVDCx16_ASAP7_75t_R g1098 ( 
.A(n_1097),
.Y(n_1098)
);

INVxp67_ASAP7_75t_L g1099 ( 
.A(n_1096),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_SL g1100 ( 
.A(n_1098),
.B(n_1095),
.Y(n_1100)
);

NOR3xp33_ASAP7_75t_L g1101 ( 
.A(n_1099),
.B(n_22),
.C(n_24),
.Y(n_1101)
);

AND2x2_ASAP7_75t_L g1102 ( 
.A(n_1100),
.B(n_24),
.Y(n_1102)
);

O2A1O1Ixp33_ASAP7_75t_SL g1103 ( 
.A1(n_1101),
.A2(n_25),
.B(n_27),
.C(n_28),
.Y(n_1103)
);

NOR2xp33_ASAP7_75t_L g1104 ( 
.A(n_1103),
.B(n_25),
.Y(n_1104)
);

NOR2xp33_ASAP7_75t_L g1105 ( 
.A(n_1102),
.B(n_28),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_1104),
.B(n_29),
.Y(n_1106)
);

AOI221xp5_ASAP7_75t_L g1107 ( 
.A1(n_1105),
.A2(n_29),
.B1(n_30),
.B2(n_31),
.C(n_32),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_1106),
.B(n_31),
.Y(n_1108)
);

OAI21xp5_ASAP7_75t_SL g1109 ( 
.A1(n_1107),
.A2(n_33),
.B(n_34),
.Y(n_1109)
);

AO22x2_ASAP7_75t_L g1110 ( 
.A1(n_1109),
.A2(n_33),
.B1(n_34),
.B2(n_35),
.Y(n_1110)
);

AOI22xp5_ASAP7_75t_L g1111 ( 
.A1(n_1108),
.A2(n_35),
.B1(n_480),
.B2(n_999),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_1109),
.Y(n_1112)
);

OAI31xp33_ASAP7_75t_SL g1113 ( 
.A1(n_1112),
.A2(n_40),
.A3(n_41),
.B(n_42),
.Y(n_1113)
);

AOI211xp5_ASAP7_75t_L g1114 ( 
.A1(n_1110),
.A2(n_44),
.B(n_45),
.C(n_46),
.Y(n_1114)
);

OAI221xp5_ASAP7_75t_L g1115 ( 
.A1(n_1111),
.A2(n_47),
.B1(n_48),
.B2(n_50),
.C(n_52),
.Y(n_1115)
);

OAI22xp33_ASAP7_75t_L g1116 ( 
.A1(n_1115),
.A2(n_493),
.B1(n_1015),
.B2(n_353),
.Y(n_1116)
);

BUFx2_ASAP7_75t_L g1117 ( 
.A(n_1113),
.Y(n_1117)
);

NOR3xp33_ASAP7_75t_SL g1118 ( 
.A(n_1117),
.B(n_1114),
.C(n_53),
.Y(n_1118)
);

NOR2x1_ASAP7_75t_L g1119 ( 
.A(n_1116),
.B(n_320),
.Y(n_1119)
);

NAND3xp33_ASAP7_75t_L g1120 ( 
.A(n_1119),
.B(n_1118),
.C(n_353),
.Y(n_1120)
);

NOR2x1_ASAP7_75t_L g1121 ( 
.A(n_1119),
.B(n_320),
.Y(n_1121)
);

NOR4xp75_ASAP7_75t_L g1122 ( 
.A(n_1120),
.B(n_56),
.C(n_57),
.D(n_59),
.Y(n_1122)
);

INVx2_ASAP7_75t_SL g1123 ( 
.A(n_1121),
.Y(n_1123)
);

XNOR2x1_ASAP7_75t_L g1124 ( 
.A(n_1123),
.B(n_62),
.Y(n_1124)
);

AOI221xp5_ASAP7_75t_L g1125 ( 
.A1(n_1122),
.A2(n_353),
.B1(n_320),
.B2(n_483),
.C(n_482),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_SL g1126 ( 
.A(n_1125),
.B(n_353),
.Y(n_1126)
);

OAI22xp5_ASAP7_75t_SL g1127 ( 
.A1(n_1124),
.A2(n_63),
.B1(n_64),
.B2(n_66),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_1126),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_1127),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_1126),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_1128),
.Y(n_1131)
);

NOR3xp33_ASAP7_75t_L g1132 ( 
.A(n_1130),
.B(n_68),
.C(n_69),
.Y(n_1132)
);

OAI211xp5_ASAP7_75t_L g1133 ( 
.A1(n_1129),
.A2(n_71),
.B(n_72),
.C(n_73),
.Y(n_1133)
);

XOR2xp5_ASAP7_75t_L g1134 ( 
.A(n_1131),
.B(n_74),
.Y(n_1134)
);

INVx2_ASAP7_75t_L g1135 ( 
.A(n_1132),
.Y(n_1135)
);

AOI22xp5_ASAP7_75t_L g1136 ( 
.A1(n_1135),
.A2(n_1133),
.B1(n_999),
.B2(n_483),
.Y(n_1136)
);

BUFx6f_ASAP7_75t_L g1137 ( 
.A(n_1134),
.Y(n_1137)
);

AOI22xp5_ASAP7_75t_SL g1138 ( 
.A1(n_1137),
.A2(n_480),
.B1(n_999),
.B2(n_483),
.Y(n_1138)
);

NOR2x1_ASAP7_75t_L g1139 ( 
.A(n_1136),
.B(n_353),
.Y(n_1139)
);

XNOR2xp5_ASAP7_75t_L g1140 ( 
.A(n_1139),
.B(n_75),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_1138),
.Y(n_1141)
);

INVxp67_ASAP7_75t_SL g1142 ( 
.A(n_1141),
.Y(n_1142)
);

OAI22xp5_ASAP7_75t_L g1143 ( 
.A1(n_1140),
.A2(n_493),
.B1(n_472),
.B2(n_470),
.Y(n_1143)
);

AOI22xp5_ASAP7_75t_L g1144 ( 
.A1(n_1142),
.A2(n_999),
.B1(n_480),
.B2(n_472),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_1143),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_1142),
.Y(n_1146)
);

AND2x2_ASAP7_75t_L g1147 ( 
.A(n_1146),
.B(n_76),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_1145),
.Y(n_1148)
);

AOI222xp33_ASAP7_75t_SL g1149 ( 
.A1(n_1144),
.A2(n_480),
.B1(n_80),
.B2(n_81),
.C1(n_84),
.C2(n_85),
.Y(n_1149)
);

INVxp67_ASAP7_75t_L g1150 ( 
.A(n_1146),
.Y(n_1150)
);

INVx2_ASAP7_75t_L g1151 ( 
.A(n_1148),
.Y(n_1151)
);

HB1xp67_ASAP7_75t_L g1152 ( 
.A(n_1150),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_1147),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_1149),
.B(n_78),
.Y(n_1154)
);

OR2x2_ASAP7_75t_L g1155 ( 
.A(n_1151),
.B(n_87),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_1152),
.Y(n_1156)
);

AOI21xp5_ASAP7_75t_L g1157 ( 
.A1(n_1153),
.A2(n_88),
.B(n_91),
.Y(n_1157)
);

OAI21xp5_ASAP7_75t_L g1158 ( 
.A1(n_1154),
.A2(n_999),
.B(n_96),
.Y(n_1158)
);

NOR2x1_ASAP7_75t_L g1159 ( 
.A(n_1151),
.B(n_93),
.Y(n_1159)
);

AOI22xp33_ASAP7_75t_L g1160 ( 
.A1(n_1151),
.A2(n_999),
.B1(n_480),
.B2(n_472),
.Y(n_1160)
);

AOI22xp33_ASAP7_75t_L g1161 ( 
.A1(n_1151),
.A2(n_470),
.B1(n_98),
.B2(n_103),
.Y(n_1161)
);

HB1xp67_ASAP7_75t_L g1162 ( 
.A(n_1152),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_1152),
.Y(n_1163)
);

AOI22xp33_ASAP7_75t_L g1164 ( 
.A1(n_1151),
.A2(n_470),
.B1(n_104),
.B2(n_106),
.Y(n_1164)
);

INVx2_ASAP7_75t_L g1165 ( 
.A(n_1151),
.Y(n_1165)
);

OAI21x1_ASAP7_75t_L g1166 ( 
.A1(n_1151),
.A2(n_97),
.B(n_107),
.Y(n_1166)
);

XNOR2xp5_ASAP7_75t_L g1167 ( 
.A(n_1162),
.B(n_108),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_1156),
.Y(n_1168)
);

NAND4xp25_ASAP7_75t_L g1169 ( 
.A(n_1163),
.B(n_109),
.C(n_110),
.D(n_112),
.Y(n_1169)
);

INVx1_ASAP7_75t_SL g1170 ( 
.A(n_1165),
.Y(n_1170)
);

OAI322xp33_ASAP7_75t_L g1171 ( 
.A1(n_1155),
.A2(n_113),
.A3(n_115),
.B1(n_116),
.B2(n_117),
.C1(n_119),
.C2(n_121),
.Y(n_1171)
);

O2A1O1Ixp33_ASAP7_75t_L g1172 ( 
.A1(n_1159),
.A2(n_122),
.B(n_123),
.C(n_124),
.Y(n_1172)
);

NAND4xp25_ASAP7_75t_L g1173 ( 
.A(n_1157),
.B(n_125),
.C(n_126),
.D(n_129),
.Y(n_1173)
);

XNOR2xp5_ASAP7_75t_L g1174 ( 
.A(n_1166),
.B(n_1161),
.Y(n_1174)
);

NAND5xp2_ASAP7_75t_L g1175 ( 
.A(n_1158),
.B(n_130),
.C(n_131),
.D(n_132),
.E(n_133),
.Y(n_1175)
);

AOI21xp5_ASAP7_75t_L g1176 ( 
.A1(n_1168),
.A2(n_1164),
.B(n_1160),
.Y(n_1176)
);

AOI221xp5_ASAP7_75t_L g1177 ( 
.A1(n_1170),
.A2(n_134),
.B1(n_135),
.B2(n_136),
.C(n_137),
.Y(n_1177)
);

AOI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_1174),
.A2(n_138),
.B(n_139),
.Y(n_1178)
);

OR2x2_ASAP7_75t_L g1179 ( 
.A(n_1175),
.B(n_140),
.Y(n_1179)
);

OAI22x1_ASAP7_75t_L g1180 ( 
.A1(n_1172),
.A2(n_142),
.B1(n_144),
.B2(n_145),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_1173),
.B(n_1167),
.Y(n_1181)
);

AOI222xp33_ASAP7_75t_SL g1182 ( 
.A1(n_1171),
.A2(n_147),
.B1(n_148),
.B2(n_149),
.C1(n_150),
.C2(n_151),
.Y(n_1182)
);

AOI22xp33_ASAP7_75t_L g1183 ( 
.A1(n_1181),
.A2(n_1169),
.B1(n_154),
.B2(n_155),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_1176),
.B(n_153),
.Y(n_1184)
);

OAI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_1179),
.A2(n_1180),
.B(n_1182),
.Y(n_1185)
);

NAND3xp33_ASAP7_75t_L g1186 ( 
.A(n_1178),
.B(n_156),
.C(n_157),
.Y(n_1186)
);

AOI21xp5_ASAP7_75t_L g1187 ( 
.A1(n_1185),
.A2(n_1177),
.B(n_159),
.Y(n_1187)
);

OR2x6_ASAP7_75t_L g1188 ( 
.A(n_1187),
.B(n_1186),
.Y(n_1188)
);

OR2x2_ASAP7_75t_L g1189 ( 
.A(n_1188),
.B(n_1183),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_1189),
.Y(n_1190)
);

AO21x2_ASAP7_75t_L g1191 ( 
.A1(n_1190),
.A2(n_1184),
.B(n_160),
.Y(n_1191)
);

AOI221xp5_ASAP7_75t_L g1192 ( 
.A1(n_1191),
.A2(n_158),
.B1(n_161),
.B2(n_162),
.C(n_163),
.Y(n_1192)
);

AOI21xp33_ASAP7_75t_SL g1193 ( 
.A1(n_1192),
.A2(n_164),
.B(n_166),
.Y(n_1193)
);

AOI21xp5_ASAP7_75t_L g1194 ( 
.A1(n_1193),
.A2(n_966),
.B(n_171),
.Y(n_1194)
);

AOI211xp5_ASAP7_75t_L g1195 ( 
.A1(n_1194),
.A2(n_169),
.B(n_174),
.C(n_175),
.Y(n_1195)
);

AOI211xp5_ASAP7_75t_L g1196 ( 
.A1(n_1195),
.A2(n_176),
.B(n_177),
.C(n_178),
.Y(n_1196)
);


endmodule