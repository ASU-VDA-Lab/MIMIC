module fake_jpeg_25203_n_101 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_101);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_101;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_SL g11 ( 
.A(n_3),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

INVx11_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx24_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_15),
.A2(n_0),
.B1(n_1),
.B2(n_4),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_24),
.A2(n_28),
.B1(n_19),
.B2(n_14),
.Y(n_45)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_25),
.B(n_33),
.Y(n_40)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_11),
.B(n_5),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_27),
.B(n_31),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g28 ( 
.A1(n_18),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_28)
);

BUFx4f_ASAP7_75t_SL g29 ( 
.A(n_23),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_29),
.Y(n_37)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_30),
.B(n_13),
.Y(n_42)
);

A2O1A1Ixp33_ASAP7_75t_L g31 ( 
.A1(n_21),
.A2(n_7),
.B(n_10),
.C(n_17),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_32),
.Y(n_34)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_36),
.B(n_41),
.Y(n_47)
);

BUFx12_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx13_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_42),
.A2(n_45),
.B1(n_19),
.B2(n_22),
.Y(n_58)
);

BUFx12_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

CKINVDCx16_ASAP7_75t_R g50 ( 
.A(n_43),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_24),
.B(n_11),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_44),
.B(n_46),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_33),
.B(n_20),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_35),
.B(n_22),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_48),
.B(n_53),
.Y(n_61)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_51),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_44),
.A2(n_30),
.B1(n_26),
.B2(n_25),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_52),
.A2(n_58),
.B1(n_39),
.B2(n_16),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_37),
.B(n_14),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_42),
.B(n_13),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_54),
.B(n_57),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_42),
.B(n_17),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_55),
.B(n_49),
.Y(n_68)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_56),
.Y(n_67)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_53),
.B(n_23),
.Y(n_60)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_60),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_51),
.B(n_23),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_63),
.B(n_64),
.Y(n_75)
);

BUFx24_ASAP7_75t_SL g64 ( 
.A(n_49),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_47),
.B(n_36),
.Y(n_66)
);

XNOR2xp5_ASAP7_75t_L g73 ( 
.A(n_66),
.B(n_65),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_SL g79 ( 
.A1(n_68),
.A2(n_70),
.B(n_50),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_69),
.A2(n_39),
.B1(n_54),
.B2(n_57),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_58),
.B(n_16),
.Y(n_70)
);

XOR2xp5_ASAP7_75t_L g71 ( 
.A(n_65),
.B(n_52),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_L g85 ( 
.A(n_71),
.B(n_78),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_73),
.B(n_76),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_74),
.A2(n_61),
.B1(n_50),
.B2(n_59),
.Y(n_80)
);

AO21x1_ASAP7_75t_L g76 ( 
.A1(n_66),
.A2(n_54),
.B(n_69),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_67),
.Y(n_77)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_77),
.Y(n_81)
);

XOR2xp5_ASAP7_75t_L g78 ( 
.A(n_62),
.B(n_56),
.Y(n_78)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_79),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_SL g88 ( 
.A1(n_80),
.A2(n_75),
.B(n_43),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_78),
.B(n_38),
.C(n_43),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_82),
.B(n_38),
.C(n_59),
.Y(n_91)
);

BUFx12_ASAP7_75t_L g83 ( 
.A(n_71),
.Y(n_83)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_83),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_86),
.A2(n_84),
.B1(n_72),
.B2(n_76),
.Y(n_87)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_87),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_88),
.B(n_90),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_81),
.B(n_85),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_91),
.B(n_82),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_93),
.B(n_83),
.Y(n_96)
);

A2O1A1Ixp33_ASAP7_75t_L g95 ( 
.A1(n_92),
.A2(n_94),
.B(n_89),
.C(n_85),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_95),
.Y(n_98)
);

INVxp33_ASAP7_75t_L g99 ( 
.A(n_96),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_93),
.B(n_91),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_99),
.B(n_97),
.C(n_83),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_100),
.B(n_98),
.Y(n_101)
);


endmodule