module fake_netlist_6_3984_n_1765 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_77, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1765);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_77;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1765;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_155;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_163;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_928;
wire n_835;
wire n_1214;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1757;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_161;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_153;
wire n_842;
wire n_1707;
wire n_1432;
wire n_156;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_154;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_683;
wire n_474;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_162;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_171;
wire n_1764;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_159;
wire n_1086;
wire n_1066;
wire n_157;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1321;
wire n_1241;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_545;
wire n_489;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_158;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

BUFx10_ASAP7_75t_L g153 ( 
.A(n_131),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_87),
.Y(n_154)
);

INVx1_ASAP7_75t_SL g155 ( 
.A(n_136),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_47),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_17),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_54),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_89),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_60),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_49),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_99),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_38),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_26),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_13),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_148),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_73),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_7),
.Y(n_168)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_108),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_93),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_111),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_3),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_85),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_114),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_18),
.Y(n_175)
);

BUFx3_ASAP7_75t_L g176 ( 
.A(n_63),
.Y(n_176)
);

BUFx10_ASAP7_75t_L g177 ( 
.A(n_19),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_8),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_33),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_21),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_45),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_47),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_48),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_101),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_119),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_84),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_19),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_121),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_128),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_117),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_97),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_110),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_127),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_28),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_8),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_75),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_62),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_49),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_15),
.Y(n_199)
);

BUFx3_ASAP7_75t_L g200 ( 
.A(n_79),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g201 ( 
.A(n_100),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_30),
.Y(n_202)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_26),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_130),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_42),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_22),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_17),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_112),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_115),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_12),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_31),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_129),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_23),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_96),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_13),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_40),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_45),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_24),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_80),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_150),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_6),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_25),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_41),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_66),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_34),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_72),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_126),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_55),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_40),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_10),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_104),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_132),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_106),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_46),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_69),
.Y(n_235)
);

BUFx2_ASAP7_75t_L g236 ( 
.A(n_6),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_71),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_134),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_32),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_50),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_9),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_146),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_57),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_27),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_120),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_50),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_35),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_7),
.Y(n_248)
);

BUFx2_ASAP7_75t_L g249 ( 
.A(n_124),
.Y(n_249)
);

BUFx8_ASAP7_75t_SL g250 ( 
.A(n_0),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_147),
.Y(n_251)
);

CKINVDCx14_ASAP7_75t_R g252 ( 
.A(n_51),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_94),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_33),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_102),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_1),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_76),
.Y(n_257)
);

INVx2_ASAP7_75t_SL g258 ( 
.A(n_95),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_116),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_78),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_46),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_27),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_34),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_107),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_149),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_15),
.Y(n_266)
);

BUFx10_ASAP7_75t_L g267 ( 
.A(n_23),
.Y(n_267)
);

CKINVDCx16_ASAP7_75t_R g268 ( 
.A(n_53),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_83),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_5),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_105),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_138),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_65),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_32),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_91),
.Y(n_275)
);

HB1xp67_ASAP7_75t_L g276 ( 
.A(n_109),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_135),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_74),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_14),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_35),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_38),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_141),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_143),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_64),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_140),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_3),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_88),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_16),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_92),
.Y(n_289)
);

INVx1_ASAP7_75t_SL g290 ( 
.A(n_52),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_59),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_82),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_68),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_67),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_42),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_48),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_122),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_30),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_118),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_58),
.Y(n_300)
);

CKINVDCx16_ASAP7_75t_R g301 ( 
.A(n_145),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_123),
.Y(n_302)
);

CKINVDCx14_ASAP7_75t_R g303 ( 
.A(n_5),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_81),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_90),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_14),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_20),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_250),
.Y(n_308)
);

HB1xp67_ASAP7_75t_L g309 ( 
.A(n_236),
.Y(n_309)
);

INVxp67_ASAP7_75t_SL g310 ( 
.A(n_276),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_189),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_178),
.Y(n_312)
);

CKINVDCx16_ASAP7_75t_R g313 ( 
.A(n_303),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_191),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_178),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_178),
.Y(n_316)
);

INVxp67_ASAP7_75t_L g317 ( 
.A(n_161),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_170),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_192),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_178),
.Y(n_320)
);

INVx1_ASAP7_75t_SL g321 ( 
.A(n_165),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_178),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_194),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_194),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_193),
.Y(n_325)
);

CKINVDCx16_ASAP7_75t_R g326 ( 
.A(n_201),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_214),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_194),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_194),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_197),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_194),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_223),
.Y(n_332)
);

INVxp67_ASAP7_75t_L g333 ( 
.A(n_175),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_204),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_223),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_223),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_223),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_223),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_209),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_203),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_203),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_203),
.Y(n_342)
);

INVxp67_ASAP7_75t_SL g343 ( 
.A(n_249),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_212),
.Y(n_344)
);

INVxp33_ASAP7_75t_L g345 ( 
.A(n_183),
.Y(n_345)
);

INVxp67_ASAP7_75t_SL g346 ( 
.A(n_176),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_219),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_230),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_230),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_234),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_220),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_234),
.Y(n_352)
);

INVxp67_ASAP7_75t_SL g353 ( 
.A(n_176),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_271),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_296),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_296),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_272),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_214),
.Y(n_358)
);

INVxp67_ASAP7_75t_L g359 ( 
.A(n_177),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_298),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_287),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_298),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_187),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_198),
.Y(n_364)
);

INVxp67_ASAP7_75t_SL g365 ( 
.A(n_200),
.Y(n_365)
);

INVxp33_ASAP7_75t_L g366 ( 
.A(n_199),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_207),
.Y(n_367)
);

BUFx2_ASAP7_75t_L g368 ( 
.A(n_156),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_294),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_211),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_227),
.Y(n_371)
);

INVxp67_ASAP7_75t_SL g372 ( 
.A(n_200),
.Y(n_372)
);

INVxp33_ASAP7_75t_L g373 ( 
.A(n_215),
.Y(n_373)
);

HB1xp67_ASAP7_75t_L g374 ( 
.A(n_156),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_228),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_268),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_231),
.Y(n_377)
);

INVxp67_ASAP7_75t_L g378 ( 
.A(n_216),
.Y(n_378)
);

INVxp33_ASAP7_75t_SL g379 ( 
.A(n_157),
.Y(n_379)
);

HB1xp67_ASAP7_75t_L g380 ( 
.A(n_157),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_312),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_312),
.Y(n_382)
);

AND2x4_ASAP7_75t_L g383 ( 
.A(n_340),
.B(n_341),
.Y(n_383)
);

AND2x2_ASAP7_75t_L g384 ( 
.A(n_346),
.B(n_252),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_315),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_311),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_314),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_319),
.Y(n_388)
);

AND2x4_ASAP7_75t_L g389 ( 
.A(n_340),
.B(n_258),
.Y(n_389)
);

INVxp67_ASAP7_75t_L g390 ( 
.A(n_380),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_327),
.Y(n_391)
);

BUFx3_ASAP7_75t_L g392 ( 
.A(n_315),
.Y(n_392)
);

HB1xp67_ASAP7_75t_L g393 ( 
.A(n_374),
.Y(n_393)
);

OA21x2_ASAP7_75t_L g394 ( 
.A1(n_327),
.A2(n_221),
.B(n_217),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_316),
.Y(n_395)
);

INVxp67_ASAP7_75t_L g396 ( 
.A(n_368),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_316),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_320),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_353),
.B(n_258),
.Y(n_399)
);

AND2x2_ASAP7_75t_L g400 ( 
.A(n_365),
.B(n_169),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_327),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_343),
.B(n_301),
.Y(n_402)
);

BUFx6f_ASAP7_75t_L g403 ( 
.A(n_358),
.Y(n_403)
);

AND2x2_ASAP7_75t_L g404 ( 
.A(n_372),
.B(n_169),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_320),
.Y(n_405)
);

NAND2xp33_ASAP7_75t_L g406 ( 
.A(n_325),
.B(n_163),
.Y(n_406)
);

AND2x2_ASAP7_75t_L g407 ( 
.A(n_341),
.B(n_342),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_322),
.Y(n_408)
);

BUFx6f_ASAP7_75t_L g409 ( 
.A(n_358),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_322),
.Y(n_410)
);

CKINVDCx16_ASAP7_75t_R g411 ( 
.A(n_313),
.Y(n_411)
);

BUFx6f_ASAP7_75t_L g412 ( 
.A(n_358),
.Y(n_412)
);

BUFx6f_ASAP7_75t_L g413 ( 
.A(n_323),
.Y(n_413)
);

BUFx2_ASAP7_75t_L g414 ( 
.A(n_376),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_323),
.Y(n_415)
);

AND2x2_ASAP7_75t_SL g416 ( 
.A(n_326),
.B(n_224),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_324),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_324),
.Y(n_418)
);

OAI21x1_ASAP7_75t_L g419 ( 
.A1(n_342),
.A2(n_233),
.B(n_224),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_328),
.B(n_158),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_328),
.Y(n_421)
);

AND2x4_ASAP7_75t_L g422 ( 
.A(n_329),
.B(n_233),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_329),
.Y(n_423)
);

CKINVDCx16_ASAP7_75t_R g424 ( 
.A(n_313),
.Y(n_424)
);

INVx3_ASAP7_75t_L g425 ( 
.A(n_331),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_331),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_332),
.Y(n_427)
);

BUFx3_ASAP7_75t_L g428 ( 
.A(n_332),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_335),
.Y(n_429)
);

CKINVDCx8_ASAP7_75t_R g430 ( 
.A(n_326),
.Y(n_430)
);

AND2x4_ASAP7_75t_L g431 ( 
.A(n_335),
.B(n_154),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_336),
.Y(n_432)
);

AND2x2_ASAP7_75t_L g433 ( 
.A(n_336),
.B(n_159),
.Y(n_433)
);

NAND2x1_ASAP7_75t_L g434 ( 
.A(n_337),
.B(n_214),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_L g435 ( 
.A1(n_310),
.A2(n_248),
.B1(n_256),
.B2(n_262),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_337),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_318),
.Y(n_437)
);

AND2x2_ASAP7_75t_L g438 ( 
.A(n_338),
.B(n_167),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_330),
.Y(n_439)
);

INVx3_ASAP7_75t_L g440 ( 
.A(n_338),
.Y(n_440)
);

XNOR2x2_ASAP7_75t_L g441 ( 
.A(n_321),
.B(n_222),
.Y(n_441)
);

AND2x2_ASAP7_75t_L g442 ( 
.A(n_348),
.B(n_171),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_363),
.Y(n_443)
);

HB1xp67_ASAP7_75t_L g444 ( 
.A(n_368),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_R g445 ( 
.A(n_334),
.B(n_235),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_418),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_394),
.Y(n_447)
);

AO22x2_ASAP7_75t_L g448 ( 
.A1(n_396),
.A2(n_306),
.B1(n_295),
.B2(n_247),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_394),
.Y(n_449)
);

INVx2_ASAP7_75t_SL g450 ( 
.A(n_384),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_SL g451 ( 
.A1(n_435),
.A2(n_369),
.B1(n_361),
.B2(n_357),
.Y(n_451)
);

INVx1_ASAP7_75t_SL g452 ( 
.A(n_437),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_394),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_384),
.B(n_339),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_394),
.Y(n_455)
);

INVx4_ASAP7_75t_L g456 ( 
.A(n_413),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_394),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_392),
.Y(n_458)
);

INVx3_ASAP7_75t_L g459 ( 
.A(n_403),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_418),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_418),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_432),
.Y(n_462)
);

BUFx4f_ASAP7_75t_L g463 ( 
.A(n_431),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_392),
.Y(n_464)
);

INVxp67_ASAP7_75t_SL g465 ( 
.A(n_392),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_428),
.Y(n_466)
);

INVx2_ASAP7_75t_SL g467 ( 
.A(n_384),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_416),
.B(n_344),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_428),
.Y(n_469)
);

NOR3xp33_ASAP7_75t_L g470 ( 
.A(n_396),
.B(n_321),
.C(n_402),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_432),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_445),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_428),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_432),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_381),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_381),
.Y(n_476)
);

NOR3xp33_ASAP7_75t_L g477 ( 
.A(n_402),
.B(n_359),
.C(n_279),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_382),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_382),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_385),
.Y(n_480)
);

INVxp33_ASAP7_75t_SL g481 ( 
.A(n_445),
.Y(n_481)
);

OR2x6_ASAP7_75t_L g482 ( 
.A(n_390),
.B(n_399),
.Y(n_482)
);

AO21x2_ASAP7_75t_L g483 ( 
.A1(n_419),
.A2(n_188),
.B(n_186),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_385),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_386),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_SL g486 ( 
.A(n_416),
.B(n_347),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_395),
.Y(n_487)
);

INVx3_ASAP7_75t_L g488 ( 
.A(n_403),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_395),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_397),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_SL g491 ( 
.A(n_416),
.B(n_351),
.Y(n_491)
);

BUFx6f_ASAP7_75t_L g492 ( 
.A(n_403),
.Y(n_492)
);

AOI22xp5_ASAP7_75t_L g493 ( 
.A1(n_406),
.A2(n_377),
.B1(n_375),
.B2(n_371),
.Y(n_493)
);

CKINVDCx16_ASAP7_75t_R g494 ( 
.A(n_411),
.Y(n_494)
);

NOR2x1p5_ASAP7_75t_L g495 ( 
.A(n_387),
.B(n_308),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_397),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_398),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_398),
.Y(n_498)
);

BUFx3_ASAP7_75t_L g499 ( 
.A(n_431),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_405),
.Y(n_500)
);

AND2x2_ASAP7_75t_SL g501 ( 
.A(n_400),
.B(n_214),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_405),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_408),
.Y(n_503)
);

INVx8_ASAP7_75t_L g504 ( 
.A(n_431),
.Y(n_504)
);

AOI22xp33_ASAP7_75t_L g505 ( 
.A1(n_400),
.A2(n_309),
.B1(n_379),
.B2(n_225),
.Y(n_505)
);

BUFx8_ASAP7_75t_SL g506 ( 
.A(n_414),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_408),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_410),
.Y(n_508)
);

INVx4_ASAP7_75t_L g509 ( 
.A(n_413),
.Y(n_509)
);

BUFx3_ASAP7_75t_L g510 ( 
.A(n_431),
.Y(n_510)
);

AOI21x1_ASAP7_75t_L g511 ( 
.A1(n_434),
.A2(n_196),
.B(n_190),
.Y(n_511)
);

OR2x6_ASAP7_75t_L g512 ( 
.A(n_390),
.B(n_317),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_410),
.Y(n_513)
);

BUFx3_ASAP7_75t_L g514 ( 
.A(n_431),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_415),
.Y(n_515)
);

INVx3_ASAP7_75t_L g516 ( 
.A(n_403),
.Y(n_516)
);

INVxp67_ASAP7_75t_L g517 ( 
.A(n_444),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_415),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_417),
.Y(n_519)
);

BUFx10_ASAP7_75t_L g520 ( 
.A(n_388),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_417),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_439),
.B(n_345),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_SL g523 ( 
.A(n_411),
.B(n_153),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_421),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_421),
.Y(n_525)
);

INVxp33_ASAP7_75t_L g526 ( 
.A(n_444),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_423),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_SL g528 ( 
.A(n_424),
.B(n_153),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_423),
.Y(n_529)
);

INVx3_ASAP7_75t_L g530 ( 
.A(n_403),
.Y(n_530)
);

OAI21xp33_ASAP7_75t_SL g531 ( 
.A1(n_399),
.A2(n_286),
.B(n_263),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_426),
.Y(n_532)
);

INVx3_ASAP7_75t_L g533 ( 
.A(n_403),
.Y(n_533)
);

AND2x4_ASAP7_75t_L g534 ( 
.A(n_400),
.B(n_363),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_426),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_427),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_420),
.B(n_366),
.Y(n_537)
);

INVx2_ASAP7_75t_SL g538 ( 
.A(n_404),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_427),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_429),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_R g541 ( 
.A(n_424),
.B(n_354),
.Y(n_541)
);

AOI22xp33_ASAP7_75t_L g542 ( 
.A1(n_404),
.A2(n_389),
.B1(n_442),
.B2(n_433),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_429),
.Y(n_543)
);

INVx3_ASAP7_75t_L g544 ( 
.A(n_403),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_436),
.Y(n_545)
);

AND2x2_ASAP7_75t_L g546 ( 
.A(n_404),
.B(n_348),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_436),
.Y(n_547)
);

INVx8_ASAP7_75t_L g548 ( 
.A(n_389),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_SL g549 ( 
.A(n_430),
.B(n_153),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_430),
.Y(n_550)
);

AOI22xp33_ASAP7_75t_L g551 ( 
.A1(n_389),
.A2(n_378),
.B1(n_317),
.B2(n_333),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_L g552 ( 
.A(n_420),
.B(n_373),
.Y(n_552)
);

INVx3_ASAP7_75t_L g553 ( 
.A(n_409),
.Y(n_553)
);

INVx3_ASAP7_75t_L g554 ( 
.A(n_409),
.Y(n_554)
);

INVx3_ASAP7_75t_L g555 ( 
.A(n_409),
.Y(n_555)
);

BUFx3_ASAP7_75t_L g556 ( 
.A(n_433),
.Y(n_556)
);

BUFx6f_ASAP7_75t_L g557 ( 
.A(n_409),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_407),
.Y(n_558)
);

NOR2xp33_ASAP7_75t_L g559 ( 
.A(n_393),
.B(n_333),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_433),
.B(n_438),
.Y(n_560)
);

INVx8_ASAP7_75t_L g561 ( 
.A(n_389),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_430),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_L g563 ( 
.A(n_393),
.B(n_378),
.Y(n_563)
);

AND2x4_ASAP7_75t_L g564 ( 
.A(n_442),
.B(n_438),
.Y(n_564)
);

AOI22xp33_ASAP7_75t_L g565 ( 
.A1(n_389),
.A2(n_214),
.B1(n_370),
.B2(n_364),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_407),
.Y(n_566)
);

BUFx6f_ASAP7_75t_L g567 ( 
.A(n_409),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_414),
.Y(n_568)
);

NOR2xp33_ASAP7_75t_L g569 ( 
.A(n_443),
.B(n_155),
.Y(n_569)
);

AND2x4_ASAP7_75t_L g570 ( 
.A(n_442),
.B(n_208),
.Y(n_570)
);

BUFx10_ASAP7_75t_L g571 ( 
.A(n_383),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_SL g572 ( 
.A(n_435),
.B(n_158),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_SL g573 ( 
.A(n_383),
.B(n_160),
.Y(n_573)
);

OR2x2_ASAP7_75t_L g574 ( 
.A(n_441),
.B(n_364),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_407),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_422),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_425),
.Y(n_577)
);

BUFx3_ASAP7_75t_L g578 ( 
.A(n_438),
.Y(n_578)
);

CKINVDCx20_ASAP7_75t_R g579 ( 
.A(n_443),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_425),
.Y(n_580)
);

BUFx2_ASAP7_75t_L g581 ( 
.A(n_441),
.Y(n_581)
);

INVx4_ASAP7_75t_L g582 ( 
.A(n_413),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_425),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_422),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_422),
.Y(n_585)
);

AOI22xp5_ASAP7_75t_L g586 ( 
.A1(n_383),
.A2(n_265),
.B1(n_185),
.B2(n_184),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_425),
.Y(n_587)
);

AOI22xp33_ASAP7_75t_L g588 ( 
.A1(n_383),
.A2(n_370),
.B1(n_367),
.B2(n_292),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_440),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_440),
.Y(n_590)
);

BUFx6f_ASAP7_75t_L g591 ( 
.A(n_409),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_SL g592 ( 
.A(n_383),
.B(n_160),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_440),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_SL g594 ( 
.A(n_501),
.B(n_290),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_501),
.B(n_538),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_501),
.B(n_422),
.Y(n_596)
);

OAI221xp5_ASAP7_75t_L g597 ( 
.A1(n_538),
.A2(n_182),
.B1(n_242),
.B2(n_245),
.C(n_289),
.Y(n_597)
);

NOR2xp67_ASAP7_75t_L g598 ( 
.A(n_472),
.B(n_238),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_558),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_SL g600 ( 
.A(n_450),
.B(n_467),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_537),
.B(n_552),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_542),
.B(n_422),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_475),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_558),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_566),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_475),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_L g607 ( 
.A(n_450),
.B(n_441),
.Y(n_607)
);

INVxp67_ASAP7_75t_SL g608 ( 
.A(n_447),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_SL g609 ( 
.A(n_564),
.B(n_226),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_SL g610 ( 
.A(n_564),
.B(n_232),
.Y(n_610)
);

BUFx6f_ASAP7_75t_L g611 ( 
.A(n_499),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_566),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_SL g613 ( 
.A(n_467),
.B(n_162),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_575),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_575),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_SL g616 ( 
.A(n_472),
.B(n_162),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_479),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_479),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_564),
.B(n_440),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_564),
.B(n_413),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_458),
.Y(n_621)
);

AOI22xp5_ASAP7_75t_L g622 ( 
.A1(n_468),
.A2(n_251),
.B1(n_282),
.B2(n_283),
.Y(n_622)
);

INVx2_ASAP7_75t_SL g623 ( 
.A(n_546),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_SL g624 ( 
.A(n_560),
.B(n_237),
.Y(n_624)
);

INVxp67_ASAP7_75t_L g625 ( 
.A(n_522),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_556),
.B(n_578),
.Y(n_626)
);

INVx2_ASAP7_75t_SL g627 ( 
.A(n_546),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_490),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_556),
.B(n_413),
.Y(n_629)
);

NAND2xp33_ASAP7_75t_L g630 ( 
.A(n_548),
.B(n_284),
.Y(n_630)
);

AOI22xp33_ASAP7_75t_L g631 ( 
.A1(n_581),
.A2(n_419),
.B1(n_299),
.B2(n_253),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_578),
.B(n_413),
.Y(n_632)
);

AND2x6_ASAP7_75t_SL g633 ( 
.A(n_559),
.B(n_563),
.Y(n_633)
);

NOR2x1p5_ASAP7_75t_L g634 ( 
.A(n_574),
.B(n_163),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_L g635 ( 
.A(n_482),
.B(n_166),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_465),
.B(n_413),
.Y(n_636)
);

AOI22xp5_ASAP7_75t_L g637 ( 
.A1(n_486),
.A2(n_285),
.B1(n_291),
.B2(n_293),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_SL g638 ( 
.A(n_499),
.B(n_243),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_458),
.B(n_255),
.Y(n_639)
);

INVxp67_ASAP7_75t_L g640 ( 
.A(n_512),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_464),
.Y(n_641)
);

NOR2xp33_ASAP7_75t_L g642 ( 
.A(n_482),
.B(n_166),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_464),
.B(n_264),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_466),
.B(n_304),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_490),
.Y(n_645)
);

INVxp33_ASAP7_75t_L g646 ( 
.A(n_526),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_466),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_496),
.Y(n_648)
);

HB1xp67_ASAP7_75t_L g649 ( 
.A(n_517),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_469),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_469),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_SL g652 ( 
.A(n_481),
.B(n_173),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_473),
.B(n_305),
.Y(n_653)
);

INVx8_ASAP7_75t_L g654 ( 
.A(n_482),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_473),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_534),
.B(n_409),
.Y(n_656)
);

AOI21xp5_ASAP7_75t_L g657 ( 
.A1(n_463),
.A2(n_434),
.B(n_419),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_534),
.B(n_412),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_SL g659 ( 
.A(n_510),
.B(n_514),
.Y(n_659)
);

OR2x2_ASAP7_75t_L g660 ( 
.A(n_512),
.B(n_367),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_496),
.Y(n_661)
);

NOR2xp33_ASAP7_75t_SL g662 ( 
.A(n_481),
.B(n_173),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_576),
.Y(n_663)
);

INVx2_ASAP7_75t_SL g664 ( 
.A(n_534),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_497),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_576),
.B(n_412),
.Y(n_666)
);

INVxp67_ASAP7_75t_L g667 ( 
.A(n_512),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_584),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_584),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_497),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_SL g671 ( 
.A(n_510),
.B(n_174),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_585),
.B(n_412),
.Y(n_672)
);

OAI22xp5_ASAP7_75t_SL g673 ( 
.A1(n_581),
.A2(n_180),
.B1(n_181),
.B2(n_179),
.Y(n_673)
);

OAI22xp33_ASAP7_75t_L g674 ( 
.A1(n_574),
.A2(n_180),
.B1(n_181),
.B2(n_179),
.Y(n_674)
);

O2A1O1Ixp33_ASAP7_75t_L g675 ( 
.A1(n_447),
.A2(n_349),
.B(n_350),
.C(n_352),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_498),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_449),
.B(n_453),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_498),
.Y(n_678)
);

AOI22xp33_ASAP7_75t_L g679 ( 
.A1(n_449),
.A2(n_266),
.B1(n_172),
.B2(n_168),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_514),
.Y(n_680)
);

AOI22xp33_ASAP7_75t_L g681 ( 
.A1(n_453),
.A2(n_266),
.B1(n_172),
.B2(n_168),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_513),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_476),
.Y(n_683)
);

INVx2_ASAP7_75t_SL g684 ( 
.A(n_482),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_476),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_513),
.Y(n_686)
);

NOR2xp33_ASAP7_75t_L g687 ( 
.A(n_454),
.B(n_174),
.Y(n_687)
);

BUFx6f_ASAP7_75t_L g688 ( 
.A(n_571),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_478),
.Y(n_689)
);

BUFx6f_ASAP7_75t_L g690 ( 
.A(n_571),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_478),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_519),
.Y(n_692)
);

NAND2xp33_ASAP7_75t_L g693 ( 
.A(n_548),
.B(n_184),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_455),
.B(n_412),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_480),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_455),
.B(n_457),
.Y(n_696)
);

INVx3_ASAP7_75t_L g697 ( 
.A(n_571),
.Y(n_697)
);

AOI21xp5_ASAP7_75t_L g698 ( 
.A1(n_463),
.A2(n_401),
.B(n_391),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_SL g699 ( 
.A(n_463),
.B(n_185),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_SL g700 ( 
.A(n_457),
.B(n_257),
.Y(n_700)
);

NOR2xp67_ASAP7_75t_SL g701 ( 
.A(n_492),
.B(n_257),
.Y(n_701)
);

BUFx5_ASAP7_75t_L g702 ( 
.A(n_480),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_484),
.B(n_412),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_484),
.Y(n_704)
);

NOR3xp33_ASAP7_75t_L g705 ( 
.A(n_491),
.B(n_195),
.C(n_202),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_487),
.B(n_412),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_487),
.B(n_412),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_489),
.Y(n_708)
);

INVx4_ASAP7_75t_L g709 ( 
.A(n_504),
.Y(n_709)
);

AOI22xp33_ASAP7_75t_L g710 ( 
.A1(n_448),
.A2(n_270),
.B1(n_261),
.B2(n_164),
.Y(n_710)
);

BUFx3_ASAP7_75t_L g711 ( 
.A(n_520),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_485),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_500),
.B(n_391),
.Y(n_713)
);

OAI221xp5_ASAP7_75t_L g714 ( 
.A1(n_531),
.A2(n_205),
.B1(n_206),
.B2(n_210),
.C(n_213),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_519),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_500),
.B(n_401),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_SL g717 ( 
.A(n_493),
.B(n_259),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_502),
.B(n_401),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_502),
.B(n_259),
.Y(n_719)
);

NOR2xp33_ASAP7_75t_L g720 ( 
.A(n_572),
.B(n_260),
.Y(n_720)
);

AND2x2_ASAP7_75t_L g721 ( 
.A(n_512),
.B(n_177),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_521),
.Y(n_722)
);

NOR2xp33_ASAP7_75t_L g723 ( 
.A(n_586),
.B(n_260),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_521),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_503),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_503),
.B(n_265),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_507),
.B(n_269),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_507),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_525),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_508),
.B(n_269),
.Y(n_730)
);

NOR2xp33_ASAP7_75t_L g731 ( 
.A(n_549),
.B(n_273),
.Y(n_731)
);

NOR2xp67_ASAP7_75t_L g732 ( 
.A(n_485),
.B(n_273),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_525),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_508),
.B(n_275),
.Y(n_734)
);

OR2x6_ASAP7_75t_L g735 ( 
.A(n_451),
.B(n_349),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_515),
.B(n_275),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_515),
.Y(n_737)
);

INVx2_ASAP7_75t_SL g738 ( 
.A(n_579),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_527),
.Y(n_739)
);

BUFx3_ASAP7_75t_L g740 ( 
.A(n_520),
.Y(n_740)
);

NAND2x1p5_ASAP7_75t_L g741 ( 
.A(n_570),
.B(n_350),
.Y(n_741)
);

AOI22xp33_ASAP7_75t_SL g742 ( 
.A1(n_550),
.A2(n_177),
.B1(n_267),
.B2(n_164),
.Y(n_742)
);

AOI22xp33_ASAP7_75t_L g743 ( 
.A1(n_448),
.A2(n_261),
.B1(n_270),
.B2(n_274),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_SL g744 ( 
.A(n_569),
.B(n_277),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_SL g745 ( 
.A(n_470),
.B(n_278),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_518),
.B(n_278),
.Y(n_746)
);

AND2x2_ASAP7_75t_L g747 ( 
.A(n_551),
.B(n_267),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_524),
.B(n_297),
.Y(n_748)
);

NOR2xp33_ASAP7_75t_L g749 ( 
.A(n_573),
.B(n_297),
.Y(n_749)
);

AND2x4_ASAP7_75t_L g750 ( 
.A(n_570),
.B(n_352),
.Y(n_750)
);

INVxp67_ASAP7_75t_L g751 ( 
.A(n_477),
.Y(n_751)
);

AND2x2_ASAP7_75t_SL g752 ( 
.A(n_494),
.B(n_362),
.Y(n_752)
);

NOR2xp33_ASAP7_75t_L g753 ( 
.A(n_592),
.B(n_300),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_527),
.Y(n_754)
);

CKINVDCx11_ASAP7_75t_R g755 ( 
.A(n_520),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_536),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_536),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_524),
.Y(n_758)
);

AOI22xp5_ASAP7_75t_L g759 ( 
.A1(n_570),
.A2(n_302),
.B1(n_229),
.B2(n_239),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_529),
.B(n_302),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_532),
.B(n_280),
.Y(n_761)
);

INVx2_ASAP7_75t_SL g762 ( 
.A(n_660),
.Y(n_762)
);

OR2x6_ASAP7_75t_L g763 ( 
.A(n_654),
.B(n_495),
.Y(n_763)
);

BUFx3_ASAP7_75t_L g764 ( 
.A(n_712),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_SL g765 ( 
.A(n_702),
.B(n_550),
.Y(n_765)
);

BUFx2_ASAP7_75t_L g766 ( 
.A(n_738),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_SL g767 ( 
.A(n_702),
.B(n_562),
.Y(n_767)
);

NOR2xp33_ASAP7_75t_L g768 ( 
.A(n_601),
.B(n_562),
.Y(n_768)
);

AOI22xp33_ASAP7_75t_L g769 ( 
.A1(n_607),
.A2(n_679),
.B1(n_681),
.B2(n_594),
.Y(n_769)
);

AOI22xp5_ASAP7_75t_L g770 ( 
.A1(n_659),
.A2(n_570),
.B1(n_548),
.B2(n_561),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_663),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_755),
.Y(n_772)
);

INVx5_ASAP7_75t_L g773 ( 
.A(n_688),
.Y(n_773)
);

BUFx6f_ASAP7_75t_L g774 ( 
.A(n_688),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_603),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_668),
.Y(n_776)
);

NOR2xp33_ASAP7_75t_L g777 ( 
.A(n_625),
.B(n_607),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_669),
.Y(n_778)
);

OR2x6_ASAP7_75t_L g779 ( 
.A(n_654),
.B(n_711),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_603),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_606),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_SL g782 ( 
.A(n_702),
.B(n_548),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_608),
.B(n_532),
.Y(n_783)
);

INVx1_ASAP7_75t_SL g784 ( 
.A(n_646),
.Y(n_784)
);

OR2x6_ASAP7_75t_SL g785 ( 
.A(n_761),
.B(n_568),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_606),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_599),
.B(n_535),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_711),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_617),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_617),
.Y(n_790)
);

INVxp67_ASAP7_75t_L g791 ( 
.A(n_649),
.Y(n_791)
);

BUFx2_ASAP7_75t_L g792 ( 
.A(n_752),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_618),
.Y(n_793)
);

INVx3_ASAP7_75t_L g794 ( 
.A(n_611),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_SL g795 ( 
.A(n_702),
.B(n_548),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_618),
.Y(n_796)
);

AND2x6_ASAP7_75t_L g797 ( 
.A(n_595),
.B(n_577),
.Y(n_797)
);

NOR2x2_ASAP7_75t_L g798 ( 
.A(n_735),
.B(n_494),
.Y(n_798)
);

HB1xp67_ASAP7_75t_L g799 ( 
.A(n_626),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_628),
.Y(n_800)
);

NOR2x2_ASAP7_75t_L g801 ( 
.A(n_735),
.B(n_541),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_628),
.Y(n_802)
);

AND2x4_ASAP7_75t_L g803 ( 
.A(n_664),
.B(n_623),
.Y(n_803)
);

BUFx4f_ASAP7_75t_SL g804 ( 
.A(n_740),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_604),
.B(n_535),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_605),
.B(n_612),
.Y(n_806)
);

INVx2_ASAP7_75t_SL g807 ( 
.A(n_634),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_614),
.B(n_543),
.Y(n_808)
);

CKINVDCx5p33_ASAP7_75t_R g809 ( 
.A(n_740),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_645),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_615),
.B(n_543),
.Y(n_811)
);

NAND2xp33_ASAP7_75t_L g812 ( 
.A(n_688),
.B(n_561),
.Y(n_812)
);

NOR2xp33_ASAP7_75t_L g813 ( 
.A(n_751),
.B(n_523),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_683),
.B(n_545),
.Y(n_814)
);

AO22x1_ASAP7_75t_L g815 ( 
.A1(n_723),
.A2(n_568),
.B1(n_274),
.B2(n_307),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_645),
.Y(n_816)
);

AND2x4_ASAP7_75t_L g817 ( 
.A(n_627),
.B(n_684),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_648),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_648),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_685),
.B(n_545),
.Y(n_820)
);

NOR2xp33_ASAP7_75t_L g821 ( 
.A(n_633),
.B(n_528),
.Y(n_821)
);

INVx3_ASAP7_75t_L g822 ( 
.A(n_611),
.Y(n_822)
);

CKINVDCx5p33_ASAP7_75t_R g823 ( 
.A(n_752),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_661),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_661),
.Y(n_825)
);

INVx3_ASAP7_75t_L g826 ( 
.A(n_611),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_665),
.Y(n_827)
);

NOR2xp33_ASAP7_75t_L g828 ( 
.A(n_687),
.B(n_600),
.Y(n_828)
);

NOR2xp33_ASAP7_75t_L g829 ( 
.A(n_687),
.B(n_505),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_SL g830 ( 
.A(n_702),
.B(n_561),
.Y(n_830)
);

INVx2_ASAP7_75t_SL g831 ( 
.A(n_721),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_665),
.Y(n_832)
);

NOR2xp33_ASAP7_75t_L g833 ( 
.A(n_640),
.B(n_452),
.Y(n_833)
);

INVx5_ASAP7_75t_L g834 ( 
.A(n_688),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_670),
.Y(n_835)
);

AND2x2_ASAP7_75t_SL g836 ( 
.A(n_631),
.B(n_565),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_689),
.B(n_561),
.Y(n_837)
);

AND2x6_ASAP7_75t_SL g838 ( 
.A(n_735),
.B(n_506),
.Y(n_838)
);

NAND3xp33_ASAP7_75t_SL g839 ( 
.A(n_720),
.B(n_307),
.C(n_218),
.Y(n_839)
);

NAND3xp33_ASAP7_75t_SL g840 ( 
.A(n_720),
.B(n_254),
.C(n_241),
.Y(n_840)
);

CKINVDCx5p33_ASAP7_75t_R g841 ( 
.A(n_654),
.Y(n_841)
);

BUFx3_ASAP7_75t_L g842 ( 
.A(n_750),
.Y(n_842)
);

INVx5_ASAP7_75t_L g843 ( 
.A(n_690),
.Y(n_843)
);

BUFx6f_ASAP7_75t_L g844 ( 
.A(n_690),
.Y(n_844)
);

AND2x2_ASAP7_75t_L g845 ( 
.A(n_747),
.B(n_448),
.Y(n_845)
);

CKINVDCx8_ASAP7_75t_R g846 ( 
.A(n_635),
.Y(n_846)
);

AND2x4_ASAP7_75t_L g847 ( 
.A(n_750),
.B(n_611),
.Y(n_847)
);

NOR2xp33_ASAP7_75t_L g848 ( 
.A(n_667),
.B(n_539),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_691),
.B(n_561),
.Y(n_849)
);

INVxp67_ASAP7_75t_SL g850 ( 
.A(n_677),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_SL g851 ( 
.A(n_702),
.B(n_577),
.Y(n_851)
);

NOR2xp33_ASAP7_75t_L g852 ( 
.A(n_662),
.B(n_539),
.Y(n_852)
);

BUFx6f_ASAP7_75t_L g853 ( 
.A(n_690),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_SL g854 ( 
.A(n_690),
.B(n_580),
.Y(n_854)
);

NAND2x1p5_ASAP7_75t_L g855 ( 
.A(n_709),
.B(n_540),
.Y(n_855)
);

BUFx3_ASAP7_75t_L g856 ( 
.A(n_741),
.Y(n_856)
);

INVx2_ASAP7_75t_SL g857 ( 
.A(n_613),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_676),
.Y(n_858)
);

NOR2x1p5_ASAP7_75t_L g859 ( 
.A(n_719),
.B(n_240),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_695),
.B(n_540),
.Y(n_860)
);

BUFx6f_ASAP7_75t_L g861 ( 
.A(n_659),
.Y(n_861)
);

OAI22xp5_ASAP7_75t_L g862 ( 
.A1(n_596),
.A2(n_588),
.B1(n_504),
.B2(n_547),
.Y(n_862)
);

OR2x2_ASAP7_75t_L g863 ( 
.A(n_616),
.B(n_495),
.Y(n_863)
);

HB1xp67_ASAP7_75t_L g864 ( 
.A(n_680),
.Y(n_864)
);

AOI22xp33_ASAP7_75t_L g865 ( 
.A1(n_679),
.A2(n_448),
.B1(n_483),
.B2(n_547),
.Y(n_865)
);

CKINVDCx20_ASAP7_75t_R g866 ( 
.A(n_652),
.Y(n_866)
);

INVx1_ASAP7_75t_SL g867 ( 
.A(n_726),
.Y(n_867)
);

AOI21xp5_ASAP7_75t_L g868 ( 
.A1(n_694),
.A2(n_504),
.B(n_509),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_704),
.B(n_580),
.Y(n_869)
);

CKINVDCx5p33_ASAP7_75t_R g870 ( 
.A(n_731),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_708),
.B(n_583),
.Y(n_871)
);

BUFx8_ASAP7_75t_L g872 ( 
.A(n_725),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_676),
.Y(n_873)
);

AOI22xp5_ASAP7_75t_L g874 ( 
.A1(n_594),
.A2(n_609),
.B1(n_610),
.B2(n_624),
.Y(n_874)
);

OAI22xp5_ASAP7_75t_SL g875 ( 
.A1(n_742),
.A2(n_244),
.B1(n_246),
.B2(n_281),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_678),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_678),
.Y(n_877)
);

BUFx6f_ASAP7_75t_L g878 ( 
.A(n_697),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_682),
.Y(n_879)
);

AND2x4_ASAP7_75t_L g880 ( 
.A(n_728),
.B(n_593),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_682),
.Y(n_881)
);

BUFx6f_ASAP7_75t_L g882 ( 
.A(n_697),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_686),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_686),
.Y(n_884)
);

OR2x2_ASAP7_75t_L g885 ( 
.A(n_745),
.B(n_483),
.Y(n_885)
);

BUFx6f_ASAP7_75t_L g886 ( 
.A(n_709),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_737),
.B(n_583),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_758),
.B(n_587),
.Y(n_888)
);

HB1xp67_ASAP7_75t_L g889 ( 
.A(n_741),
.Y(n_889)
);

INVx3_ASAP7_75t_L g890 ( 
.A(n_692),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_692),
.Y(n_891)
);

OR2x6_ASAP7_75t_L g892 ( 
.A(n_732),
.B(n_504),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_715),
.Y(n_893)
);

BUFx2_ASAP7_75t_L g894 ( 
.A(n_727),
.Y(n_894)
);

BUFx3_ASAP7_75t_L g895 ( 
.A(n_621),
.Y(n_895)
);

INVx2_ASAP7_75t_SL g896 ( 
.A(n_730),
.Y(n_896)
);

AOI22xp33_ASAP7_75t_L g897 ( 
.A1(n_681),
.A2(n_483),
.B1(n_593),
.B2(n_590),
.Y(n_897)
);

AND2x6_ASAP7_75t_SL g898 ( 
.A(n_723),
.B(n_355),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_715),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_SL g900 ( 
.A(n_619),
.B(n_620),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_722),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_722),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_SL g903 ( 
.A(n_696),
.B(n_656),
.Y(n_903)
);

INVx2_ASAP7_75t_SL g904 ( 
.A(n_734),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_724),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_724),
.Y(n_906)
);

A2O1A1Ixp33_ASAP7_75t_SL g907 ( 
.A1(n_701),
.A2(n_714),
.B(n_675),
.C(n_749),
.Y(n_907)
);

NOR2xp33_ASAP7_75t_L g908 ( 
.A(n_731),
.B(n_587),
.Y(n_908)
);

AND2x2_ASAP7_75t_L g909 ( 
.A(n_635),
.B(n_267),
.Y(n_909)
);

AOI22xp5_ASAP7_75t_L g910 ( 
.A1(n_609),
.A2(n_610),
.B1(n_624),
.B2(n_753),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_641),
.B(n_589),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_647),
.B(n_589),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_729),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_729),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_SL g915 ( 
.A(n_658),
.B(n_590),
.Y(n_915)
);

BUFx3_ASAP7_75t_L g916 ( 
.A(n_642),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_733),
.Y(n_917)
);

INVx2_ASAP7_75t_L g918 ( 
.A(n_733),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_650),
.B(n_651),
.Y(n_919)
);

CKINVDCx5p33_ASAP7_75t_R g920 ( 
.A(n_642),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_739),
.Y(n_921)
);

INVx3_ASAP7_75t_L g922 ( 
.A(n_739),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_754),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_754),
.Y(n_924)
);

INVxp67_ASAP7_75t_L g925 ( 
.A(n_736),
.Y(n_925)
);

NOR2xp33_ASAP7_75t_L g926 ( 
.A(n_744),
.B(n_288),
.Y(n_926)
);

AOI22xp33_ASAP7_75t_L g927 ( 
.A1(n_631),
.A2(n_461),
.B1(n_462),
.B2(n_471),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_SL g928 ( 
.A(n_602),
.B(n_459),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_756),
.Y(n_929)
);

BUFx2_ASAP7_75t_L g930 ( 
.A(n_746),
.Y(n_930)
);

AOI21xp5_ASAP7_75t_L g931 ( 
.A1(n_629),
.A2(n_504),
.B(n_582),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_756),
.Y(n_932)
);

AND3x2_ASAP7_75t_SL g933 ( 
.A(n_710),
.B(n_0),
.C(n_1),
.Y(n_933)
);

CKINVDCx5p33_ASAP7_75t_R g934 ( 
.A(n_717),
.Y(n_934)
);

AOI22xp33_ASAP7_75t_L g935 ( 
.A1(n_710),
.A2(n_743),
.B1(n_700),
.B2(n_673),
.Y(n_935)
);

AND2x4_ASAP7_75t_L g936 ( 
.A(n_655),
.B(n_355),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_757),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_SL g938 ( 
.A(n_757),
.B(n_459),
.Y(n_938)
);

INVx4_ASAP7_75t_L g939 ( 
.A(n_598),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_749),
.B(n_459),
.Y(n_940)
);

INVxp67_ASAP7_75t_L g941 ( 
.A(n_748),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_SL g942 ( 
.A(n_632),
.B(n_488),
.Y(n_942)
);

INVx2_ASAP7_75t_L g943 ( 
.A(n_703),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_753),
.B(n_488),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_706),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_SL g946 ( 
.A(n_657),
.B(n_488),
.Y(n_946)
);

NAND2xp33_ASAP7_75t_SL g947 ( 
.A(n_870),
.B(n_743),
.Y(n_947)
);

OAI22xp33_ASAP7_75t_L g948 ( 
.A1(n_829),
.A2(n_777),
.B1(n_910),
.B2(n_850),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_850),
.B(n_760),
.Y(n_949)
);

NAND3xp33_ASAP7_75t_L g950 ( 
.A(n_829),
.B(n_705),
.C(n_622),
.Y(n_950)
);

HB1xp67_ASAP7_75t_L g951 ( 
.A(n_784),
.Y(n_951)
);

O2A1O1Ixp33_ASAP7_75t_L g952 ( 
.A1(n_777),
.A2(n_597),
.B(n_671),
.C(n_700),
.Y(n_952)
);

NOR2xp33_ASAP7_75t_L g953 ( 
.A(n_768),
.B(n_674),
.Y(n_953)
);

AND2x4_ASAP7_75t_L g954 ( 
.A(n_847),
.B(n_671),
.Y(n_954)
);

NOR2xp33_ASAP7_75t_L g955 ( 
.A(n_768),
.B(n_759),
.Y(n_955)
);

CKINVDCx5p33_ASAP7_75t_R g956 ( 
.A(n_764),
.Y(n_956)
);

AOI22xp33_ASAP7_75t_L g957 ( 
.A1(n_769),
.A2(n_638),
.B1(n_644),
.B2(n_639),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_828),
.B(n_699),
.Y(n_958)
);

INVx3_ASAP7_75t_L g959 ( 
.A(n_774),
.Y(n_959)
);

O2A1O1Ixp33_ASAP7_75t_L g960 ( 
.A1(n_839),
.A2(n_638),
.B(n_699),
.C(n_653),
.Y(n_960)
);

AOI21xp5_ASAP7_75t_L g961 ( 
.A1(n_946),
.A2(n_630),
.B(n_636),
.Y(n_961)
);

AOI21xp5_ASAP7_75t_L g962 ( 
.A1(n_946),
.A2(n_693),
.B(n_672),
.Y(n_962)
);

INVx2_ASAP7_75t_L g963 ( 
.A(n_890),
.Y(n_963)
);

AOI21xp5_ASAP7_75t_L g964 ( 
.A1(n_868),
.A2(n_666),
.B(n_698),
.Y(n_964)
);

INVx3_ASAP7_75t_L g965 ( 
.A(n_774),
.Y(n_965)
);

NOR2xp33_ASAP7_75t_L g966 ( 
.A(n_925),
.B(n_637),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_SL g967 ( 
.A(n_867),
.B(n_643),
.Y(n_967)
);

A2O1A1Ixp33_ASAP7_75t_SL g968 ( 
.A1(n_852),
.A2(n_530),
.B(n_516),
.C(n_533),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_SL g969 ( 
.A(n_828),
.B(n_707),
.Y(n_969)
);

O2A1O1Ixp5_ASAP7_75t_L g970 ( 
.A1(n_940),
.A2(n_718),
.B(n_716),
.C(n_713),
.Y(n_970)
);

AOI21xp5_ASAP7_75t_L g971 ( 
.A1(n_903),
.A2(n_456),
.B(n_582),
.Y(n_971)
);

CKINVDCx6p67_ASAP7_75t_R g972 ( 
.A(n_763),
.Y(n_972)
);

AOI21xp5_ASAP7_75t_L g973 ( 
.A1(n_903),
.A2(n_456),
.B(n_582),
.Y(n_973)
);

NAND3xp33_ASAP7_75t_L g974 ( 
.A(n_769),
.B(n_356),
.C(n_360),
.Y(n_974)
);

CKINVDCx14_ASAP7_75t_R g975 ( 
.A(n_772),
.Y(n_975)
);

AND2x2_ASAP7_75t_L g976 ( 
.A(n_792),
.B(n_356),
.Y(n_976)
);

AOI22xp33_ASAP7_75t_L g977 ( 
.A1(n_935),
.A2(n_462),
.B1(n_471),
.B2(n_446),
.Y(n_977)
);

BUFx6f_ASAP7_75t_L g978 ( 
.A(n_774),
.Y(n_978)
);

BUFx2_ASAP7_75t_L g979 ( 
.A(n_766),
.Y(n_979)
);

AOI22xp33_ASAP7_75t_L g980 ( 
.A1(n_935),
.A2(n_446),
.B1(n_460),
.B2(n_461),
.Y(n_980)
);

NOR2xp33_ASAP7_75t_L g981 ( 
.A(n_925),
.B(n_516),
.Y(n_981)
);

OR2x6_ASAP7_75t_L g982 ( 
.A(n_779),
.B(n_456),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_799),
.B(n_530),
.Y(n_983)
);

HB1xp67_ASAP7_75t_L g984 ( 
.A(n_799),
.Y(n_984)
);

AOI21xp5_ASAP7_75t_L g985 ( 
.A1(n_773),
.A2(n_509),
.B(n_567),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_941),
.B(n_530),
.Y(n_986)
);

INVx2_ASAP7_75t_L g987 ( 
.A(n_890),
.Y(n_987)
);

BUFx2_ASAP7_75t_L g988 ( 
.A(n_791),
.Y(n_988)
);

AOI21xp5_ASAP7_75t_L g989 ( 
.A1(n_773),
.A2(n_509),
.B(n_567),
.Y(n_989)
);

BUFx12f_ASAP7_75t_L g990 ( 
.A(n_872),
.Y(n_990)
);

A2O1A1Ixp33_ASAP7_75t_L g991 ( 
.A1(n_874),
.A2(n_926),
.B(n_941),
.C(n_813),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_771),
.Y(n_992)
);

AOI22xp33_ASAP7_75t_L g993 ( 
.A1(n_836),
.A2(n_460),
.B1(n_474),
.B2(n_360),
.Y(n_993)
);

BUFx6f_ASAP7_75t_L g994 ( 
.A(n_774),
.Y(n_994)
);

AOI22xp5_ASAP7_75t_L g995 ( 
.A1(n_840),
.A2(n_544),
.B1(n_533),
.B2(n_553),
.Y(n_995)
);

O2A1O1Ixp5_ASAP7_75t_L g996 ( 
.A1(n_944),
.A2(n_511),
.B(n_474),
.C(n_553),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_896),
.B(n_904),
.Y(n_997)
);

HB1xp67_ASAP7_75t_L g998 ( 
.A(n_791),
.Y(n_998)
);

O2A1O1Ixp33_ASAP7_75t_L g999 ( 
.A1(n_840),
.A2(n_554),
.B(n_555),
.C(n_9),
.Y(n_999)
);

INVx2_ASAP7_75t_L g1000 ( 
.A(n_922),
.Y(n_1000)
);

OAI22xp5_ASAP7_75t_L g1001 ( 
.A1(n_836),
.A2(n_555),
.B1(n_554),
.B2(n_557),
.Y(n_1001)
);

CKINVDCx20_ASAP7_75t_R g1002 ( 
.A(n_804),
.Y(n_1002)
);

INVx5_ASAP7_75t_L g1003 ( 
.A(n_886),
.Y(n_1003)
);

AOI21xp5_ASAP7_75t_L g1004 ( 
.A1(n_773),
.A2(n_591),
.B(n_567),
.Y(n_1004)
);

O2A1O1Ixp33_ASAP7_75t_L g1005 ( 
.A1(n_926),
.A2(n_2),
.B(n_4),
.C(n_10),
.Y(n_1005)
);

INVx2_ASAP7_75t_L g1006 ( 
.A(n_922),
.Y(n_1006)
);

OR2x6_ASAP7_75t_SL g1007 ( 
.A(n_920),
.B(n_788),
.Y(n_1007)
);

AND2x2_ASAP7_75t_L g1008 ( 
.A(n_845),
.B(n_2),
.Y(n_1008)
);

OAI22xp5_ASAP7_75t_L g1009 ( 
.A1(n_908),
.A2(n_591),
.B1(n_567),
.B2(n_557),
.Y(n_1009)
);

AOI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_834),
.A2(n_591),
.B(n_557),
.Y(n_1010)
);

BUFx6f_ASAP7_75t_L g1011 ( 
.A(n_844),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_776),
.Y(n_1012)
);

NOR2xp33_ASAP7_75t_L g1013 ( 
.A(n_894),
.B(n_4),
.Y(n_1013)
);

NAND3xp33_ASAP7_75t_L g1014 ( 
.A(n_815),
.B(n_557),
.C(n_492),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_SL g1015 ( 
.A(n_930),
.B(n_557),
.Y(n_1015)
);

A2O1A1Ixp33_ASAP7_75t_L g1016 ( 
.A1(n_852),
.A2(n_492),
.B(n_511),
.C(n_16),
.Y(n_1016)
);

NAND2xp33_ASAP7_75t_L g1017 ( 
.A(n_886),
.B(n_492),
.Y(n_1017)
);

A2O1A1Ixp33_ASAP7_75t_L g1018 ( 
.A1(n_908),
.A2(n_11),
.B(n_12),
.C(n_18),
.Y(n_1018)
);

O2A1O1Ixp33_ASAP7_75t_L g1019 ( 
.A1(n_907),
.A2(n_11),
.B(n_20),
.C(n_21),
.Y(n_1019)
);

INVx2_ASAP7_75t_L g1020 ( 
.A(n_775),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_806),
.B(n_22),
.Y(n_1021)
);

OAI22xp5_ASAP7_75t_L g1022 ( 
.A1(n_861),
.A2(n_77),
.B1(n_151),
.B2(n_144),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_778),
.B(n_24),
.Y(n_1023)
);

OAI22xp5_ASAP7_75t_L g1024 ( 
.A1(n_861),
.A2(n_70),
.B1(n_142),
.B2(n_139),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_786),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_787),
.B(n_25),
.Y(n_1026)
);

BUFx2_ASAP7_75t_L g1027 ( 
.A(n_823),
.Y(n_1027)
);

INVx2_ASAP7_75t_L g1028 ( 
.A(n_780),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_805),
.B(n_28),
.Y(n_1029)
);

INVx1_ASAP7_75t_SL g1030 ( 
.A(n_809),
.Y(n_1030)
);

A2O1A1Ixp33_ASAP7_75t_L g1031 ( 
.A1(n_857),
.A2(n_29),
.B(n_31),
.C(n_36),
.Y(n_1031)
);

CKINVDCx5p33_ASAP7_75t_R g1032 ( 
.A(n_838),
.Y(n_1032)
);

AOI21x1_ASAP7_75t_L g1033 ( 
.A1(n_854),
.A2(n_928),
.B(n_900),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_SL g1034 ( 
.A(n_834),
.B(n_86),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_789),
.Y(n_1035)
);

INVx2_ASAP7_75t_L g1036 ( 
.A(n_781),
.Y(n_1036)
);

OAI21xp5_ASAP7_75t_L g1037 ( 
.A1(n_885),
.A2(n_98),
.B(n_137),
.Y(n_1037)
);

CKINVDCx5p33_ASAP7_75t_R g1038 ( 
.A(n_841),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_808),
.B(n_29),
.Y(n_1039)
);

NOR2xp33_ASAP7_75t_L g1040 ( 
.A(n_916),
.B(n_36),
.Y(n_1040)
);

AOI21xp5_ASAP7_75t_L g1041 ( 
.A1(n_834),
.A2(n_843),
.B(n_812),
.Y(n_1041)
);

OAI22xp5_ASAP7_75t_L g1042 ( 
.A1(n_861),
.A2(n_783),
.B1(n_767),
.B2(n_765),
.Y(n_1042)
);

INVx2_ASAP7_75t_L g1043 ( 
.A(n_790),
.Y(n_1043)
);

INVx2_ASAP7_75t_L g1044 ( 
.A(n_793),
.Y(n_1044)
);

AOI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_843),
.A2(n_103),
.B(n_133),
.Y(n_1045)
);

BUFx3_ASAP7_75t_L g1046 ( 
.A(n_804),
.Y(n_1046)
);

NOR2xp33_ASAP7_75t_L g1047 ( 
.A(n_846),
.B(n_37),
.Y(n_1047)
);

OAI21xp33_ASAP7_75t_SL g1048 ( 
.A1(n_814),
.A2(n_37),
.B(n_39),
.Y(n_1048)
);

INVx2_ASAP7_75t_L g1049 ( 
.A(n_802),
.Y(n_1049)
);

O2A1O1Ixp33_ASAP7_75t_L g1050 ( 
.A1(n_811),
.A2(n_39),
.B(n_41),
.C(n_43),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_796),
.Y(n_1051)
);

BUFx2_ASAP7_75t_L g1052 ( 
.A(n_762),
.Y(n_1052)
);

AOI21xp5_ASAP7_75t_L g1053 ( 
.A1(n_843),
.A2(n_113),
.B(n_125),
.Y(n_1053)
);

AOI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_843),
.A2(n_56),
.B(n_61),
.Y(n_1054)
);

NAND2xp33_ASAP7_75t_SL g1055 ( 
.A(n_934),
.B(n_43),
.Y(n_1055)
);

AOI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_782),
.A2(n_152),
.B(n_44),
.Y(n_1056)
);

OR2x2_ASAP7_75t_L g1057 ( 
.A(n_833),
.B(n_44),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_820),
.B(n_848),
.Y(n_1058)
);

OAI22xp5_ASAP7_75t_L g1059 ( 
.A1(n_861),
.A2(n_767),
.B1(n_770),
.B2(n_895),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_848),
.B(n_943),
.Y(n_1060)
);

INVx2_ASAP7_75t_L g1061 ( 
.A(n_816),
.Y(n_1061)
);

A2O1A1Ixp33_ASAP7_75t_SL g1062 ( 
.A1(n_821),
.A2(n_822),
.B(n_794),
.C(n_826),
.Y(n_1062)
);

AOI21xp5_ASAP7_75t_L g1063 ( 
.A1(n_782),
.A2(n_795),
.B(n_830),
.Y(n_1063)
);

AOI21x1_ASAP7_75t_L g1064 ( 
.A1(n_942),
.A2(n_851),
.B(n_915),
.Y(n_1064)
);

AO22x1_ASAP7_75t_L g1065 ( 
.A1(n_821),
.A2(n_872),
.B1(n_933),
.B2(n_833),
.Y(n_1065)
);

OAI21x1_ASAP7_75t_L g1066 ( 
.A1(n_931),
.A2(n_915),
.B(n_942),
.Y(n_1066)
);

OAI22xp5_ASAP7_75t_L g1067 ( 
.A1(n_895),
.A2(n_889),
.B1(n_919),
.B2(n_856),
.Y(n_1067)
);

AOI21xp5_ASAP7_75t_L g1068 ( 
.A1(n_795),
.A2(n_830),
.B(n_837),
.Y(n_1068)
);

AOI22xp5_ASAP7_75t_L g1069 ( 
.A1(n_831),
.A2(n_866),
.B1(n_803),
.B2(n_859),
.Y(n_1069)
);

A2O1A1Ixp33_ASAP7_75t_L g1070 ( 
.A1(n_909),
.A2(n_860),
.B(n_865),
.C(n_849),
.Y(n_1070)
);

HB1xp67_ASAP7_75t_L g1071 ( 
.A(n_864),
.Y(n_1071)
);

O2A1O1Ixp33_ASAP7_75t_L g1072 ( 
.A1(n_864),
.A2(n_807),
.B(n_863),
.C(n_869),
.Y(n_1072)
);

INVx2_ASAP7_75t_L g1073 ( 
.A(n_818),
.Y(n_1073)
);

OAI22xp5_ASAP7_75t_L g1074 ( 
.A1(n_889),
.A2(n_897),
.B1(n_862),
.B2(n_886),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_800),
.Y(n_1075)
);

AOI21xp5_ASAP7_75t_L g1076 ( 
.A1(n_851),
.A2(n_945),
.B(n_855),
.Y(n_1076)
);

A2O1A1Ixp33_ASAP7_75t_L g1077 ( 
.A1(n_865),
.A2(n_803),
.B(n_880),
.C(n_897),
.Y(n_1077)
);

A2O1A1Ixp33_ASAP7_75t_L g1078 ( 
.A1(n_880),
.A2(n_817),
.B(n_887),
.C(n_888),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_SL g1079 ( 
.A(n_844),
.B(n_853),
.Y(n_1079)
);

AOI21xp5_ASAP7_75t_L g1080 ( 
.A1(n_855),
.A2(n_938),
.B(n_871),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_936),
.B(n_939),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_992),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_1012),
.Y(n_1083)
);

AO21x2_ASAP7_75t_L g1084 ( 
.A1(n_968),
.A2(n_912),
.B(n_911),
.Y(n_1084)
);

NOR2xp33_ASAP7_75t_L g1085 ( 
.A(n_955),
.B(n_953),
.Y(n_1085)
);

A2O1A1Ixp33_ASAP7_75t_L g1086 ( 
.A1(n_955),
.A2(n_817),
.B(n_936),
.C(n_842),
.Y(n_1086)
);

NOR2x1_ASAP7_75t_SL g1087 ( 
.A(n_1003),
.B(n_853),
.Y(n_1087)
);

INVx3_ASAP7_75t_L g1088 ( 
.A(n_1003),
.Y(n_1088)
);

AOI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_961),
.A2(n_892),
.B(n_882),
.Y(n_1089)
);

AOI22xp5_ASAP7_75t_L g1090 ( 
.A1(n_953),
.A2(n_875),
.B1(n_763),
.B2(n_779),
.Y(n_1090)
);

A2O1A1Ixp33_ASAP7_75t_L g1091 ( 
.A1(n_991),
.A2(n_877),
.B(n_917),
.C(n_914),
.Y(n_1091)
);

OAI21x1_ASAP7_75t_L g1092 ( 
.A1(n_964),
.A2(n_873),
.B(n_932),
.Y(n_1092)
);

OAI21xp5_ASAP7_75t_L g1093 ( 
.A1(n_1070),
.A2(n_927),
.B(n_797),
.Y(n_1093)
);

CKINVDCx8_ASAP7_75t_R g1094 ( 
.A(n_956),
.Y(n_1094)
);

AO31x2_ASAP7_75t_L g1095 ( 
.A1(n_1074),
.A2(n_905),
.A3(n_902),
.B(n_929),
.Y(n_1095)
);

OAI21x1_ASAP7_75t_L g1096 ( 
.A1(n_1066),
.A2(n_879),
.B(n_923),
.Y(n_1096)
);

OAI21x1_ASAP7_75t_SL g1097 ( 
.A1(n_1037),
.A2(n_937),
.B(n_893),
.Y(n_1097)
);

AOI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_962),
.A2(n_949),
.B(n_1068),
.Y(n_1098)
);

OAI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_958),
.A2(n_927),
.B(n_797),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_948),
.B(n_901),
.Y(n_1100)
);

AOI22xp5_ASAP7_75t_L g1101 ( 
.A1(n_947),
.A2(n_763),
.B1(n_779),
.B2(n_822),
.Y(n_1101)
);

OAI21x1_ASAP7_75t_L g1102 ( 
.A1(n_1064),
.A2(n_835),
.B(n_913),
.Y(n_1102)
);

OAI21x1_ASAP7_75t_L g1103 ( 
.A1(n_1033),
.A2(n_891),
.B(n_884),
.Y(n_1103)
);

OAI21x1_ASAP7_75t_L g1104 ( 
.A1(n_1076),
.A2(n_827),
.B(n_883),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_948),
.B(n_881),
.Y(n_1105)
);

CKINVDCx5p33_ASAP7_75t_R g1106 ( 
.A(n_1038),
.Y(n_1106)
);

OAI21x1_ASAP7_75t_SL g1107 ( 
.A1(n_1056),
.A2(n_858),
.B(n_924),
.Y(n_1107)
);

OAI21x1_ASAP7_75t_L g1108 ( 
.A1(n_971),
.A2(n_973),
.B(n_1080),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_1025),
.Y(n_1109)
);

INVx2_ASAP7_75t_L g1110 ( 
.A(n_1020),
.Y(n_1110)
);

OA21x2_ASAP7_75t_L g1111 ( 
.A1(n_996),
.A2(n_810),
.B(n_921),
.Y(n_1111)
);

AOI221x1_ASAP7_75t_L g1112 ( 
.A1(n_950),
.A2(n_933),
.B1(n_825),
.B2(n_824),
.C(n_826),
.Y(n_1112)
);

AOI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_1058),
.A2(n_892),
.B(n_882),
.Y(n_1113)
);

NOR2xp67_ASAP7_75t_R g1114 ( 
.A(n_1046),
.B(n_882),
.Y(n_1114)
);

NAND2xp33_ASAP7_75t_R g1115 ( 
.A(n_979),
.B(n_794),
.Y(n_1115)
);

OAI22xp5_ASAP7_75t_L g1116 ( 
.A1(n_1077),
.A2(n_878),
.B1(n_785),
.B2(n_876),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_1060),
.B(n_918),
.Y(n_1117)
);

BUFx2_ASAP7_75t_L g1118 ( 
.A(n_951),
.Y(n_1118)
);

AOI21xp5_ASAP7_75t_L g1119 ( 
.A1(n_1078),
.A2(n_878),
.B(n_906),
.Y(n_1119)
);

AND3x4_ASAP7_75t_L g1120 ( 
.A(n_1007),
.B(n_798),
.C(n_801),
.Y(n_1120)
);

AND2x4_ASAP7_75t_L g1121 ( 
.A(n_954),
.B(n_878),
.Y(n_1121)
);

BUFx3_ASAP7_75t_L g1122 ( 
.A(n_1002),
.Y(n_1122)
);

OAI22xp5_ASAP7_75t_L g1123 ( 
.A1(n_966),
.A2(n_878),
.B1(n_819),
.B2(n_832),
.Y(n_1123)
);

OAI22x1_ASAP7_75t_L g1124 ( 
.A1(n_1047),
.A2(n_1069),
.B1(n_1040),
.B2(n_966),
.Y(n_1124)
);

CKINVDCx11_ASAP7_75t_R g1125 ( 
.A(n_990),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_969),
.B(n_899),
.Y(n_1126)
);

INVxp67_ASAP7_75t_L g1127 ( 
.A(n_951),
.Y(n_1127)
);

NAND2xp33_ASAP7_75t_R g1128 ( 
.A(n_1027),
.B(n_898),
.Y(n_1128)
);

BUFx3_ASAP7_75t_L g1129 ( 
.A(n_988),
.Y(n_1129)
);

AOI21xp5_ASAP7_75t_L g1130 ( 
.A1(n_1003),
.A2(n_797),
.B(n_1042),
.Y(n_1130)
);

BUFx2_ASAP7_75t_L g1131 ( 
.A(n_1052),
.Y(n_1131)
);

OAI21x1_ASAP7_75t_SL g1132 ( 
.A1(n_1005),
.A2(n_797),
.B(n_1041),
.Y(n_1132)
);

NOR2xp33_ASAP7_75t_L g1133 ( 
.A(n_997),
.B(n_797),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_SL g1134 ( 
.A(n_998),
.B(n_1072),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_981),
.B(n_986),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_981),
.B(n_954),
.Y(n_1136)
);

AOI21xp5_ASAP7_75t_L g1137 ( 
.A1(n_1059),
.A2(n_970),
.B(n_1009),
.Y(n_1137)
);

AO21x2_ASAP7_75t_L g1138 ( 
.A1(n_1016),
.A2(n_960),
.B(n_1014),
.Y(n_1138)
);

AOI221x1_ASAP7_75t_L g1139 ( 
.A1(n_1018),
.A2(n_1055),
.B1(n_1031),
.B2(n_974),
.C(n_1067),
.Y(n_1139)
);

OAI21x1_ASAP7_75t_L g1140 ( 
.A1(n_996),
.A2(n_1001),
.B(n_970),
.Y(n_1140)
);

CKINVDCx11_ASAP7_75t_R g1141 ( 
.A(n_1030),
.Y(n_1141)
);

OAI221xp5_ASAP7_75t_L g1142 ( 
.A1(n_952),
.A2(n_1057),
.B1(n_1048),
.B2(n_1047),
.C(n_1013),
.Y(n_1142)
);

O2A1O1Ixp33_ASAP7_75t_L g1143 ( 
.A1(n_1019),
.A2(n_967),
.B(n_999),
.C(n_1050),
.Y(n_1143)
);

AOI211x1_ASAP7_75t_L g1144 ( 
.A1(n_1065),
.A2(n_1023),
.B(n_1008),
.C(n_1021),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_1035),
.B(n_1075),
.Y(n_1145)
);

OR2x2_ASAP7_75t_L g1146 ( 
.A(n_976),
.B(n_998),
.Y(n_1146)
);

NAND2x1_ASAP7_75t_L g1147 ( 
.A(n_978),
.B(n_1011),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_1051),
.B(n_984),
.Y(n_1148)
);

AOI21xp5_ASAP7_75t_L g1149 ( 
.A1(n_957),
.A2(n_1081),
.B(n_989),
.Y(n_1149)
);

NOR2xp33_ASAP7_75t_L g1150 ( 
.A(n_984),
.B(n_1071),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_957),
.B(n_1061),
.Y(n_1151)
);

OAI21x1_ASAP7_75t_L g1152 ( 
.A1(n_985),
.A2(n_1004),
.B(n_1010),
.Y(n_1152)
);

O2A1O1Ixp5_ASAP7_75t_L g1153 ( 
.A1(n_1026),
.A2(n_1039),
.B(n_1029),
.C(n_1015),
.Y(n_1153)
);

CKINVDCx20_ASAP7_75t_R g1154 ( 
.A(n_975),
.Y(n_1154)
);

INVx4_ASAP7_75t_L g1155 ( 
.A(n_978),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_1028),
.B(n_1036),
.Y(n_1156)
);

INVx3_ASAP7_75t_L g1157 ( 
.A(n_978),
.Y(n_1157)
);

HB1xp67_ASAP7_75t_L g1158 ( 
.A(n_1071),
.Y(n_1158)
);

O2A1O1Ixp33_ASAP7_75t_L g1159 ( 
.A1(n_1013),
.A2(n_1062),
.B(n_1022),
.C(n_1024),
.Y(n_1159)
);

BUFx2_ASAP7_75t_L g1160 ( 
.A(n_978),
.Y(n_1160)
);

BUFx2_ASAP7_75t_L g1161 ( 
.A(n_994),
.Y(n_1161)
);

NAND3x1_ASAP7_75t_L g1162 ( 
.A(n_1032),
.B(n_972),
.C(n_959),
.Y(n_1162)
);

OAI21x1_ASAP7_75t_L g1163 ( 
.A1(n_977),
.A2(n_980),
.B(n_993),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_L g1164 ( 
.A(n_1043),
.B(n_1044),
.Y(n_1164)
);

INVx2_ASAP7_75t_L g1165 ( 
.A(n_1049),
.Y(n_1165)
);

AOI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_1079),
.A2(n_983),
.B(n_1034),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_1073),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_993),
.B(n_963),
.Y(n_1168)
);

INVx5_ASAP7_75t_L g1169 ( 
.A(n_994),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_987),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_1000),
.Y(n_1171)
);

AOI22xp33_ASAP7_75t_SL g1172 ( 
.A1(n_994),
.A2(n_1011),
.B1(n_959),
.B2(n_965),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_1006),
.B(n_965),
.Y(n_1173)
);

NAND3x1_ASAP7_75t_L g1174 ( 
.A(n_1045),
.B(n_1053),
.C(n_1054),
.Y(n_1174)
);

OAI21x1_ASAP7_75t_L g1175 ( 
.A1(n_995),
.A2(n_982),
.B(n_1011),
.Y(n_1175)
);

OR2x2_ASAP7_75t_L g1176 ( 
.A(n_982),
.B(n_994),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_1011),
.B(n_948),
.Y(n_1177)
);

AOI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_1017),
.A2(n_961),
.B(n_812),
.Y(n_1178)
);

OAI21x1_ASAP7_75t_L g1179 ( 
.A1(n_964),
.A2(n_1066),
.B(n_1063),
.Y(n_1179)
);

OR2x2_ASAP7_75t_L g1180 ( 
.A(n_951),
.B(n_452),
.Y(n_1180)
);

AO21x2_ASAP7_75t_L g1181 ( 
.A1(n_968),
.A2(n_948),
.B(n_961),
.Y(n_1181)
);

O2A1O1Ixp5_ASAP7_75t_L g1182 ( 
.A1(n_953),
.A2(n_829),
.B(n_955),
.C(n_948),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_948),
.B(n_777),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_948),
.B(n_777),
.Y(n_1184)
);

OA21x2_ASAP7_75t_L g1185 ( 
.A1(n_1066),
.A2(n_1070),
.B(n_996),
.Y(n_1185)
);

OAI21xp5_ASAP7_75t_L g1186 ( 
.A1(n_991),
.A2(n_829),
.B(n_1070),
.Y(n_1186)
);

AOI21xp5_ASAP7_75t_SL g1187 ( 
.A1(n_1077),
.A2(n_709),
.B(n_886),
.Y(n_1187)
);

AO21x2_ASAP7_75t_L g1188 ( 
.A1(n_968),
.A2(n_948),
.B(n_961),
.Y(n_1188)
);

NAND2xp33_ASAP7_75t_L g1189 ( 
.A(n_991),
.B(n_870),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_992),
.Y(n_1190)
);

OAI21xp5_ASAP7_75t_SL g1191 ( 
.A1(n_953),
.A2(n_829),
.B(n_435),
.Y(n_1191)
);

AOI21xp5_ASAP7_75t_L g1192 ( 
.A1(n_1017),
.A2(n_961),
.B(n_812),
.Y(n_1192)
);

BUFx2_ASAP7_75t_L g1193 ( 
.A(n_951),
.Y(n_1193)
);

INVx3_ASAP7_75t_L g1194 ( 
.A(n_1003),
.Y(n_1194)
);

AO31x2_ASAP7_75t_L g1195 ( 
.A1(n_1074),
.A2(n_1042),
.A3(n_1070),
.B(n_1016),
.Y(n_1195)
);

AOI31xp67_ASAP7_75t_L g1196 ( 
.A1(n_969),
.A2(n_910),
.A3(n_874),
.B(n_700),
.Y(n_1196)
);

CKINVDCx5p33_ASAP7_75t_R g1197 ( 
.A(n_956),
.Y(n_1197)
);

OAI21x1_ASAP7_75t_L g1198 ( 
.A1(n_964),
.A2(n_1066),
.B(n_1063),
.Y(n_1198)
);

AOI21xp5_ASAP7_75t_L g1199 ( 
.A1(n_1017),
.A2(n_961),
.B(n_812),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_L g1200 ( 
.A(n_948),
.B(n_777),
.Y(n_1200)
);

OA22x2_ASAP7_75t_L g1201 ( 
.A1(n_1069),
.A2(n_581),
.B1(n_870),
.B2(n_435),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_948),
.B(n_777),
.Y(n_1202)
);

NAND3x1_ASAP7_75t_L g1203 ( 
.A(n_953),
.B(n_1047),
.C(n_829),
.Y(n_1203)
);

NOR2xp67_ASAP7_75t_R g1204 ( 
.A(n_1046),
.B(n_711),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_992),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_948),
.B(n_777),
.Y(n_1206)
);

INVx3_ASAP7_75t_L g1207 ( 
.A(n_1003),
.Y(n_1207)
);

OAI21x1_ASAP7_75t_SL g1208 ( 
.A1(n_1037),
.A2(n_1056),
.B(n_1005),
.Y(n_1208)
);

NOR2xp33_ASAP7_75t_L g1209 ( 
.A(n_955),
.B(n_768),
.Y(n_1209)
);

NAND2xp33_ASAP7_75t_L g1210 ( 
.A(n_991),
.B(n_870),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_SL g1211 ( 
.A(n_948),
.B(n_870),
.Y(n_1211)
);

AND2x2_ASAP7_75t_L g1212 ( 
.A(n_976),
.B(n_777),
.Y(n_1212)
);

INVx2_ASAP7_75t_SL g1213 ( 
.A(n_951),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_948),
.B(n_777),
.Y(n_1214)
);

OAI21x1_ASAP7_75t_L g1215 ( 
.A1(n_964),
.A2(n_1066),
.B(n_1063),
.Y(n_1215)
);

INVx2_ASAP7_75t_L g1216 ( 
.A(n_992),
.Y(n_1216)
);

OR2x2_ASAP7_75t_L g1217 ( 
.A(n_951),
.B(n_452),
.Y(n_1217)
);

NAND3xp33_ASAP7_75t_SL g1218 ( 
.A(n_955),
.B(n_870),
.C(n_829),
.Y(n_1218)
);

OAI21x1_ASAP7_75t_L g1219 ( 
.A1(n_964),
.A2(n_1066),
.B(n_1063),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_SL g1220 ( 
.A(n_948),
.B(n_870),
.Y(n_1220)
);

AO21x2_ASAP7_75t_L g1221 ( 
.A1(n_1137),
.A2(n_1186),
.B(n_1098),
.Y(n_1221)
);

NOR2xp33_ASAP7_75t_L g1222 ( 
.A(n_1085),
.B(n_1209),
.Y(n_1222)
);

OAI21x1_ASAP7_75t_L g1223 ( 
.A1(n_1092),
.A2(n_1096),
.B(n_1179),
.Y(n_1223)
);

AND2x4_ASAP7_75t_L g1224 ( 
.A(n_1121),
.B(n_1086),
.Y(n_1224)
);

INVx2_ASAP7_75t_L g1225 ( 
.A(n_1111),
.Y(n_1225)
);

BUFx2_ASAP7_75t_L g1226 ( 
.A(n_1129),
.Y(n_1226)
);

OAI21x1_ASAP7_75t_L g1227 ( 
.A1(n_1198),
.A2(n_1219),
.B(n_1215),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1216),
.Y(n_1228)
);

OAI21x1_ASAP7_75t_L g1229 ( 
.A1(n_1089),
.A2(n_1104),
.B(n_1152),
.Y(n_1229)
);

OA21x2_ASAP7_75t_L g1230 ( 
.A1(n_1140),
.A2(n_1186),
.B(n_1093),
.Y(n_1230)
);

BUFx6f_ASAP7_75t_L g1231 ( 
.A(n_1169),
.Y(n_1231)
);

INVx2_ASAP7_75t_L g1232 ( 
.A(n_1111),
.Y(n_1232)
);

OAI21x1_ASAP7_75t_L g1233 ( 
.A1(n_1108),
.A2(n_1192),
.B(n_1178),
.Y(n_1233)
);

AO21x2_ASAP7_75t_L g1234 ( 
.A1(n_1208),
.A2(n_1130),
.B(n_1132),
.Y(n_1234)
);

INVx2_ASAP7_75t_L g1235 ( 
.A(n_1102),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1082),
.Y(n_1236)
);

INVx2_ASAP7_75t_L g1237 ( 
.A(n_1103),
.Y(n_1237)
);

INVx1_ASAP7_75t_SL g1238 ( 
.A(n_1180),
.Y(n_1238)
);

INVx2_ASAP7_75t_L g1239 ( 
.A(n_1083),
.Y(n_1239)
);

OAI22xp33_ASAP7_75t_L g1240 ( 
.A1(n_1191),
.A2(n_1218),
.B1(n_1201),
.B2(n_1200),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_1190),
.Y(n_1241)
);

OAI22xp5_ASAP7_75t_L g1242 ( 
.A1(n_1203),
.A2(n_1220),
.B1(n_1211),
.B2(n_1142),
.Y(n_1242)
);

BUFx8_ASAP7_75t_L g1243 ( 
.A(n_1131),
.Y(n_1243)
);

AOI22xp33_ASAP7_75t_L g1244 ( 
.A1(n_1142),
.A2(n_1200),
.B1(n_1214),
.B2(n_1183),
.Y(n_1244)
);

AOI21xp5_ASAP7_75t_L g1245 ( 
.A1(n_1199),
.A2(n_1187),
.B(n_1093),
.Y(n_1245)
);

AND2x4_ASAP7_75t_L g1246 ( 
.A(n_1121),
.B(n_1176),
.Y(n_1246)
);

INVx5_ASAP7_75t_L g1247 ( 
.A(n_1169),
.Y(n_1247)
);

AO31x2_ASAP7_75t_L g1248 ( 
.A1(n_1112),
.A2(n_1149),
.A3(n_1091),
.B(n_1139),
.Y(n_1248)
);

BUFx6f_ASAP7_75t_L g1249 ( 
.A(n_1169),
.Y(n_1249)
);

BUFx6f_ASAP7_75t_L g1250 ( 
.A(n_1169),
.Y(n_1250)
);

AOI222xp33_ASAP7_75t_L g1251 ( 
.A1(n_1124),
.A2(n_1212),
.B1(n_1214),
.B2(n_1202),
.C1(n_1183),
.C2(n_1184),
.Y(n_1251)
);

NOR2x1_ASAP7_75t_SL g1252 ( 
.A(n_1134),
.B(n_1116),
.Y(n_1252)
);

OAI21x1_ASAP7_75t_L g1253 ( 
.A1(n_1174),
.A2(n_1175),
.B(n_1119),
.Y(n_1253)
);

INVxp67_ASAP7_75t_L g1254 ( 
.A(n_1150),
.Y(n_1254)
);

INVx2_ASAP7_75t_SL g1255 ( 
.A(n_1197),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1205),
.Y(n_1256)
);

INVx2_ASAP7_75t_L g1257 ( 
.A(n_1109),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1145),
.Y(n_1258)
);

INVx2_ASAP7_75t_SL g1259 ( 
.A(n_1106),
.Y(n_1259)
);

OAI21x1_ASAP7_75t_L g1260 ( 
.A1(n_1113),
.A2(n_1097),
.B(n_1107),
.Y(n_1260)
);

OAI21xp5_ASAP7_75t_L g1261 ( 
.A1(n_1182),
.A2(n_1153),
.B(n_1206),
.Y(n_1261)
);

AO21x2_ASAP7_75t_L g1262 ( 
.A1(n_1181),
.A2(n_1188),
.B(n_1138),
.Y(n_1262)
);

INVx2_ASAP7_75t_SL g1263 ( 
.A(n_1118),
.Y(n_1263)
);

AOI21x1_ASAP7_75t_L g1264 ( 
.A1(n_1116),
.A2(n_1105),
.B(n_1100),
.Y(n_1264)
);

CKINVDCx20_ASAP7_75t_R g1265 ( 
.A(n_1154),
.Y(n_1265)
);

INVx2_ASAP7_75t_L g1266 ( 
.A(n_1126),
.Y(n_1266)
);

AOI21xp5_ASAP7_75t_L g1267 ( 
.A1(n_1189),
.A2(n_1210),
.B(n_1099),
.Y(n_1267)
);

AOI22xp33_ASAP7_75t_SL g1268 ( 
.A1(n_1201),
.A2(n_1184),
.B1(n_1206),
.B2(n_1202),
.Y(n_1268)
);

INVx2_ASAP7_75t_L g1269 ( 
.A(n_1126),
.Y(n_1269)
);

AO21x1_ASAP7_75t_L g1270 ( 
.A1(n_1143),
.A2(n_1159),
.B(n_1135),
.Y(n_1270)
);

OAI21x1_ASAP7_75t_L g1271 ( 
.A1(n_1185),
.A2(n_1166),
.B(n_1163),
.Y(n_1271)
);

NOR2x1_ASAP7_75t_R g1272 ( 
.A(n_1125),
.B(n_1141),
.Y(n_1272)
);

BUFx3_ASAP7_75t_L g1273 ( 
.A(n_1193),
.Y(n_1273)
);

CKINVDCx20_ASAP7_75t_R g1274 ( 
.A(n_1094),
.Y(n_1274)
);

OA21x2_ASAP7_75t_L g1275 ( 
.A1(n_1100),
.A2(n_1105),
.B(n_1177),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_L g1276 ( 
.A(n_1146),
.B(n_1117),
.Y(n_1276)
);

OAI21x1_ASAP7_75t_L g1277 ( 
.A1(n_1151),
.A2(n_1123),
.B(n_1177),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1145),
.Y(n_1278)
);

AOI21xp5_ASAP7_75t_L g1279 ( 
.A1(n_1138),
.A2(n_1188),
.B(n_1181),
.Y(n_1279)
);

O2A1O1Ixp33_ASAP7_75t_L g1280 ( 
.A1(n_1127),
.A2(n_1136),
.B(n_1213),
.C(n_1217),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1148),
.Y(n_1281)
);

AOI22xp5_ASAP7_75t_L g1282 ( 
.A1(n_1128),
.A2(n_1090),
.B1(n_1120),
.B2(n_1101),
.Y(n_1282)
);

BUFx2_ASAP7_75t_R g1283 ( 
.A(n_1122),
.Y(n_1283)
);

BUFx6f_ASAP7_75t_L g1284 ( 
.A(n_1147),
.Y(n_1284)
);

OA21x2_ASAP7_75t_L g1285 ( 
.A1(n_1168),
.A2(n_1117),
.B(n_1133),
.Y(n_1285)
);

HB1xp67_ASAP7_75t_L g1286 ( 
.A(n_1158),
.Y(n_1286)
);

OAI22xp5_ASAP7_75t_L g1287 ( 
.A1(n_1144),
.A2(n_1148),
.B1(n_1167),
.B2(n_1162),
.Y(n_1287)
);

OAI21x1_ASAP7_75t_SL g1288 ( 
.A1(n_1087),
.A2(n_1173),
.B(n_1156),
.Y(n_1288)
);

OAI21x1_ASAP7_75t_L g1289 ( 
.A1(n_1173),
.A2(n_1164),
.B(n_1156),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1164),
.Y(n_1290)
);

INVx1_ASAP7_75t_SL g1291 ( 
.A(n_1160),
.Y(n_1291)
);

OAI21xp5_ASAP7_75t_L g1292 ( 
.A1(n_1196),
.A2(n_1165),
.B(n_1110),
.Y(n_1292)
);

OAI21x1_ASAP7_75t_L g1293 ( 
.A1(n_1157),
.A2(n_1207),
.B(n_1088),
.Y(n_1293)
);

OAI22xp5_ASAP7_75t_L g1294 ( 
.A1(n_1172),
.A2(n_1171),
.B1(n_1170),
.B2(n_1194),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1161),
.Y(n_1295)
);

CKINVDCx11_ASAP7_75t_R g1296 ( 
.A(n_1155),
.Y(n_1296)
);

OAI21x1_ASAP7_75t_L g1297 ( 
.A1(n_1157),
.A2(n_1207),
.B(n_1088),
.Y(n_1297)
);

CKINVDCx5p33_ASAP7_75t_R g1298 ( 
.A(n_1115),
.Y(n_1298)
);

BUFx2_ASAP7_75t_L g1299 ( 
.A(n_1155),
.Y(n_1299)
);

INVxp67_ASAP7_75t_L g1300 ( 
.A(n_1114),
.Y(n_1300)
);

BUFx6f_ASAP7_75t_L g1301 ( 
.A(n_1084),
.Y(n_1301)
);

AND2x4_ASAP7_75t_L g1302 ( 
.A(n_1195),
.B(n_1095),
.Y(n_1302)
);

INVx2_ASAP7_75t_L g1303 ( 
.A(n_1195),
.Y(n_1303)
);

BUFx12f_ASAP7_75t_L g1304 ( 
.A(n_1204),
.Y(n_1304)
);

NAND2x1p5_ASAP7_75t_L g1305 ( 
.A(n_1195),
.B(n_1003),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1216),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1216),
.Y(n_1307)
);

NOR2xp33_ASAP7_75t_L g1308 ( 
.A(n_1085),
.B(n_1209),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1216),
.Y(n_1309)
);

INVx2_ASAP7_75t_L g1310 ( 
.A(n_1111),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_L g1311 ( 
.A(n_1209),
.B(n_1085),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1216),
.Y(n_1312)
);

INVx2_ASAP7_75t_L g1313 ( 
.A(n_1111),
.Y(n_1313)
);

OAI221xp5_ASAP7_75t_L g1314 ( 
.A1(n_1191),
.A2(n_829),
.B1(n_1085),
.B2(n_1209),
.C(n_601),
.Y(n_1314)
);

OAI21xp5_ASAP7_75t_L g1315 ( 
.A1(n_1209),
.A2(n_1085),
.B(n_829),
.Y(n_1315)
);

INVxp67_ASAP7_75t_SL g1316 ( 
.A(n_1163),
.Y(n_1316)
);

NOR2xp33_ASAP7_75t_SL g1317 ( 
.A(n_1094),
.B(n_712),
.Y(n_1317)
);

NAND2x1p5_ASAP7_75t_L g1318 ( 
.A(n_1169),
.B(n_1003),
.Y(n_1318)
);

INVx6_ASAP7_75t_L g1319 ( 
.A(n_1169),
.Y(n_1319)
);

HB1xp67_ASAP7_75t_L g1320 ( 
.A(n_1158),
.Y(n_1320)
);

OAI21x1_ASAP7_75t_L g1321 ( 
.A1(n_1092),
.A2(n_1096),
.B(n_1179),
.Y(n_1321)
);

NOR2xp67_ASAP7_75t_SL g1322 ( 
.A(n_1094),
.B(n_711),
.Y(n_1322)
);

OR2x2_ASAP7_75t_L g1323 ( 
.A(n_1146),
.B(n_1212),
.Y(n_1323)
);

CKINVDCx5p33_ASAP7_75t_R g1324 ( 
.A(n_1141),
.Y(n_1324)
);

OR2x2_ASAP7_75t_L g1325 ( 
.A(n_1146),
.B(n_1212),
.Y(n_1325)
);

INVx2_ASAP7_75t_L g1326 ( 
.A(n_1111),
.Y(n_1326)
);

INVx2_ASAP7_75t_L g1327 ( 
.A(n_1111),
.Y(n_1327)
);

AND2x6_ASAP7_75t_L g1328 ( 
.A(n_1177),
.B(n_1100),
.Y(n_1328)
);

AO21x2_ASAP7_75t_L g1329 ( 
.A1(n_1137),
.A2(n_1186),
.B(n_1098),
.Y(n_1329)
);

AND2x4_ASAP7_75t_L g1330 ( 
.A(n_1121),
.B(n_954),
.Y(n_1330)
);

OAI21x1_ASAP7_75t_L g1331 ( 
.A1(n_1092),
.A2(n_1198),
.B(n_1179),
.Y(n_1331)
);

OR2x2_ASAP7_75t_L g1332 ( 
.A(n_1146),
.B(n_1212),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_L g1333 ( 
.A(n_1209),
.B(n_1085),
.Y(n_1333)
);

BUFx2_ASAP7_75t_L g1334 ( 
.A(n_1129),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1216),
.Y(n_1335)
);

OAI21x1_ASAP7_75t_L g1336 ( 
.A1(n_1092),
.A2(n_1096),
.B(n_1179),
.Y(n_1336)
);

OAI222xp33_ASAP7_75t_L g1337 ( 
.A1(n_1085),
.A2(n_769),
.B1(n_935),
.B2(n_1209),
.C1(n_1220),
.C2(n_1211),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_L g1338 ( 
.A(n_1209),
.B(n_1085),
.Y(n_1338)
);

O2A1O1Ixp33_ASAP7_75t_SL g1339 ( 
.A1(n_1183),
.A2(n_991),
.B(n_1018),
.C(n_1214),
.Y(n_1339)
);

OAI21x1_ASAP7_75t_SL g1340 ( 
.A1(n_1208),
.A2(n_1132),
.B(n_1019),
.Y(n_1340)
);

O2A1O1Ixp33_ASAP7_75t_L g1341 ( 
.A1(n_1085),
.A2(n_1209),
.B(n_829),
.C(n_1191),
.Y(n_1341)
);

NAND3xp33_ASAP7_75t_L g1342 ( 
.A(n_1209),
.B(n_829),
.C(n_1085),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_SL g1343 ( 
.A(n_1085),
.B(n_1209),
.Y(n_1343)
);

OAI21x1_ASAP7_75t_L g1344 ( 
.A1(n_1092),
.A2(n_1096),
.B(n_1179),
.Y(n_1344)
);

INVx4_ASAP7_75t_L g1345 ( 
.A(n_1169),
.Y(n_1345)
);

AOI22xp33_ASAP7_75t_L g1346 ( 
.A1(n_1085),
.A2(n_1209),
.B1(n_829),
.B2(n_1218),
.Y(n_1346)
);

OAI22xp33_ASAP7_75t_L g1347 ( 
.A1(n_1085),
.A2(n_1191),
.B1(n_1209),
.B2(n_870),
.Y(n_1347)
);

INVx2_ASAP7_75t_L g1348 ( 
.A(n_1111),
.Y(n_1348)
);

BUFx3_ASAP7_75t_L g1349 ( 
.A(n_1118),
.Y(n_1349)
);

BUFx6f_ASAP7_75t_L g1350 ( 
.A(n_1169),
.Y(n_1350)
);

OA21x2_ASAP7_75t_L g1351 ( 
.A1(n_1137),
.A2(n_1140),
.B(n_1186),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1239),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_L g1353 ( 
.A(n_1244),
.B(n_1275),
.Y(n_1353)
);

AND2x4_ASAP7_75t_L g1354 ( 
.A(n_1246),
.B(n_1273),
.Y(n_1354)
);

O2A1O1Ixp5_ASAP7_75t_L g1355 ( 
.A1(n_1337),
.A2(n_1315),
.B(n_1267),
.C(n_1242),
.Y(n_1355)
);

AOI21x1_ASAP7_75t_SL g1356 ( 
.A1(n_1311),
.A2(n_1338),
.B(n_1333),
.Y(n_1356)
);

BUFx6f_ASAP7_75t_L g1357 ( 
.A(n_1296),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_L g1358 ( 
.A(n_1244),
.B(n_1275),
.Y(n_1358)
);

AOI211xp5_ASAP7_75t_L g1359 ( 
.A1(n_1347),
.A2(n_1314),
.B(n_1341),
.C(n_1240),
.Y(n_1359)
);

OA21x2_ASAP7_75t_L g1360 ( 
.A1(n_1279),
.A2(n_1271),
.B(n_1261),
.Y(n_1360)
);

AND2x2_ASAP7_75t_SL g1361 ( 
.A(n_1346),
.B(n_1222),
.Y(n_1361)
);

OAI22xp5_ASAP7_75t_L g1362 ( 
.A1(n_1222),
.A2(n_1308),
.B1(n_1342),
.B2(n_1346),
.Y(n_1362)
);

AND2x2_ASAP7_75t_L g1363 ( 
.A(n_1246),
.B(n_1323),
.Y(n_1363)
);

AND2x2_ASAP7_75t_L g1364 ( 
.A(n_1246),
.B(n_1325),
.Y(n_1364)
);

AND2x2_ASAP7_75t_L g1365 ( 
.A(n_1332),
.B(n_1308),
.Y(n_1365)
);

AOI21xp5_ASAP7_75t_SL g1366 ( 
.A1(n_1318),
.A2(n_1343),
.B(n_1245),
.Y(n_1366)
);

NAND2xp5_ASAP7_75t_L g1367 ( 
.A(n_1275),
.B(n_1328),
.Y(n_1367)
);

AOI221xp5_ASAP7_75t_L g1368 ( 
.A1(n_1337),
.A2(n_1347),
.B1(n_1240),
.B2(n_1343),
.C(n_1339),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_L g1369 ( 
.A(n_1328),
.B(n_1281),
.Y(n_1369)
);

CKINVDCx20_ASAP7_75t_R g1370 ( 
.A(n_1274),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1328),
.B(n_1258),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_L g1372 ( 
.A(n_1328),
.B(n_1278),
.Y(n_1372)
);

CKINVDCx5p33_ASAP7_75t_R g1373 ( 
.A(n_1324),
.Y(n_1373)
);

CKINVDCx5p33_ASAP7_75t_R g1374 ( 
.A(n_1324),
.Y(n_1374)
);

O2A1O1Ixp33_ASAP7_75t_L g1375 ( 
.A1(n_1339),
.A2(n_1287),
.B(n_1280),
.C(n_1340),
.Y(n_1375)
);

INVxp33_ASAP7_75t_L g1376 ( 
.A(n_1317),
.Y(n_1376)
);

O2A1O1Ixp5_ASAP7_75t_L g1377 ( 
.A1(n_1270),
.A2(n_1264),
.B(n_1294),
.C(n_1302),
.Y(n_1377)
);

AND2x2_ASAP7_75t_L g1378 ( 
.A(n_1330),
.B(n_1268),
.Y(n_1378)
);

INVx1_ASAP7_75t_SL g1379 ( 
.A(n_1238),
.Y(n_1379)
);

NOR2xp33_ASAP7_75t_L g1380 ( 
.A(n_1298),
.B(n_1226),
.Y(n_1380)
);

AND2x2_ASAP7_75t_L g1381 ( 
.A(n_1330),
.B(n_1268),
.Y(n_1381)
);

NOR2xp67_ASAP7_75t_L g1382 ( 
.A(n_1259),
.B(n_1255),
.Y(n_1382)
);

HB1xp67_ASAP7_75t_L g1383 ( 
.A(n_1286),
.Y(n_1383)
);

INVx2_ASAP7_75t_L g1384 ( 
.A(n_1257),
.Y(n_1384)
);

OA21x2_ASAP7_75t_L g1385 ( 
.A1(n_1223),
.A2(n_1321),
.B(n_1336),
.Y(n_1385)
);

CKINVDCx20_ASAP7_75t_R g1386 ( 
.A(n_1274),
.Y(n_1386)
);

OAI22xp5_ASAP7_75t_L g1387 ( 
.A1(n_1298),
.A2(n_1282),
.B1(n_1254),
.B2(n_1276),
.Y(n_1387)
);

AOI221x1_ASAP7_75t_SL g1388 ( 
.A1(n_1236),
.A2(n_1241),
.B1(n_1256),
.B2(n_1312),
.C(n_1309),
.Y(n_1388)
);

NOR2xp67_ASAP7_75t_L g1389 ( 
.A(n_1304),
.B(n_1254),
.Y(n_1389)
);

INVx2_ASAP7_75t_L g1390 ( 
.A(n_1228),
.Y(n_1390)
);

OAI22xp5_ASAP7_75t_L g1391 ( 
.A1(n_1286),
.A2(n_1320),
.B1(n_1306),
.B2(n_1307),
.Y(n_1391)
);

AOI21xp5_ASAP7_75t_L g1392 ( 
.A1(n_1221),
.A2(n_1329),
.B(n_1233),
.Y(n_1392)
);

AOI21x1_ASAP7_75t_SL g1393 ( 
.A1(n_1302),
.A2(n_1224),
.B(n_1320),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1335),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1266),
.Y(n_1395)
);

AND2x4_ASAP7_75t_L g1396 ( 
.A(n_1273),
.B(n_1349),
.Y(n_1396)
);

AND2x4_ASAP7_75t_L g1397 ( 
.A(n_1349),
.B(n_1224),
.Y(n_1397)
);

HB1xp67_ASAP7_75t_L g1398 ( 
.A(n_1263),
.Y(n_1398)
);

O2A1O1Ixp33_ASAP7_75t_L g1399 ( 
.A1(n_1251),
.A2(n_1300),
.B(n_1288),
.C(n_1291),
.Y(n_1399)
);

INVx2_ASAP7_75t_SL g1400 ( 
.A(n_1243),
.Y(n_1400)
);

OAI22xp5_ASAP7_75t_SL g1401 ( 
.A1(n_1265),
.A2(n_1304),
.B1(n_1300),
.B2(n_1334),
.Y(n_1401)
);

NAND2xp5_ASAP7_75t_L g1402 ( 
.A(n_1328),
.B(n_1266),
.Y(n_1402)
);

AND2x2_ASAP7_75t_L g1403 ( 
.A(n_1330),
.B(n_1295),
.Y(n_1403)
);

CKINVDCx20_ASAP7_75t_R g1404 ( 
.A(n_1265),
.Y(n_1404)
);

BUFx5_ASAP7_75t_L g1405 ( 
.A(n_1302),
.Y(n_1405)
);

AND2x4_ASAP7_75t_L g1406 ( 
.A(n_1224),
.B(n_1299),
.Y(n_1406)
);

AND2x2_ASAP7_75t_L g1407 ( 
.A(n_1269),
.B(n_1290),
.Y(n_1407)
);

OAI22xp5_ASAP7_75t_L g1408 ( 
.A1(n_1247),
.A2(n_1269),
.B1(n_1319),
.B2(n_1303),
.Y(n_1408)
);

AOI21xp5_ASAP7_75t_L g1409 ( 
.A1(n_1329),
.A2(n_1252),
.B(n_1253),
.Y(n_1409)
);

O2A1O1Ixp33_ASAP7_75t_L g1410 ( 
.A1(n_1292),
.A2(n_1305),
.B(n_1316),
.C(n_1303),
.Y(n_1410)
);

AOI221xp5_ASAP7_75t_L g1411 ( 
.A1(n_1322),
.A2(n_1316),
.B1(n_1234),
.B2(n_1262),
.C(n_1305),
.Y(n_1411)
);

OAI22xp5_ASAP7_75t_L g1412 ( 
.A1(n_1247),
.A2(n_1319),
.B1(n_1283),
.B2(n_1318),
.Y(n_1412)
);

AOI21xp5_ASAP7_75t_L g1413 ( 
.A1(n_1229),
.A2(n_1285),
.B(n_1260),
.Y(n_1413)
);

AND2x2_ASAP7_75t_L g1414 ( 
.A(n_1289),
.B(n_1285),
.Y(n_1414)
);

NOR2xp67_ASAP7_75t_L g1415 ( 
.A(n_1345),
.B(n_1284),
.Y(n_1415)
);

AND2x2_ASAP7_75t_L g1416 ( 
.A(n_1285),
.B(n_1277),
.Y(n_1416)
);

INVx2_ASAP7_75t_L g1417 ( 
.A(n_1293),
.Y(n_1417)
);

AND2x2_ASAP7_75t_L g1418 ( 
.A(n_1297),
.B(n_1296),
.Y(n_1418)
);

NAND2xp5_ASAP7_75t_L g1419 ( 
.A(n_1248),
.B(n_1230),
.Y(n_1419)
);

O2A1O1Ixp5_ASAP7_75t_L g1420 ( 
.A1(n_1235),
.A2(n_1237),
.B(n_1348),
.C(n_1327),
.Y(n_1420)
);

O2A1O1Ixp33_ASAP7_75t_L g1421 ( 
.A1(n_1234),
.A2(n_1237),
.B(n_1235),
.C(n_1262),
.Y(n_1421)
);

INVx3_ASAP7_75t_SL g1422 ( 
.A(n_1231),
.Y(n_1422)
);

OAI22xp5_ASAP7_75t_L g1423 ( 
.A1(n_1231),
.A2(n_1350),
.B1(n_1250),
.B2(n_1249),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1225),
.Y(n_1424)
);

OAI22xp5_ASAP7_75t_L g1425 ( 
.A1(n_1231),
.A2(n_1250),
.B1(n_1249),
.B2(n_1350),
.Y(n_1425)
);

CKINVDCx16_ASAP7_75t_R g1426 ( 
.A(n_1272),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1232),
.Y(n_1427)
);

AOI21xp5_ASAP7_75t_L g1428 ( 
.A1(n_1351),
.A2(n_1230),
.B(n_1331),
.Y(n_1428)
);

INVxp67_ASAP7_75t_L g1429 ( 
.A(n_1243),
.Y(n_1429)
);

CKINVDCx5p33_ASAP7_75t_R g1430 ( 
.A(n_1243),
.Y(n_1430)
);

HB1xp67_ASAP7_75t_L g1431 ( 
.A(n_1231),
.Y(n_1431)
);

AND2x2_ASAP7_75t_L g1432 ( 
.A(n_1284),
.B(n_1350),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1232),
.Y(n_1433)
);

O2A1O1Ixp33_ASAP7_75t_L g1434 ( 
.A1(n_1351),
.A2(n_1310),
.B(n_1327),
.C(n_1326),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_L g1435 ( 
.A(n_1248),
.B(n_1310),
.Y(n_1435)
);

AOI21xp5_ASAP7_75t_L g1436 ( 
.A1(n_1331),
.A2(n_1227),
.B(n_1344),
.Y(n_1436)
);

AND2x2_ASAP7_75t_L g1437 ( 
.A(n_1284),
.B(n_1249),
.Y(n_1437)
);

OAI22xp5_ASAP7_75t_L g1438 ( 
.A1(n_1250),
.A2(n_1284),
.B1(n_1313),
.B2(n_1326),
.Y(n_1438)
);

OR2x2_ASAP7_75t_L g1439 ( 
.A(n_1248),
.B(n_1348),
.Y(n_1439)
);

OR2x2_ASAP7_75t_L g1440 ( 
.A(n_1301),
.B(n_1323),
.Y(n_1440)
);

AND2x4_ASAP7_75t_L g1441 ( 
.A(n_1301),
.B(n_1246),
.Y(n_1441)
);

OA21x2_ASAP7_75t_L g1442 ( 
.A1(n_1279),
.A2(n_1271),
.B(n_1137),
.Y(n_1442)
);

NAND2xp5_ASAP7_75t_L g1443 ( 
.A(n_1244),
.B(n_1275),
.Y(n_1443)
);

NAND2x1_ASAP7_75t_L g1444 ( 
.A(n_1288),
.B(n_1319),
.Y(n_1444)
);

AOI21x1_ASAP7_75t_SL g1445 ( 
.A1(n_1311),
.A2(n_1338),
.B(n_1333),
.Y(n_1445)
);

INVxp33_ASAP7_75t_SL g1446 ( 
.A(n_1317),
.Y(n_1446)
);

O2A1O1Ixp33_ASAP7_75t_L g1447 ( 
.A1(n_1314),
.A2(n_1085),
.B(n_1209),
.C(n_1341),
.Y(n_1447)
);

O2A1O1Ixp5_ASAP7_75t_L g1448 ( 
.A1(n_1337),
.A2(n_1209),
.B(n_1085),
.C(n_1186),
.Y(n_1448)
);

HB1xp67_ASAP7_75t_L g1449 ( 
.A(n_1286),
.Y(n_1449)
);

OR2x2_ASAP7_75t_L g1450 ( 
.A(n_1367),
.B(n_1353),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1424),
.Y(n_1451)
);

AND2x4_ASAP7_75t_L g1452 ( 
.A(n_1417),
.B(n_1416),
.Y(n_1452)
);

AND2x2_ASAP7_75t_L g1453 ( 
.A(n_1414),
.B(n_1367),
.Y(n_1453)
);

AO21x2_ASAP7_75t_L g1454 ( 
.A1(n_1392),
.A2(n_1428),
.B(n_1413),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1427),
.Y(n_1455)
);

INVxp67_ASAP7_75t_L g1456 ( 
.A(n_1383),
.Y(n_1456)
);

INVx2_ASAP7_75t_L g1457 ( 
.A(n_1420),
.Y(n_1457)
);

OR2x2_ASAP7_75t_L g1458 ( 
.A(n_1353),
.B(n_1358),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1433),
.Y(n_1459)
);

INVx2_ASAP7_75t_L g1460 ( 
.A(n_1439),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1352),
.Y(n_1461)
);

AOI21xp5_ASAP7_75t_SL g1462 ( 
.A1(n_1447),
.A2(n_1368),
.B(n_1362),
.Y(n_1462)
);

INVx1_ASAP7_75t_SL g1463 ( 
.A(n_1440),
.Y(n_1463)
);

NAND2xp5_ASAP7_75t_L g1464 ( 
.A(n_1369),
.B(n_1371),
.Y(n_1464)
);

AOI22xp33_ASAP7_75t_L g1465 ( 
.A1(n_1361),
.A2(n_1362),
.B1(n_1387),
.B2(n_1378),
.Y(n_1465)
);

OA21x2_ASAP7_75t_L g1466 ( 
.A1(n_1419),
.A2(n_1377),
.B(n_1409),
.Y(n_1466)
);

OAI22xp5_ASAP7_75t_L g1467 ( 
.A1(n_1359),
.A2(n_1387),
.B1(n_1379),
.B2(n_1365),
.Y(n_1467)
);

OAI21x1_ASAP7_75t_L g1468 ( 
.A1(n_1436),
.A2(n_1421),
.B(n_1434),
.Y(n_1468)
);

OR2x6_ASAP7_75t_L g1469 ( 
.A(n_1366),
.B(n_1410),
.Y(n_1469)
);

HB1xp67_ASAP7_75t_L g1470 ( 
.A(n_1435),
.Y(n_1470)
);

AND2x2_ASAP7_75t_L g1471 ( 
.A(n_1435),
.B(n_1405),
.Y(n_1471)
);

BUFx2_ASAP7_75t_L g1472 ( 
.A(n_1405),
.Y(n_1472)
);

BUFx2_ASAP7_75t_L g1473 ( 
.A(n_1402),
.Y(n_1473)
);

OAI22xp33_ASAP7_75t_L g1474 ( 
.A1(n_1357),
.A2(n_1443),
.B1(n_1358),
.B2(n_1376),
.Y(n_1474)
);

OR2x2_ASAP7_75t_L g1475 ( 
.A(n_1443),
.B(n_1402),
.Y(n_1475)
);

HB1xp67_ASAP7_75t_L g1476 ( 
.A(n_1438),
.Y(n_1476)
);

OAI21xp5_ASAP7_75t_L g1477 ( 
.A1(n_1448),
.A2(n_1355),
.B(n_1375),
.Y(n_1477)
);

AND2x4_ASAP7_75t_L g1478 ( 
.A(n_1371),
.B(n_1372),
.Y(n_1478)
);

AOI221xp5_ASAP7_75t_L g1479 ( 
.A1(n_1399),
.A2(n_1388),
.B1(n_1391),
.B2(n_1398),
.C(n_1449),
.Y(n_1479)
);

INVx2_ASAP7_75t_L g1480 ( 
.A(n_1384),
.Y(n_1480)
);

AO21x2_ASAP7_75t_L g1481 ( 
.A1(n_1438),
.A2(n_1408),
.B(n_1369),
.Y(n_1481)
);

BUFx3_ASAP7_75t_L g1482 ( 
.A(n_1418),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1395),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1394),
.Y(n_1484)
);

OA21x2_ASAP7_75t_L g1485 ( 
.A1(n_1411),
.A2(n_1390),
.B(n_1381),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1407),
.Y(n_1486)
);

INVx2_ASAP7_75t_L g1487 ( 
.A(n_1385),
.Y(n_1487)
);

INVx1_ASAP7_75t_SL g1488 ( 
.A(n_1403),
.Y(n_1488)
);

HB1xp67_ASAP7_75t_L g1489 ( 
.A(n_1360),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1442),
.Y(n_1490)
);

HB1xp67_ASAP7_75t_L g1491 ( 
.A(n_1411),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1441),
.Y(n_1492)
);

AO21x2_ASAP7_75t_L g1493 ( 
.A1(n_1423),
.A2(n_1425),
.B(n_1412),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_L g1494 ( 
.A(n_1406),
.B(n_1397),
.Y(n_1494)
);

AO21x2_ASAP7_75t_L g1495 ( 
.A1(n_1412),
.A2(n_1415),
.B(n_1406),
.Y(n_1495)
);

OR2x2_ASAP7_75t_L g1496 ( 
.A(n_1397),
.B(n_1364),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1363),
.B(n_1354),
.Y(n_1497)
);

AND2x2_ASAP7_75t_L g1498 ( 
.A(n_1354),
.B(n_1396),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_L g1499 ( 
.A(n_1431),
.B(n_1396),
.Y(n_1499)
);

INVxp67_ASAP7_75t_L g1500 ( 
.A(n_1432),
.Y(n_1500)
);

NAND2xp5_ASAP7_75t_L g1501 ( 
.A(n_1458),
.B(n_1444),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_L g1502 ( 
.A(n_1458),
.B(n_1389),
.Y(n_1502)
);

INVxp67_ASAP7_75t_SL g1503 ( 
.A(n_1470),
.Y(n_1503)
);

AND2x2_ASAP7_75t_L g1504 ( 
.A(n_1453),
.B(n_1437),
.Y(n_1504)
);

AND2x2_ASAP7_75t_L g1505 ( 
.A(n_1453),
.B(n_1380),
.Y(n_1505)
);

AND2x2_ASAP7_75t_L g1506 ( 
.A(n_1453),
.B(n_1357),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1478),
.B(n_1471),
.Y(n_1507)
);

AND2x2_ASAP7_75t_L g1508 ( 
.A(n_1478),
.B(n_1357),
.Y(n_1508)
);

AND2x2_ASAP7_75t_L g1509 ( 
.A(n_1478),
.B(n_1400),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1461),
.Y(n_1510)
);

AND2x2_ASAP7_75t_L g1511 ( 
.A(n_1478),
.B(n_1429),
.Y(n_1511)
);

OR2x2_ASAP7_75t_L g1512 ( 
.A(n_1450),
.B(n_1422),
.Y(n_1512)
);

NAND2xp5_ASAP7_75t_L g1513 ( 
.A(n_1475),
.B(n_1382),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1461),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1475),
.B(n_1446),
.Y(n_1515)
);

INVx2_ASAP7_75t_L g1516 ( 
.A(n_1487),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_L g1517 ( 
.A(n_1450),
.B(n_1401),
.Y(n_1517)
);

INVx2_ASAP7_75t_L g1518 ( 
.A(n_1487),
.Y(n_1518)
);

HB1xp67_ASAP7_75t_L g1519 ( 
.A(n_1470),
.Y(n_1519)
);

AND2x2_ASAP7_75t_L g1520 ( 
.A(n_1478),
.B(n_1393),
.Y(n_1520)
);

NAND2xp5_ASAP7_75t_L g1521 ( 
.A(n_1464),
.B(n_1473),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1471),
.B(n_1430),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_SL g1523 ( 
.A(n_1477),
.B(n_1374),
.Y(n_1523)
);

AND2x2_ASAP7_75t_L g1524 ( 
.A(n_1471),
.B(n_1426),
.Y(n_1524)
);

OR2x2_ASAP7_75t_L g1525 ( 
.A(n_1460),
.B(n_1464),
.Y(n_1525)
);

INVx5_ASAP7_75t_L g1526 ( 
.A(n_1469),
.Y(n_1526)
);

INVx2_ASAP7_75t_SL g1527 ( 
.A(n_1452),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1491),
.B(n_1356),
.Y(n_1528)
);

OA21x2_ASAP7_75t_L g1529 ( 
.A1(n_1468),
.A2(n_1445),
.B(n_1373),
.Y(n_1529)
);

CKINVDCx20_ASAP7_75t_R g1530 ( 
.A(n_1482),
.Y(n_1530)
);

OAI31xp33_ASAP7_75t_L g1531 ( 
.A1(n_1523),
.A2(n_1467),
.A3(n_1465),
.B(n_1474),
.Y(n_1531)
);

OAI211xp5_ASAP7_75t_SL g1532 ( 
.A1(n_1528),
.A2(n_1462),
.B(n_1523),
.C(n_1517),
.Y(n_1532)
);

OAI211xp5_ASAP7_75t_L g1533 ( 
.A1(n_1528),
.A2(n_1477),
.B(n_1491),
.C(n_1479),
.Y(n_1533)
);

OAI22xp5_ASAP7_75t_L g1534 ( 
.A1(n_1530),
.A2(n_1467),
.B1(n_1469),
.B2(n_1479),
.Y(n_1534)
);

BUFx10_ASAP7_75t_L g1535 ( 
.A(n_1510),
.Y(n_1535)
);

AOI33xp33_ASAP7_75t_L g1536 ( 
.A1(n_1505),
.A2(n_1474),
.A3(n_1484),
.B1(n_1486),
.B2(n_1488),
.B3(n_1463),
.Y(n_1536)
);

AOI222xp33_ASAP7_75t_SL g1537 ( 
.A1(n_1519),
.A2(n_1456),
.B1(n_1463),
.B2(n_1484),
.C1(n_1488),
.C2(n_1486),
.Y(n_1537)
);

AOI22xp33_ASAP7_75t_L g1538 ( 
.A1(n_1511),
.A2(n_1469),
.B1(n_1482),
.B2(n_1493),
.Y(n_1538)
);

AOI33xp33_ASAP7_75t_L g1539 ( 
.A1(n_1505),
.A2(n_1483),
.A3(n_1457),
.B1(n_1459),
.B2(n_1451),
.B3(n_1455),
.Y(n_1539)
);

OR2x2_ASAP7_75t_L g1540 ( 
.A(n_1521),
.B(n_1460),
.Y(n_1540)
);

AND2x2_ASAP7_75t_L g1541 ( 
.A(n_1507),
.B(n_1485),
.Y(n_1541)
);

AOI221xp5_ASAP7_75t_L g1542 ( 
.A1(n_1517),
.A2(n_1456),
.B1(n_1476),
.B2(n_1500),
.C(n_1499),
.Y(n_1542)
);

NAND2xp33_ASAP7_75t_SL g1543 ( 
.A(n_1530),
.B(n_1404),
.Y(n_1543)
);

INVx2_ASAP7_75t_L g1544 ( 
.A(n_1516),
.Y(n_1544)
);

OAI211xp5_ASAP7_75t_L g1545 ( 
.A1(n_1513),
.A2(n_1476),
.B(n_1485),
.C(n_1466),
.Y(n_1545)
);

NAND2xp5_ASAP7_75t_L g1546 ( 
.A(n_1521),
.B(n_1500),
.Y(n_1546)
);

OAI22xp5_ASAP7_75t_L g1547 ( 
.A1(n_1513),
.A2(n_1469),
.B1(n_1496),
.B2(n_1482),
.Y(n_1547)
);

AND2x2_ASAP7_75t_L g1548 ( 
.A(n_1507),
.B(n_1485),
.Y(n_1548)
);

OR2x2_ASAP7_75t_L g1549 ( 
.A(n_1525),
.B(n_1485),
.Y(n_1549)
);

INVx4_ASAP7_75t_SL g1550 ( 
.A(n_1520),
.Y(n_1550)
);

BUFx2_ASAP7_75t_L g1551 ( 
.A(n_1519),
.Y(n_1551)
);

AOI221xp5_ASAP7_75t_L g1552 ( 
.A1(n_1515),
.A2(n_1501),
.B1(n_1502),
.B2(n_1505),
.C(n_1520),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1507),
.B(n_1485),
.Y(n_1553)
);

AOI22xp33_ASAP7_75t_L g1554 ( 
.A1(n_1511),
.A2(n_1469),
.B1(n_1493),
.B2(n_1495),
.Y(n_1554)
);

AOI22xp33_ASAP7_75t_L g1555 ( 
.A1(n_1511),
.A2(n_1469),
.B1(n_1493),
.B2(n_1495),
.Y(n_1555)
);

OAI33xp33_ASAP7_75t_L g1556 ( 
.A1(n_1501),
.A2(n_1483),
.A3(n_1499),
.B1(n_1451),
.B2(n_1459),
.B3(n_1455),
.Y(n_1556)
);

BUFx3_ASAP7_75t_L g1557 ( 
.A(n_1508),
.Y(n_1557)
);

AO21x2_ASAP7_75t_L g1558 ( 
.A1(n_1518),
.A2(n_1490),
.B(n_1489),
.Y(n_1558)
);

OAI33xp33_ASAP7_75t_L g1559 ( 
.A1(n_1515),
.A2(n_1492),
.A3(n_1490),
.B1(n_1457),
.B2(n_1494),
.B3(n_1480),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1504),
.B(n_1472),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1510),
.Y(n_1561)
);

NAND5xp2_ASAP7_75t_L g1562 ( 
.A(n_1524),
.B(n_1492),
.C(n_1498),
.D(n_1494),
.E(n_1472),
.Y(n_1562)
);

OR2x2_ASAP7_75t_L g1563 ( 
.A(n_1525),
.B(n_1481),
.Y(n_1563)
);

AND3x1_ASAP7_75t_L g1564 ( 
.A(n_1524),
.B(n_1498),
.C(n_1497),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1514),
.Y(n_1565)
);

INVx2_ASAP7_75t_L g1566 ( 
.A(n_1558),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1561),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1561),
.Y(n_1568)
);

AND2x2_ASAP7_75t_L g1569 ( 
.A(n_1541),
.B(n_1527),
.Y(n_1569)
);

NAND3xp33_ASAP7_75t_SL g1570 ( 
.A(n_1531),
.B(n_1502),
.C(n_1524),
.Y(n_1570)
);

INVx1_ASAP7_75t_SL g1571 ( 
.A(n_1551),
.Y(n_1571)
);

BUFx2_ASAP7_75t_L g1572 ( 
.A(n_1550),
.Y(n_1572)
);

INVx1_ASAP7_75t_SL g1573 ( 
.A(n_1551),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1565),
.Y(n_1574)
);

INVxp67_ASAP7_75t_SL g1575 ( 
.A(n_1549),
.Y(n_1575)
);

BUFx2_ASAP7_75t_L g1576 ( 
.A(n_1550),
.Y(n_1576)
);

INVx2_ASAP7_75t_L g1577 ( 
.A(n_1558),
.Y(n_1577)
);

INVx2_ASAP7_75t_L g1578 ( 
.A(n_1544),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_L g1579 ( 
.A(n_1539),
.B(n_1503),
.Y(n_1579)
);

NOR2xp33_ASAP7_75t_L g1580 ( 
.A(n_1532),
.B(n_1522),
.Y(n_1580)
);

INVx4_ASAP7_75t_SL g1581 ( 
.A(n_1557),
.Y(n_1581)
);

INVxp67_ASAP7_75t_L g1582 ( 
.A(n_1537),
.Y(n_1582)
);

OAI21xp33_ASAP7_75t_L g1583 ( 
.A1(n_1533),
.A2(n_1520),
.B(n_1512),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1563),
.B(n_1504),
.Y(n_1584)
);

BUFx2_ASAP7_75t_L g1585 ( 
.A(n_1550),
.Y(n_1585)
);

AO21x2_ASAP7_75t_L g1586 ( 
.A1(n_1545),
.A2(n_1454),
.B(n_1489),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1535),
.Y(n_1587)
);

NOR2xp67_ASAP7_75t_L g1588 ( 
.A(n_1562),
.B(n_1526),
.Y(n_1588)
);

INVx3_ASAP7_75t_L g1589 ( 
.A(n_1535),
.Y(n_1589)
);

INVx4_ASAP7_75t_SL g1590 ( 
.A(n_1557),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1572),
.B(n_1550),
.Y(n_1591)
);

BUFx6f_ASAP7_75t_L g1592 ( 
.A(n_1572),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1567),
.Y(n_1593)
);

OR2x2_ASAP7_75t_L g1594 ( 
.A(n_1579),
.B(n_1563),
.Y(n_1594)
);

INVx2_ASAP7_75t_L g1595 ( 
.A(n_1578),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1567),
.Y(n_1596)
);

NOR2xp33_ASAP7_75t_L g1597 ( 
.A(n_1580),
.B(n_1543),
.Y(n_1597)
);

NAND3xp33_ASAP7_75t_L g1598 ( 
.A(n_1582),
.B(n_1531),
.C(n_1534),
.Y(n_1598)
);

AOI21xp5_ASAP7_75t_L g1599 ( 
.A1(n_1570),
.A2(n_1555),
.B(n_1554),
.Y(n_1599)
);

NAND2x1p5_ASAP7_75t_L g1600 ( 
.A(n_1572),
.B(n_1526),
.Y(n_1600)
);

AND2x2_ASAP7_75t_L g1601 ( 
.A(n_1576),
.B(n_1550),
.Y(n_1601)
);

INVx1_ASAP7_75t_SL g1602 ( 
.A(n_1576),
.Y(n_1602)
);

AOI221xp5_ASAP7_75t_L g1603 ( 
.A1(n_1570),
.A2(n_1559),
.B1(n_1542),
.B2(n_1552),
.C(n_1556),
.Y(n_1603)
);

BUFx3_ASAP7_75t_L g1604 ( 
.A(n_1576),
.Y(n_1604)
);

AOI22xp33_ASAP7_75t_L g1605 ( 
.A1(n_1583),
.A2(n_1526),
.B1(n_1538),
.B2(n_1547),
.Y(n_1605)
);

AND2x2_ASAP7_75t_L g1606 ( 
.A(n_1585),
.B(n_1564),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1582),
.B(n_1536),
.Y(n_1607)
);

AND2x2_ASAP7_75t_L g1608 ( 
.A(n_1585),
.B(n_1564),
.Y(n_1608)
);

HB1xp67_ASAP7_75t_L g1609 ( 
.A(n_1571),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1568),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_L g1611 ( 
.A(n_1583),
.B(n_1506),
.Y(n_1611)
);

OR2x2_ASAP7_75t_L g1612 ( 
.A(n_1579),
.B(n_1549),
.Y(n_1612)
);

OR2x2_ASAP7_75t_L g1613 ( 
.A(n_1584),
.B(n_1540),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1568),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_L g1615 ( 
.A(n_1580),
.B(n_1506),
.Y(n_1615)
);

INVx1_ASAP7_75t_SL g1616 ( 
.A(n_1585),
.Y(n_1616)
);

OR2x2_ASAP7_75t_L g1617 ( 
.A(n_1571),
.B(n_1540),
.Y(n_1617)
);

AND2x2_ASAP7_75t_L g1618 ( 
.A(n_1581),
.B(n_1548),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1581),
.B(n_1553),
.Y(n_1619)
);

NOR3xp33_ASAP7_75t_SL g1620 ( 
.A(n_1587),
.B(n_1546),
.C(n_1514),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_SL g1621 ( 
.A(n_1588),
.B(n_1526),
.Y(n_1621)
);

INVx2_ASAP7_75t_L g1622 ( 
.A(n_1578),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_L g1623 ( 
.A(n_1573),
.B(n_1553),
.Y(n_1623)
);

AND2x4_ASAP7_75t_L g1624 ( 
.A(n_1581),
.B(n_1590),
.Y(n_1624)
);

INVx3_ASAP7_75t_L g1625 ( 
.A(n_1589),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1574),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1581),
.B(n_1557),
.Y(n_1627)
);

HB1xp67_ASAP7_75t_L g1628 ( 
.A(n_1573),
.Y(n_1628)
);

NAND4xp25_ASAP7_75t_SL g1629 ( 
.A(n_1569),
.B(n_1537),
.C(n_1522),
.D(n_1508),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1593),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_L g1631 ( 
.A(n_1607),
.B(n_1560),
.Y(n_1631)
);

INVx1_ASAP7_75t_SL g1632 ( 
.A(n_1591),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_L g1633 ( 
.A(n_1598),
.B(n_1560),
.Y(n_1633)
);

NAND2x1p5_ASAP7_75t_L g1634 ( 
.A(n_1624),
.B(n_1526),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1593),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_L g1636 ( 
.A(n_1598),
.B(n_1603),
.Y(n_1636)
);

AND2x2_ASAP7_75t_L g1637 ( 
.A(n_1591),
.B(n_1581),
.Y(n_1637)
);

AND2x2_ASAP7_75t_L g1638 ( 
.A(n_1601),
.B(n_1581),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1601),
.B(n_1590),
.Y(n_1639)
);

NAND2x1_ASAP7_75t_L g1640 ( 
.A(n_1624),
.B(n_1588),
.Y(n_1640)
);

INVx2_ASAP7_75t_L g1641 ( 
.A(n_1592),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1596),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1596),
.Y(n_1643)
);

OR2x2_ASAP7_75t_L g1644 ( 
.A(n_1594),
.B(n_1612),
.Y(n_1644)
);

OR2x2_ASAP7_75t_L g1645 ( 
.A(n_1594),
.B(n_1575),
.Y(n_1645)
);

AND2x2_ASAP7_75t_L g1646 ( 
.A(n_1606),
.B(n_1608),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1610),
.Y(n_1647)
);

NOR2xp67_ASAP7_75t_L g1648 ( 
.A(n_1624),
.B(n_1629),
.Y(n_1648)
);

OR2x2_ASAP7_75t_L g1649 ( 
.A(n_1612),
.B(n_1575),
.Y(n_1649)
);

INVx3_ASAP7_75t_L g1650 ( 
.A(n_1592),
.Y(n_1650)
);

OR2x2_ASAP7_75t_L g1651 ( 
.A(n_1617),
.B(n_1574),
.Y(n_1651)
);

OAI22xp5_ASAP7_75t_L g1652 ( 
.A1(n_1599),
.A2(n_1526),
.B1(n_1520),
.B2(n_1529),
.Y(n_1652)
);

INVx2_ASAP7_75t_L g1653 ( 
.A(n_1592),
.Y(n_1653)
);

AND2x2_ASAP7_75t_L g1654 ( 
.A(n_1606),
.B(n_1590),
.Y(n_1654)
);

NAND2xp5_ASAP7_75t_L g1655 ( 
.A(n_1609),
.B(n_1508),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1608),
.B(n_1590),
.Y(n_1656)
);

AND2x4_ASAP7_75t_L g1657 ( 
.A(n_1604),
.B(n_1590),
.Y(n_1657)
);

INVx2_ASAP7_75t_L g1658 ( 
.A(n_1592),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1627),
.B(n_1590),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1610),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_L g1661 ( 
.A(n_1628),
.B(n_1509),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1614),
.Y(n_1662)
);

AND2x2_ASAP7_75t_L g1663 ( 
.A(n_1627),
.B(n_1569),
.Y(n_1663)
);

AOI21xp5_ASAP7_75t_L g1664 ( 
.A1(n_1597),
.A2(n_1586),
.B(n_1526),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1630),
.Y(n_1665)
);

OR2x2_ASAP7_75t_L g1666 ( 
.A(n_1644),
.B(n_1617),
.Y(n_1666)
);

INVx2_ASAP7_75t_L g1667 ( 
.A(n_1650),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_L g1668 ( 
.A(n_1632),
.B(n_1620),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1630),
.Y(n_1669)
);

HB1xp67_ASAP7_75t_L g1670 ( 
.A(n_1650),
.Y(n_1670)
);

INVx3_ASAP7_75t_SL g1671 ( 
.A(n_1650),
.Y(n_1671)
);

OR2x6_ASAP7_75t_L g1672 ( 
.A(n_1641),
.B(n_1592),
.Y(n_1672)
);

AND2x2_ASAP7_75t_L g1673 ( 
.A(n_1646),
.B(n_1604),
.Y(n_1673)
);

INVx3_ASAP7_75t_L g1674 ( 
.A(n_1640),
.Y(n_1674)
);

BUFx3_ASAP7_75t_L g1675 ( 
.A(n_1641),
.Y(n_1675)
);

HB1xp67_ASAP7_75t_L g1676 ( 
.A(n_1653),
.Y(n_1676)
);

AOI22xp33_ASAP7_75t_L g1677 ( 
.A1(n_1636),
.A2(n_1605),
.B1(n_1526),
.B2(n_1621),
.Y(n_1677)
);

OR2x6_ASAP7_75t_L g1678 ( 
.A(n_1653),
.B(n_1600),
.Y(n_1678)
);

AO22x1_ASAP7_75t_L g1679 ( 
.A1(n_1657),
.A2(n_1602),
.B1(n_1616),
.B2(n_1618),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1635),
.Y(n_1680)
);

INVx3_ASAP7_75t_L g1681 ( 
.A(n_1640),
.Y(n_1681)
);

BUFx2_ASAP7_75t_L g1682 ( 
.A(n_1657),
.Y(n_1682)
);

NAND2xp5_ASAP7_75t_L g1683 ( 
.A(n_1633),
.B(n_1646),
.Y(n_1683)
);

OR2x2_ASAP7_75t_L g1684 ( 
.A(n_1644),
.B(n_1613),
.Y(n_1684)
);

AND2x2_ASAP7_75t_L g1685 ( 
.A(n_1637),
.B(n_1600),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1635),
.Y(n_1686)
);

INVx1_ASAP7_75t_SL g1687 ( 
.A(n_1637),
.Y(n_1687)
);

NOR2xp33_ASAP7_75t_L g1688 ( 
.A(n_1631),
.B(n_1615),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1642),
.Y(n_1689)
);

INVx2_ASAP7_75t_L g1690 ( 
.A(n_1672),
.Y(n_1690)
);

AND2x2_ASAP7_75t_L g1691 ( 
.A(n_1673),
.B(n_1638),
.Y(n_1691)
);

XOR2x2_ASAP7_75t_L g1692 ( 
.A(n_1683),
.B(n_1648),
.Y(n_1692)
);

INVxp67_ASAP7_75t_L g1693 ( 
.A(n_1673),
.Y(n_1693)
);

AOI21xp5_ASAP7_75t_L g1694 ( 
.A1(n_1679),
.A2(n_1668),
.B(n_1648),
.Y(n_1694)
);

NOR2xp33_ASAP7_75t_L g1695 ( 
.A(n_1687),
.B(n_1659),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1676),
.Y(n_1696)
);

OAI22xp5_ASAP7_75t_L g1697 ( 
.A1(n_1666),
.A2(n_1611),
.B1(n_1638),
.B2(n_1639),
.Y(n_1697)
);

OR2x2_ASAP7_75t_L g1698 ( 
.A(n_1666),
.B(n_1655),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1689),
.Y(n_1699)
);

OAI21xp33_ASAP7_75t_L g1700 ( 
.A1(n_1688),
.A2(n_1639),
.B(n_1656),
.Y(n_1700)
);

AND2x2_ASAP7_75t_L g1701 ( 
.A(n_1685),
.B(n_1659),
.Y(n_1701)
);

AOI31xp33_ASAP7_75t_L g1702 ( 
.A1(n_1685),
.A2(n_1656),
.A3(n_1654),
.B(n_1657),
.Y(n_1702)
);

BUFx3_ASAP7_75t_L g1703 ( 
.A(n_1682),
.Y(n_1703)
);

INVxp67_ASAP7_75t_L g1704 ( 
.A(n_1682),
.Y(n_1704)
);

AOI21xp5_ASAP7_75t_L g1705 ( 
.A1(n_1679),
.A2(n_1664),
.B(n_1652),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1689),
.Y(n_1706)
);

AND2x2_ASAP7_75t_L g1707 ( 
.A(n_1671),
.B(n_1654),
.Y(n_1707)
);

AOI222xp33_ASAP7_75t_L g1708 ( 
.A1(n_1677),
.A2(n_1657),
.B1(n_1658),
.B2(n_1643),
.C1(n_1660),
.C2(n_1662),
.Y(n_1708)
);

AND2x2_ASAP7_75t_L g1709 ( 
.A(n_1691),
.B(n_1663),
.Y(n_1709)
);

HB1xp67_ASAP7_75t_L g1710 ( 
.A(n_1703),
.Y(n_1710)
);

INVx2_ASAP7_75t_L g1711 ( 
.A(n_1703),
.Y(n_1711)
);

AND2x2_ASAP7_75t_L g1712 ( 
.A(n_1691),
.B(n_1663),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_L g1713 ( 
.A(n_1693),
.B(n_1675),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_L g1714 ( 
.A(n_1704),
.B(n_1675),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_1695),
.B(n_1707),
.Y(n_1715)
);

NAND2x1p5_ASAP7_75t_L g1716 ( 
.A(n_1707),
.B(n_1674),
.Y(n_1716)
);

NAND2xp5_ASAP7_75t_L g1717 ( 
.A(n_1695),
.B(n_1670),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_L g1718 ( 
.A(n_1696),
.B(n_1667),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_L g1719 ( 
.A(n_1701),
.B(n_1667),
.Y(n_1719)
);

NAND3xp33_ASAP7_75t_SL g1720 ( 
.A(n_1716),
.B(n_1694),
.C(n_1708),
.Y(n_1720)
);

OAI22xp5_ASAP7_75t_L g1721 ( 
.A1(n_1715),
.A2(n_1702),
.B1(n_1698),
.B2(n_1684),
.Y(n_1721)
);

AOI221xp5_ASAP7_75t_L g1722 ( 
.A1(n_1717),
.A2(n_1700),
.B1(n_1697),
.B2(n_1705),
.C(n_1690),
.Y(n_1722)
);

NOR2x1_ASAP7_75t_L g1723 ( 
.A(n_1714),
.B(n_1690),
.Y(n_1723)
);

NAND3xp33_ASAP7_75t_L g1724 ( 
.A(n_1710),
.B(n_1672),
.C(n_1658),
.Y(n_1724)
);

NAND5xp2_ASAP7_75t_SL g1725 ( 
.A(n_1709),
.B(n_1692),
.C(n_1671),
.D(n_1672),
.E(n_1618),
.Y(n_1725)
);

AOI322xp5_ASAP7_75t_L g1726 ( 
.A1(n_1714),
.A2(n_1706),
.A3(n_1699),
.B1(n_1692),
.B2(n_1686),
.C1(n_1665),
.C2(n_1680),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1718),
.Y(n_1727)
);

NAND2xp5_ASAP7_75t_SL g1728 ( 
.A(n_1711),
.B(n_1684),
.Y(n_1728)
);

NOR2x1_ASAP7_75t_L g1729 ( 
.A(n_1713),
.B(n_1672),
.Y(n_1729)
);

AOI31xp33_ASAP7_75t_L g1730 ( 
.A1(n_1719),
.A2(n_1712),
.A3(n_1634),
.B(n_1600),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1723),
.Y(n_1731)
);

AOI22xp5_ASAP7_75t_L g1732 ( 
.A1(n_1720),
.A2(n_1671),
.B1(n_1681),
.B2(n_1674),
.Y(n_1732)
);

AO22x1_ASAP7_75t_L g1733 ( 
.A1(n_1729),
.A2(n_1681),
.B1(n_1674),
.B2(n_1686),
.Y(n_1733)
);

AOI21xp33_ASAP7_75t_L g1734 ( 
.A1(n_1721),
.A2(n_1681),
.B(n_1678),
.Y(n_1734)
);

NOR3xp33_ASAP7_75t_L g1735 ( 
.A(n_1728),
.B(n_1680),
.C(n_1669),
.Y(n_1735)
);

AND2x2_ASAP7_75t_L g1736 ( 
.A(n_1732),
.B(n_1727),
.Y(n_1736)
);

AND2x2_ASAP7_75t_L g1737 ( 
.A(n_1731),
.B(n_1722),
.Y(n_1737)
);

BUFx2_ASAP7_75t_L g1738 ( 
.A(n_1733),
.Y(n_1738)
);

INVxp67_ASAP7_75t_L g1739 ( 
.A(n_1734),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1735),
.Y(n_1740)
);

OR2x2_ASAP7_75t_L g1741 ( 
.A(n_1731),
.B(n_1724),
.Y(n_1741)
);

XOR2xp5_ASAP7_75t_L g1742 ( 
.A(n_1741),
.B(n_1725),
.Y(n_1742)
);

AOI31xp33_ASAP7_75t_L g1743 ( 
.A1(n_1737),
.A2(n_1634),
.A3(n_1726),
.B(n_1669),
.Y(n_1743)
);

AOI221xp5_ASAP7_75t_L g1744 ( 
.A1(n_1740),
.A2(n_1730),
.B1(n_1665),
.B2(n_1662),
.C(n_1642),
.Y(n_1744)
);

INVxp33_ASAP7_75t_L g1745 ( 
.A(n_1736),
.Y(n_1745)
);

XNOR2xp5_ASAP7_75t_L g1746 ( 
.A(n_1736),
.B(n_1370),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1746),
.Y(n_1747)
);

NAND2xp5_ASAP7_75t_SL g1748 ( 
.A(n_1743),
.B(n_1738),
.Y(n_1748)
);

NOR2xp33_ASAP7_75t_L g1749 ( 
.A(n_1745),
.B(n_1739),
.Y(n_1749)
);

AND3x4_ASAP7_75t_L g1750 ( 
.A(n_1748),
.B(n_1742),
.C(n_1739),
.Y(n_1750)
);

AOI322xp5_ASAP7_75t_L g1751 ( 
.A1(n_1750),
.A2(n_1749),
.A3(n_1747),
.B1(n_1744),
.B2(n_1660),
.C1(n_1647),
.C2(n_1643),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1751),
.Y(n_1752)
);

INVx2_ASAP7_75t_L g1753 ( 
.A(n_1752),
.Y(n_1753)
);

OAI21xp5_ASAP7_75t_L g1754 ( 
.A1(n_1753),
.A2(n_1678),
.B(n_1634),
.Y(n_1754)
);

OAI22x1_ASAP7_75t_L g1755 ( 
.A1(n_1754),
.A2(n_1647),
.B1(n_1645),
.B2(n_1649),
.Y(n_1755)
);

AOI22xp5_ASAP7_75t_SL g1756 ( 
.A1(n_1754),
.A2(n_1386),
.B1(n_1625),
.B2(n_1619),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1756),
.Y(n_1757)
);

AO221x2_ASAP7_75t_L g1758 ( 
.A1(n_1755),
.A2(n_1678),
.B1(n_1622),
.B2(n_1595),
.C(n_1661),
.Y(n_1758)
);

NAND3xp33_ASAP7_75t_L g1759 ( 
.A(n_1757),
.B(n_1678),
.C(n_1645),
.Y(n_1759)
);

NOR2xp33_ASAP7_75t_L g1760 ( 
.A(n_1758),
.B(n_1649),
.Y(n_1760)
);

AOI322xp5_ASAP7_75t_L g1761 ( 
.A1(n_1760),
.A2(n_1625),
.A3(n_1619),
.B1(n_1622),
.B2(n_1595),
.C1(n_1614),
.C2(n_1626),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1759),
.Y(n_1762)
);

AOI22xp5_ASAP7_75t_L g1763 ( 
.A1(n_1762),
.A2(n_1625),
.B1(n_1651),
.B2(n_1626),
.Y(n_1763)
);

OAI22xp33_ASAP7_75t_L g1764 ( 
.A1(n_1761),
.A2(n_1651),
.B1(n_1623),
.B2(n_1613),
.Y(n_1764)
);

AOI211xp5_ASAP7_75t_L g1765 ( 
.A1(n_1764),
.A2(n_1763),
.B(n_1566),
.C(n_1577),
.Y(n_1765)
);


endmodule