module fake_jpeg_29322_n_282 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_282);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_282;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_165;
wire n_78;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_259;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_260;
wire n_112;
wire n_199;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_13),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_18),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_17),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_15),
.Y(n_22)
);

BUFx16f_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_5),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_12),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_16),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_9),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_4),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

INVx13_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_4),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_41),
.Y(n_42)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_42),
.Y(n_98)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_41),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_43),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_21),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_44),
.B(n_51),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_45),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_26),
.Y(n_47)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_47),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_48),
.Y(n_91)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_49),
.Y(n_95)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_26),
.Y(n_50)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_50),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_21),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_25),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_52),
.Y(n_80)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_29),
.Y(n_53)
);

BUFx2_ASAP7_75t_L g64 ( 
.A(n_53),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_25),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_54),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_21),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_55),
.B(n_61),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_25),
.Y(n_56)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_56),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_23),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_57),
.B(n_39),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_25),
.Y(n_58)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_58),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_32),
.Y(n_59)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_59),
.Y(n_79)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_60),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_32),
.Y(n_61)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_29),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_62),
.B(n_63),
.Y(n_72)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_33),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_59),
.A2(n_32),
.B1(n_26),
.B2(n_28),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_66),
.A2(n_75),
.B1(n_96),
.B2(n_99),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_47),
.B(n_40),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_68),
.B(n_70),
.Y(n_129)
);

NAND2x1p5_ASAP7_75t_L g69 ( 
.A(n_49),
.B(n_23),
.Y(n_69)
);

OR2x4_ASAP7_75t_L g118 ( 
.A(n_69),
.B(n_2),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_61),
.B(n_40),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_45),
.B(n_19),
.Y(n_73)
);

NAND3xp33_ASAP7_75t_L g109 ( 
.A(n_73),
.B(n_76),
.C(n_17),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_42),
.A2(n_28),
.B1(n_29),
.B2(n_23),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_45),
.B(n_19),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_43),
.B(n_37),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_77),
.B(n_92),
.Y(n_135)
);

OAI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_52),
.A2(n_28),
.B1(n_23),
.B2(n_34),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_82),
.A2(n_87),
.B1(n_3),
.B2(n_7),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_53),
.B(n_20),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_83),
.B(n_86),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_62),
.B(n_20),
.Y(n_86)
);

OAI22xp33_ASAP7_75t_L g87 ( 
.A1(n_54),
.A2(n_24),
.B1(n_38),
.B2(n_34),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_46),
.B(n_22),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_90),
.B(n_97),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_58),
.B(n_30),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_56),
.B(n_30),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_94),
.B(n_1),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_48),
.A2(n_29),
.B1(n_38),
.B2(n_24),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_60),
.B(n_35),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_47),
.A2(n_37),
.B1(n_36),
.B2(n_27),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_47),
.A2(n_36),
.B1(n_27),
.B2(n_35),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_100),
.A2(n_101),
.B1(n_3),
.B2(n_4),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_47),
.A2(n_31),
.B1(n_22),
.B2(n_39),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_60),
.B(n_31),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_102),
.B(n_103),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_77),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_104),
.A2(n_131),
.B1(n_112),
.B2(n_107),
.Y(n_142)
);

XNOR2x1_ASAP7_75t_L g106 ( 
.A(n_68),
.B(n_70),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_106),
.B(n_115),
.C(n_112),
.Y(n_159)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_84),
.Y(n_108)
);

INVx4_ASAP7_75t_SL g136 ( 
.A(n_108),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_109),
.B(n_128),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_65),
.Y(n_110)
);

OR2x2_ASAP7_75t_L g143 ( 
.A(n_110),
.B(n_118),
.Y(n_143)
);

BUFx2_ASAP7_75t_L g111 ( 
.A(n_98),
.Y(n_111)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_111),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_112),
.B(n_115),
.Y(n_164)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_69),
.B(n_94),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_80),
.Y(n_116)
);

INVx6_ASAP7_75t_L g138 ( 
.A(n_116),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_72),
.B(n_13),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_117),
.B(n_120),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_119),
.A2(n_7),
.B(n_8),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_81),
.B(n_14),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_67),
.B(n_92),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_121),
.B(n_124),
.Y(n_162)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_95),
.Y(n_122)
);

INVx1_ASAP7_75t_SL g163 ( 
.A(n_122),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_64),
.Y(n_123)
);

OR2x2_ASAP7_75t_L g155 ( 
.A(n_123),
.B(n_125),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_93),
.B(n_12),
.Y(n_124)
);

AO22x2_ASAP7_75t_L g125 ( 
.A1(n_69),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_84),
.Y(n_126)
);

INVx13_ASAP7_75t_L g137 ( 
.A(n_126),
.Y(n_137)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_88),
.Y(n_127)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_127),
.Y(n_139)
);

CKINVDCx12_ASAP7_75t_R g128 ( 
.A(n_64),
.Y(n_128)
);

A2O1A1Ixp33_ASAP7_75t_L g130 ( 
.A1(n_87),
.A2(n_11),
.B(n_5),
.C(n_6),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_130),
.B(n_7),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_79),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_132),
.B(n_133),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_95),
.B(n_11),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_88),
.Y(n_134)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_134),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_135),
.B(n_93),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_140),
.B(n_145),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_142),
.A2(n_160),
.B1(n_91),
.B2(n_126),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_135),
.B(n_74),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_127),
.Y(n_146)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_146),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_147),
.A2(n_155),
.B1(n_161),
.B2(n_165),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_129),
.B(n_74),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_149),
.B(n_156),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_110),
.B(n_71),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_151),
.B(n_153),
.Y(n_190)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_134),
.Y(n_152)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_152),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_114),
.B(n_71),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_129),
.B(n_89),
.Y(n_156)
);

INVx6_ASAP7_75t_L g157 ( 
.A(n_116),
.Y(n_157)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_157),
.Y(n_170)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_122),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_159),
.B(n_113),
.C(n_123),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_115),
.A2(n_106),
.B1(n_131),
.B2(n_104),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_161),
.A2(n_125),
.B(n_130),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_125),
.B(n_78),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_165),
.B(n_80),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_155),
.A2(n_118),
.B(n_125),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_166),
.B(n_172),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_169),
.B(n_174),
.Y(n_195)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_160),
.B(n_125),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g197 ( 
.A(n_171),
.B(n_178),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_149),
.B(n_105),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_156),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_139),
.Y(n_175)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_175),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_142),
.A2(n_78),
.B1(n_89),
.B2(n_132),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_176),
.A2(n_136),
.B1(n_163),
.B2(n_144),
.Y(n_205)
);

OAI32xp33_ASAP7_75t_L g193 ( 
.A1(n_179),
.A2(n_146),
.A3(n_152),
.B1(n_141),
.B2(n_164),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_180),
.B(n_189),
.C(n_147),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_154),
.B(n_108),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_181),
.B(n_148),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_150),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_182),
.B(n_183),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_162),
.B(n_9),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_145),
.B(n_111),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_184),
.B(n_186),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_140),
.A2(n_85),
.B1(n_91),
.B2(n_98),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_185),
.A2(n_187),
.B1(n_163),
.B2(n_138),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_159),
.B(n_85),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_164),
.B(n_10),
.Y(n_188)
);

OAI21xp33_ASAP7_75t_L g208 ( 
.A1(n_188),
.A2(n_144),
.B(n_138),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_164),
.B(n_10),
.C(n_143),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_139),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_191),
.Y(n_200)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_192),
.Y(n_214)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_193),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_182),
.B(n_143),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_198),
.B(n_206),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_SL g226 ( 
.A(n_201),
.B(n_189),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_186),
.B(n_141),
.C(n_158),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_203),
.B(n_184),
.C(n_171),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_190),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_204),
.B(n_205),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_183),
.B(n_136),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_191),
.Y(n_207)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_207),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_208),
.B(n_185),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_172),
.B(n_180),
.Y(n_209)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_209),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_210),
.A2(n_212),
.B1(n_176),
.B2(n_170),
.Y(n_222)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_167),
.Y(n_211)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_211),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_187),
.A2(n_137),
.B1(n_157),
.B2(n_178),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_196),
.A2(n_169),
.B(n_166),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_213),
.A2(n_177),
.B(n_173),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_197),
.A2(n_171),
.B(n_179),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_216),
.A2(n_223),
.B(n_224),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_200),
.B(n_174),
.Y(n_218)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_218),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_222),
.A2(n_227),
.B1(n_193),
.B2(n_211),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_197),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_225),
.B(n_226),
.C(n_201),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_212),
.A2(n_195),
.B1(n_210),
.B2(n_196),
.Y(n_227)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_194),
.Y(n_229)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_229),
.Y(n_234)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_194),
.Y(n_230)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_230),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_218),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_231),
.B(n_228),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_224),
.A2(n_197),
.B(n_200),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_232),
.A2(n_235),
.B(n_239),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_236),
.B(n_237),
.C(n_241),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_226),
.B(n_202),
.C(n_203),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_213),
.A2(n_177),
.B(n_204),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_225),
.B(n_202),
.C(n_173),
.Y(n_241)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_242),
.Y(n_244)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_230),
.Y(n_243)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_243),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_245),
.B(n_247),
.Y(n_256)
);

BUFx12f_ASAP7_75t_SL g247 ( 
.A(n_239),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_232),
.A2(n_217),
.B(n_238),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_248),
.B(n_251),
.Y(n_261)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_233),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_237),
.B(n_227),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_252),
.B(n_241),
.Y(n_257)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_240),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_253),
.A2(n_254),
.B1(n_220),
.B2(n_215),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_234),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_255),
.B(n_257),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_SL g258 ( 
.A(n_252),
.B(n_249),
.Y(n_258)
);

OAI221xp5_ASAP7_75t_L g263 ( 
.A1(n_258),
.A2(n_262),
.B1(n_247),
.B2(n_249),
.C(n_221),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_244),
.A2(n_221),
.B1(n_242),
.B2(n_215),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_259),
.A2(n_223),
.B1(n_246),
.B2(n_216),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_250),
.B(n_236),
.C(n_219),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_260),
.A2(n_254),
.B(n_188),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_250),
.B(n_235),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_263),
.A2(n_266),
.B(n_199),
.Y(n_271)
);

INVx1_ASAP7_75t_SL g265 ( 
.A(n_256),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_265),
.B(n_267),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_261),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_268),
.B(n_258),
.Y(n_270)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_270),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_L g275 ( 
.A1(n_271),
.A2(n_167),
.B(n_168),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_265),
.A2(n_264),
.B(n_262),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_272),
.A2(n_273),
.B(n_214),
.Y(n_274)
);

MAJx2_ASAP7_75t_L g273 ( 
.A(n_265),
.B(n_260),
.C(n_257),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_274),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_275),
.A2(n_269),
.B(n_168),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_278),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_279),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_280),
.A2(n_277),
.B(n_276),
.Y(n_281)
);

BUFx24_ASAP7_75t_SL g282 ( 
.A(n_281),
.Y(n_282)
);


endmodule