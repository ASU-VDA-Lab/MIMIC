module fake_aes_3967_n_805 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_97, n_80, n_107, n_60, n_41, n_35, n_94, n_65, n_9, n_10, n_103, n_19, n_87, n_104, n_98, n_74, n_7, n_29, n_45, n_85, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_16, n_13, n_113, n_95, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_111, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_112, n_55, n_12, n_86, n_75, n_105, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_110, n_66, n_1, n_82, n_106, n_15, n_61, n_21, n_99, n_109, n_93, n_51, n_96, n_39, n_805);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_97;
input n_80;
input n_107;
input n_60;
input n_41;
input n_35;
input n_94;
input n_65;
input n_9;
input n_10;
input n_103;
input n_19;
input n_87;
input n_104;
input n_98;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_16;
input n_13;
input n_113;
input n_95;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_111;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_112;
input n_55;
input n_12;
input n_86;
input n_75;
input n_105;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_110;
input n_66;
input n_1;
input n_82;
input n_106;
input n_15;
input n_61;
input n_21;
input n_99;
input n_109;
input n_93;
input n_51;
input n_96;
input n_39;
output n_805;
wire n_117;
wire n_663;
wire n_707;
wire n_791;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_801;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_523;
wire n_229;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_252;
wire n_152;
wire n_637;
wire n_802;
wire n_353;
wire n_564;
wire n_779;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_762;
wire n_672;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_400;
wire n_787;
wire n_296;
wire n_157;
wire n_765;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_789;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_476;
wire n_227;
wire n_384;
wire n_434;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_777;
wire n_732;
wire n_752;
wire n_199;
wire n_351;
wire n_401;
wire n_461;
wire n_305;
wire n_599;
wire n_724;
wire n_228;
wire n_786;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_773;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_764;
wire n_314;
wire n_237;
wire n_181;
wire n_769;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_798;
wire n_241;
wire n_575;
wire n_711;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_767;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_490;
wire n_247;
wire n_648;
wire n_613;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_735;
wire n_696;
wire n_771;
wire n_784;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_746;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_803;
wire n_299;
wire n_338;
wire n_699;
wire n_519;
wire n_729;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_747;
wire n_635;
wire n_731;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_760;
wire n_751;
wire n_800;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_788;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_450;
wire n_579;
wire n_776;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_649;
wire n_526;
wire n_276;
wire n_320;
wire n_768;
wire n_797;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_666;
wire n_621;
wire n_799;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_754;
wire n_775;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_733;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_790;
wire n_761;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_396;
wire n_168;
wire n_804;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_723;
wire n_597;
wire n_749;
wire n_225;
wire n_535;
wire n_530;
wire n_737;
wire n_778;
wire n_220;
wire n_358;
wire n_795;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_782;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_734;
wire n_524;
wire n_121;
wire n_584;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_180;
wire n_441;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_766;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_774;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_722;
wire n_618;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_785;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_793;
wire n_182;
wire n_492;
wire n_592;
wire n_753;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_742;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_759;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_736;
wire n_194;
wire n_287;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_781;
wire n_421;
wire n_175;
wire n_709;
wire n_739;
wire n_145;
wire n_740;
wire n_483;
wire n_408;
wire n_772;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
BUFx3_ASAP7_75t_L g114 ( .A(n_49), .Y(n_114) );
CKINVDCx5p33_ASAP7_75t_R g115 ( .A(n_19), .Y(n_115) );
HB1xp67_ASAP7_75t_L g116 ( .A(n_110), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_79), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_81), .Y(n_118) );
CKINVDCx5p33_ASAP7_75t_R g119 ( .A(n_2), .Y(n_119) );
CKINVDCx5p33_ASAP7_75t_R g120 ( .A(n_13), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_50), .Y(n_121) );
BUFx6f_ASAP7_75t_L g122 ( .A(n_36), .Y(n_122) );
CKINVDCx5p33_ASAP7_75t_R g123 ( .A(n_63), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_105), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_31), .Y(n_125) );
CKINVDCx5p33_ASAP7_75t_R g126 ( .A(n_88), .Y(n_126) );
CKINVDCx5p33_ASAP7_75t_R g127 ( .A(n_47), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_9), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_111), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_59), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_97), .Y(n_131) );
INVx2_ASAP7_75t_L g132 ( .A(n_112), .Y(n_132) );
CKINVDCx5p33_ASAP7_75t_R g133 ( .A(n_90), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_68), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_38), .Y(n_135) );
CKINVDCx5p33_ASAP7_75t_R g136 ( .A(n_41), .Y(n_136) );
INVx2_ASAP7_75t_L g137 ( .A(n_87), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_39), .Y(n_138) );
CKINVDCx5p33_ASAP7_75t_R g139 ( .A(n_19), .Y(n_139) );
CKINVDCx5p33_ASAP7_75t_R g140 ( .A(n_12), .Y(n_140) );
NOR2xp67_ASAP7_75t_L g141 ( .A(n_107), .B(n_16), .Y(n_141) );
CKINVDCx5p33_ASAP7_75t_R g142 ( .A(n_17), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_0), .Y(n_143) );
CKINVDCx5p33_ASAP7_75t_R g144 ( .A(n_53), .Y(n_144) );
CKINVDCx5p33_ASAP7_75t_R g145 ( .A(n_80), .Y(n_145) );
BUFx10_ASAP7_75t_L g146 ( .A(n_104), .Y(n_146) );
INVx2_ASAP7_75t_SL g147 ( .A(n_34), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_45), .Y(n_148) );
HB1xp67_ASAP7_75t_L g149 ( .A(n_65), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_85), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_8), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_10), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_52), .Y(n_153) );
CKINVDCx20_ASAP7_75t_R g154 ( .A(n_76), .Y(n_154) );
CKINVDCx5p33_ASAP7_75t_R g155 ( .A(n_11), .Y(n_155) );
CKINVDCx5p33_ASAP7_75t_R g156 ( .A(n_91), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_18), .Y(n_157) );
INVx2_ASAP7_75t_L g158 ( .A(n_60), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_62), .Y(n_159) );
CKINVDCx5p33_ASAP7_75t_R g160 ( .A(n_56), .Y(n_160) );
CKINVDCx5p33_ASAP7_75t_R g161 ( .A(n_46), .Y(n_161) );
INVx2_ASAP7_75t_L g162 ( .A(n_122), .Y(n_162) );
BUFx8_ASAP7_75t_L g163 ( .A(n_147), .Y(n_163) );
INVx2_ASAP7_75t_L g164 ( .A(n_122), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_116), .B(n_0), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_117), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_118), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_121), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_124), .Y(n_169) );
AND2x4_ASAP7_75t_L g170 ( .A(n_147), .B(n_1), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_125), .Y(n_171) );
BUFx6f_ASAP7_75t_L g172 ( .A(n_122), .Y(n_172) );
OAI21x1_ASAP7_75t_L g173 ( .A1(n_132), .A2(n_51), .B(n_109), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_129), .Y(n_174) );
INVx3_ASAP7_75t_L g175 ( .A(n_146), .Y(n_175) );
OA21x2_ASAP7_75t_L g176 ( .A1(n_132), .A2(n_48), .B(n_108), .Y(n_176) );
INVx2_ASAP7_75t_L g177 ( .A(n_122), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_130), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_131), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_149), .B(n_1), .Y(n_180) );
INVx2_ASAP7_75t_L g181 ( .A(n_122), .Y(n_181) );
INVx3_ASAP7_75t_L g182 ( .A(n_146), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_128), .B(n_2), .Y(n_183) );
OR2x6_ASAP7_75t_L g184 ( .A(n_165), .B(n_143), .Y(n_184) );
INVx2_ASAP7_75t_SL g185 ( .A(n_175), .Y(n_185) );
NAND3xp33_ASAP7_75t_L g186 ( .A(n_165), .B(n_142), .C(n_115), .Y(n_186) );
INVx2_ASAP7_75t_L g187 ( .A(n_162), .Y(n_187) );
INVx2_ASAP7_75t_L g188 ( .A(n_162), .Y(n_188) );
INVx2_ASAP7_75t_L g189 ( .A(n_162), .Y(n_189) );
AND3x1_ASAP7_75t_L g190 ( .A(n_175), .B(n_152), .C(n_151), .Y(n_190) );
BUFx3_ASAP7_75t_L g191 ( .A(n_170), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_170), .Y(n_192) );
AND2x4_ASAP7_75t_L g193 ( .A(n_175), .B(n_157), .Y(n_193) );
BUFx6f_ASAP7_75t_L g194 ( .A(n_172), .Y(n_194) );
INVx2_ASAP7_75t_L g195 ( .A(n_164), .Y(n_195) );
INVx2_ASAP7_75t_L g196 ( .A(n_164), .Y(n_196) );
INVx2_ASAP7_75t_L g197 ( .A(n_164), .Y(n_197) );
AND2x6_ASAP7_75t_L g198 ( .A(n_170), .B(n_114), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_170), .Y(n_199) );
BUFx6f_ASAP7_75t_L g200 ( .A(n_172), .Y(n_200) );
NAND2xp5_ASAP7_75t_SL g201 ( .A(n_175), .B(n_146), .Y(n_201) );
INVx3_ASAP7_75t_L g202 ( .A(n_173), .Y(n_202) );
INVx2_ASAP7_75t_L g203 ( .A(n_177), .Y(n_203) );
INVx2_ASAP7_75t_L g204 ( .A(n_177), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_177), .Y(n_205) );
INVx1_ASAP7_75t_L g206 ( .A(n_181), .Y(n_206) );
OR2x6_ASAP7_75t_L g207 ( .A(n_180), .B(n_141), .Y(n_207) );
INVx2_ASAP7_75t_L g208 ( .A(n_181), .Y(n_208) );
CKINVDCx6p67_ASAP7_75t_R g209 ( .A(n_180), .Y(n_209) );
INVx2_ASAP7_75t_L g210 ( .A(n_181), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_182), .B(n_115), .Y(n_211) );
INVx1_ASAP7_75t_L g212 ( .A(n_173), .Y(n_212) );
INVx2_ASAP7_75t_L g213 ( .A(n_172), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_173), .Y(n_214) );
AOI22xp33_ASAP7_75t_L g215 ( .A1(n_166), .A2(n_140), .B1(n_119), .B2(n_142), .Y(n_215) );
AOI222xp33_ASAP7_75t_L g216 ( .A1(n_215), .A2(n_186), .B1(n_183), .B2(n_168), .C1(n_169), .C2(n_171), .Y(n_216) );
OR2x6_ASAP7_75t_L g217 ( .A(n_184), .B(n_182), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_192), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_211), .B(n_182), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_184), .B(n_182), .Y(n_220) );
INVx1_ASAP7_75t_L g221 ( .A(n_192), .Y(n_221) );
BUFx6f_ASAP7_75t_SL g222 ( .A(n_198), .Y(n_222) );
NAND2xp5_ASAP7_75t_SL g223 ( .A(n_199), .B(n_163), .Y(n_223) );
O2A1O1Ixp5_ASAP7_75t_L g224 ( .A1(n_202), .A2(n_174), .B(n_179), .C(n_178), .Y(n_224) );
NOR2xp67_ASAP7_75t_L g225 ( .A(n_201), .B(n_166), .Y(n_225) );
NAND2xp5_ASAP7_75t_SL g226 ( .A(n_199), .B(n_163), .Y(n_226) );
AND2x2_ASAP7_75t_L g227 ( .A(n_184), .B(n_167), .Y(n_227) );
NOR2xp67_ASAP7_75t_L g228 ( .A(n_193), .B(n_167), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_184), .B(n_163), .Y(n_229) );
NOR2xp33_ASAP7_75t_SL g230 ( .A(n_209), .B(n_154), .Y(n_230) );
AOI22xp33_ASAP7_75t_L g231 ( .A1(n_198), .A2(n_171), .B1(n_179), .B2(n_178), .Y(n_231) );
INVxp67_ASAP7_75t_L g232 ( .A(n_190), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_193), .B(n_163), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_193), .B(n_168), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_193), .Y(n_235) );
HB1xp67_ASAP7_75t_L g236 ( .A(n_209), .Y(n_236) );
AND2x2_ASAP7_75t_L g237 ( .A(n_191), .B(n_169), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_185), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_185), .B(n_174), .Y(n_239) );
AND2x2_ASAP7_75t_SL g240 ( .A(n_190), .B(n_176), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_191), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_198), .B(n_123), .Y(n_242) );
NOR2xp33_ASAP7_75t_L g243 ( .A(n_207), .B(n_183), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_212), .Y(n_244) );
NOR2xp33_ASAP7_75t_L g245 ( .A(n_207), .B(n_123), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_198), .B(n_144), .Y(n_246) );
A2O1A1Ixp33_ASAP7_75t_L g247 ( .A1(n_212), .A2(n_135), .B(n_148), .C(n_150), .Y(n_247) );
NOR2xp33_ASAP7_75t_L g248 ( .A(n_207), .B(n_144), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_198), .B(n_145), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_207), .Y(n_250) );
AND2x2_ASAP7_75t_L g251 ( .A(n_198), .B(n_119), .Y(n_251) );
OAI22xp33_ASAP7_75t_L g252 ( .A1(n_214), .A2(n_140), .B1(n_120), .B2(n_155), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_198), .B(n_145), .Y(n_253) );
AND2x6_ASAP7_75t_SL g254 ( .A(n_214), .B(n_134), .Y(n_254) );
BUFx3_ASAP7_75t_L g255 ( .A(n_202), .Y(n_255) );
INVx2_ASAP7_75t_SL g256 ( .A(n_202), .Y(n_256) );
AOI22xp5_ASAP7_75t_L g257 ( .A1(n_205), .A2(n_155), .B1(n_120), .B2(n_139), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_205), .B(n_156), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_206), .B(n_156), .Y(n_259) );
AOI21xp5_ASAP7_75t_L g260 ( .A1(n_244), .A2(n_176), .B(n_206), .Y(n_260) );
AOI21xp5_ASAP7_75t_L g261 ( .A1(n_244), .A2(n_176), .B(n_210), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_227), .B(n_160), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_227), .B(n_160), .Y(n_263) );
A2O1A1Ixp33_ASAP7_75t_L g264 ( .A1(n_218), .A2(n_138), .B(n_153), .C(n_159), .Y(n_264) );
AOI21xp5_ASAP7_75t_L g265 ( .A1(n_223), .A2(n_176), .B(n_210), .Y(n_265) );
INVx3_ASAP7_75t_L g266 ( .A(n_235), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_243), .B(n_161), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_216), .B(n_161), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_228), .B(n_126), .Y(n_269) );
AOI21xp5_ASAP7_75t_L g270 ( .A1(n_223), .A2(n_176), .B(n_208), .Y(n_270) );
INVx4_ASAP7_75t_L g271 ( .A(n_217), .Y(n_271) );
AOI22xp33_ASAP7_75t_L g272 ( .A1(n_251), .A2(n_114), .B1(n_137), .B2(n_158), .Y(n_272) );
NAND2xp5_ASAP7_75t_SL g273 ( .A(n_229), .B(n_127), .Y(n_273) );
INVx3_ASAP7_75t_L g274 ( .A(n_222), .Y(n_274) );
AOI21x1_ASAP7_75t_L g275 ( .A1(n_226), .A2(n_213), .B(n_208), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_237), .B(n_133), .Y(n_276) );
AOI21xp5_ASAP7_75t_L g277 ( .A1(n_226), .A2(n_256), .B(n_233), .Y(n_277) );
HB1xp67_ASAP7_75t_L g278 ( .A(n_217), .Y(n_278) );
OAI21xp33_ASAP7_75t_L g279 ( .A1(n_257), .A2(n_136), .B(n_158), .Y(n_279) );
AO21x1_ASAP7_75t_L g280 ( .A1(n_218), .A2(n_137), .B(n_204), .Y(n_280) );
OAI22xp5_ASAP7_75t_L g281 ( .A1(n_217), .A2(n_195), .B1(n_204), .B2(n_203), .Y(n_281) );
OR2x6_ASAP7_75t_L g282 ( .A(n_217), .B(n_172), .Y(n_282) );
OR2x6_ASAP7_75t_L g283 ( .A(n_236), .B(n_172), .Y(n_283) );
AOI21xp5_ASAP7_75t_L g284 ( .A1(n_256), .A2(n_195), .B(n_203), .Y(n_284) );
NOR2xp67_ASAP7_75t_R g285 ( .A(n_221), .B(n_187), .Y(n_285) );
AOI22xp5_ASAP7_75t_L g286 ( .A1(n_232), .A2(n_187), .B1(n_197), .B2(n_196), .Y(n_286) );
AOI21xp33_ASAP7_75t_L g287 ( .A1(n_245), .A2(n_188), .B(n_189), .Y(n_287) );
AOI21xp5_ASAP7_75t_L g288 ( .A1(n_221), .A2(n_188), .B(n_197), .Y(n_288) );
NOR2xp33_ASAP7_75t_L g289 ( .A(n_250), .B(n_3), .Y(n_289) );
OAI21x1_ASAP7_75t_L g290 ( .A1(n_224), .A2(n_213), .B(n_196), .Y(n_290) );
AOI21xp5_ASAP7_75t_L g291 ( .A1(n_255), .A2(n_189), .B(n_194), .Y(n_291) );
BUFx2_ASAP7_75t_L g292 ( .A(n_251), .Y(n_292) );
OAI22xp5_ASAP7_75t_L g293 ( .A1(n_231), .A2(n_172), .B1(n_4), .B2(n_5), .Y(n_293) );
NAND2xp5_ASAP7_75t_SL g294 ( .A(n_252), .B(n_194), .Y(n_294) );
O2A1O1Ixp33_ASAP7_75t_L g295 ( .A1(n_247), .A2(n_3), .B(n_4), .C(n_5), .Y(n_295) );
BUFx6f_ASAP7_75t_L g296 ( .A(n_255), .Y(n_296) );
NOR2xp33_ASAP7_75t_L g297 ( .A(n_248), .B(n_6), .Y(n_297) );
OR2x2_ASAP7_75t_L g298 ( .A(n_262), .B(n_220), .Y(n_298) );
NOR2xp33_ASAP7_75t_L g299 ( .A(n_263), .B(n_234), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_292), .B(n_237), .Y(n_300) );
AO22x2_ASAP7_75t_L g301 ( .A1(n_271), .A2(n_254), .B1(n_230), .B2(n_240), .Y(n_301) );
AOI221xp5_ASAP7_75t_SL g302 ( .A1(n_264), .A2(n_268), .B1(n_247), .B2(n_279), .C(n_272), .Y(n_302) );
CKINVDCx20_ASAP7_75t_R g303 ( .A(n_271), .Y(n_303) );
INVx5_ASAP7_75t_L g304 ( .A(n_282), .Y(n_304) );
BUFx3_ASAP7_75t_L g305 ( .A(n_282), .Y(n_305) );
OAI21x1_ASAP7_75t_L g306 ( .A1(n_275), .A2(n_238), .B(n_241), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_278), .B(n_225), .Y(n_307) );
INVxp67_ASAP7_75t_L g308 ( .A(n_289), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_297), .B(n_219), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_267), .B(n_239), .Y(n_310) );
AOI21x1_ASAP7_75t_L g311 ( .A1(n_261), .A2(n_259), .B(n_258), .Y(n_311) );
AOI21xp5_ASAP7_75t_L g312 ( .A1(n_277), .A2(n_240), .B(n_249), .Y(n_312) );
AO31x2_ASAP7_75t_L g313 ( .A1(n_280), .A2(n_253), .A3(n_246), .B(n_242), .Y(n_313) );
AND2x4_ASAP7_75t_L g314 ( .A(n_282), .B(n_222), .Y(n_314) );
OAI22xp5_ASAP7_75t_L g315 ( .A1(n_281), .A2(n_222), .B1(n_7), .B2(n_8), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_276), .B(n_6), .Y(n_316) );
OAI21x1_ASAP7_75t_L g317 ( .A1(n_265), .A2(n_200), .B(n_194), .Y(n_317) );
AOI21xp5_ASAP7_75t_L g318 ( .A1(n_270), .A2(n_200), .B(n_194), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_266), .Y(n_319) );
NOR2xp33_ASAP7_75t_L g320 ( .A(n_273), .B(n_7), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_266), .Y(n_321) );
INVx2_ASAP7_75t_L g322 ( .A(n_290), .Y(n_322) );
AOI21x1_ASAP7_75t_L g323 ( .A1(n_260), .A2(n_200), .B(n_194), .Y(n_323) );
OAI21x1_ASAP7_75t_L g324 ( .A1(n_291), .A2(n_200), .B(n_58), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_269), .B(n_9), .Y(n_325) );
AO21x2_ASAP7_75t_L g326 ( .A1(n_322), .A2(n_294), .B(n_295), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_299), .B(n_285), .Y(n_327) );
AOI21x1_ASAP7_75t_L g328 ( .A1(n_323), .A2(n_284), .B(n_288), .Y(n_328) );
OAI22xp5_ASAP7_75t_L g329 ( .A1(n_301), .A2(n_283), .B1(n_293), .B2(n_296), .Y(n_329) );
INVx3_ASAP7_75t_L g330 ( .A(n_304), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_319), .Y(n_331) );
INVx2_ASAP7_75t_L g332 ( .A(n_322), .Y(n_332) );
OAI21x1_ASAP7_75t_L g333 ( .A1(n_317), .A2(n_274), .B(n_285), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_321), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_300), .Y(n_335) );
BUFx2_ASAP7_75t_SL g336 ( .A(n_304), .Y(n_336) );
INVx3_ASAP7_75t_L g337 ( .A(n_304), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_299), .B(n_286), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_316), .Y(n_339) );
AND2x4_ASAP7_75t_L g340 ( .A(n_314), .B(n_274), .Y(n_340) );
INVx3_ASAP7_75t_L g341 ( .A(n_304), .Y(n_341) );
OAI21x1_ASAP7_75t_L g342 ( .A1(n_317), .A2(n_296), .B(n_287), .Y(n_342) );
NOR2xp33_ASAP7_75t_L g343 ( .A(n_308), .B(n_283), .Y(n_343) );
OA21x2_ASAP7_75t_L g344 ( .A1(n_318), .A2(n_296), .B(n_200), .Y(n_344) );
AOI22xp5_ASAP7_75t_L g345 ( .A1(n_301), .A2(n_283), .B1(n_11), .B2(n_12), .Y(n_345) );
AND2x4_ASAP7_75t_L g346 ( .A(n_314), .B(n_64), .Y(n_346) );
INVx4_ASAP7_75t_L g347 ( .A(n_314), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_310), .B(n_10), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_298), .B(n_13), .Y(n_349) );
INVx2_ASAP7_75t_L g350 ( .A(n_332), .Y(n_350) );
BUFx3_ASAP7_75t_L g351 ( .A(n_330), .Y(n_351) );
INVx3_ASAP7_75t_L g352 ( .A(n_347), .Y(n_352) );
OAI21x1_ASAP7_75t_L g353 ( .A1(n_342), .A2(n_324), .B(n_311), .Y(n_353) );
INVx2_ASAP7_75t_L g354 ( .A(n_332), .Y(n_354) );
OA21x2_ASAP7_75t_L g355 ( .A1(n_342), .A2(n_324), .B(n_312), .Y(n_355) );
AO21x2_ASAP7_75t_L g356 ( .A1(n_328), .A2(n_325), .B(n_309), .Y(n_356) );
OAI21x1_ASAP7_75t_L g357 ( .A1(n_333), .A2(n_306), .B(n_315), .Y(n_357) );
HB1xp67_ASAP7_75t_L g358 ( .A(n_332), .Y(n_358) );
AND2x2_ASAP7_75t_L g359 ( .A(n_339), .B(n_301), .Y(n_359) );
OAI21x1_ASAP7_75t_L g360 ( .A1(n_333), .A2(n_307), .B(n_320), .Y(n_360) );
HB1xp67_ASAP7_75t_L g361 ( .A(n_327), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_331), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_331), .Y(n_363) );
BUFx2_ASAP7_75t_L g364 ( .A(n_330), .Y(n_364) );
AND2x2_ASAP7_75t_L g365 ( .A(n_339), .B(n_313), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_334), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_334), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_335), .Y(n_368) );
AND2x2_ASAP7_75t_L g369 ( .A(n_345), .B(n_313), .Y(n_369) );
INVx3_ASAP7_75t_L g370 ( .A(n_347), .Y(n_370) );
HB1xp67_ASAP7_75t_L g371 ( .A(n_327), .Y(n_371) );
INVx2_ASAP7_75t_L g372 ( .A(n_344), .Y(n_372) );
INVx2_ASAP7_75t_L g373 ( .A(n_344), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_335), .Y(n_374) );
INVx2_ASAP7_75t_L g375 ( .A(n_344), .Y(n_375) );
INVx2_ASAP7_75t_SL g376 ( .A(n_330), .Y(n_376) );
INVx2_ASAP7_75t_L g377 ( .A(n_344), .Y(n_377) );
OA21x2_ASAP7_75t_L g378 ( .A1(n_333), .A2(n_302), .B(n_320), .Y(n_378) );
HB1xp67_ASAP7_75t_L g379 ( .A(n_330), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_358), .Y(n_380) );
AND2x2_ASAP7_75t_L g381 ( .A(n_365), .B(n_345), .Y(n_381) );
NAND3xp33_ASAP7_75t_L g382 ( .A(n_365), .B(n_348), .C(n_349), .Y(n_382) );
AOI22xp5_ASAP7_75t_L g383 ( .A1(n_359), .A2(n_338), .B1(n_348), .B2(n_303), .Y(n_383) );
AND2x2_ASAP7_75t_L g384 ( .A(n_365), .B(n_326), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_368), .B(n_338), .Y(n_385) );
AND2x2_ASAP7_75t_L g386 ( .A(n_358), .B(n_326), .Y(n_386) );
INVx3_ASAP7_75t_L g387 ( .A(n_372), .Y(n_387) );
HB1xp67_ASAP7_75t_L g388 ( .A(n_379), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_363), .Y(n_389) );
AND2x2_ASAP7_75t_L g390 ( .A(n_359), .B(n_326), .Y(n_390) );
NAND2x1p5_ASAP7_75t_L g391 ( .A(n_352), .B(n_346), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_363), .Y(n_392) );
HB1xp67_ASAP7_75t_L g393 ( .A(n_379), .Y(n_393) );
NOR4xp25_ASAP7_75t_SL g394 ( .A(n_364), .B(n_336), .C(n_329), .D(n_346), .Y(n_394) );
BUFx3_ASAP7_75t_L g395 ( .A(n_351), .Y(n_395) );
INVx2_ASAP7_75t_L g396 ( .A(n_350), .Y(n_396) );
INVxp67_ASAP7_75t_SL g397 ( .A(n_350), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_368), .B(n_349), .Y(n_398) );
INVx2_ASAP7_75t_L g399 ( .A(n_350), .Y(n_399) );
AND2x2_ASAP7_75t_L g400 ( .A(n_359), .B(n_326), .Y(n_400) );
AND2x2_ASAP7_75t_L g401 ( .A(n_369), .B(n_346), .Y(n_401) );
CKINVDCx5p33_ASAP7_75t_R g402 ( .A(n_351), .Y(n_402) );
INVx2_ASAP7_75t_L g403 ( .A(n_350), .Y(n_403) );
AND2x2_ASAP7_75t_L g404 ( .A(n_369), .B(n_346), .Y(n_404) );
BUFx2_ASAP7_75t_L g405 ( .A(n_364), .Y(n_405) );
HB1xp67_ASAP7_75t_L g406 ( .A(n_374), .Y(n_406) );
BUFx5_ASAP7_75t_L g407 ( .A(n_351), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_363), .Y(n_408) );
INVx8_ASAP7_75t_L g409 ( .A(n_352), .Y(n_409) );
AND2x2_ASAP7_75t_L g410 ( .A(n_369), .B(n_347), .Y(n_410) );
AOI22xp33_ASAP7_75t_SL g411 ( .A1(n_352), .A2(n_347), .B1(n_336), .B2(n_329), .Y(n_411) );
AND2x2_ASAP7_75t_L g412 ( .A(n_366), .B(n_337), .Y(n_412) );
INVx2_ASAP7_75t_L g413 ( .A(n_354), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_374), .B(n_337), .Y(n_414) );
INVx2_ASAP7_75t_L g415 ( .A(n_354), .Y(n_415) );
AND2x2_ASAP7_75t_L g416 ( .A(n_366), .B(n_337), .Y(n_416) );
AND2x4_ASAP7_75t_L g417 ( .A(n_372), .B(n_373), .Y(n_417) );
AND2x4_ASAP7_75t_L g418 ( .A(n_372), .B(n_337), .Y(n_418) );
INVxp67_ASAP7_75t_L g419 ( .A(n_364), .Y(n_419) );
AND2x2_ASAP7_75t_L g420 ( .A(n_366), .B(n_341), .Y(n_420) );
INVx2_ASAP7_75t_L g421 ( .A(n_354), .Y(n_421) );
AND2x2_ASAP7_75t_L g422 ( .A(n_362), .B(n_341), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_354), .Y(n_423) );
OAI22xp5_ASAP7_75t_L g424 ( .A1(n_361), .A2(n_303), .B1(n_341), .B2(n_305), .Y(n_424) );
AND2x2_ASAP7_75t_L g425 ( .A(n_362), .B(n_341), .Y(n_425) );
NOR2xp33_ASAP7_75t_L g426 ( .A(n_367), .B(n_343), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_367), .B(n_340), .Y(n_427) );
OAI222xp33_ASAP7_75t_L g428 ( .A1(n_376), .A2(n_340), .B1(n_305), .B2(n_328), .C1(n_17), .C2(n_18), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_361), .B(n_340), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_389), .B(n_371), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_389), .Y(n_431) );
AND2x2_ASAP7_75t_L g432 ( .A(n_384), .B(n_371), .Y(n_432) );
AND2x2_ASAP7_75t_L g433 ( .A(n_384), .B(n_372), .Y(n_433) );
BUFx2_ASAP7_75t_L g434 ( .A(n_418), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_392), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_426), .B(n_376), .Y(n_436) );
OR2x2_ASAP7_75t_L g437 ( .A(n_380), .B(n_373), .Y(n_437) );
AND2x4_ASAP7_75t_L g438 ( .A(n_418), .B(n_373), .Y(n_438) );
INVx3_ASAP7_75t_L g439 ( .A(n_387), .Y(n_439) );
NOR2x1_ASAP7_75t_L g440 ( .A(n_424), .B(n_351), .Y(n_440) );
OR2x2_ASAP7_75t_L g441 ( .A(n_380), .B(n_373), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_390), .B(n_375), .Y(n_442) );
OR2x2_ASAP7_75t_L g443 ( .A(n_388), .B(n_375), .Y(n_443) );
INVx2_ASAP7_75t_L g444 ( .A(n_396), .Y(n_444) );
AND2x2_ASAP7_75t_L g445 ( .A(n_390), .B(n_375), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_406), .B(n_376), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_385), .B(n_352), .Y(n_447) );
INVxp67_ASAP7_75t_L g448 ( .A(n_393), .Y(n_448) );
INVx1_ASAP7_75t_SL g449 ( .A(n_402), .Y(n_449) );
CKINVDCx5p33_ASAP7_75t_R g450 ( .A(n_409), .Y(n_450) );
INVx2_ASAP7_75t_L g451 ( .A(n_396), .Y(n_451) );
OR2x2_ASAP7_75t_L g452 ( .A(n_405), .B(n_375), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_392), .B(n_352), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_408), .Y(n_454) );
AND2x2_ASAP7_75t_L g455 ( .A(n_400), .B(n_377), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_408), .Y(n_456) );
AND2x2_ASAP7_75t_L g457 ( .A(n_400), .B(n_377), .Y(n_457) );
HB1xp67_ASAP7_75t_L g458 ( .A(n_405), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_423), .Y(n_459) );
INVx2_ASAP7_75t_L g460 ( .A(n_396), .Y(n_460) );
INVx1_ASAP7_75t_SL g461 ( .A(n_418), .Y(n_461) );
AND2x2_ASAP7_75t_L g462 ( .A(n_401), .B(n_377), .Y(n_462) );
INVxp33_ASAP7_75t_L g463 ( .A(n_391), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_422), .B(n_370), .Y(n_464) );
AND2x2_ASAP7_75t_L g465 ( .A(n_401), .B(n_377), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_423), .Y(n_466) );
AND2x2_ASAP7_75t_L g467 ( .A(n_404), .B(n_360), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_422), .B(n_370), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_399), .Y(n_469) );
AND2x2_ASAP7_75t_L g470 ( .A(n_404), .B(n_360), .Y(n_470) );
INVx2_ASAP7_75t_L g471 ( .A(n_399), .Y(n_471) );
HB1xp67_ASAP7_75t_L g472 ( .A(n_419), .Y(n_472) );
INVx2_ASAP7_75t_L g473 ( .A(n_399), .Y(n_473) );
AND2x2_ASAP7_75t_L g474 ( .A(n_410), .B(n_360), .Y(n_474) );
AND2x2_ASAP7_75t_L g475 ( .A(n_410), .B(n_378), .Y(n_475) );
AND2x2_ASAP7_75t_L g476 ( .A(n_381), .B(n_378), .Y(n_476) );
INVx2_ASAP7_75t_L g477 ( .A(n_403), .Y(n_477) );
AND2x2_ASAP7_75t_L g478 ( .A(n_381), .B(n_378), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_425), .B(n_370), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_403), .Y(n_480) );
AND2x4_ASAP7_75t_L g481 ( .A(n_418), .B(n_353), .Y(n_481) );
AND2x2_ASAP7_75t_L g482 ( .A(n_417), .B(n_378), .Y(n_482) );
AND2x2_ASAP7_75t_L g483 ( .A(n_417), .B(n_378), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_403), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_413), .Y(n_485) );
AND2x2_ASAP7_75t_L g486 ( .A(n_417), .B(n_378), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_413), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_413), .Y(n_488) );
AND2x4_ASAP7_75t_L g489 ( .A(n_417), .B(n_353), .Y(n_489) );
AND2x2_ASAP7_75t_L g490 ( .A(n_387), .B(n_356), .Y(n_490) );
AND2x2_ASAP7_75t_L g491 ( .A(n_387), .B(n_356), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_425), .B(n_370), .Y(n_492) );
INVx2_ASAP7_75t_L g493 ( .A(n_415), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_415), .Y(n_494) );
INVx2_ASAP7_75t_L g495 ( .A(n_415), .Y(n_495) );
INVx2_ASAP7_75t_L g496 ( .A(n_421), .Y(n_496) );
INVx2_ASAP7_75t_L g497 ( .A(n_421), .Y(n_497) );
AND2x2_ASAP7_75t_L g498 ( .A(n_387), .B(n_356), .Y(n_498) );
BUFx3_ASAP7_75t_L g499 ( .A(n_409), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_421), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_412), .B(n_370), .Y(n_501) );
AND2x2_ASAP7_75t_L g502 ( .A(n_397), .B(n_356), .Y(n_502) );
OR2x2_ASAP7_75t_L g503 ( .A(n_429), .B(n_356), .Y(n_503) );
AND2x2_ASAP7_75t_L g504 ( .A(n_386), .B(n_412), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_431), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_431), .Y(n_506) );
INVx2_ASAP7_75t_SL g507 ( .A(n_443), .Y(n_507) );
INVx1_ASAP7_75t_SL g508 ( .A(n_449), .Y(n_508) );
BUFx2_ASAP7_75t_L g509 ( .A(n_450), .Y(n_509) );
OR2x2_ASAP7_75t_L g510 ( .A(n_432), .B(n_416), .Y(n_510) );
OR2x2_ASAP7_75t_L g511 ( .A(n_432), .B(n_416), .Y(n_511) );
INVx2_ASAP7_75t_L g512 ( .A(n_444), .Y(n_512) );
INVxp67_ASAP7_75t_L g513 ( .A(n_458), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_435), .Y(n_514) );
NOR2x1_ASAP7_75t_L g515 ( .A(n_499), .B(n_424), .Y(n_515) );
OR2x2_ASAP7_75t_L g516 ( .A(n_504), .B(n_420), .Y(n_516) );
AND2x2_ASAP7_75t_L g517 ( .A(n_504), .B(n_420), .Y(n_517) );
INVx2_ASAP7_75t_L g518 ( .A(n_444), .Y(n_518) );
OR2x2_ASAP7_75t_L g519 ( .A(n_433), .B(n_395), .Y(n_519) );
NOR2xp33_ASAP7_75t_L g520 ( .A(n_448), .B(n_383), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_435), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_433), .B(n_383), .Y(n_522) );
INVx2_ASAP7_75t_L g523 ( .A(n_444), .Y(n_523) );
AND2x2_ASAP7_75t_L g524 ( .A(n_462), .B(n_395), .Y(n_524) );
NOR2x1p5_ASAP7_75t_L g525 ( .A(n_499), .B(n_395), .Y(n_525) );
AND2x2_ASAP7_75t_L g526 ( .A(n_462), .B(n_465), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_476), .B(n_382), .Y(n_527) );
INVx2_ASAP7_75t_SL g528 ( .A(n_443), .Y(n_528) );
INVxp67_ASAP7_75t_L g529 ( .A(n_440), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_476), .B(n_382), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_454), .Y(n_531) );
OR2x2_ASAP7_75t_L g532 ( .A(n_442), .B(n_427), .Y(n_532) );
OR2x2_ASAP7_75t_L g533 ( .A(n_442), .B(n_414), .Y(n_533) );
AND2x2_ASAP7_75t_L g534 ( .A(n_475), .B(n_386), .Y(n_534) );
AND2x2_ASAP7_75t_L g535 ( .A(n_475), .B(n_407), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_454), .Y(n_536) );
HB1xp67_ASAP7_75t_L g537 ( .A(n_452), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_478), .B(n_398), .Y(n_538) );
AND2x2_ASAP7_75t_L g539 ( .A(n_465), .B(n_407), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_456), .Y(n_540) );
OR2x2_ASAP7_75t_L g541 ( .A(n_445), .B(n_407), .Y(n_541) );
AOI22xp33_ASAP7_75t_L g542 ( .A1(n_436), .A2(n_411), .B1(n_391), .B2(n_340), .Y(n_542) );
INVx2_ASAP7_75t_L g543 ( .A(n_451), .Y(n_543) );
AND2x2_ASAP7_75t_L g544 ( .A(n_445), .B(n_407), .Y(n_544) );
NOR2xp33_ASAP7_75t_L g545 ( .A(n_449), .B(n_428), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_478), .B(n_407), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_456), .Y(n_547) );
AND2x2_ASAP7_75t_L g548 ( .A(n_455), .B(n_407), .Y(n_548) );
BUFx2_ASAP7_75t_L g549 ( .A(n_499), .Y(n_549) );
INVx2_ASAP7_75t_L g550 ( .A(n_451), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_455), .B(n_407), .Y(n_551) );
NAND2xp5_ASAP7_75t_SL g552 ( .A(n_440), .B(n_407), .Y(n_552) );
OR2x2_ASAP7_75t_L g553 ( .A(n_457), .B(n_407), .Y(n_553) );
INVx2_ASAP7_75t_L g554 ( .A(n_451), .Y(n_554) );
NOR2x1_ASAP7_75t_L g555 ( .A(n_446), .B(n_409), .Y(n_555) );
OR2x2_ASAP7_75t_L g556 ( .A(n_457), .B(n_391), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_430), .B(n_409), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_430), .B(n_409), .Y(n_558) );
BUFx3_ASAP7_75t_L g559 ( .A(n_434), .Y(n_559) );
AND2x2_ASAP7_75t_L g560 ( .A(n_434), .B(n_394), .Y(n_560) );
OR2x2_ASAP7_75t_L g561 ( .A(n_437), .B(n_355), .Y(n_561) );
AND2x2_ASAP7_75t_L g562 ( .A(n_472), .B(n_394), .Y(n_562) );
INVx2_ASAP7_75t_L g563 ( .A(n_460), .Y(n_563) );
HB1xp67_ASAP7_75t_L g564 ( .A(n_452), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_459), .Y(n_565) );
AND2x2_ASAP7_75t_L g566 ( .A(n_474), .B(n_355), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_459), .Y(n_567) );
INVx1_ASAP7_75t_SL g568 ( .A(n_461), .Y(n_568) );
INVx3_ASAP7_75t_SL g569 ( .A(n_438), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_466), .Y(n_570) );
AND2x2_ASAP7_75t_L g571 ( .A(n_474), .B(n_355), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_466), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_453), .Y(n_573) );
INVx2_ASAP7_75t_L g574 ( .A(n_460), .Y(n_574) );
AND2x4_ASAP7_75t_L g575 ( .A(n_489), .B(n_353), .Y(n_575) );
INVx2_ASAP7_75t_L g576 ( .A(n_460), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_447), .B(n_355), .Y(n_577) );
NOR2xp33_ASAP7_75t_L g578 ( .A(n_503), .B(n_14), .Y(n_578) );
AND2x4_ASAP7_75t_L g579 ( .A(n_489), .B(n_357), .Y(n_579) );
AND2x4_ASAP7_75t_L g580 ( .A(n_489), .B(n_357), .Y(n_580) );
INVx2_ASAP7_75t_L g581 ( .A(n_471), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_437), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_441), .Y(n_583) );
AND2x2_ASAP7_75t_L g584 ( .A(n_467), .B(n_355), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_503), .B(n_355), .Y(n_585) );
NOR2xp67_ASAP7_75t_L g586 ( .A(n_439), .B(n_14), .Y(n_586) );
INVx2_ASAP7_75t_SL g587 ( .A(n_441), .Y(n_587) );
INVx2_ASAP7_75t_L g588 ( .A(n_471), .Y(n_588) );
INVx2_ASAP7_75t_L g589 ( .A(n_471), .Y(n_589) );
OR2x2_ASAP7_75t_L g590 ( .A(n_501), .B(n_15), .Y(n_590) );
AND2x2_ASAP7_75t_L g591 ( .A(n_467), .B(n_357), .Y(n_591) );
INVx1_ASAP7_75t_SL g592 ( .A(n_461), .Y(n_592) );
INVx2_ASAP7_75t_L g593 ( .A(n_473), .Y(n_593) );
AND2x2_ASAP7_75t_L g594 ( .A(n_470), .B(n_15), .Y(n_594) );
AND2x2_ASAP7_75t_L g595 ( .A(n_526), .B(n_470), .Y(n_595) );
AND2x4_ASAP7_75t_L g596 ( .A(n_525), .B(n_575), .Y(n_596) );
INVx2_ASAP7_75t_L g597 ( .A(n_507), .Y(n_597) );
INVx1_ASAP7_75t_SL g598 ( .A(n_569), .Y(n_598) );
NOR2xp33_ASAP7_75t_L g599 ( .A(n_508), .B(n_463), .Y(n_599) );
INVxp67_ASAP7_75t_L g600 ( .A(n_545), .Y(n_600) );
AND2x2_ASAP7_75t_L g601 ( .A(n_534), .B(n_482), .Y(n_601) );
OR2x2_ASAP7_75t_L g602 ( .A(n_587), .B(n_464), .Y(n_602) );
NAND2xp5_ASAP7_75t_SL g603 ( .A(n_515), .B(n_489), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_527), .B(n_502), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_565), .Y(n_605) );
OAI21xp5_ASAP7_75t_L g606 ( .A1(n_586), .A2(n_502), .B(n_490), .Y(n_606) );
HB1xp67_ASAP7_75t_L g607 ( .A(n_537), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_567), .Y(n_608) );
NAND2x1p5_ASAP7_75t_L g609 ( .A(n_549), .B(n_439), .Y(n_609) );
NOR2xp33_ASAP7_75t_L g610 ( .A(n_509), .B(n_468), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_570), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_572), .Y(n_612) );
OR2x2_ASAP7_75t_L g613 ( .A(n_587), .B(n_479), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_530), .B(n_482), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_505), .Y(n_615) );
AND2x4_ASAP7_75t_L g616 ( .A(n_575), .B(n_481), .Y(n_616) );
INVx2_ASAP7_75t_L g617 ( .A(n_507), .Y(n_617) );
NOR2xp33_ASAP7_75t_L g618 ( .A(n_520), .B(n_492), .Y(n_618) );
INVx2_ASAP7_75t_L g619 ( .A(n_528), .Y(n_619) );
AND2x2_ASAP7_75t_L g620 ( .A(n_534), .B(n_483), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_506), .Y(n_621) );
INVxp33_ASAP7_75t_L g622 ( .A(n_555), .Y(n_622) );
INVx3_ASAP7_75t_L g623 ( .A(n_569), .Y(n_623) );
AND2x4_ASAP7_75t_L g624 ( .A(n_575), .B(n_481), .Y(n_624) );
AOI322xp5_ASAP7_75t_L g625 ( .A1(n_545), .A2(n_486), .A3(n_483), .B1(n_498), .B2(n_490), .C1(n_491), .C2(n_481), .Y(n_625) );
NOR2xp33_ASAP7_75t_L g626 ( .A(n_520), .B(n_16), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_582), .B(n_486), .Y(n_627) );
NAND2x1_ASAP7_75t_L g628 ( .A(n_528), .B(n_439), .Y(n_628) );
INVx2_ASAP7_75t_SL g629 ( .A(n_519), .Y(n_629) );
AND2x2_ASAP7_75t_L g630 ( .A(n_517), .B(n_438), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_583), .B(n_491), .Y(n_631) );
INVx2_ASAP7_75t_L g632 ( .A(n_537), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_573), .B(n_498), .Y(n_633) );
NAND2x1p5_ASAP7_75t_L g634 ( .A(n_552), .B(n_439), .Y(n_634) );
AND2x2_ASAP7_75t_L g635 ( .A(n_524), .B(n_438), .Y(n_635) );
NOR2xp33_ASAP7_75t_L g636 ( .A(n_590), .B(n_20), .Y(n_636) );
NOR2xp67_ASAP7_75t_L g637 ( .A(n_529), .B(n_438), .Y(n_637) );
INVx2_ASAP7_75t_L g638 ( .A(n_564), .Y(n_638) );
INVx2_ASAP7_75t_SL g639 ( .A(n_516), .Y(n_639) );
BUFx2_ASAP7_75t_L g640 ( .A(n_564), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_538), .B(n_469), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_585), .B(n_469), .Y(n_642) );
INVxp67_ASAP7_75t_L g643 ( .A(n_562), .Y(n_643) );
AND2x2_ASAP7_75t_L g644 ( .A(n_535), .B(n_481), .Y(n_644) );
AND2x2_ASAP7_75t_L g645 ( .A(n_535), .B(n_480), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_514), .Y(n_646) );
NAND2x1_ASAP7_75t_L g647 ( .A(n_579), .B(n_480), .Y(n_647) );
HB1xp67_ASAP7_75t_L g648 ( .A(n_513), .Y(n_648) );
AND2x2_ASAP7_75t_L g649 ( .A(n_544), .B(n_484), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_521), .Y(n_650) );
AND2x2_ASAP7_75t_L g651 ( .A(n_548), .B(n_484), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_531), .Y(n_652) );
AND2x2_ASAP7_75t_L g653 ( .A(n_539), .B(n_485), .Y(n_653) );
HB1xp67_ASAP7_75t_L g654 ( .A(n_513), .Y(n_654) );
AND2x2_ASAP7_75t_L g655 ( .A(n_510), .B(n_485), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_536), .Y(n_656) );
OR2x6_ASAP7_75t_L g657 ( .A(n_552), .B(n_493), .Y(n_657) );
INVx1_ASAP7_75t_SL g658 ( .A(n_559), .Y(n_658) );
INVx1_ASAP7_75t_L g659 ( .A(n_540), .Y(n_659) );
AND2x2_ASAP7_75t_L g660 ( .A(n_511), .B(n_487), .Y(n_660) );
AND2x4_ASAP7_75t_L g661 ( .A(n_579), .B(n_500), .Y(n_661) );
AND2x2_ASAP7_75t_L g662 ( .A(n_559), .B(n_487), .Y(n_662) );
INVx2_ASAP7_75t_L g663 ( .A(n_512), .Y(n_663) );
INVx2_ASAP7_75t_L g664 ( .A(n_512), .Y(n_664) );
AND2x4_ASAP7_75t_L g665 ( .A(n_579), .B(n_500), .Y(n_665) );
NOR2xp33_ASAP7_75t_L g666 ( .A(n_578), .B(n_20), .Y(n_666) );
AOI32xp33_ASAP7_75t_SL g667 ( .A1(n_578), .A2(n_494), .A3(n_488), .B1(n_23), .B2(n_24), .Y(n_667) );
INVx2_ASAP7_75t_L g668 ( .A(n_518), .Y(n_668) );
CKINVDCx16_ASAP7_75t_R g669 ( .A(n_594), .Y(n_669) );
AOI21xp5_ASAP7_75t_L g670 ( .A1(n_529), .A2(n_497), .B(n_496), .Y(n_670) );
AND2x2_ASAP7_75t_L g671 ( .A(n_532), .B(n_488), .Y(n_671) );
AND2x2_ASAP7_75t_L g672 ( .A(n_533), .B(n_494), .Y(n_672) );
OAI21xp5_ASAP7_75t_L g673 ( .A1(n_542), .A2(n_497), .B(n_496), .Y(n_673) );
OR2x2_ASAP7_75t_L g674 ( .A(n_541), .B(n_497), .Y(n_674) );
OR2x2_ASAP7_75t_L g675 ( .A(n_553), .B(n_496), .Y(n_675) );
OR2x2_ASAP7_75t_L g676 ( .A(n_546), .B(n_495), .Y(n_676) );
AND2x2_ASAP7_75t_L g677 ( .A(n_598), .B(n_566), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_625), .B(n_571), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_604), .B(n_584), .Y(n_679) );
AOI33xp33_ASAP7_75t_L g680 ( .A1(n_598), .A2(n_542), .A3(n_591), .B1(n_580), .B2(n_560), .B3(n_568), .Y(n_680) );
A2O1A1Ixp33_ASAP7_75t_L g681 ( .A1(n_622), .A2(n_558), .B(n_557), .C(n_580), .Y(n_681) );
NOR2xp33_ASAP7_75t_L g682 ( .A(n_600), .B(n_522), .Y(n_682) );
INVx2_ASAP7_75t_SL g683 ( .A(n_629), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_600), .B(n_591), .Y(n_684) );
AOI22xp5_ASAP7_75t_L g685 ( .A1(n_626), .A2(n_580), .B1(n_551), .B2(n_547), .Y(n_685) );
INVx1_ASAP7_75t_L g686 ( .A(n_648), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_648), .B(n_577), .Y(n_687) );
INVx2_ASAP7_75t_L g688 ( .A(n_640), .Y(n_688) );
INVx1_ASAP7_75t_L g689 ( .A(n_654), .Y(n_689) );
AOI322xp5_ASAP7_75t_L g690 ( .A1(n_669), .A2(n_592), .A3(n_554), .B1(n_589), .B2(n_588), .C1(n_581), .C2(n_576), .Y(n_690) );
INVx1_ASAP7_75t_L g691 ( .A(n_654), .Y(n_691) );
INVx1_ASAP7_75t_L g692 ( .A(n_607), .Y(n_692) );
OAI222xp33_ASAP7_75t_L g693 ( .A1(n_643), .A2(n_556), .B1(n_561), .B2(n_588), .C1(n_581), .C2(n_576), .Y(n_693) );
NOR2xp33_ASAP7_75t_L g694 ( .A(n_618), .B(n_593), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_604), .B(n_593), .Y(n_695) );
AND2x2_ASAP7_75t_L g696 ( .A(n_644), .B(n_589), .Y(n_696) );
HB1xp67_ASAP7_75t_L g697 ( .A(n_607), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_614), .B(n_574), .Y(n_698) );
INVx1_ASAP7_75t_L g699 ( .A(n_641), .Y(n_699) );
INVx1_ASAP7_75t_L g700 ( .A(n_641), .Y(n_700) );
OAI22xp33_ASAP7_75t_L g701 ( .A1(n_623), .A2(n_574), .B1(n_563), .B2(n_554), .Y(n_701) );
AOI21xp33_ASAP7_75t_L g702 ( .A1(n_636), .A2(n_563), .B(n_550), .Y(n_702) );
INVx1_ASAP7_75t_L g703 ( .A(n_605), .Y(n_703) );
O2A1O1Ixp33_ASAP7_75t_L g704 ( .A1(n_643), .A2(n_550), .B(n_543), .C(n_523), .Y(n_704) );
INVx1_ASAP7_75t_L g705 ( .A(n_608), .Y(n_705) );
OAI22xp5_ASAP7_75t_L g706 ( .A1(n_623), .A2(n_543), .B1(n_523), .B2(n_518), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_642), .B(n_495), .Y(n_707) );
AND2x2_ASAP7_75t_L g708 ( .A(n_595), .B(n_495), .Y(n_708) );
AND2x2_ASAP7_75t_L g709 ( .A(n_601), .B(n_493), .Y(n_709) );
INVxp67_ASAP7_75t_L g710 ( .A(n_599), .Y(n_710) );
OAI32xp33_ASAP7_75t_L g711 ( .A1(n_658), .A2(n_493), .A3(n_477), .B1(n_473), .B2(n_313), .Y(n_711) );
INVx2_ASAP7_75t_SL g712 ( .A(n_635), .Y(n_712) );
AOI221xp5_ASAP7_75t_L g713 ( .A1(n_666), .A2(n_477), .B1(n_473), .B2(n_313), .C(n_26), .Y(n_713) );
OR4x1_ASAP7_75t_L g714 ( .A(n_647), .B(n_477), .C(n_22), .D(n_25), .Y(n_714) );
AOI22xp5_ASAP7_75t_L g715 ( .A1(n_610), .A2(n_21), .B1(n_27), .B2(n_28), .Y(n_715) );
INVx1_ASAP7_75t_L g716 ( .A(n_611), .Y(n_716) );
INVx1_ASAP7_75t_L g717 ( .A(n_612), .Y(n_717) );
INVx1_ASAP7_75t_L g718 ( .A(n_615), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_614), .B(n_113), .Y(n_719) );
INVx1_ASAP7_75t_L g720 ( .A(n_621), .Y(n_720) );
INVx1_ASAP7_75t_L g721 ( .A(n_646), .Y(n_721) );
OR2x2_ASAP7_75t_L g722 ( .A(n_627), .B(n_29), .Y(n_722) );
AOI32xp33_ASAP7_75t_L g723 ( .A1(n_596), .A2(n_106), .A3(n_32), .B1(n_33), .B2(n_35), .Y(n_723) );
INVx1_ASAP7_75t_L g724 ( .A(n_650), .Y(n_724) );
INVx1_ASAP7_75t_L g725 ( .A(n_652), .Y(n_725) );
OAI221xp5_ASAP7_75t_L g726 ( .A1(n_673), .A2(n_30), .B1(n_37), .B2(n_40), .C(n_42), .Y(n_726) );
INVx1_ASAP7_75t_L g727 ( .A(n_656), .Y(n_727) );
INVx1_ASAP7_75t_L g728 ( .A(n_659), .Y(n_728) );
NOR2xp67_ASAP7_75t_L g729 ( .A(n_596), .B(n_43), .Y(n_729) );
INVx1_ASAP7_75t_L g730 ( .A(n_631), .Y(n_730) );
OAI22xp33_ASAP7_75t_L g731 ( .A1(n_678), .A2(n_637), .B1(n_628), .B2(n_603), .Y(n_731) );
AOI21xp5_ASAP7_75t_SL g732 ( .A1(n_681), .A2(n_606), .B(n_673), .Y(n_732) );
OAI211xp5_ASAP7_75t_L g733 ( .A1(n_690), .A2(n_606), .B(n_658), .C(n_670), .Y(n_733) );
AOI321xp33_ASAP7_75t_L g734 ( .A1(n_678), .A2(n_665), .A3(n_661), .B1(n_670), .B2(n_624), .C(n_616), .Y(n_734) );
OAI22xp5_ASAP7_75t_L g735 ( .A1(n_683), .A2(n_616), .B1(n_624), .B2(n_639), .Y(n_735) );
AOI21xp5_ASAP7_75t_L g736 ( .A1(n_693), .A2(n_657), .B(n_642), .Y(n_736) );
AOI22xp5_ASAP7_75t_L g737 ( .A1(n_682), .A2(n_661), .B1(n_665), .B2(n_631), .Y(n_737) );
NAND3xp33_ASAP7_75t_L g738 ( .A(n_680), .B(n_638), .C(n_632), .Y(n_738) );
AOI22xp5_ASAP7_75t_L g739 ( .A1(n_685), .A2(n_633), .B1(n_671), .B2(n_672), .Y(n_739) );
INVx1_ASAP7_75t_L g740 ( .A(n_699), .Y(n_740) );
AOI21xp5_ASAP7_75t_L g741 ( .A1(n_704), .A2(n_657), .B(n_609), .Y(n_741) );
AOI22xp5_ASAP7_75t_L g742 ( .A1(n_710), .A2(n_633), .B1(n_645), .B2(n_627), .Y(n_742) );
AOI21xp5_ASAP7_75t_L g743 ( .A1(n_706), .A2(n_657), .B(n_609), .Y(n_743) );
OAI21xp5_ASAP7_75t_L g744 ( .A1(n_729), .A2(n_634), .B(n_667), .Y(n_744) );
AOI21xp33_ASAP7_75t_SL g745 ( .A1(n_723), .A2(n_634), .B(n_597), .Y(n_745) );
NAND2xp5_ASAP7_75t_L g746 ( .A(n_700), .B(n_660), .Y(n_746) );
AOI221xp5_ASAP7_75t_L g747 ( .A1(n_702), .A2(n_617), .B1(n_619), .B2(n_655), .C(n_653), .Y(n_747) );
OAI22xp5_ASAP7_75t_L g748 ( .A1(n_712), .A2(n_602), .B1(n_613), .B2(n_620), .Y(n_748) );
NAND2xp5_ASAP7_75t_L g749 ( .A(n_730), .B(n_649), .Y(n_749) );
AOI211x1_ASAP7_75t_L g750 ( .A1(n_702), .A2(n_630), .B(n_651), .C(n_662), .Y(n_750) );
AOI21xp5_ASAP7_75t_L g751 ( .A1(n_706), .A2(n_675), .B(n_674), .Y(n_751) );
AOI22xp5_ASAP7_75t_L g752 ( .A1(n_694), .A2(n_676), .B1(n_668), .B2(n_664), .Y(n_752) );
OAI221xp5_ASAP7_75t_L g753 ( .A1(n_684), .A2(n_663), .B1(n_54), .B2(n_55), .C(n_57), .Y(n_753) );
AOI221xp5_ASAP7_75t_SL g754 ( .A1(n_701), .A2(n_44), .B1(n_61), .B2(n_66), .C(n_67), .Y(n_754) );
INVx1_ASAP7_75t_L g755 ( .A(n_686), .Y(n_755) );
AOI21xp5_ASAP7_75t_L g756 ( .A1(n_707), .A2(n_69), .B(n_70), .Y(n_756) );
INVx2_ASAP7_75t_L g757 ( .A(n_697), .Y(n_757) );
INVx1_ASAP7_75t_L g758 ( .A(n_689), .Y(n_758) );
OAI21xp5_ASAP7_75t_SL g759 ( .A1(n_713), .A2(n_71), .B(n_72), .Y(n_759) );
OA22x2_ASAP7_75t_L g760 ( .A1(n_677), .A2(n_73), .B1(n_74), .B2(n_75), .Y(n_760) );
AOI221xp5_ASAP7_75t_L g761 ( .A1(n_711), .A2(n_77), .B1(n_78), .B2(n_82), .C(n_83), .Y(n_761) );
A2O1A1Ixp33_ASAP7_75t_L g762 ( .A1(n_734), .A2(n_688), .B(n_679), .C(n_687), .Y(n_762) );
OAI221xp5_ASAP7_75t_L g763 ( .A1(n_732), .A2(n_691), .B1(n_692), .B2(n_728), .C(n_725), .Y(n_763) );
NOR2xp33_ASAP7_75t_L g764 ( .A(n_735), .B(n_679), .Y(n_764) );
NAND2xp5_ASAP7_75t_L g765 ( .A(n_740), .B(n_703), .Y(n_765) );
AOI21xp5_ASAP7_75t_L g766 ( .A1(n_741), .A2(n_707), .B(n_698), .Y(n_766) );
AOI22xp5_ASAP7_75t_L g767 ( .A1(n_731), .A2(n_727), .B1(n_724), .B2(n_721), .Y(n_767) );
NAND3xp33_ASAP7_75t_L g768 ( .A(n_733), .B(n_719), .C(n_722), .Y(n_768) );
NAND3xp33_ASAP7_75t_L g769 ( .A(n_750), .B(n_726), .C(n_720), .Y(n_769) );
NOR3xp33_ASAP7_75t_SL g770 ( .A(n_759), .B(n_714), .C(n_695), .Y(n_770) );
AOI21xp5_ASAP7_75t_L g771 ( .A1(n_743), .A2(n_718), .B(n_717), .Y(n_771) );
OAI32xp33_ASAP7_75t_L g772 ( .A1(n_738), .A2(n_716), .A3(n_705), .B1(n_709), .B2(n_696), .Y(n_772) );
NOR2x1_ASAP7_75t_L g773 ( .A(n_744), .B(n_708), .Y(n_773) );
NAND2xp5_ASAP7_75t_L g774 ( .A(n_742), .B(n_715), .Y(n_774) );
NOR2xp33_ASAP7_75t_SL g775 ( .A(n_753), .B(n_84), .Y(n_775) );
O2A1O1Ixp33_ASAP7_75t_L g776 ( .A1(n_745), .A2(n_86), .B(n_89), .C(n_92), .Y(n_776) );
O2A1O1Ixp33_ASAP7_75t_L g777 ( .A1(n_759), .A2(n_93), .B(n_94), .C(n_95), .Y(n_777) );
NAND2xp5_ASAP7_75t_L g778 ( .A(n_764), .B(n_747), .Y(n_778) );
AOI21xp5_ASAP7_75t_L g779 ( .A1(n_776), .A2(n_736), .B(n_760), .Y(n_779) );
NAND2xp5_ASAP7_75t_SL g780 ( .A(n_771), .B(n_754), .Y(n_780) );
XNOR2x1_ASAP7_75t_L g781 ( .A(n_773), .B(n_737), .Y(n_781) );
INVx2_ASAP7_75t_L g782 ( .A(n_765), .Y(n_782) );
NOR2xp33_ASAP7_75t_L g783 ( .A(n_763), .B(n_757), .Y(n_783) );
AOI211x1_ASAP7_75t_L g784 ( .A1(n_772), .A2(n_751), .B(n_748), .C(n_758), .Y(n_784) );
NOR2x1_ASAP7_75t_L g785 ( .A(n_777), .B(n_756), .Y(n_785) );
NAND4xp75_ASAP7_75t_L g786 ( .A(n_784), .B(n_767), .C(n_770), .D(n_774), .Y(n_786) );
NOR3xp33_ASAP7_75t_L g787 ( .A(n_780), .B(n_769), .C(n_768), .Y(n_787) );
HB1xp67_ASAP7_75t_L g788 ( .A(n_782), .Y(n_788) );
NOR3xp33_ASAP7_75t_L g789 ( .A(n_785), .B(n_762), .C(n_761), .Y(n_789) );
INVx1_ASAP7_75t_L g790 ( .A(n_778), .Y(n_790) );
NAND2x1p5_ASAP7_75t_L g791 ( .A(n_790), .B(n_779), .Y(n_791) );
NOR3xp33_ASAP7_75t_L g792 ( .A(n_786), .B(n_783), .C(n_766), .Y(n_792) );
INVx2_ASAP7_75t_L g793 ( .A(n_788), .Y(n_793) );
XOR2x2_ASAP7_75t_L g794 ( .A(n_791), .B(n_787), .Y(n_794) );
OAI22xp5_ASAP7_75t_SL g795 ( .A1(n_793), .A2(n_789), .B1(n_781), .B2(n_739), .Y(n_795) );
INVx1_ASAP7_75t_L g796 ( .A(n_794), .Y(n_796) );
INVx2_ASAP7_75t_L g797 ( .A(n_795), .Y(n_797) );
NAND2xp5_ASAP7_75t_SL g798 ( .A(n_797), .B(n_792), .Y(n_798) );
OAI22xp5_ASAP7_75t_L g799 ( .A1(n_796), .A2(n_755), .B1(n_752), .B2(n_749), .Y(n_799) );
NAND2xp5_ASAP7_75t_L g800 ( .A(n_798), .B(n_775), .Y(n_800) );
INVx1_ASAP7_75t_L g801 ( .A(n_799), .Y(n_801) );
AOI22xp5_ASAP7_75t_L g802 ( .A1(n_801), .A2(n_800), .B1(n_746), .B2(n_99), .Y(n_802) );
AOI22xp5_ASAP7_75t_L g803 ( .A1(n_802), .A2(n_96), .B1(n_98), .B2(n_100), .Y(n_803) );
OR2x6_ASAP7_75t_L g804 ( .A(n_803), .B(n_101), .Y(n_804) );
AOI21xp5_ASAP7_75t_L g805 ( .A1(n_804), .A2(n_102), .B(n_103), .Y(n_805) );
endmodule