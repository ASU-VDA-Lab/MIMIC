module fake_netlist_5_2545_n_1998 (n_137, n_210, n_168, n_164, n_191, n_91, n_208, n_82, n_122, n_194, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_65, n_78, n_74, n_144, n_207, n_114, n_57, n_96, n_37, n_189, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_197, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_195, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_203, n_205, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_202, n_130, n_157, n_29, n_79, n_193, n_131, n_151, n_47, n_173, n_192, n_25, n_53, n_160, n_198, n_188, n_190, n_8, n_201, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_55, n_196, n_99, n_2, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_200, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_209, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_199, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_206, n_171, n_153, n_7, n_15, n_145, n_48, n_204, n_50, n_52, n_88, n_110, n_1998);

input n_137;
input n_210;
input n_168;
input n_164;
input n_191;
input n_91;
input n_208;
input n_82;
input n_122;
input n_194;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_65;
input n_78;
input n_74;
input n_144;
input n_207;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_197;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_195;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_203;
input n_205;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_202;
input n_130;
input n_157;
input n_29;
input n_79;
input n_193;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_25;
input n_53;
input n_160;
input n_198;
input n_188;
input n_190;
input n_8;
input n_201;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_196;
input n_99;
input n_2;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_200;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_209;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_199;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_206;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_204;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1998;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_1021;
wire n_1960;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1947;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_1580;
wire n_674;
wire n_417;
wire n_1939;
wire n_1806;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1860;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_1896;
wire n_929;
wire n_1124;
wire n_1818;
wire n_902;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_1845;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_1949;
wire n_343;
wire n_1449;
wire n_308;
wire n_1946;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_1948;
wire n_1984;
wire n_264;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_339;
wire n_1146;
wire n_882;
wire n_243;
wire n_1097;
wire n_1036;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_580;
wire n_290;
wire n_1040;
wire n_1872;
wire n_1852;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_1931;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1880;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_446;
wire n_1863;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1986;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1971;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_1950;
wire n_907;
wire n_1447;
wire n_1377;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1926;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_1819;
wire n_476;
wire n_1527;
wire n_534;
wire n_1882;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_561;
wire n_1319;
wire n_1825;
wire n_1951;
wire n_1883;
wire n_1906;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_352;
wire n_1884;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1891;
wire n_1481;
wire n_1942;
wire n_434;
wire n_1978;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_1810;
wire n_1888;
wire n_759;
wire n_1892;
wire n_806;
wire n_1997;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1963;
wire n_1571;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_1925;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1798;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_1916;
wire n_293;
wire n_677;
wire n_372;
wire n_244;
wire n_1333;
wire n_1121;
wire n_433;
wire n_604;
wire n_314;
wire n_368;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_624;
wire n_252;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1994;
wire n_1231;
wire n_739;
wire n_1406;
wire n_1279;
wire n_1195;
wire n_1837;
wire n_1839;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_1832;
wire n_259;
wire n_448;
wire n_1851;
wire n_758;
wire n_999;
wire n_1933;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_1874;
wire n_563;
wire n_1987;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_1964;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1923;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_1989;
wire n_396;
wire n_1887;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1959;
wire n_1758;
wire n_1574;
wire n_473;
wire n_1921;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_1820;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_1870;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1980;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1927;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_1965;
wire n_239;
wire n_630;
wire n_1902;
wire n_1941;
wire n_1913;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1875;
wire n_1982;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_261;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_1849;
wire n_729;
wire n_1131;
wire n_1084;
wire n_1961;
wire n_970;
wire n_1935;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_1821;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_1893;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_1958;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1954;
wire n_1608;
wire n_983;
wire n_1844;
wire n_280;
wire n_1305;
wire n_873;
wire n_1826;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_1974;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1966;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_1953;
wire n_1938;
wire n_820;
wire n_1200;
wire n_1911;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_1967;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_1932;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1992;
wire n_1643;
wire n_883;
wire n_1983;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1400;
wire n_1342;
wire n_900;
wire n_856;
wire n_1793;
wire n_1976;
wire n_918;
wire n_942;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1977;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1735;
wire n_1697;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_1881;
wire n_988;
wire n_1940;
wire n_814;
wire n_1549;
wire n_1934;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1824;
wire n_1917;
wire n_1219;
wire n_1204;
wire n_1814;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1848;
wire n_1928;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_584;
wire n_336;
wire n_681;
wire n_1638;
wire n_1786;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1895;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1929;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_1968;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_1970;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_1737;
wire n_1904;
wire n_1993;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1957;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_1899;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1835;
wire n_1440;
wire n_421;
wire n_1988;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_232;
wire n_1915;
wire n_1109;
wire n_895;
wire n_1310;
wire n_1803;
wire n_427;
wire n_1399;
wire n_1543;
wire n_1991;
wire n_1979;
wire n_791;
wire n_732;
wire n_1533;
wire n_808;
wire n_797;
wire n_1025;
wire n_1930;
wire n_1955;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1972;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_1855;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_1985;
wire n_1898;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_1890;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1944;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_1981;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1952;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1922;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_1867;
wire n_1945;
wire n_481;
wire n_1675;
wire n_1924;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_1995;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_1813;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_428;
wire n_379;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_1973;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_1873;
wire n_1411;
wire n_221;
wire n_622;
wire n_1962;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_1842;
wire n_871;
wire n_598;
wire n_685;
wire n_928;
wire n_608;
wire n_1367;
wire n_1943;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1858;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_384;
wire n_1404;
wire n_1794;
wire n_1315;
wire n_277;
wire n_1061;
wire n_1910;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_844;
wire n_471;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_1975;
wire n_273;
wire n_1937;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_1914;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_1936;
wire n_1956;
wire n_437;
wire n_1642;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_1918;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_1879;
wire n_597;
wire n_1996;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1969;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_1089;
wire n_927;
wire n_1990;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_202),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_130),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_175),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_88),
.Y(n_214)
);

HB1xp67_ASAP7_75t_L g215 ( 
.A(n_132),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_65),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_210),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_181),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_122),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_188),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_42),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_92),
.Y(n_222)
);

INVx1_ASAP7_75t_SL g223 ( 
.A(n_86),
.Y(n_223)
);

BUFx10_ASAP7_75t_L g224 ( 
.A(n_100),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_136),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_15),
.Y(n_226)
);

BUFx10_ASAP7_75t_L g227 ( 
.A(n_145),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_140),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_4),
.Y(n_229)
);

HB1xp67_ASAP7_75t_L g230 ( 
.A(n_38),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_190),
.Y(n_231)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_90),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_38),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_79),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_9),
.Y(n_235)
);

BUFx3_ASAP7_75t_L g236 ( 
.A(n_7),
.Y(n_236)
);

INVx2_ASAP7_75t_SL g237 ( 
.A(n_117),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_115),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_32),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_71),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_157),
.Y(n_241)
);

BUFx2_ASAP7_75t_SL g242 ( 
.A(n_147),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_83),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_2),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_124),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_168),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_13),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_180),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_81),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_131),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_151),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_114),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_158),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_8),
.Y(n_254)
);

CKINVDCx16_ASAP7_75t_R g255 ( 
.A(n_142),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_120),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_7),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_155),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_194),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_118),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_126),
.Y(n_261)
);

BUFx3_ASAP7_75t_L g262 ( 
.A(n_0),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_112),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_85),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_108),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_143),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_80),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_148),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_39),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_22),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_17),
.Y(n_271)
);

CKINVDCx16_ASAP7_75t_R g272 ( 
.A(n_27),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_75),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_14),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_149),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_36),
.Y(n_276)
);

BUFx3_ASAP7_75t_L g277 ( 
.A(n_2),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_102),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_141),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_97),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_94),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_199),
.Y(n_282)
);

BUFx10_ASAP7_75t_L g283 ( 
.A(n_89),
.Y(n_283)
);

BUFx6f_ASAP7_75t_L g284 ( 
.A(n_183),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_54),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_26),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_134),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_163),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_139),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_95),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_44),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_176),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_64),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_70),
.Y(n_294)
);

BUFx6f_ASAP7_75t_L g295 ( 
.A(n_61),
.Y(n_295)
);

INVx2_ASAP7_75t_SL g296 ( 
.A(n_186),
.Y(n_296)
);

INVx1_ASAP7_75t_SL g297 ( 
.A(n_192),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_125),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_57),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_51),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_0),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_32),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_121),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_93),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_154),
.Y(n_305)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_128),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_169),
.Y(n_307)
);

INVx2_ASAP7_75t_SL g308 ( 
.A(n_104),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_144),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_113),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_166),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_61),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_28),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_161),
.Y(n_314)
);

BUFx8_ASAP7_75t_SL g315 ( 
.A(n_31),
.Y(n_315)
);

INVx1_ASAP7_75t_SL g316 ( 
.A(n_96),
.Y(n_316)
);

INVx1_ASAP7_75t_SL g317 ( 
.A(n_12),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_82),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_174),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_135),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_23),
.Y(n_321)
);

BUFx6f_ASAP7_75t_L g322 ( 
.A(n_162),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_184),
.Y(n_323)
);

INVx1_ASAP7_75t_SL g324 ( 
.A(n_153),
.Y(n_324)
);

CKINVDCx16_ASAP7_75t_R g325 ( 
.A(n_110),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_12),
.Y(n_326)
);

BUFx5_ASAP7_75t_L g327 ( 
.A(n_106),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_98),
.Y(n_328)
);

INVx2_ASAP7_75t_SL g329 ( 
.A(n_57),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_50),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_193),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_49),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_44),
.Y(n_333)
);

INVx1_ASAP7_75t_SL g334 ( 
.A(n_8),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_127),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_189),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_209),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_66),
.Y(n_338)
);

INVx1_ASAP7_75t_SL g339 ( 
.A(n_206),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_19),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_195),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_21),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_63),
.Y(n_343)
);

BUFx3_ASAP7_75t_L g344 ( 
.A(n_22),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_107),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_63),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_196),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_200),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_146),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_198),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_40),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_156),
.Y(n_352)
);

INVx1_ASAP7_75t_SL g353 ( 
.A(n_170),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_203),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_46),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_28),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_103),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_201),
.Y(n_358)
);

INVxp67_ASAP7_75t_L g359 ( 
.A(n_51),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_187),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_5),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_197),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_4),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_205),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_84),
.Y(n_365)
);

BUFx10_ASAP7_75t_L g366 ( 
.A(n_171),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_159),
.Y(n_367)
);

BUFx10_ASAP7_75t_L g368 ( 
.A(n_152),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_1),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_101),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_178),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_59),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_16),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_9),
.Y(n_374)
);

CKINVDCx6p67_ASAP7_75t_R g375 ( 
.A(n_160),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_55),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_177),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_47),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_150),
.Y(n_379)
);

BUFx3_ASAP7_75t_L g380 ( 
.A(n_40),
.Y(n_380)
);

INVx2_ASAP7_75t_SL g381 ( 
.A(n_49),
.Y(n_381)
);

INVx1_ASAP7_75t_SL g382 ( 
.A(n_207),
.Y(n_382)
);

BUFx3_ASAP7_75t_L g383 ( 
.A(n_27),
.Y(n_383)
);

BUFx2_ASAP7_75t_L g384 ( 
.A(n_47),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_55),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_58),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_72),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_179),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_182),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_25),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_33),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_1),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_53),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_3),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_25),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_164),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_34),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_56),
.Y(n_398)
);

BUFx3_ASAP7_75t_L g399 ( 
.A(n_69),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_31),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_34),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_23),
.Y(n_402)
);

BUFx3_ASAP7_75t_L g403 ( 
.A(n_204),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_48),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_109),
.Y(n_405)
);

BUFx2_ASAP7_75t_L g406 ( 
.A(n_13),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_67),
.Y(n_407)
);

BUFx3_ASAP7_75t_L g408 ( 
.A(n_21),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_129),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_111),
.Y(n_410)
);

BUFx3_ASAP7_75t_L g411 ( 
.A(n_35),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_185),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_17),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_20),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_133),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_64),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_68),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_236),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_212),
.Y(n_419)
);

AND2x2_ASAP7_75t_L g420 ( 
.A(n_384),
.B(n_3),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_236),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_217),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_315),
.Y(n_423)
);

INVxp67_ASAP7_75t_L g424 ( 
.A(n_406),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_229),
.B(n_5),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_262),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_262),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_277),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_253),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_272),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_292),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_257),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_305),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_295),
.Y(n_434)
);

INVxp33_ASAP7_75t_SL g435 ( 
.A(n_230),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_269),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_270),
.Y(n_437)
);

INVxp67_ASAP7_75t_SL g438 ( 
.A(n_215),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_295),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_271),
.Y(n_440)
);

NOR2xp67_ASAP7_75t_L g441 ( 
.A(n_359),
.B(n_6),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_274),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_286),
.Y(n_443)
);

INVxp67_ASAP7_75t_L g444 ( 
.A(n_276),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_348),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_412),
.Y(n_446)
);

INVxp67_ASAP7_75t_SL g447 ( 
.A(n_399),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_291),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_295),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_299),
.Y(n_450)
);

INVxp33_ASAP7_75t_L g451 ( 
.A(n_285),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_295),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_277),
.Y(n_453)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_255),
.Y(n_454)
);

INVxp67_ASAP7_75t_SL g455 ( 
.A(n_399),
.Y(n_455)
);

HB1xp67_ASAP7_75t_L g456 ( 
.A(n_221),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_344),
.Y(n_457)
);

INVxp67_ASAP7_75t_L g458 ( 
.A(n_293),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_344),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_380),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_295),
.Y(n_461)
);

INVxp33_ASAP7_75t_SL g462 ( 
.A(n_221),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_237),
.B(n_6),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_380),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_383),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_383),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_408),
.Y(n_467)
);

INVxp67_ASAP7_75t_SL g468 ( 
.A(n_403),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_408),
.Y(n_469)
);

HB1xp67_ASAP7_75t_L g470 ( 
.A(n_226),
.Y(n_470)
);

CKINVDCx20_ASAP7_75t_R g471 ( 
.A(n_325),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_392),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_300),
.Y(n_473)
);

BUFx2_ASAP7_75t_L g474 ( 
.A(n_411),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_301),
.Y(n_475)
);

INVxp67_ASAP7_75t_SL g476 ( 
.A(n_403),
.Y(n_476)
);

CKINVDCx20_ASAP7_75t_R g477 ( 
.A(n_258),
.Y(n_477)
);

INVxp67_ASAP7_75t_SL g478 ( 
.A(n_411),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_302),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_343),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_346),
.Y(n_481)
);

HB1xp67_ASAP7_75t_L g482 ( 
.A(n_226),
.Y(n_482)
);

NAND2xp33_ASAP7_75t_R g483 ( 
.A(n_211),
.B(n_10),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_237),
.B(n_10),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_296),
.B(n_11),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_313),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_321),
.Y(n_487)
);

CKINVDCx20_ASAP7_75t_R g488 ( 
.A(n_259),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_326),
.Y(n_489)
);

CKINVDCx20_ASAP7_75t_R g490 ( 
.A(n_260),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_296),
.B(n_11),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_330),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_308),
.B(n_14),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_308),
.B(n_219),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_351),
.Y(n_495)
);

INVxp33_ASAP7_75t_SL g496 ( 
.A(n_233),
.Y(n_496)
);

INVx1_ASAP7_75t_SL g497 ( 
.A(n_244),
.Y(n_497)
);

HB1xp67_ASAP7_75t_L g498 ( 
.A(n_233),
.Y(n_498)
);

CKINVDCx16_ASAP7_75t_R g499 ( 
.A(n_224),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_392),
.Y(n_500)
);

CKINVDCx16_ASAP7_75t_R g501 ( 
.A(n_224),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_393),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_356),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_393),
.Y(n_504)
);

INVxp33_ASAP7_75t_L g505 ( 
.A(n_361),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_332),
.Y(n_506)
);

CKINVDCx16_ASAP7_75t_R g507 ( 
.A(n_224),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_219),
.B(n_15),
.Y(n_508)
);

INVxp67_ASAP7_75t_SL g509 ( 
.A(n_216),
.Y(n_509)
);

INVxp33_ASAP7_75t_SL g510 ( 
.A(n_235),
.Y(n_510)
);

NAND2xp33_ASAP7_75t_R g511 ( 
.A(n_211),
.B(n_16),
.Y(n_511)
);

CKINVDCx16_ASAP7_75t_R g512 ( 
.A(n_227),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_333),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_363),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_369),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_395),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_400),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_401),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_402),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_404),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_329),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_329),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_381),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_381),
.Y(n_524)
);

CKINVDCx20_ASAP7_75t_R g525 ( 
.A(n_261),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_SL g526 ( 
.A(n_499),
.B(n_227),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_447),
.B(n_232),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_455),
.B(n_232),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_434),
.Y(n_529)
);

NOR2xp67_ASAP7_75t_L g530 ( 
.A(n_432),
.B(n_220),
.Y(n_530)
);

XOR2x2_ASAP7_75t_SL g531 ( 
.A(n_463),
.B(n_247),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_461),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_477),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_434),
.Y(n_534)
);

AND2x6_ASAP7_75t_L g535 ( 
.A(n_420),
.B(n_213),
.Y(n_535)
);

CKINVDCx11_ASAP7_75t_R g536 ( 
.A(n_419),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_461),
.Y(n_537)
);

CKINVDCx20_ASAP7_75t_R g538 ( 
.A(n_422),
.Y(n_538)
);

AND2x2_ASAP7_75t_L g539 ( 
.A(n_478),
.B(n_227),
.Y(n_539)
);

AND2x2_ASAP7_75t_L g540 ( 
.A(n_468),
.B(n_283),
.Y(n_540)
);

INVx3_ASAP7_75t_L g541 ( 
.A(n_439),
.Y(n_541)
);

INVx4_ASAP7_75t_L g542 ( 
.A(n_432),
.Y(n_542)
);

BUFx8_ASAP7_75t_L g543 ( 
.A(n_420),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_439),
.Y(n_544)
);

BUFx6f_ASAP7_75t_L g545 ( 
.A(n_449),
.Y(n_545)
);

AND2x2_ASAP7_75t_L g546 ( 
.A(n_476),
.B(n_283),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_449),
.Y(n_547)
);

CKINVDCx20_ASAP7_75t_R g548 ( 
.A(n_429),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_452),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_488),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_490),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_452),
.Y(n_552)
);

BUFx6f_ASAP7_75t_L g553 ( 
.A(n_472),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_519),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_480),
.Y(n_555)
);

AND2x2_ASAP7_75t_L g556 ( 
.A(n_418),
.B(n_283),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_525),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_481),
.Y(n_558)
);

BUFx2_ASAP7_75t_L g559 ( 
.A(n_430),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_454),
.Y(n_560)
);

BUFx2_ASAP7_75t_L g561 ( 
.A(n_430),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_495),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_472),
.Y(n_563)
);

BUFx8_ASAP7_75t_L g564 ( 
.A(n_474),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_R g565 ( 
.A(n_436),
.B(n_263),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_471),
.Y(n_566)
);

CKINVDCx20_ASAP7_75t_R g567 ( 
.A(n_431),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_500),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_433),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_519),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_503),
.Y(n_571)
);

BUFx6f_ASAP7_75t_L g572 ( 
.A(n_500),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_445),
.Y(n_573)
);

BUFx6f_ASAP7_75t_L g574 ( 
.A(n_502),
.Y(n_574)
);

CKINVDCx20_ASAP7_75t_R g575 ( 
.A(n_446),
.Y(n_575)
);

BUFx6f_ASAP7_75t_L g576 ( 
.A(n_502),
.Y(n_576)
);

CKINVDCx20_ASAP7_75t_R g577 ( 
.A(n_497),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_514),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_504),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_520),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_509),
.B(n_240),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_504),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_520),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_R g584 ( 
.A(n_436),
.B(n_264),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_515),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_516),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_517),
.Y(n_587)
);

OR2x2_ASAP7_75t_L g588 ( 
.A(n_474),
.B(n_317),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_518),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_521),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_521),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_423),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_423),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_522),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_421),
.Y(n_595)
);

NOR2xp33_ASAP7_75t_L g596 ( 
.A(n_462),
.B(n_223),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_522),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_426),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_437),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_427),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_523),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_437),
.Y(n_602)
);

NAND2xp33_ASAP7_75t_L g603 ( 
.A(n_440),
.B(n_235),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_438),
.B(n_494),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_440),
.Y(n_605)
);

BUFx6f_ASAP7_75t_L g606 ( 
.A(n_485),
.Y(n_606)
);

NOR2xp67_ASAP7_75t_L g607 ( 
.A(n_442),
.B(n_225),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_442),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_428),
.Y(n_609)
);

CKINVDCx20_ASAP7_75t_R g610 ( 
.A(n_501),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_453),
.Y(n_611)
);

AOI22xp33_ASAP7_75t_L g612 ( 
.A1(n_606),
.A2(n_508),
.B1(n_491),
.B2(n_493),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_532),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_606),
.B(n_484),
.Y(n_614)
);

BUFx2_ASAP7_75t_L g615 ( 
.A(n_577),
.Y(n_615)
);

AND2x2_ASAP7_75t_L g616 ( 
.A(n_540),
.B(n_457),
.Y(n_616)
);

INVx4_ASAP7_75t_L g617 ( 
.A(n_545),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_606),
.B(n_443),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_537),
.Y(n_619)
);

BUFx6f_ASAP7_75t_L g620 ( 
.A(n_545),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_537),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_598),
.Y(n_622)
);

AND2x4_ASAP7_75t_L g623 ( 
.A(n_606),
.B(n_459),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_SL g624 ( 
.A(n_606),
.B(n_240),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_552),
.Y(n_625)
);

AOI22xp33_ASAP7_75t_L g626 ( 
.A1(n_581),
.A2(n_435),
.B1(n_424),
.B2(n_496),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_552),
.Y(n_627)
);

AND2x2_ASAP7_75t_SL g628 ( 
.A(n_596),
.B(n_256),
.Y(n_628)
);

BUFx3_ASAP7_75t_L g629 ( 
.A(n_600),
.Y(n_629)
);

INVx1_ASAP7_75t_SL g630 ( 
.A(n_588),
.Y(n_630)
);

AOI22xp33_ASAP7_75t_L g631 ( 
.A1(n_535),
.A2(n_510),
.B1(n_289),
.B2(n_306),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_SL g632 ( 
.A(n_530),
.B(n_256),
.Y(n_632)
);

INVx5_ASAP7_75t_L g633 ( 
.A(n_535),
.Y(n_633)
);

OR2x2_ASAP7_75t_L g634 ( 
.A(n_588),
.B(n_456),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_604),
.B(n_443),
.Y(n_635)
);

NOR2xp33_ASAP7_75t_L g636 ( 
.A(n_603),
.B(n_448),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_607),
.B(n_448),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_555),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_541),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_558),
.Y(n_640)
);

INVx6_ASAP7_75t_L g641 ( 
.A(n_564),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_541),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_562),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_571),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_SL g645 ( 
.A(n_531),
.B(n_289),
.Y(n_645)
);

NOR2xp33_ASAP7_75t_L g646 ( 
.A(n_542),
.B(n_450),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_578),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_SL g648 ( 
.A(n_531),
.B(n_306),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_595),
.Y(n_649)
);

INVx3_ASAP7_75t_L g650 ( 
.A(n_545),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_540),
.B(n_450),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_546),
.B(n_473),
.Y(n_652)
);

AND2x4_ASAP7_75t_L g653 ( 
.A(n_595),
.B(n_460),
.Y(n_653)
);

AND2x2_ASAP7_75t_L g654 ( 
.A(n_546),
.B(n_464),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_535),
.B(n_473),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_609),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_609),
.Y(n_657)
);

NOR2xp33_ASAP7_75t_L g658 ( 
.A(n_542),
.B(n_475),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_541),
.Y(n_659)
);

HB1xp67_ASAP7_75t_L g660 ( 
.A(n_539),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_611),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_611),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_585),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_SL g664 ( 
.A(n_542),
.B(n_539),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_535),
.B(n_475),
.Y(n_665)
);

OR2x2_ASAP7_75t_L g666 ( 
.A(n_527),
.B(n_470),
.Y(n_666)
);

INVx4_ASAP7_75t_L g667 ( 
.A(n_545),
.Y(n_667)
);

INVxp67_ASAP7_75t_SL g668 ( 
.A(n_545),
.Y(n_668)
);

NAND2xp33_ASAP7_75t_L g669 ( 
.A(n_535),
.B(n_213),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_SL g670 ( 
.A(n_528),
.B(n_362),
.Y(n_670)
);

AOI22xp33_ASAP7_75t_L g671 ( 
.A1(n_535),
.A2(n_362),
.B1(n_377),
.B2(n_441),
.Y(n_671)
);

INVx4_ASAP7_75t_L g672 ( 
.A(n_535),
.Y(n_672)
);

INVx5_ASAP7_75t_L g673 ( 
.A(n_553),
.Y(n_673)
);

INVx3_ASAP7_75t_L g674 ( 
.A(n_553),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_586),
.Y(n_675)
);

NAND3xp33_ASAP7_75t_L g676 ( 
.A(n_556),
.B(n_486),
.C(n_479),
.Y(n_676)
);

INVx6_ASAP7_75t_L g677 ( 
.A(n_564),
.Y(n_677)
);

NOR2xp33_ASAP7_75t_L g678 ( 
.A(n_526),
.B(n_479),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_586),
.Y(n_679)
);

OR2x6_ASAP7_75t_L g680 ( 
.A(n_556),
.B(n_242),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_544),
.Y(n_681)
);

NAND2xp33_ASAP7_75t_R g682 ( 
.A(n_599),
.B(n_486),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_589),
.Y(n_683)
);

INVx4_ASAP7_75t_SL g684 ( 
.A(n_553),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_529),
.B(n_487),
.Y(n_685)
);

OAI22xp33_ASAP7_75t_L g686 ( 
.A1(n_599),
.A2(n_512),
.B1(n_507),
.B2(n_483),
.Y(n_686)
);

OR2x2_ASAP7_75t_L g687 ( 
.A(n_559),
.B(n_482),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_544),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_534),
.B(n_487),
.Y(n_689)
);

BUFx4f_ASAP7_75t_L g690 ( 
.A(n_553),
.Y(n_690)
);

INVxp67_ASAP7_75t_L g691 ( 
.A(n_559),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_589),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_547),
.B(n_489),
.Y(n_693)
);

INVx3_ASAP7_75t_L g694 ( 
.A(n_553),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_547),
.Y(n_695)
);

AND2x6_ASAP7_75t_L g696 ( 
.A(n_554),
.B(n_377),
.Y(n_696)
);

AND2x2_ASAP7_75t_L g697 ( 
.A(n_554),
.B(n_465),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_570),
.Y(n_698)
);

BUFx10_ASAP7_75t_L g699 ( 
.A(n_592),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_SL g700 ( 
.A(n_565),
.B(n_213),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_SL g701 ( 
.A(n_584),
.B(n_213),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_570),
.Y(n_702)
);

AND2x2_ASAP7_75t_L g703 ( 
.A(n_580),
.B(n_466),
.Y(n_703)
);

INVx3_ASAP7_75t_L g704 ( 
.A(n_572),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_580),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_549),
.Y(n_706)
);

NOR2xp33_ASAP7_75t_L g707 ( 
.A(n_602),
.B(n_489),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_549),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_572),
.Y(n_709)
);

INVx5_ASAP7_75t_L g710 ( 
.A(n_572),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_572),
.B(n_492),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_583),
.Y(n_712)
);

AOI22xp33_ASAP7_75t_L g713 ( 
.A1(n_583),
.A2(n_498),
.B1(n_458),
.B2(n_444),
.Y(n_713)
);

INVx4_ASAP7_75t_L g714 ( 
.A(n_572),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_587),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_587),
.Y(n_716)
);

INVx5_ASAP7_75t_L g717 ( 
.A(n_574),
.Y(n_717)
);

OR2x2_ASAP7_75t_L g718 ( 
.A(n_561),
.B(n_492),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_574),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_590),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_SL g721 ( 
.A(n_543),
.B(n_213),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_574),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_SL g723 ( 
.A(n_543),
.B(n_284),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_590),
.Y(n_724)
);

NOR2xp33_ASAP7_75t_L g725 ( 
.A(n_602),
.B(n_506),
.Y(n_725)
);

INVx4_ASAP7_75t_L g726 ( 
.A(n_574),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_SL g727 ( 
.A(n_543),
.B(n_284),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_574),
.Y(n_728)
);

BUFx6f_ASAP7_75t_L g729 ( 
.A(n_576),
.Y(n_729)
);

INVx3_ASAP7_75t_L g730 ( 
.A(n_576),
.Y(n_730)
);

INVx1_ASAP7_75t_SL g731 ( 
.A(n_561),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_SL g732 ( 
.A(n_605),
.B(n_284),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_SL g733 ( 
.A(n_605),
.B(n_284),
.Y(n_733)
);

OR2x6_ASAP7_75t_L g734 ( 
.A(n_591),
.B(n_467),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_591),
.Y(n_735)
);

INVx3_ASAP7_75t_L g736 ( 
.A(n_576),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_594),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_594),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_597),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_576),
.Y(n_740)
);

BUFx3_ASAP7_75t_L g741 ( 
.A(n_576),
.Y(n_741)
);

NOR2xp33_ASAP7_75t_L g742 ( 
.A(n_608),
.B(n_506),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_597),
.Y(n_743)
);

AND2x4_ASAP7_75t_L g744 ( 
.A(n_601),
.B(n_469),
.Y(n_744)
);

AND2x2_ASAP7_75t_L g745 ( 
.A(n_563),
.B(n_568),
.Y(n_745)
);

NOR2xp33_ASAP7_75t_L g746 ( 
.A(n_608),
.B(n_513),
.Y(n_746)
);

BUFx3_ASAP7_75t_L g747 ( 
.A(n_601),
.Y(n_747)
);

NOR2xp33_ASAP7_75t_L g748 ( 
.A(n_563),
.B(n_513),
.Y(n_748)
);

BUFx10_ASAP7_75t_L g749 ( 
.A(n_592),
.Y(n_749)
);

INVx2_ASAP7_75t_SL g750 ( 
.A(n_564),
.Y(n_750)
);

AND2x2_ASAP7_75t_SL g751 ( 
.A(n_568),
.B(n_284),
.Y(n_751)
);

INVx4_ASAP7_75t_L g752 ( 
.A(n_579),
.Y(n_752)
);

BUFx8_ASAP7_75t_SL g753 ( 
.A(n_538),
.Y(n_753)
);

OAI21xp33_ASAP7_75t_SL g754 ( 
.A1(n_579),
.A2(n_524),
.B(n_523),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_582),
.Y(n_755)
);

NOR2xp33_ASAP7_75t_L g756 ( 
.A(n_582),
.B(n_451),
.Y(n_756)
);

INVxp67_ASAP7_75t_SL g757 ( 
.A(n_548),
.Y(n_757)
);

BUFx2_ASAP7_75t_L g758 ( 
.A(n_560),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_593),
.Y(n_759)
);

OR2x6_ASAP7_75t_L g760 ( 
.A(n_536),
.B(n_524),
.Y(n_760)
);

NOR2xp33_ASAP7_75t_L g761 ( 
.A(n_593),
.B(n_505),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_533),
.Y(n_762)
);

AOI22xp33_ASAP7_75t_L g763 ( 
.A1(n_628),
.A2(n_334),
.B1(n_397),
.B2(n_322),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_613),
.Y(n_764)
);

INVx8_ASAP7_75t_L g765 ( 
.A(n_680),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_SL g766 ( 
.A(n_628),
.B(n_322),
.Y(n_766)
);

OAI22xp5_ASAP7_75t_L g767 ( 
.A1(n_612),
.A2(n_382),
.B1(n_297),
.B2(n_316),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_614),
.B(n_246),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_649),
.Y(n_769)
);

AND2x2_ASAP7_75t_L g770 ( 
.A(n_630),
.B(n_533),
.Y(n_770)
);

BUFx3_ASAP7_75t_L g771 ( 
.A(n_623),
.Y(n_771)
);

OR2x2_ASAP7_75t_L g772 ( 
.A(n_634),
.B(n_560),
.Y(n_772)
);

NOR2xp67_ASAP7_75t_L g773 ( 
.A(n_676),
.B(n_550),
.Y(n_773)
);

AOI22xp33_ASAP7_75t_L g774 ( 
.A1(n_645),
.A2(n_322),
.B1(n_327),
.B2(n_417),
.Y(n_774)
);

BUFx6f_ASAP7_75t_L g775 ( 
.A(n_623),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_656),
.Y(n_776)
);

NOR2xp33_ASAP7_75t_SL g777 ( 
.A(n_641),
.B(n_550),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_623),
.B(n_248),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_618),
.B(n_249),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_SL g780 ( 
.A(n_633),
.B(n_322),
.Y(n_780)
);

NOR2xp67_ASAP7_75t_SL g781 ( 
.A(n_633),
.B(n_322),
.Y(n_781)
);

NOR2xp33_ASAP7_75t_L g782 ( 
.A(n_635),
.B(n_324),
.Y(n_782)
);

NOR2xp33_ASAP7_75t_L g783 ( 
.A(n_651),
.B(n_339),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_698),
.B(n_265),
.Y(n_784)
);

AND2x6_ASAP7_75t_L g785 ( 
.A(n_616),
.B(n_275),
.Y(n_785)
);

AOI22xp33_ASAP7_75t_L g786 ( 
.A1(n_645),
.A2(n_327),
.B1(n_338),
.B2(n_294),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_SL g787 ( 
.A(n_633),
.B(n_327),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_702),
.B(n_278),
.Y(n_788)
);

AOI22xp33_ASAP7_75t_L g789 ( 
.A1(n_648),
.A2(n_327),
.B1(n_303),
.B2(n_350),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_SL g790 ( 
.A(n_633),
.B(n_327),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_619),
.Y(n_791)
);

BUFx10_ASAP7_75t_L g792 ( 
.A(n_707),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_621),
.Y(n_793)
);

O2A1O1Ixp5_ASAP7_75t_L g794 ( 
.A1(n_624),
.A2(n_357),
.B(n_388),
.C(n_349),
.Y(n_794)
);

NOR2xp33_ASAP7_75t_L g795 ( 
.A(n_652),
.B(n_353),
.Y(n_795)
);

INVx1_ASAP7_75t_SL g796 ( 
.A(n_731),
.Y(n_796)
);

NOR2xp33_ASAP7_75t_L g797 ( 
.A(n_666),
.B(n_214),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_SL g798 ( 
.A(n_633),
.B(n_327),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_SL g799 ( 
.A(n_672),
.B(n_327),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_657),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_705),
.B(n_282),
.Y(n_801)
);

HB1xp67_ASAP7_75t_L g802 ( 
.A(n_660),
.Y(n_802)
);

OR2x6_ASAP7_75t_L g803 ( 
.A(n_641),
.B(n_567),
.Y(n_803)
);

INVxp33_ASAP7_75t_L g804 ( 
.A(n_761),
.Y(n_804)
);

BUFx2_ASAP7_75t_L g805 ( 
.A(n_615),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_SL g806 ( 
.A(n_672),
.B(n_327),
.Y(n_806)
);

OR2x2_ASAP7_75t_L g807 ( 
.A(n_687),
.B(n_566),
.Y(n_807)
);

NOR2xp33_ASAP7_75t_L g808 ( 
.A(n_664),
.B(n_214),
.Y(n_808)
);

A2O1A1Ixp33_ASAP7_75t_L g809 ( 
.A1(n_648),
.A2(n_288),
.B(n_323),
.C(n_319),
.Y(n_809)
);

AOI22xp33_ASAP7_75t_L g810 ( 
.A1(n_751),
.A2(n_314),
.B1(n_345),
.B2(n_347),
.Y(n_810)
);

NOR2xp33_ASAP7_75t_L g811 ( 
.A(n_664),
.B(n_218),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_661),
.Y(n_812)
);

NOR3xp33_ASAP7_75t_L g813 ( 
.A(n_686),
.B(n_566),
.C(n_557),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_712),
.B(n_290),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_SL g815 ( 
.A(n_672),
.B(n_307),
.Y(n_815)
);

AOI22xp33_ASAP7_75t_L g816 ( 
.A1(n_751),
.A2(n_311),
.B1(n_371),
.B2(n_396),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_662),
.Y(n_817)
);

OR2x6_ASAP7_75t_L g818 ( 
.A(n_641),
.B(n_575),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_752),
.B(n_266),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_752),
.B(n_267),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_663),
.Y(n_821)
);

NOR2x1p5_ASAP7_75t_L g822 ( 
.A(n_718),
.B(n_551),
.Y(n_822)
);

INVx4_ASAP7_75t_L g823 ( 
.A(n_729),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_752),
.B(n_268),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_SL g825 ( 
.A(n_655),
.B(n_273),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_753),
.Y(n_826)
);

NOR2xp33_ASAP7_75t_L g827 ( 
.A(n_693),
.B(n_218),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_748),
.B(n_279),
.Y(n_828)
);

AND2x2_ASAP7_75t_L g829 ( 
.A(n_756),
.B(n_551),
.Y(n_829)
);

OAI221xp5_ASAP7_75t_L g830 ( 
.A1(n_670),
.A2(n_511),
.B1(n_342),
.B2(n_355),
.C(n_340),
.Y(n_830)
);

NAND2x1_ASAP7_75t_L g831 ( 
.A(n_714),
.B(n_73),
.Y(n_831)
);

AOI22xp33_ASAP7_75t_L g832 ( 
.A1(n_631),
.A2(n_312),
.B1(n_239),
.B2(n_416),
.Y(n_832)
);

AND2x2_ASAP7_75t_L g833 ( 
.A(n_616),
.B(n_654),
.Y(n_833)
);

AND2x2_ASAP7_75t_L g834 ( 
.A(n_654),
.B(n_557),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_747),
.B(n_280),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_SL g836 ( 
.A(n_665),
.B(n_281),
.Y(n_836)
);

BUFx6f_ASAP7_75t_L g837 ( 
.A(n_629),
.Y(n_837)
);

INVxp67_ASAP7_75t_SL g838 ( 
.A(n_729),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_747),
.B(n_287),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_675),
.B(n_298),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_679),
.Y(n_841)
);

AOI22xp33_ASAP7_75t_L g842 ( 
.A1(n_670),
.A2(n_696),
.B1(n_671),
.B2(n_624),
.Y(n_842)
);

BUFx3_ASAP7_75t_L g843 ( 
.A(n_629),
.Y(n_843)
);

AOI21xp5_ASAP7_75t_L g844 ( 
.A1(n_668),
.A2(n_690),
.B(n_711),
.Y(n_844)
);

AND2x4_ASAP7_75t_L g845 ( 
.A(n_683),
.B(n_222),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_692),
.B(n_304),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_SL g847 ( 
.A(n_636),
.B(n_318),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_745),
.B(n_320),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_639),
.Y(n_849)
);

NOR2xp33_ASAP7_75t_L g850 ( 
.A(n_685),
.B(n_222),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_745),
.B(n_328),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_638),
.B(n_640),
.Y(n_852)
);

AND2x4_ASAP7_75t_SL g853 ( 
.A(n_699),
.B(n_610),
.Y(n_853)
);

INVx2_ASAP7_75t_L g854 ( 
.A(n_642),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_643),
.B(n_331),
.Y(n_855)
);

OAI22xp33_ASAP7_75t_L g856 ( 
.A1(n_680),
.A2(n_239),
.B1(n_416),
.B2(n_254),
.Y(n_856)
);

BUFx3_ASAP7_75t_L g857 ( 
.A(n_653),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_644),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_647),
.B(n_335),
.Y(n_859)
);

AOI22xp5_ASAP7_75t_L g860 ( 
.A1(n_678),
.A2(n_354),
.B1(n_336),
.B2(n_337),
.Y(n_860)
);

NOR2xp33_ASAP7_75t_L g861 ( 
.A(n_689),
.B(n_228),
.Y(n_861)
);

AND2x2_ASAP7_75t_L g862 ( 
.A(n_725),
.B(n_569),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_622),
.B(n_341),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_697),
.Y(n_864)
);

OAI22xp5_ASAP7_75t_L g865 ( 
.A1(n_680),
.A2(n_231),
.B1(n_415),
.B2(n_234),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_659),
.Y(n_866)
);

INVx2_ASAP7_75t_L g867 ( 
.A(n_625),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_681),
.B(n_352),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_697),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_SL g870 ( 
.A(n_646),
.B(n_358),
.Y(n_870)
);

HB1xp67_ASAP7_75t_L g871 ( 
.A(n_734),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_703),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_703),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_SL g874 ( 
.A(n_658),
.B(n_360),
.Y(n_874)
);

INVx2_ASAP7_75t_L g875 ( 
.A(n_625),
.Y(n_875)
);

NOR2xp33_ASAP7_75t_L g876 ( 
.A(n_732),
.B(n_228),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_627),
.Y(n_877)
);

NOR2xp33_ASAP7_75t_L g878 ( 
.A(n_732),
.B(n_231),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_688),
.B(n_364),
.Y(n_879)
);

NAND2xp33_ASAP7_75t_L g880 ( 
.A(n_696),
.B(n_365),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_715),
.Y(n_881)
);

NOR2xp33_ASAP7_75t_SL g882 ( 
.A(n_677),
.B(n_569),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_688),
.B(n_367),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_SL g884 ( 
.A(n_637),
.B(n_370),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_SL g885 ( 
.A(n_695),
.B(n_234),
.Y(n_885)
);

NOR2xp33_ASAP7_75t_L g886 ( 
.A(n_733),
.B(n_238),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_716),
.Y(n_887)
);

NOR2xp67_ASAP7_75t_SL g888 ( 
.A(n_721),
.B(n_238),
.Y(n_888)
);

NAND2x1_ASAP7_75t_L g889 ( 
.A(n_714),
.B(n_74),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_744),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_695),
.B(n_241),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_744),
.Y(n_892)
);

NAND2xp33_ASAP7_75t_SL g893 ( 
.A(n_721),
.B(n_254),
.Y(n_893)
);

NOR2xp33_ASAP7_75t_L g894 ( 
.A(n_733),
.B(n_241),
.Y(n_894)
);

OR2x6_ASAP7_75t_L g895 ( 
.A(n_677),
.B(n_573),
.Y(n_895)
);

AND2x4_ASAP7_75t_L g896 ( 
.A(n_653),
.B(n_243),
.Y(n_896)
);

AOI22x1_ASAP7_75t_L g897 ( 
.A1(n_706),
.A2(n_379),
.B1(n_245),
.B2(n_415),
.Y(n_897)
);

OAI22xp33_ASAP7_75t_L g898 ( 
.A1(n_680),
.A2(n_312),
.B1(n_372),
.B2(n_414),
.Y(n_898)
);

CKINVDCx5p33_ASAP7_75t_R g899 ( 
.A(n_753),
.Y(n_899)
);

AOI21xp5_ASAP7_75t_L g900 ( 
.A1(n_690),
.A2(n_245),
.B(n_250),
.Y(n_900)
);

INVx3_ASAP7_75t_L g901 ( 
.A(n_744),
.Y(n_901)
);

INVx2_ASAP7_75t_SL g902 ( 
.A(n_653),
.Y(n_902)
);

AOI22xp5_ASAP7_75t_L g903 ( 
.A1(n_723),
.A2(n_250),
.B1(n_251),
.B2(n_252),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_SL g904 ( 
.A(n_708),
.B(n_251),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_708),
.B(n_252),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_720),
.B(n_309),
.Y(n_906)
);

OR2x2_ASAP7_75t_L g907 ( 
.A(n_626),
.B(n_573),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_724),
.B(n_309),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_735),
.B(n_310),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_737),
.Y(n_910)
);

AOI22xp5_ASAP7_75t_L g911 ( 
.A1(n_723),
.A2(n_387),
.B1(n_379),
.B2(n_310),
.Y(n_911)
);

INVx2_ASAP7_75t_L g912 ( 
.A(n_627),
.Y(n_912)
);

NOR2xp33_ASAP7_75t_L g913 ( 
.A(n_742),
.B(n_387),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_738),
.B(n_389),
.Y(n_914)
);

INVx4_ASAP7_75t_L g915 ( 
.A(n_729),
.Y(n_915)
);

NOR2xp33_ASAP7_75t_L g916 ( 
.A(n_746),
.B(n_389),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_739),
.Y(n_917)
);

NOR2x1p5_ASAP7_75t_L g918 ( 
.A(n_759),
.B(n_375),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_743),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_755),
.B(n_405),
.Y(n_920)
);

INVx2_ASAP7_75t_SL g921 ( 
.A(n_734),
.Y(n_921)
);

AOI21xp5_ASAP7_75t_L g922 ( 
.A1(n_844),
.A2(n_690),
.B(n_714),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_782),
.B(n_700),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_782),
.B(n_783),
.Y(n_924)
);

AOI21xp5_ASAP7_75t_L g925 ( 
.A1(n_815),
.A2(n_726),
.B(n_669),
.Y(n_925)
);

INVx2_ASAP7_75t_L g926 ( 
.A(n_849),
.Y(n_926)
);

NOR3xp33_ASAP7_75t_L g927 ( 
.A(n_913),
.B(n_691),
.C(n_758),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_890),
.Y(n_928)
);

AOI22xp5_ASAP7_75t_L g929 ( 
.A1(n_783),
.A2(n_795),
.B1(n_785),
.B2(n_808),
.Y(n_929)
);

OAI21xp5_ASAP7_75t_L g930 ( 
.A1(n_766),
.A2(n_669),
.B(n_632),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_795),
.B(n_700),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_913),
.B(n_701),
.Y(n_932)
);

INVx3_ASAP7_75t_L g933 ( 
.A(n_775),
.Y(n_933)
);

AOI21xp5_ASAP7_75t_L g934 ( 
.A1(n_815),
.A2(n_726),
.B(n_667),
.Y(n_934)
);

AND2x4_ASAP7_75t_L g935 ( 
.A(n_843),
.B(n_734),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_916),
.B(n_701),
.Y(n_936)
);

OAI22xp5_ASAP7_75t_L g937 ( 
.A1(n_810),
.A2(n_727),
.B1(n_759),
.B2(n_713),
.Y(n_937)
);

OAI21xp5_ASAP7_75t_L g938 ( 
.A1(n_766),
.A2(n_632),
.B(n_709),
.Y(n_938)
);

AND2x2_ASAP7_75t_SL g939 ( 
.A(n_853),
.B(n_762),
.Y(n_939)
);

A2O1A1Ixp33_ASAP7_75t_L g940 ( 
.A1(n_808),
.A2(n_727),
.B(n_754),
.C(n_762),
.Y(n_940)
);

A2O1A1Ixp33_ASAP7_75t_L g941 ( 
.A1(n_811),
.A2(n_750),
.B(n_709),
.C(n_728),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_833),
.B(n_719),
.Y(n_942)
);

AND2x2_ASAP7_75t_L g943 ( 
.A(n_834),
.B(n_797),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_892),
.Y(n_944)
);

AOI22xp5_ASAP7_75t_L g945 ( 
.A1(n_785),
.A2(n_682),
.B1(n_696),
.B2(n_734),
.Y(n_945)
);

AND2x2_ASAP7_75t_L g946 ( 
.A(n_797),
.B(n_699),
.Y(n_946)
);

AOI21xp5_ASAP7_75t_L g947 ( 
.A1(n_823),
.A2(n_915),
.B(n_838),
.Y(n_947)
);

AOI21xp5_ASAP7_75t_L g948 ( 
.A1(n_823),
.A2(n_667),
.B(n_617),
.Y(n_948)
);

AOI21xp5_ASAP7_75t_L g949 ( 
.A1(n_915),
.A2(n_741),
.B(n_620),
.Y(n_949)
);

OAI22xp5_ASAP7_75t_L g950 ( 
.A1(n_810),
.A2(n_816),
.B1(n_763),
.B2(n_767),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_916),
.B(n_741),
.Y(n_951)
);

AOI21xp5_ASAP7_75t_L g952 ( 
.A1(n_799),
.A2(n_620),
.B(n_719),
.Y(n_952)
);

INVx3_ASAP7_75t_SL g953 ( 
.A(n_895),
.Y(n_953)
);

AOI21xp5_ASAP7_75t_L g954 ( 
.A1(n_799),
.A2(n_620),
.B(n_722),
.Y(n_954)
);

AOI21xp5_ASAP7_75t_L g955 ( 
.A1(n_806),
.A2(n_620),
.B(n_722),
.Y(n_955)
);

AOI21x1_ASAP7_75t_L g956 ( 
.A1(n_806),
.A2(n_740),
.B(n_728),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_827),
.B(n_674),
.Y(n_957)
);

NOR2xp33_ASAP7_75t_L g958 ( 
.A(n_804),
.B(n_757),
.Y(n_958)
);

INVx3_ASAP7_75t_L g959 ( 
.A(n_775),
.Y(n_959)
);

AOI21xp5_ASAP7_75t_L g960 ( 
.A1(n_819),
.A2(n_740),
.B(n_673),
.Y(n_960)
);

NOR2xp33_ASAP7_75t_L g961 ( 
.A(n_796),
.B(n_699),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_827),
.B(n_674),
.Y(n_962)
);

INVx3_ASAP7_75t_L g963 ( 
.A(n_775),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_SL g964 ( 
.A(n_837),
.B(n_749),
.Y(n_964)
);

O2A1O1Ixp33_ASAP7_75t_L g965 ( 
.A1(n_809),
.A2(n_704),
.B(n_694),
.C(n_736),
.Y(n_965)
);

OAI21xp5_ASAP7_75t_L g966 ( 
.A1(n_842),
.A2(n_696),
.B(n_694),
.Y(n_966)
);

INVx3_ASAP7_75t_L g967 ( 
.A(n_775),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_SL g968 ( 
.A(n_837),
.B(n_749),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_SL g969 ( 
.A(n_837),
.B(n_749),
.Y(n_969)
);

BUFx12f_ASAP7_75t_L g970 ( 
.A(n_803),
.Y(n_970)
);

BUFx3_ASAP7_75t_L g971 ( 
.A(n_805),
.Y(n_971)
);

AOI21xp5_ASAP7_75t_L g972 ( 
.A1(n_820),
.A2(n_710),
.B(n_673),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_850),
.B(n_861),
.Y(n_973)
);

A2O1A1Ixp33_ASAP7_75t_L g974 ( 
.A1(n_811),
.A2(n_750),
.B(n_736),
.C(n_730),
.Y(n_974)
);

O2A1O1Ixp33_ASAP7_75t_SL g975 ( 
.A1(n_847),
.A2(n_836),
.B(n_825),
.C(n_787),
.Y(n_975)
);

AOI21xp5_ASAP7_75t_L g976 ( 
.A1(n_824),
.A2(n_673),
.B(n_710),
.Y(n_976)
);

AOI22xp33_ASAP7_75t_L g977 ( 
.A1(n_786),
.A2(n_696),
.B1(n_736),
.B2(n_730),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_SL g978 ( 
.A(n_837),
.B(n_405),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_850),
.B(n_674),
.Y(n_979)
);

AOI21xp5_ASAP7_75t_L g980 ( 
.A1(n_768),
.A2(n_852),
.B(n_836),
.Y(n_980)
);

OAI21xp5_ASAP7_75t_L g981 ( 
.A1(n_842),
.A2(n_696),
.B(n_730),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_861),
.B(n_694),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_828),
.B(n_704),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_779),
.B(n_704),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_901),
.B(n_650),
.Y(n_985)
);

AOI21xp5_ASAP7_75t_L g986 ( 
.A1(n_825),
.A2(n_673),
.B(n_717),
.Y(n_986)
);

AOI21xp5_ASAP7_75t_L g987 ( 
.A1(n_835),
.A2(n_673),
.B(n_717),
.Y(n_987)
);

AOI21xp5_ASAP7_75t_L g988 ( 
.A1(n_839),
.A2(n_717),
.B(n_710),
.Y(n_988)
);

NOR2xp33_ASAP7_75t_L g989 ( 
.A(n_829),
.B(n_677),
.Y(n_989)
);

AOI21xp5_ASAP7_75t_L g990 ( 
.A1(n_778),
.A2(n_717),
.B(n_710),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_901),
.Y(n_991)
);

AOI21x1_ASAP7_75t_L g992 ( 
.A1(n_780),
.A2(n_684),
.B(n_650),
.Y(n_992)
);

INVx2_ASAP7_75t_L g993 ( 
.A(n_854),
.Y(n_993)
);

AOI21x1_ASAP7_75t_L g994 ( 
.A1(n_780),
.A2(n_684),
.B(n_650),
.Y(n_994)
);

OAI21xp33_ASAP7_75t_L g995 ( 
.A1(n_763),
.A2(n_425),
.B(n_390),
.Y(n_995)
);

AOI21x1_ASAP7_75t_L g996 ( 
.A1(n_787),
.A2(n_684),
.B(n_717),
.Y(n_996)
);

AOI21xp5_ASAP7_75t_L g997 ( 
.A1(n_848),
.A2(n_851),
.B(n_771),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_769),
.B(n_407),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_776),
.B(n_800),
.Y(n_999)
);

NAND3xp33_ASAP7_75t_SL g1000 ( 
.A(n_907),
.B(n_386),
.C(n_374),
.Y(n_1000)
);

O2A1O1Ixp33_ASAP7_75t_SL g1001 ( 
.A1(n_847),
.A2(n_425),
.B(n_375),
.C(n_368),
.Y(n_1001)
);

O2A1O1Ixp5_ASAP7_75t_L g1002 ( 
.A1(n_870),
.A2(n_366),
.B(n_368),
.C(n_409),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_812),
.Y(n_1003)
);

OAI21xp33_ASAP7_75t_L g1004 ( 
.A1(n_832),
.A2(n_386),
.B(n_414),
.Y(n_1004)
);

AND2x4_ASAP7_75t_L g1005 ( 
.A(n_843),
.B(n_760),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_817),
.B(n_410),
.Y(n_1006)
);

OAI321xp33_ASAP7_75t_L g1007 ( 
.A1(n_856),
.A2(n_760),
.A3(n_413),
.B1(n_398),
.B2(n_394),
.C(n_391),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_821),
.B(n_378),
.Y(n_1008)
);

O2A1O1Ixp33_ASAP7_75t_L g1009 ( 
.A1(n_864),
.A2(n_760),
.B(n_366),
.C(n_368),
.Y(n_1009)
);

AND2x2_ASAP7_75t_L g1010 ( 
.A(n_770),
.B(n_760),
.Y(n_1010)
);

AOI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_868),
.A2(n_413),
.B(n_398),
.Y(n_1011)
);

AO21x1_ASAP7_75t_L g1012 ( 
.A1(n_876),
.A2(n_886),
.B(n_878),
.Y(n_1012)
);

AOI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_879),
.A2(n_394),
.B(n_391),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_841),
.Y(n_1014)
);

AOI21xp5_ASAP7_75t_L g1015 ( 
.A1(n_883),
.A2(n_390),
.B(n_385),
.Y(n_1015)
);

AOI21x1_ASAP7_75t_L g1016 ( 
.A1(n_790),
.A2(n_366),
.B(n_76),
.Y(n_1016)
);

AOI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_880),
.A2(n_378),
.B(n_376),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_816),
.B(n_376),
.Y(n_1018)
);

AND2x6_ASAP7_75t_SL g1019 ( 
.A(n_803),
.B(n_374),
.Y(n_1019)
);

AOI21x1_ASAP7_75t_L g1020 ( 
.A1(n_790),
.A2(n_137),
.B(n_78),
.Y(n_1020)
);

AOI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_840),
.A2(n_373),
.B(n_372),
.Y(n_1021)
);

AOI21x1_ASAP7_75t_L g1022 ( 
.A1(n_798),
.A2(n_123),
.B(n_208),
.Y(n_1022)
);

OAI22xp5_ASAP7_75t_L g1023 ( 
.A1(n_774),
.A2(n_373),
.B1(n_19),
.B2(n_20),
.Y(n_1023)
);

AOI21x1_ASAP7_75t_L g1024 ( 
.A1(n_798),
.A2(n_191),
.B(n_173),
.Y(n_1024)
);

AND2x2_ASAP7_75t_L g1025 ( 
.A(n_802),
.B(n_18),
.Y(n_1025)
);

INVx3_ASAP7_75t_L g1026 ( 
.A(n_857),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_876),
.B(n_18),
.Y(n_1027)
);

AOI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_846),
.A2(n_172),
.B(n_167),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_878),
.B(n_24),
.Y(n_1029)
);

AOI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_866),
.A2(n_165),
.B(n_138),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_SL g1031 ( 
.A(n_857),
.B(n_902),
.Y(n_1031)
);

OAI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_786),
.A2(n_119),
.B(n_116),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_886),
.B(n_24),
.Y(n_1033)
);

OAI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_789),
.A2(n_105),
.B(n_99),
.Y(n_1034)
);

AND2x4_ASAP7_75t_L g1035 ( 
.A(n_921),
.B(n_91),
.Y(n_1035)
);

AOI21xp5_ASAP7_75t_L g1036 ( 
.A1(n_855),
.A2(n_87),
.B(n_77),
.Y(n_1036)
);

OAI21xp5_ASAP7_75t_L g1037 ( 
.A1(n_789),
.A2(n_774),
.B(n_869),
.Y(n_1037)
);

AOI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_859),
.A2(n_26),
.B(n_29),
.Y(n_1038)
);

BUFx6f_ASAP7_75t_L g1039 ( 
.A(n_831),
.Y(n_1039)
);

NOR2x1p5_ASAP7_75t_SL g1040 ( 
.A(n_867),
.B(n_29),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_894),
.B(n_30),
.Y(n_1041)
);

NOR2xp67_ASAP7_75t_L g1042 ( 
.A(n_772),
.B(n_30),
.Y(n_1042)
);

INVx5_ASAP7_75t_L g1043 ( 
.A(n_785),
.Y(n_1043)
);

AOI21x1_ASAP7_75t_L g1044 ( 
.A1(n_884),
.A2(n_33),
.B(n_35),
.Y(n_1044)
);

OAI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_872),
.A2(n_36),
.B(n_37),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_873),
.B(n_39),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_SL g1047 ( 
.A(n_894),
.B(n_41),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_785),
.B(n_41),
.Y(n_1048)
);

AOI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_863),
.A2(n_42),
.B(n_43),
.Y(n_1049)
);

O2A1O1Ixp33_ASAP7_75t_L g1050 ( 
.A1(n_885),
.A2(n_43),
.B(n_45),
.C(n_46),
.Y(n_1050)
);

INVx2_ASAP7_75t_L g1051 ( 
.A(n_764),
.Y(n_1051)
);

AOI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_884),
.A2(n_45),
.B(n_48),
.Y(n_1052)
);

NOR3xp33_ASAP7_75t_L g1053 ( 
.A(n_862),
.B(n_50),
.C(n_52),
.Y(n_1053)
);

NOR2xp67_ASAP7_75t_L g1054 ( 
.A(n_807),
.B(n_830),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_910),
.Y(n_1055)
);

AOI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_875),
.A2(n_52),
.B(n_53),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_SL g1057 ( 
.A(n_856),
.B(n_54),
.Y(n_1057)
);

AOI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_877),
.A2(n_56),
.B(n_58),
.Y(n_1058)
);

AOI22xp5_ASAP7_75t_L g1059 ( 
.A1(n_785),
.A2(n_59),
.B1(n_60),
.B2(n_62),
.Y(n_1059)
);

OAI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_794),
.A2(n_60),
.B(n_62),
.Y(n_1060)
);

O2A1O1Ixp5_ASAP7_75t_L g1061 ( 
.A1(n_870),
.A2(n_874),
.B(n_888),
.C(n_814),
.Y(n_1061)
);

NOR3xp33_ASAP7_75t_L g1062 ( 
.A(n_813),
.B(n_898),
.C(n_865),
.Y(n_1062)
);

AND2x6_ASAP7_75t_L g1063 ( 
.A(n_858),
.B(n_896),
.Y(n_1063)
);

AOI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_912),
.A2(n_791),
.B(n_793),
.Y(n_1064)
);

O2A1O1Ixp33_ASAP7_75t_L g1065 ( 
.A1(n_885),
.A2(n_904),
.B(n_874),
.C(n_802),
.Y(n_1065)
);

O2A1O1Ixp33_ASAP7_75t_L g1066 ( 
.A1(n_904),
.A2(n_788),
.B(n_801),
.C(n_784),
.Y(n_1066)
);

INVx3_ASAP7_75t_L g1067 ( 
.A(n_917),
.Y(n_1067)
);

BUFx6f_ASAP7_75t_L g1068 ( 
.A(n_889),
.Y(n_1068)
);

AND2x2_ASAP7_75t_L g1069 ( 
.A(n_792),
.B(n_896),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_881),
.B(n_887),
.Y(n_1070)
);

O2A1O1Ixp33_ASAP7_75t_L g1071 ( 
.A1(n_891),
.A2(n_905),
.B(n_898),
.C(n_871),
.Y(n_1071)
);

AOI21xp5_ASAP7_75t_L g1072 ( 
.A1(n_919),
.A2(n_920),
.B(n_914),
.Y(n_1072)
);

INVx1_ASAP7_75t_SL g1073 ( 
.A(n_803),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_871),
.Y(n_1074)
);

AO22x1_ASAP7_75t_L g1075 ( 
.A1(n_845),
.A2(n_909),
.B1(n_908),
.B2(n_906),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_845),
.B(n_860),
.Y(n_1076)
);

INVx4_ASAP7_75t_L g1077 ( 
.A(n_765),
.Y(n_1077)
);

NOR2xp33_ASAP7_75t_L g1078 ( 
.A(n_792),
.B(n_911),
.Y(n_1078)
);

NOR2xp33_ASAP7_75t_L g1079 ( 
.A(n_903),
.B(n_777),
.Y(n_1079)
);

INVx3_ASAP7_75t_L g1080 ( 
.A(n_765),
.Y(n_1080)
);

OAI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_900),
.A2(n_832),
.B(n_893),
.Y(n_1081)
);

INVx2_ASAP7_75t_L g1082 ( 
.A(n_897),
.Y(n_1082)
);

BUFx4f_ASAP7_75t_L g1083 ( 
.A(n_818),
.Y(n_1083)
);

AOI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_765),
.A2(n_773),
.B(n_781),
.Y(n_1084)
);

AOI22xp5_ASAP7_75t_L g1085 ( 
.A1(n_822),
.A2(n_918),
.B1(n_882),
.B2(n_895),
.Y(n_1085)
);

AOI21xp5_ASAP7_75t_L g1086 ( 
.A1(n_818),
.A2(n_895),
.B(n_826),
.Y(n_1086)
);

BUFx8_ASAP7_75t_SL g1087 ( 
.A(n_899),
.Y(n_1087)
);

AND2x4_ASAP7_75t_L g1088 ( 
.A(n_818),
.B(n_843),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_782),
.B(n_833),
.Y(n_1089)
);

NAND2x1p5_ASAP7_75t_L g1090 ( 
.A(n_775),
.B(n_771),
.Y(n_1090)
);

OAI21xp5_ASAP7_75t_L g1091 ( 
.A1(n_766),
.A2(n_806),
.B(n_799),
.Y(n_1091)
);

CKINVDCx16_ASAP7_75t_R g1092 ( 
.A(n_882),
.Y(n_1092)
);

AOI21xp5_ASAP7_75t_L g1093 ( 
.A1(n_844),
.A2(n_690),
.B(n_672),
.Y(n_1093)
);

NAND2x1p5_ASAP7_75t_L g1094 ( 
.A(n_775),
.B(n_771),
.Y(n_1094)
);

HB1xp67_ASAP7_75t_L g1095 ( 
.A(n_796),
.Y(n_1095)
);

AOI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_844),
.A2(n_690),
.B(n_672),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_SL g1097 ( 
.A(n_837),
.B(n_628),
.Y(n_1097)
);

NOR2xp33_ASAP7_75t_L g1098 ( 
.A(n_804),
.B(n_782),
.Y(n_1098)
);

OAI22xp5_ASAP7_75t_L g1099 ( 
.A1(n_810),
.A2(n_816),
.B1(n_763),
.B2(n_628),
.Y(n_1099)
);

OAI22xp5_ASAP7_75t_L g1100 ( 
.A1(n_810),
.A2(n_816),
.B1(n_763),
.B2(n_628),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_782),
.B(n_783),
.Y(n_1101)
);

OAI22xp5_ASAP7_75t_L g1102 ( 
.A1(n_810),
.A2(n_816),
.B1(n_763),
.B2(n_628),
.Y(n_1102)
);

AOI21xp33_ASAP7_75t_L g1103 ( 
.A1(n_924),
.A2(n_1101),
.B(n_973),
.Y(n_1103)
);

AOI21x1_ASAP7_75t_L g1104 ( 
.A1(n_957),
.A2(n_962),
.B(n_979),
.Y(n_1104)
);

AOI21x1_ASAP7_75t_L g1105 ( 
.A1(n_982),
.A2(n_980),
.B(n_922),
.Y(n_1105)
);

OAI21x1_ASAP7_75t_L g1106 ( 
.A1(n_956),
.A2(n_1096),
.B(n_1093),
.Y(n_1106)
);

BUFx4f_ASAP7_75t_SL g1107 ( 
.A(n_970),
.Y(n_1107)
);

BUFx6f_ASAP7_75t_L g1108 ( 
.A(n_935),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_1089),
.B(n_1098),
.Y(n_1109)
);

AOI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_983),
.A2(n_997),
.B(n_975),
.Y(n_1110)
);

OAI22xp5_ASAP7_75t_L g1111 ( 
.A1(n_1099),
.A2(n_1102),
.B1(n_1100),
.B2(n_950),
.Y(n_1111)
);

OAI21xp5_ASAP7_75t_L g1112 ( 
.A1(n_1099),
.A2(n_1102),
.B(n_1100),
.Y(n_1112)
);

AOI21x1_ASAP7_75t_L g1113 ( 
.A1(n_951),
.A2(n_1075),
.B(n_960),
.Y(n_1113)
);

OAI21x1_ASAP7_75t_L g1114 ( 
.A1(n_952),
.A2(n_955),
.B(n_954),
.Y(n_1114)
);

NAND2x1_ASAP7_75t_L g1115 ( 
.A(n_933),
.B(n_959),
.Y(n_1115)
);

A2O1A1Ixp33_ASAP7_75t_L g1116 ( 
.A1(n_929),
.A2(n_950),
.B(n_923),
.C(n_1065),
.Y(n_1116)
);

OAI21x1_ASAP7_75t_L g1117 ( 
.A1(n_996),
.A2(n_994),
.B(n_992),
.Y(n_1117)
);

BUFx12f_ASAP7_75t_L g1118 ( 
.A(n_1019),
.Y(n_1118)
);

AO31x2_ASAP7_75t_L g1119 ( 
.A1(n_1012),
.A2(n_941),
.A3(n_974),
.B(n_940),
.Y(n_1119)
);

OAI21x1_ASAP7_75t_L g1120 ( 
.A1(n_948),
.A2(n_981),
.B(n_966),
.Y(n_1120)
);

AOI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_1091),
.A2(n_981),
.B(n_966),
.Y(n_1121)
);

OAI21x1_ASAP7_75t_L g1122 ( 
.A1(n_972),
.A2(n_976),
.B(n_965),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_1089),
.B(n_931),
.Y(n_1123)
);

OAI21x1_ASAP7_75t_SL g1124 ( 
.A1(n_1045),
.A2(n_1034),
.B(n_1032),
.Y(n_1124)
);

OAI21x1_ASAP7_75t_L g1125 ( 
.A1(n_986),
.A2(n_934),
.B(n_987),
.Y(n_1125)
);

AOI21x1_ASAP7_75t_L g1126 ( 
.A1(n_984),
.A2(n_985),
.B(n_1072),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_SL g1127 ( 
.A(n_943),
.B(n_946),
.Y(n_1127)
);

OR2x6_ASAP7_75t_L g1128 ( 
.A(n_971),
.B(n_1088),
.Y(n_1128)
);

OAI21xp5_ASAP7_75t_L g1129 ( 
.A1(n_1091),
.A2(n_1037),
.B(n_930),
.Y(n_1129)
);

OAI21x1_ASAP7_75t_L g1130 ( 
.A1(n_988),
.A2(n_949),
.B(n_1064),
.Y(n_1130)
);

INVx2_ASAP7_75t_L g1131 ( 
.A(n_928),
.Y(n_1131)
);

NAND3xp33_ASAP7_75t_L g1132 ( 
.A(n_1027),
.B(n_1033),
.C(n_1029),
.Y(n_1132)
);

AOI21xp5_ASAP7_75t_L g1133 ( 
.A1(n_925),
.A2(n_932),
.B(n_936),
.Y(n_1133)
);

OAI21x1_ASAP7_75t_L g1134 ( 
.A1(n_990),
.A2(n_938),
.B(n_947),
.Y(n_1134)
);

AO31x2_ASAP7_75t_L g1135 ( 
.A1(n_1082),
.A2(n_1041),
.A3(n_937),
.B(n_1048),
.Y(n_1135)
);

AOI21xp5_ASAP7_75t_L g1136 ( 
.A1(n_1043),
.A2(n_1097),
.B(n_1066),
.Y(n_1136)
);

OAI21xp5_ASAP7_75t_L g1137 ( 
.A1(n_1037),
.A2(n_930),
.B(n_938),
.Y(n_1137)
);

INVx2_ASAP7_75t_L g1138 ( 
.A(n_944),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_1003),
.Y(n_1139)
);

AND2x2_ASAP7_75t_L g1140 ( 
.A(n_958),
.B(n_927),
.Y(n_1140)
);

A2O1A1Ixp33_ASAP7_75t_L g1141 ( 
.A1(n_1079),
.A2(n_1071),
.B(n_1081),
.C(n_937),
.Y(n_1141)
);

INVx8_ASAP7_75t_L g1142 ( 
.A(n_1063),
.Y(n_1142)
);

NAND2x1p5_ASAP7_75t_L g1143 ( 
.A(n_1077),
.B(n_1080),
.Y(n_1143)
);

OAI21x1_ASAP7_75t_L g1144 ( 
.A1(n_942),
.A2(n_1024),
.B(n_1020),
.Y(n_1144)
);

INVx3_ASAP7_75t_L g1145 ( 
.A(n_933),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_942),
.B(n_999),
.Y(n_1146)
);

OAI21xp5_ASAP7_75t_L g1147 ( 
.A1(n_1081),
.A2(n_1061),
.B(n_1032),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_1014),
.B(n_1055),
.Y(n_1148)
);

AOI21xp5_ASAP7_75t_L g1149 ( 
.A1(n_1043),
.A2(n_1076),
.B(n_1034),
.Y(n_1149)
);

AND3x1_ASAP7_75t_SL g1150 ( 
.A(n_1074),
.B(n_1007),
.C(n_995),
.Y(n_1150)
);

AND2x2_ASAP7_75t_L g1151 ( 
.A(n_961),
.B(n_1069),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_1070),
.B(n_1046),
.Y(n_1152)
);

OAI21x1_ASAP7_75t_L g1153 ( 
.A1(n_1022),
.A2(n_1084),
.B(n_1016),
.Y(n_1153)
);

OAI21x1_ASAP7_75t_L g1154 ( 
.A1(n_1090),
.A2(n_1094),
.B(n_926),
.Y(n_1154)
);

NOR2xp67_ASAP7_75t_L g1155 ( 
.A(n_1026),
.B(n_1080),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_SL g1156 ( 
.A(n_1054),
.B(n_935),
.Y(n_1156)
);

BUFx2_ASAP7_75t_L g1157 ( 
.A(n_1088),
.Y(n_1157)
);

AOI21x1_ASAP7_75t_L g1158 ( 
.A1(n_991),
.A2(n_1031),
.B(n_978),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_1051),
.Y(n_1159)
);

OAI21x1_ASAP7_75t_L g1160 ( 
.A1(n_1090),
.A2(n_1094),
.B(n_993),
.Y(n_1160)
);

A2O1A1Ixp33_ASAP7_75t_L g1161 ( 
.A1(n_1062),
.A2(n_1078),
.B(n_1018),
.C(n_1047),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_SL g1162 ( 
.A(n_1092),
.B(n_1026),
.Y(n_1162)
);

OR2x6_ASAP7_75t_L g1163 ( 
.A(n_1086),
.B(n_1005),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_L g1164 ( 
.A(n_1046),
.B(n_1067),
.Y(n_1164)
);

BUFx6f_ASAP7_75t_L g1165 ( 
.A(n_1077),
.Y(n_1165)
);

BUFx12f_ASAP7_75t_L g1166 ( 
.A(n_1005),
.Y(n_1166)
);

INVx2_ASAP7_75t_SL g1167 ( 
.A(n_1025),
.Y(n_1167)
);

AOI21xp5_ASAP7_75t_L g1168 ( 
.A1(n_1043),
.A2(n_977),
.B(n_1039),
.Y(n_1168)
);

OR2x6_ASAP7_75t_L g1169 ( 
.A(n_1010),
.B(n_1035),
.Y(n_1169)
);

INVxp67_ASAP7_75t_SL g1170 ( 
.A(n_959),
.Y(n_1170)
);

OAI22xp5_ASAP7_75t_L g1171 ( 
.A1(n_1023),
.A2(n_1045),
.B1(n_1057),
.B2(n_1043),
.Y(n_1171)
);

AND2x2_ASAP7_75t_L g1172 ( 
.A(n_989),
.B(n_939),
.Y(n_1172)
);

NOR2x1_ASAP7_75t_SL g1173 ( 
.A(n_1039),
.B(n_1068),
.Y(n_1173)
);

AOI21xp5_ASAP7_75t_L g1174 ( 
.A1(n_1039),
.A2(n_1068),
.B(n_967),
.Y(n_1174)
);

BUFx6f_ASAP7_75t_L g1175 ( 
.A(n_1035),
.Y(n_1175)
);

A2O1A1Ixp33_ASAP7_75t_L g1176 ( 
.A1(n_1052),
.A2(n_945),
.B(n_1050),
.C(n_1017),
.Y(n_1176)
);

A2O1A1Ixp33_ASAP7_75t_L g1177 ( 
.A1(n_1004),
.A2(n_1021),
.B(n_1049),
.C(n_1038),
.Y(n_1177)
);

INVx2_ASAP7_75t_SL g1178 ( 
.A(n_1073),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_SL g1179 ( 
.A(n_963),
.B(n_967),
.Y(n_1179)
);

AOI21x1_ASAP7_75t_L g1180 ( 
.A1(n_964),
.A2(n_968),
.B(n_969),
.Y(n_1180)
);

OAI21x1_ASAP7_75t_L g1181 ( 
.A1(n_963),
.A2(n_1030),
.B(n_1028),
.Y(n_1181)
);

OAI21x1_ASAP7_75t_L g1182 ( 
.A1(n_1036),
.A2(n_1044),
.B(n_1056),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_998),
.B(n_1006),
.Y(n_1183)
);

BUFx5_ASAP7_75t_L g1184 ( 
.A(n_1063),
.Y(n_1184)
);

OAI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_1048),
.A2(n_1002),
.B(n_1060),
.Y(n_1185)
);

INVx2_ASAP7_75t_L g1186 ( 
.A(n_1068),
.Y(n_1186)
);

OAI21x1_ASAP7_75t_L g1187 ( 
.A1(n_1058),
.A2(n_1060),
.B(n_1008),
.Y(n_1187)
);

INVx3_ASAP7_75t_L g1188 ( 
.A(n_1063),
.Y(n_1188)
);

NOR2x1_ASAP7_75t_L g1189 ( 
.A(n_1000),
.B(n_1042),
.Y(n_1189)
);

AO31x2_ASAP7_75t_L g1190 ( 
.A1(n_1023),
.A2(n_1015),
.A3(n_1013),
.B(n_1011),
.Y(n_1190)
);

INVx2_ASAP7_75t_SL g1191 ( 
.A(n_1083),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_1063),
.B(n_1053),
.Y(n_1192)
);

AOI21x1_ASAP7_75t_L g1193 ( 
.A1(n_1040),
.A2(n_1063),
.B(n_1001),
.Y(n_1193)
);

OAI21x1_ASAP7_75t_L g1194 ( 
.A1(n_1059),
.A2(n_1009),
.B(n_1085),
.Y(n_1194)
);

AND2x4_ASAP7_75t_L g1195 ( 
.A(n_1083),
.B(n_953),
.Y(n_1195)
);

AND2x2_ASAP7_75t_L g1196 ( 
.A(n_1087),
.B(n_1098),
.Y(n_1196)
);

OAI21xp5_ASAP7_75t_L g1197 ( 
.A1(n_924),
.A2(n_1101),
.B(n_1100),
.Y(n_1197)
);

OR2x2_ASAP7_75t_L g1198 ( 
.A(n_1089),
.B(n_630),
.Y(n_1198)
);

OAI21xp5_ASAP7_75t_L g1199 ( 
.A1(n_924),
.A2(n_1101),
.B(n_1100),
.Y(n_1199)
);

AOI21xp33_ASAP7_75t_L g1200 ( 
.A1(n_924),
.A2(n_1101),
.B(n_973),
.Y(n_1200)
);

NOR2xp33_ASAP7_75t_L g1201 ( 
.A(n_1098),
.B(n_924),
.Y(n_1201)
);

OA21x2_ASAP7_75t_L g1202 ( 
.A1(n_938),
.A2(n_981),
.B(n_966),
.Y(n_1202)
);

AND2x2_ASAP7_75t_L g1203 ( 
.A(n_1098),
.B(n_943),
.Y(n_1203)
);

AOI221xp5_ASAP7_75t_SL g1204 ( 
.A1(n_950),
.A2(n_1100),
.B1(n_1102),
.B2(n_1099),
.C(n_1101),
.Y(n_1204)
);

AOI21xp5_ASAP7_75t_L g1205 ( 
.A1(n_980),
.A2(n_672),
.B(n_1093),
.Y(n_1205)
);

OAI22xp5_ASAP7_75t_L g1206 ( 
.A1(n_1099),
.A2(n_1102),
.B1(n_1100),
.B2(n_1101),
.Y(n_1206)
);

AOI21xp5_ASAP7_75t_L g1207 ( 
.A1(n_980),
.A2(n_672),
.B(n_1093),
.Y(n_1207)
);

NOR2xp67_ASAP7_75t_L g1208 ( 
.A(n_929),
.B(n_1026),
.Y(n_1208)
);

OR2x2_ASAP7_75t_L g1209 ( 
.A(n_1089),
.B(n_630),
.Y(n_1209)
);

OAI21x1_ASAP7_75t_L g1210 ( 
.A1(n_956),
.A2(n_922),
.B(n_1093),
.Y(n_1210)
);

OR2x2_ASAP7_75t_L g1211 ( 
.A(n_1089),
.B(n_630),
.Y(n_1211)
);

AND2x6_ASAP7_75t_L g1212 ( 
.A(n_929),
.B(n_945),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_924),
.B(n_1101),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_924),
.B(n_1101),
.Y(n_1214)
);

BUFx6f_ASAP7_75t_L g1215 ( 
.A(n_935),
.Y(n_1215)
);

OAI22x1_ASAP7_75t_L g1216 ( 
.A1(n_1057),
.A2(n_1098),
.B1(n_1101),
.B2(n_924),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_924),
.B(n_1101),
.Y(n_1217)
);

OAI21x1_ASAP7_75t_L g1218 ( 
.A1(n_956),
.A2(n_922),
.B(n_1093),
.Y(n_1218)
);

AND2x4_ASAP7_75t_L g1219 ( 
.A(n_1077),
.B(n_935),
.Y(n_1219)
);

OAI21xp5_ASAP7_75t_L g1220 ( 
.A1(n_924),
.A2(n_1101),
.B(n_1100),
.Y(n_1220)
);

OAI21xp5_ASAP7_75t_L g1221 ( 
.A1(n_924),
.A2(n_1101),
.B(n_1100),
.Y(n_1221)
);

OAI21x1_ASAP7_75t_SL g1222 ( 
.A1(n_1045),
.A2(n_1034),
.B(n_1032),
.Y(n_1222)
);

AOI21xp5_ASAP7_75t_L g1223 ( 
.A1(n_980),
.A2(n_672),
.B(n_1093),
.Y(n_1223)
);

BUFx2_ASAP7_75t_L g1224 ( 
.A(n_1095),
.Y(n_1224)
);

OAI21xp5_ASAP7_75t_L g1225 ( 
.A1(n_924),
.A2(n_1101),
.B(n_1100),
.Y(n_1225)
);

AOI221x1_ASAP7_75t_L g1226 ( 
.A1(n_924),
.A2(n_1101),
.B1(n_1099),
.B2(n_1102),
.C(n_1100),
.Y(n_1226)
);

AND2x4_ASAP7_75t_L g1227 ( 
.A(n_1077),
.B(n_935),
.Y(n_1227)
);

OAI21xp5_ASAP7_75t_L g1228 ( 
.A1(n_924),
.A2(n_1101),
.B(n_1100),
.Y(n_1228)
);

OAI21xp5_ASAP7_75t_L g1229 ( 
.A1(n_924),
.A2(n_1101),
.B(n_1100),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_L g1230 ( 
.A(n_924),
.B(n_1101),
.Y(n_1230)
);

INVxp67_ASAP7_75t_L g1231 ( 
.A(n_1095),
.Y(n_1231)
);

HB1xp67_ASAP7_75t_L g1232 ( 
.A(n_1095),
.Y(n_1232)
);

INVx5_ASAP7_75t_L g1233 ( 
.A(n_970),
.Y(n_1233)
);

NAND2x1p5_ASAP7_75t_L g1234 ( 
.A(n_1077),
.B(n_1080),
.Y(n_1234)
);

BUFx6f_ASAP7_75t_L g1235 ( 
.A(n_935),
.Y(n_1235)
);

A2O1A1Ixp33_ASAP7_75t_L g1236 ( 
.A1(n_924),
.A2(n_1101),
.B(n_973),
.C(n_929),
.Y(n_1236)
);

AOI21x1_ASAP7_75t_L g1237 ( 
.A1(n_957),
.A2(n_962),
.B(n_979),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_924),
.B(n_1101),
.Y(n_1238)
);

NOR2xp33_ASAP7_75t_L g1239 ( 
.A(n_1098),
.B(n_924),
.Y(n_1239)
);

O2A1O1Ixp5_ASAP7_75t_L g1240 ( 
.A1(n_924),
.A2(n_1101),
.B(n_973),
.C(n_1012),
.Y(n_1240)
);

BUFx8_ASAP7_75t_SL g1241 ( 
.A(n_1087),
.Y(n_1241)
);

AOI21xp5_ASAP7_75t_L g1242 ( 
.A1(n_980),
.A2(n_672),
.B(n_1093),
.Y(n_1242)
);

BUFx4f_ASAP7_75t_L g1243 ( 
.A(n_953),
.Y(n_1243)
);

INVx5_ASAP7_75t_L g1244 ( 
.A(n_970),
.Y(n_1244)
);

OAI22x1_ASAP7_75t_L g1245 ( 
.A1(n_1057),
.A2(n_1098),
.B1(n_1101),
.B2(n_924),
.Y(n_1245)
);

AOI21xp5_ASAP7_75t_L g1246 ( 
.A1(n_980),
.A2(n_672),
.B(n_1093),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1003),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_L g1248 ( 
.A(n_924),
.B(n_1101),
.Y(n_1248)
);

OAI21x1_ASAP7_75t_L g1249 ( 
.A1(n_956),
.A2(n_922),
.B(n_1093),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_L g1250 ( 
.A(n_924),
.B(n_1101),
.Y(n_1250)
);

BUFx6f_ASAP7_75t_L g1251 ( 
.A(n_935),
.Y(n_1251)
);

AOI21x1_ASAP7_75t_L g1252 ( 
.A1(n_957),
.A2(n_962),
.B(n_979),
.Y(n_1252)
);

NAND3xp33_ASAP7_75t_L g1253 ( 
.A(n_924),
.B(n_1101),
.C(n_973),
.Y(n_1253)
);

NOR2x1_ASAP7_75t_L g1254 ( 
.A(n_961),
.B(n_895),
.Y(n_1254)
);

OAI22xp5_ASAP7_75t_L g1255 ( 
.A1(n_1099),
.A2(n_1102),
.B1(n_1100),
.B2(n_1101),
.Y(n_1255)
);

AOI21xp5_ASAP7_75t_L g1256 ( 
.A1(n_980),
.A2(n_672),
.B(n_1093),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_SL g1257 ( 
.A(n_924),
.B(n_1101),
.Y(n_1257)
);

AOI21x1_ASAP7_75t_L g1258 ( 
.A1(n_957),
.A2(n_962),
.B(n_979),
.Y(n_1258)
);

NOR3xp33_ASAP7_75t_L g1259 ( 
.A(n_1201),
.B(n_1239),
.C(n_1127),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_L g1260 ( 
.A(n_1213),
.B(n_1214),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1139),
.Y(n_1261)
);

AOI21xp5_ASAP7_75t_L g1262 ( 
.A1(n_1133),
.A2(n_1110),
.B(n_1147),
.Y(n_1262)
);

OAI21xp5_ASAP7_75t_L g1263 ( 
.A1(n_1141),
.A2(n_1255),
.B(n_1206),
.Y(n_1263)
);

INVx5_ASAP7_75t_L g1264 ( 
.A(n_1165),
.Y(n_1264)
);

BUFx6f_ASAP7_75t_L g1265 ( 
.A(n_1165),
.Y(n_1265)
);

OAI22xp5_ASAP7_75t_L g1266 ( 
.A1(n_1112),
.A2(n_1111),
.B1(n_1206),
.B2(n_1255),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_L g1267 ( 
.A(n_1217),
.B(n_1230),
.Y(n_1267)
);

AND2x4_ASAP7_75t_L g1268 ( 
.A(n_1219),
.B(n_1227),
.Y(n_1268)
);

HB1xp67_ASAP7_75t_L g1269 ( 
.A(n_1232),
.Y(n_1269)
);

CKINVDCx16_ASAP7_75t_R g1270 ( 
.A(n_1166),
.Y(n_1270)
);

INVx2_ASAP7_75t_SL g1271 ( 
.A(n_1224),
.Y(n_1271)
);

CKINVDCx20_ASAP7_75t_R g1272 ( 
.A(n_1241),
.Y(n_1272)
);

AOI21xp5_ASAP7_75t_L g1273 ( 
.A1(n_1205),
.A2(n_1223),
.B(n_1207),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_SL g1274 ( 
.A(n_1140),
.B(n_1198),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_L g1275 ( 
.A(n_1238),
.B(n_1248),
.Y(n_1275)
);

AOI21xp33_ASAP7_75t_SL g1276 ( 
.A1(n_1162),
.A2(n_1211),
.B(n_1209),
.Y(n_1276)
);

CKINVDCx5p33_ASAP7_75t_R g1277 ( 
.A(n_1128),
.Y(n_1277)
);

NOR2xp33_ASAP7_75t_R g1278 ( 
.A(n_1243),
.B(n_1107),
.Y(n_1278)
);

AOI21xp5_ASAP7_75t_L g1279 ( 
.A1(n_1242),
.A2(n_1256),
.B(n_1246),
.Y(n_1279)
);

AOI21xp5_ASAP7_75t_L g1280 ( 
.A1(n_1168),
.A2(n_1136),
.B(n_1173),
.Y(n_1280)
);

BUFx12f_ASAP7_75t_L g1281 ( 
.A(n_1128),
.Y(n_1281)
);

AOI22xp5_ASAP7_75t_L g1282 ( 
.A1(n_1111),
.A2(n_1203),
.B1(n_1204),
.B2(n_1112),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_L g1283 ( 
.A(n_1250),
.B(n_1109),
.Y(n_1283)
);

BUFx2_ASAP7_75t_SL g1284 ( 
.A(n_1165),
.Y(n_1284)
);

BUFx3_ASAP7_75t_L g1285 ( 
.A(n_1128),
.Y(n_1285)
);

AND2x6_ASAP7_75t_L g1286 ( 
.A(n_1188),
.B(n_1175),
.Y(n_1286)
);

INVx3_ASAP7_75t_L g1287 ( 
.A(n_1142),
.Y(n_1287)
);

OR2x2_ASAP7_75t_L g1288 ( 
.A(n_1257),
.B(n_1253),
.Y(n_1288)
);

OAI21x1_ASAP7_75t_L g1289 ( 
.A1(n_1117),
.A2(n_1106),
.B(n_1210),
.Y(n_1289)
);

INVxp67_ASAP7_75t_L g1290 ( 
.A(n_1178),
.Y(n_1290)
);

BUFx8_ASAP7_75t_L g1291 ( 
.A(n_1157),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_L g1292 ( 
.A(n_1123),
.B(n_1103),
.Y(n_1292)
);

INVx3_ASAP7_75t_L g1293 ( 
.A(n_1142),
.Y(n_1293)
);

INVx3_ASAP7_75t_L g1294 ( 
.A(n_1142),
.Y(n_1294)
);

AND2x2_ASAP7_75t_L g1295 ( 
.A(n_1172),
.B(n_1151),
.Y(n_1295)
);

NOR2xp33_ASAP7_75t_L g1296 ( 
.A(n_1200),
.B(n_1183),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1247),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1148),
.Y(n_1298)
);

AOI21xp5_ASAP7_75t_L g1299 ( 
.A1(n_1124),
.A2(n_1222),
.B(n_1116),
.Y(n_1299)
);

NAND2x2_ASAP7_75t_L g1300 ( 
.A(n_1191),
.B(n_1167),
.Y(n_1300)
);

AND2x4_ASAP7_75t_L g1301 ( 
.A(n_1219),
.B(n_1227),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1138),
.Y(n_1302)
);

BUFx6f_ASAP7_75t_L g1303 ( 
.A(n_1108),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_L g1304 ( 
.A(n_1253),
.B(n_1152),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1146),
.B(n_1197),
.Y(n_1305)
);

BUFx2_ASAP7_75t_L g1306 ( 
.A(n_1231),
.Y(n_1306)
);

BUFx2_ASAP7_75t_L g1307 ( 
.A(n_1169),
.Y(n_1307)
);

HB1xp67_ASAP7_75t_L g1308 ( 
.A(n_1169),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1159),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_L g1310 ( 
.A(n_1197),
.B(n_1199),
.Y(n_1310)
);

INVx5_ASAP7_75t_L g1311 ( 
.A(n_1188),
.Y(n_1311)
);

AO21x1_ASAP7_75t_L g1312 ( 
.A1(n_1199),
.A2(n_1229),
.B(n_1228),
.Y(n_1312)
);

A2O1A1Ixp33_ASAP7_75t_L g1313 ( 
.A1(n_1161),
.A2(n_1229),
.B(n_1225),
.C(n_1228),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_L g1314 ( 
.A(n_1220),
.B(n_1221),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_L g1315 ( 
.A(n_1220),
.B(n_1221),
.Y(n_1315)
);

OAI22xp5_ASAP7_75t_SL g1316 ( 
.A1(n_1171),
.A2(n_1225),
.B1(n_1118),
.B2(n_1216),
.Y(n_1316)
);

BUFx4_ASAP7_75t_SL g1317 ( 
.A(n_1163),
.Y(n_1317)
);

A2O1A1Ixp33_ASAP7_75t_L g1318 ( 
.A1(n_1236),
.A2(n_1240),
.B(n_1132),
.C(n_1204),
.Y(n_1318)
);

OAI22xp5_ASAP7_75t_L g1319 ( 
.A1(n_1171),
.A2(n_1121),
.B1(n_1129),
.B2(n_1132),
.Y(n_1319)
);

OAI22xp5_ASAP7_75t_L g1320 ( 
.A1(n_1129),
.A2(n_1169),
.B1(n_1175),
.B2(n_1137),
.Y(n_1320)
);

AOI21xp5_ASAP7_75t_L g1321 ( 
.A1(n_1176),
.A2(n_1137),
.B(n_1174),
.Y(n_1321)
);

INVx4_ASAP7_75t_SL g1322 ( 
.A(n_1195),
.Y(n_1322)
);

AND2x2_ASAP7_75t_L g1323 ( 
.A(n_1245),
.B(n_1108),
.Y(n_1323)
);

AND2x2_ASAP7_75t_L g1324 ( 
.A(n_1215),
.B(n_1235),
.Y(n_1324)
);

CKINVDCx8_ASAP7_75t_R g1325 ( 
.A(n_1233),
.Y(n_1325)
);

O2A1O1Ixp33_ASAP7_75t_L g1326 ( 
.A1(n_1177),
.A2(n_1156),
.B(n_1192),
.C(n_1185),
.Y(n_1326)
);

AND2x2_ASAP7_75t_L g1327 ( 
.A(n_1215),
.B(n_1251),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_L g1328 ( 
.A(n_1164),
.B(n_1226),
.Y(n_1328)
);

BUFx6f_ASAP7_75t_L g1329 ( 
.A(n_1235),
.Y(n_1329)
);

NOR2xp33_ASAP7_75t_L g1330 ( 
.A(n_1175),
.B(n_1196),
.Y(n_1330)
);

NOR2xp67_ASAP7_75t_SL g1331 ( 
.A(n_1233),
.B(n_1244),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1170),
.Y(n_1332)
);

AND2x4_ASAP7_75t_L g1333 ( 
.A(n_1235),
.B(n_1251),
.Y(n_1333)
);

INVx1_ASAP7_75t_SL g1334 ( 
.A(n_1251),
.Y(n_1334)
);

INVx1_ASAP7_75t_SL g1335 ( 
.A(n_1195),
.Y(n_1335)
);

BUFx2_ASAP7_75t_L g1336 ( 
.A(n_1163),
.Y(n_1336)
);

INVx3_ASAP7_75t_L g1337 ( 
.A(n_1145),
.Y(n_1337)
);

AND2x4_ASAP7_75t_L g1338 ( 
.A(n_1163),
.B(n_1233),
.Y(n_1338)
);

AOI21xp5_ASAP7_75t_L g1339 ( 
.A1(n_1181),
.A2(n_1218),
.B(n_1249),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_L g1340 ( 
.A(n_1208),
.B(n_1189),
.Y(n_1340)
);

NAND2xp5_ASAP7_75t_L g1341 ( 
.A(n_1208),
.B(n_1212),
.Y(n_1341)
);

BUFx2_ASAP7_75t_L g1342 ( 
.A(n_1254),
.Y(n_1342)
);

CKINVDCx5p33_ASAP7_75t_R g1343 ( 
.A(n_1244),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_L g1344 ( 
.A(n_1212),
.B(n_1135),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_L g1345 ( 
.A(n_1212),
.B(n_1135),
.Y(n_1345)
);

NOR2xp33_ASAP7_75t_L g1346 ( 
.A(n_1179),
.B(n_1180),
.Y(n_1346)
);

OA21x2_ASAP7_75t_L g1347 ( 
.A1(n_1120),
.A2(n_1134),
.B(n_1122),
.Y(n_1347)
);

BUFx6f_ASAP7_75t_L g1348 ( 
.A(n_1143),
.Y(n_1348)
);

AOI21xp5_ASAP7_75t_L g1349 ( 
.A1(n_1125),
.A2(n_1187),
.B(n_1130),
.Y(n_1349)
);

OAI21xp33_ASAP7_75t_L g1350 ( 
.A1(n_1194),
.A2(n_1158),
.B(n_1150),
.Y(n_1350)
);

AND2x4_ASAP7_75t_L g1351 ( 
.A(n_1244),
.B(n_1155),
.Y(n_1351)
);

NAND2xp33_ASAP7_75t_L g1352 ( 
.A(n_1184),
.B(n_1234),
.Y(n_1352)
);

INVx3_ASAP7_75t_L g1353 ( 
.A(n_1115),
.Y(n_1353)
);

AOI22xp33_ASAP7_75t_L g1354 ( 
.A1(n_1212),
.A2(n_1202),
.B1(n_1186),
.B2(n_1155),
.Y(n_1354)
);

BUFx6f_ASAP7_75t_L g1355 ( 
.A(n_1154),
.Y(n_1355)
);

AOI21xp5_ASAP7_75t_L g1356 ( 
.A1(n_1202),
.A2(n_1153),
.B(n_1182),
.Y(n_1356)
);

O2A1O1Ixp5_ASAP7_75t_SL g1357 ( 
.A1(n_1113),
.A2(n_1135),
.B(n_1105),
.C(n_1119),
.Y(n_1357)
);

CKINVDCx20_ASAP7_75t_R g1358 ( 
.A(n_1184),
.Y(n_1358)
);

AOI22xp33_ASAP7_75t_L g1359 ( 
.A1(n_1184),
.A2(n_1160),
.B1(n_1144),
.B2(n_1114),
.Y(n_1359)
);

BUFx2_ASAP7_75t_L g1360 ( 
.A(n_1190),
.Y(n_1360)
);

AOI21xp5_ASAP7_75t_L g1361 ( 
.A1(n_1104),
.A2(n_1258),
.B(n_1252),
.Y(n_1361)
);

INVx3_ASAP7_75t_L g1362 ( 
.A(n_1184),
.Y(n_1362)
);

AOI21xp5_ASAP7_75t_L g1363 ( 
.A1(n_1237),
.A2(n_1126),
.B(n_1184),
.Y(n_1363)
);

AOI21xp5_ASAP7_75t_L g1364 ( 
.A1(n_1119),
.A2(n_1193),
.B(n_1190),
.Y(n_1364)
);

OAI22xp5_ASAP7_75t_L g1365 ( 
.A1(n_1112),
.A2(n_1100),
.B1(n_1102),
.B2(n_1099),
.Y(n_1365)
);

AND2x4_ASAP7_75t_L g1366 ( 
.A(n_1219),
.B(n_1227),
.Y(n_1366)
);

BUFx4f_ASAP7_75t_L g1367 ( 
.A(n_1195),
.Y(n_1367)
);

AND2x4_ASAP7_75t_L g1368 ( 
.A(n_1219),
.B(n_1227),
.Y(n_1368)
);

CKINVDCx20_ASAP7_75t_R g1369 ( 
.A(n_1241),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1201),
.B(n_1239),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1139),
.Y(n_1371)
);

AND2x2_ASAP7_75t_L g1372 ( 
.A(n_1203),
.B(n_943),
.Y(n_1372)
);

OAI21xp5_ASAP7_75t_L g1373 ( 
.A1(n_1141),
.A2(n_1255),
.B(n_1206),
.Y(n_1373)
);

AND2x2_ASAP7_75t_L g1374 ( 
.A(n_1203),
.B(n_943),
.Y(n_1374)
);

AOI21xp5_ASAP7_75t_L g1375 ( 
.A1(n_1133),
.A2(n_1110),
.B(n_1147),
.Y(n_1375)
);

AOI21xp5_ASAP7_75t_L g1376 ( 
.A1(n_1133),
.A2(n_1110),
.B(n_1147),
.Y(n_1376)
);

INVx2_ASAP7_75t_L g1377 ( 
.A(n_1131),
.Y(n_1377)
);

AOI22xp5_ASAP7_75t_L g1378 ( 
.A1(n_1111),
.A2(n_1099),
.B1(n_1102),
.B2(n_1100),
.Y(n_1378)
);

AOI22xp5_ASAP7_75t_L g1379 ( 
.A1(n_1111),
.A2(n_1099),
.B1(n_1102),
.B2(n_1100),
.Y(n_1379)
);

BUFx6f_ASAP7_75t_L g1380 ( 
.A(n_1165),
.Y(n_1380)
);

AOI21xp5_ASAP7_75t_L g1381 ( 
.A1(n_1133),
.A2(n_1110),
.B(n_1147),
.Y(n_1381)
);

AOI21x1_ASAP7_75t_L g1382 ( 
.A1(n_1149),
.A2(n_1136),
.B(n_1113),
.Y(n_1382)
);

AND2x4_ASAP7_75t_L g1383 ( 
.A(n_1219),
.B(n_1227),
.Y(n_1383)
);

O2A1O1Ixp33_ASAP7_75t_L g1384 ( 
.A1(n_1161),
.A2(n_1101),
.B(n_924),
.C(n_973),
.Y(n_1384)
);

NAND2x1p5_ASAP7_75t_L g1385 ( 
.A(n_1165),
.B(n_1219),
.Y(n_1385)
);

AOI21xp5_ASAP7_75t_L g1386 ( 
.A1(n_1133),
.A2(n_1110),
.B(n_1147),
.Y(n_1386)
);

AND2x4_ASAP7_75t_L g1387 ( 
.A(n_1219),
.B(n_1227),
.Y(n_1387)
);

OAI22xp33_ASAP7_75t_L g1388 ( 
.A1(n_1213),
.A2(n_924),
.B1(n_1101),
.B2(n_973),
.Y(n_1388)
);

INVx3_ASAP7_75t_L g1389 ( 
.A(n_1142),
.Y(n_1389)
);

NAND2xp5_ASAP7_75t_L g1390 ( 
.A(n_1213),
.B(n_1214),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_1213),
.B(n_1214),
.Y(n_1391)
);

BUFx2_ASAP7_75t_L g1392 ( 
.A(n_1224),
.Y(n_1392)
);

BUFx2_ASAP7_75t_L g1393 ( 
.A(n_1224),
.Y(n_1393)
);

AND2x4_ASAP7_75t_L g1394 ( 
.A(n_1219),
.B(n_1227),
.Y(n_1394)
);

CKINVDCx11_ASAP7_75t_R g1395 ( 
.A(n_1118),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1139),
.Y(n_1396)
);

AND2x2_ASAP7_75t_L g1397 ( 
.A(n_1203),
.B(n_943),
.Y(n_1397)
);

AOI21xp5_ASAP7_75t_L g1398 ( 
.A1(n_1133),
.A2(n_1110),
.B(n_1147),
.Y(n_1398)
);

BUFx6f_ASAP7_75t_L g1399 ( 
.A(n_1165),
.Y(n_1399)
);

HB1xp67_ASAP7_75t_L g1400 ( 
.A(n_1232),
.Y(n_1400)
);

AND2x2_ASAP7_75t_L g1401 ( 
.A(n_1203),
.B(n_943),
.Y(n_1401)
);

INVx3_ASAP7_75t_L g1402 ( 
.A(n_1142),
.Y(n_1402)
);

AOI21x1_ASAP7_75t_L g1403 ( 
.A1(n_1149),
.A2(n_1136),
.B(n_1113),
.Y(n_1403)
);

AND2x4_ASAP7_75t_L g1404 ( 
.A(n_1219),
.B(n_1227),
.Y(n_1404)
);

INVx5_ASAP7_75t_L g1405 ( 
.A(n_1165),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_L g1406 ( 
.A(n_1201),
.B(n_1239),
.Y(n_1406)
);

BUFx2_ASAP7_75t_L g1407 ( 
.A(n_1224),
.Y(n_1407)
);

OAI21x1_ASAP7_75t_SL g1408 ( 
.A1(n_1124),
.A2(n_1222),
.B(n_1193),
.Y(n_1408)
);

NOR2xp33_ASAP7_75t_L g1409 ( 
.A(n_1370),
.B(n_1406),
.Y(n_1409)
);

INVx6_ASAP7_75t_L g1410 ( 
.A(n_1264),
.Y(n_1410)
);

INVx2_ASAP7_75t_L g1411 ( 
.A(n_1297),
.Y(n_1411)
);

NAND2x1p5_ASAP7_75t_L g1412 ( 
.A(n_1264),
.B(n_1405),
.Y(n_1412)
);

BUFx6f_ASAP7_75t_L g1413 ( 
.A(n_1268),
.Y(n_1413)
);

BUFx6f_ASAP7_75t_L g1414 ( 
.A(n_1268),
.Y(n_1414)
);

AOI22xp33_ASAP7_75t_L g1415 ( 
.A1(n_1365),
.A2(n_1266),
.B1(n_1379),
.B2(n_1378),
.Y(n_1415)
);

AOI22xp33_ASAP7_75t_SL g1416 ( 
.A1(n_1365),
.A2(n_1266),
.B1(n_1316),
.B2(n_1263),
.Y(n_1416)
);

INVx2_ASAP7_75t_SL g1417 ( 
.A(n_1291),
.Y(n_1417)
);

INVx2_ASAP7_75t_L g1418 ( 
.A(n_1371),
.Y(n_1418)
);

NAND2x1p5_ASAP7_75t_L g1419 ( 
.A(n_1264),
.B(n_1405),
.Y(n_1419)
);

AOI22xp33_ASAP7_75t_L g1420 ( 
.A1(n_1378),
.A2(n_1379),
.B1(n_1373),
.B2(n_1263),
.Y(n_1420)
);

OAI22xp33_ASAP7_75t_L g1421 ( 
.A1(n_1275),
.A2(n_1390),
.B1(n_1391),
.B2(n_1267),
.Y(n_1421)
);

HB1xp67_ASAP7_75t_L g1422 ( 
.A(n_1269),
.Y(n_1422)
);

BUFx4f_ASAP7_75t_L g1423 ( 
.A(n_1301),
.Y(n_1423)
);

OAI22xp5_ASAP7_75t_L g1424 ( 
.A1(n_1260),
.A2(n_1275),
.B1(n_1390),
.B2(n_1391),
.Y(n_1424)
);

INVx11_ASAP7_75t_L g1425 ( 
.A(n_1291),
.Y(n_1425)
);

BUFx2_ASAP7_75t_L g1426 ( 
.A(n_1392),
.Y(n_1426)
);

OAI21x1_ASAP7_75t_L g1427 ( 
.A1(n_1289),
.A2(n_1363),
.B(n_1356),
.Y(n_1427)
);

CKINVDCx8_ASAP7_75t_R g1428 ( 
.A(n_1284),
.Y(n_1428)
);

OAI22xp5_ASAP7_75t_L g1429 ( 
.A1(n_1283),
.A2(n_1296),
.B1(n_1313),
.B2(n_1340),
.Y(n_1429)
);

AO21x2_ASAP7_75t_L g1430 ( 
.A1(n_1339),
.A2(n_1361),
.B(n_1349),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1396),
.Y(n_1431)
);

NAND2x1p5_ASAP7_75t_L g1432 ( 
.A(n_1405),
.B(n_1338),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1302),
.Y(n_1433)
);

INVx4_ASAP7_75t_L g1434 ( 
.A(n_1265),
.Y(n_1434)
);

BUFx2_ASAP7_75t_SL g1435 ( 
.A(n_1325),
.Y(n_1435)
);

OAI22xp33_ASAP7_75t_L g1436 ( 
.A1(n_1282),
.A2(n_1373),
.B1(n_1310),
.B2(n_1315),
.Y(n_1436)
);

BUFx2_ASAP7_75t_L g1437 ( 
.A(n_1393),
.Y(n_1437)
);

AND2x4_ASAP7_75t_L g1438 ( 
.A(n_1287),
.B(n_1293),
.Y(n_1438)
);

OAI21x1_ASAP7_75t_L g1439 ( 
.A1(n_1273),
.A2(n_1279),
.B(n_1382),
.Y(n_1439)
);

BUFx3_ASAP7_75t_L g1440 ( 
.A(n_1367),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1309),
.Y(n_1441)
);

AOI22xp33_ASAP7_75t_L g1442 ( 
.A1(n_1259),
.A2(n_1316),
.B1(n_1312),
.B2(n_1388),
.Y(n_1442)
);

AOI21x1_ASAP7_75t_L g1443 ( 
.A1(n_1280),
.A2(n_1403),
.B(n_1321),
.Y(n_1443)
);

OAI22xp5_ASAP7_75t_SL g1444 ( 
.A1(n_1330),
.A2(n_1335),
.B1(n_1270),
.B2(n_1277),
.Y(n_1444)
);

AOI22xp33_ASAP7_75t_L g1445 ( 
.A1(n_1310),
.A2(n_1315),
.B1(n_1314),
.B2(n_1319),
.Y(n_1445)
);

AOI21xp5_ASAP7_75t_L g1446 ( 
.A1(n_1262),
.A2(n_1376),
.B(n_1398),
.Y(n_1446)
);

BUFx3_ASAP7_75t_L g1447 ( 
.A(n_1367),
.Y(n_1447)
);

INVxp67_ASAP7_75t_L g1448 ( 
.A(n_1400),
.Y(n_1448)
);

HB1xp67_ASAP7_75t_L g1449 ( 
.A(n_1407),
.Y(n_1449)
);

INVx2_ASAP7_75t_L g1450 ( 
.A(n_1377),
.Y(n_1450)
);

AOI22xp33_ASAP7_75t_L g1451 ( 
.A1(n_1314),
.A2(n_1319),
.B1(n_1282),
.B2(n_1274),
.Y(n_1451)
);

AOI22xp33_ASAP7_75t_L g1452 ( 
.A1(n_1292),
.A2(n_1304),
.B1(n_1299),
.B2(n_1401),
.Y(n_1452)
);

CKINVDCx5p33_ASAP7_75t_R g1453 ( 
.A(n_1272),
.Y(n_1453)
);

BUFx6f_ASAP7_75t_L g1454 ( 
.A(n_1301),
.Y(n_1454)
);

AOI22xp33_ASAP7_75t_L g1455 ( 
.A1(n_1292),
.A2(n_1397),
.B1(n_1374),
.B2(n_1372),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1298),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1288),
.Y(n_1457)
);

HB1xp67_ASAP7_75t_L g1458 ( 
.A(n_1306),
.Y(n_1458)
);

AOI22xp33_ASAP7_75t_SL g1459 ( 
.A1(n_1295),
.A2(n_1342),
.B1(n_1336),
.B2(n_1358),
.Y(n_1459)
);

OAI22xp5_ASAP7_75t_L g1460 ( 
.A1(n_1341),
.A2(n_1276),
.B1(n_1305),
.B2(n_1335),
.Y(n_1460)
);

BUFx12f_ASAP7_75t_L g1461 ( 
.A(n_1395),
.Y(n_1461)
);

HB1xp67_ASAP7_75t_SL g1462 ( 
.A(n_1343),
.Y(n_1462)
);

OAI22xp5_ASAP7_75t_L g1463 ( 
.A1(n_1305),
.A2(n_1271),
.B1(n_1384),
.B2(n_1354),
.Y(n_1463)
);

OAI21xp5_ASAP7_75t_L g1464 ( 
.A1(n_1326),
.A2(n_1318),
.B(n_1386),
.Y(n_1464)
);

AOI22xp33_ASAP7_75t_L g1465 ( 
.A1(n_1323),
.A2(n_1320),
.B1(n_1350),
.B2(n_1307),
.Y(n_1465)
);

NAND2x1p5_ASAP7_75t_L g1466 ( 
.A(n_1293),
.B(n_1402),
.Y(n_1466)
);

AND2x2_ASAP7_75t_L g1467 ( 
.A(n_1366),
.B(n_1387),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1332),
.Y(n_1468)
);

OA21x2_ASAP7_75t_L g1469 ( 
.A1(n_1364),
.A2(n_1381),
.B(n_1375),
.Y(n_1469)
);

AOI22xp33_ASAP7_75t_L g1470 ( 
.A1(n_1320),
.A2(n_1350),
.B1(n_1308),
.B2(n_1328),
.Y(n_1470)
);

CKINVDCx11_ASAP7_75t_R g1471 ( 
.A(n_1369),
.Y(n_1471)
);

HB1xp67_ASAP7_75t_L g1472 ( 
.A(n_1290),
.Y(n_1472)
);

BUFx8_ASAP7_75t_L g1473 ( 
.A(n_1281),
.Y(n_1473)
);

BUFx2_ASAP7_75t_L g1474 ( 
.A(n_1324),
.Y(n_1474)
);

OAI21xp33_ASAP7_75t_L g1475 ( 
.A1(n_1344),
.A2(n_1345),
.B(n_1346),
.Y(n_1475)
);

INVxp67_ASAP7_75t_SL g1476 ( 
.A(n_1337),
.Y(n_1476)
);

INVxp67_ASAP7_75t_L g1477 ( 
.A(n_1327),
.Y(n_1477)
);

BUFx3_ASAP7_75t_L g1478 ( 
.A(n_1366),
.Y(n_1478)
);

OAI22xp5_ASAP7_75t_L g1479 ( 
.A1(n_1300),
.A2(n_1285),
.B1(n_1345),
.B2(n_1334),
.Y(n_1479)
);

AND2x2_ASAP7_75t_L g1480 ( 
.A(n_1368),
.B(n_1394),
.Y(n_1480)
);

AOI22xp33_ASAP7_75t_L g1481 ( 
.A1(n_1360),
.A2(n_1408),
.B1(n_1368),
.B2(n_1383),
.Y(n_1481)
);

INVx8_ASAP7_75t_L g1482 ( 
.A(n_1286),
.Y(n_1482)
);

AOI22xp33_ASAP7_75t_SL g1483 ( 
.A1(n_1278),
.A2(n_1351),
.B1(n_1317),
.B2(n_1387),
.Y(n_1483)
);

OR2x6_ASAP7_75t_L g1484 ( 
.A(n_1294),
.B(n_1389),
.Y(n_1484)
);

OA21x2_ASAP7_75t_L g1485 ( 
.A1(n_1359),
.A2(n_1357),
.B(n_1347),
.Y(n_1485)
);

INVx2_ASAP7_75t_SL g1486 ( 
.A(n_1380),
.Y(n_1486)
);

INVxp33_ASAP7_75t_L g1487 ( 
.A(n_1383),
.Y(n_1487)
);

BUFx12f_ASAP7_75t_L g1488 ( 
.A(n_1380),
.Y(n_1488)
);

OA21x2_ASAP7_75t_L g1489 ( 
.A1(n_1355),
.A2(n_1334),
.B(n_1333),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1303),
.Y(n_1490)
);

CKINVDCx20_ASAP7_75t_R g1491 ( 
.A(n_1322),
.Y(n_1491)
);

INVx2_ASAP7_75t_L g1492 ( 
.A(n_1311),
.Y(n_1492)
);

OAI22xp5_ASAP7_75t_L g1493 ( 
.A1(n_1385),
.A2(n_1404),
.B1(n_1394),
.B2(n_1348),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1303),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1303),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1329),
.Y(n_1496)
);

OAI21x1_ASAP7_75t_L g1497 ( 
.A1(n_1362),
.A2(n_1294),
.B(n_1402),
.Y(n_1497)
);

BUFx12f_ASAP7_75t_L g1498 ( 
.A(n_1399),
.Y(n_1498)
);

BUFx3_ASAP7_75t_L g1499 ( 
.A(n_1404),
.Y(n_1499)
);

INVxp67_ASAP7_75t_L g1500 ( 
.A(n_1331),
.Y(n_1500)
);

INVx2_ASAP7_75t_L g1501 ( 
.A(n_1355),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1353),
.Y(n_1502)
);

HB1xp67_ASAP7_75t_L g1503 ( 
.A(n_1399),
.Y(n_1503)
);

INVx1_ASAP7_75t_SL g1504 ( 
.A(n_1322),
.Y(n_1504)
);

AOI22xp5_ASAP7_75t_SL g1505 ( 
.A1(n_1286),
.A2(n_1348),
.B1(n_1399),
.B2(n_1353),
.Y(n_1505)
);

AOI21x1_ASAP7_75t_L g1506 ( 
.A1(n_1355),
.A2(n_1352),
.B(n_1362),
.Y(n_1506)
);

AOI22xp33_ASAP7_75t_L g1507 ( 
.A1(n_1286),
.A2(n_1365),
.B1(n_1101),
.B2(n_924),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1348),
.Y(n_1508)
);

INVxp67_ASAP7_75t_L g1509 ( 
.A(n_1269),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1261),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1261),
.Y(n_1511)
);

BUFx3_ASAP7_75t_L g1512 ( 
.A(n_1264),
.Y(n_1512)
);

OR2x2_ASAP7_75t_L g1513 ( 
.A(n_1295),
.B(n_1274),
.Y(n_1513)
);

CKINVDCx11_ASAP7_75t_R g1514 ( 
.A(n_1272),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1261),
.Y(n_1515)
);

NAND2xp5_ASAP7_75t_L g1516 ( 
.A(n_1370),
.B(n_1201),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1261),
.Y(n_1517)
);

BUFx6f_ASAP7_75t_L g1518 ( 
.A(n_1268),
.Y(n_1518)
);

AOI22xp33_ASAP7_75t_L g1519 ( 
.A1(n_1365),
.A2(n_1101),
.B1(n_924),
.B2(n_1112),
.Y(n_1519)
);

INVx2_ASAP7_75t_SL g1520 ( 
.A(n_1291),
.Y(n_1520)
);

BUFx3_ASAP7_75t_L g1521 ( 
.A(n_1264),
.Y(n_1521)
);

CKINVDCx14_ASAP7_75t_R g1522 ( 
.A(n_1278),
.Y(n_1522)
);

AOI22xp33_ASAP7_75t_L g1523 ( 
.A1(n_1365),
.A2(n_1101),
.B1(n_924),
.B2(n_1112),
.Y(n_1523)
);

AOI22xp33_ASAP7_75t_L g1524 ( 
.A1(n_1365),
.A2(n_1101),
.B1(n_924),
.B2(n_1112),
.Y(n_1524)
);

AOI22xp33_ASAP7_75t_SL g1525 ( 
.A1(n_1365),
.A2(n_1100),
.B1(n_1102),
.B2(n_1099),
.Y(n_1525)
);

HB1xp67_ASAP7_75t_L g1526 ( 
.A(n_1269),
.Y(n_1526)
);

AND2x2_ASAP7_75t_L g1527 ( 
.A(n_1372),
.B(n_1374),
.Y(n_1527)
);

AOI22xp33_ASAP7_75t_SL g1528 ( 
.A1(n_1365),
.A2(n_1100),
.B1(n_1102),
.B2(n_1099),
.Y(n_1528)
);

BUFx8_ASAP7_75t_L g1529 ( 
.A(n_1392),
.Y(n_1529)
);

AOI22xp33_ASAP7_75t_L g1530 ( 
.A1(n_1365),
.A2(n_1101),
.B1(n_924),
.B2(n_1112),
.Y(n_1530)
);

INVx3_ASAP7_75t_L g1531 ( 
.A(n_1265),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_L g1532 ( 
.A(n_1370),
.B(n_1201),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1261),
.Y(n_1533)
);

AND2x2_ASAP7_75t_L g1534 ( 
.A(n_1372),
.B(n_1374),
.Y(n_1534)
);

INVx8_ASAP7_75t_L g1535 ( 
.A(n_1264),
.Y(n_1535)
);

AND2x2_ASAP7_75t_L g1536 ( 
.A(n_1372),
.B(n_1374),
.Y(n_1536)
);

CKINVDCx11_ASAP7_75t_R g1537 ( 
.A(n_1272),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1261),
.Y(n_1538)
);

BUFx3_ASAP7_75t_L g1539 ( 
.A(n_1264),
.Y(n_1539)
);

AOI21x1_ASAP7_75t_L g1540 ( 
.A1(n_1363),
.A2(n_1149),
.B(n_1356),
.Y(n_1540)
);

OAI22xp33_ASAP7_75t_L g1541 ( 
.A1(n_1370),
.A2(n_1099),
.B1(n_1102),
.B2(n_1100),
.Y(n_1541)
);

AOI22xp33_ASAP7_75t_L g1542 ( 
.A1(n_1365),
.A2(n_1101),
.B1(n_924),
.B2(n_1112),
.Y(n_1542)
);

INVx2_ASAP7_75t_SL g1543 ( 
.A(n_1291),
.Y(n_1543)
);

AND2x2_ASAP7_75t_L g1544 ( 
.A(n_1416),
.B(n_1445),
.Y(n_1544)
);

OAI21x1_ASAP7_75t_L g1545 ( 
.A1(n_1427),
.A2(n_1540),
.B(n_1443),
.Y(n_1545)
);

AOI21x1_ASAP7_75t_L g1546 ( 
.A1(n_1446),
.A2(n_1429),
.B(n_1506),
.Y(n_1546)
);

HB1xp67_ASAP7_75t_L g1547 ( 
.A(n_1422),
.Y(n_1547)
);

OR2x2_ASAP7_75t_L g1548 ( 
.A(n_1445),
.B(n_1451),
.Y(n_1548)
);

INVxp67_ASAP7_75t_L g1549 ( 
.A(n_1472),
.Y(n_1549)
);

BUFx2_ASAP7_75t_L g1550 ( 
.A(n_1457),
.Y(n_1550)
);

AOI222xp33_ASAP7_75t_L g1551 ( 
.A1(n_1415),
.A2(n_1420),
.B1(n_1542),
.B2(n_1523),
.C1(n_1524),
.C2(n_1519),
.Y(n_1551)
);

NAND3xp33_ASAP7_75t_L g1552 ( 
.A(n_1519),
.B(n_1524),
.C(n_1523),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1411),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1424),
.B(n_1409),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1418),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1409),
.B(n_1516),
.Y(n_1556)
);

HB1xp67_ASAP7_75t_L g1557 ( 
.A(n_1526),
.Y(n_1557)
);

OAI21x1_ASAP7_75t_L g1558 ( 
.A1(n_1439),
.A2(n_1464),
.B(n_1497),
.Y(n_1558)
);

OR2x6_ASAP7_75t_L g1559 ( 
.A(n_1439),
.B(n_1482),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1525),
.B(n_1528),
.Y(n_1560)
);

BUFx2_ASAP7_75t_L g1561 ( 
.A(n_1489),
.Y(n_1561)
);

INVx8_ASAP7_75t_L g1562 ( 
.A(n_1482),
.Y(n_1562)
);

INVx4_ASAP7_75t_SL g1563 ( 
.A(n_1484),
.Y(n_1563)
);

OR2x2_ASAP7_75t_L g1564 ( 
.A(n_1451),
.B(n_1475),
.Y(n_1564)
);

OA21x2_ASAP7_75t_L g1565 ( 
.A1(n_1470),
.A2(n_1442),
.B(n_1415),
.Y(n_1565)
);

INVxp67_ASAP7_75t_L g1566 ( 
.A(n_1458),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1420),
.B(n_1452),
.Y(n_1567)
);

INVx2_ASAP7_75t_SL g1568 ( 
.A(n_1410),
.Y(n_1568)
);

OAI21x1_ASAP7_75t_L g1569 ( 
.A1(n_1469),
.A2(n_1501),
.B(n_1485),
.Y(n_1569)
);

BUFx2_ASAP7_75t_L g1570 ( 
.A(n_1489),
.Y(n_1570)
);

HB1xp67_ASAP7_75t_L g1571 ( 
.A(n_1449),
.Y(n_1571)
);

AOI22xp5_ASAP7_75t_L g1572 ( 
.A1(n_1530),
.A2(n_1542),
.B1(n_1541),
.B2(n_1532),
.Y(n_1572)
);

CKINVDCx14_ASAP7_75t_R g1573 ( 
.A(n_1522),
.Y(n_1573)
);

BUFx3_ASAP7_75t_L g1574 ( 
.A(n_1529),
.Y(n_1574)
);

INVx3_ASAP7_75t_L g1575 ( 
.A(n_1489),
.Y(n_1575)
);

HB1xp67_ASAP7_75t_L g1576 ( 
.A(n_1513),
.Y(n_1576)
);

AO31x2_ASAP7_75t_L g1577 ( 
.A1(n_1463),
.A2(n_1460),
.A3(n_1515),
.B(n_1538),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1431),
.Y(n_1578)
);

OAI21x1_ASAP7_75t_L g1579 ( 
.A1(n_1469),
.A2(n_1485),
.B(n_1481),
.Y(n_1579)
);

INVx2_ASAP7_75t_L g1580 ( 
.A(n_1510),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1452),
.B(n_1470),
.Y(n_1581)
);

AND2x2_ASAP7_75t_L g1582 ( 
.A(n_1455),
.B(n_1465),
.Y(n_1582)
);

INVx2_ASAP7_75t_L g1583 ( 
.A(n_1511),
.Y(n_1583)
);

INVxp67_ASAP7_75t_SL g1584 ( 
.A(n_1421),
.Y(n_1584)
);

OR2x2_ASAP7_75t_L g1585 ( 
.A(n_1436),
.B(n_1455),
.Y(n_1585)
);

OR2x2_ASAP7_75t_L g1586 ( 
.A(n_1436),
.B(n_1465),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1442),
.B(n_1527),
.Y(n_1587)
);

HB1xp67_ASAP7_75t_L g1588 ( 
.A(n_1456),
.Y(n_1588)
);

INVx2_ASAP7_75t_L g1589 ( 
.A(n_1517),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1533),
.Y(n_1590)
);

BUFx3_ASAP7_75t_L g1591 ( 
.A(n_1529),
.Y(n_1591)
);

OA21x2_ASAP7_75t_L g1592 ( 
.A1(n_1530),
.A2(n_1507),
.B(n_1481),
.Y(n_1592)
);

OR2x2_ASAP7_75t_L g1593 ( 
.A(n_1421),
.B(n_1469),
.Y(n_1593)
);

INVx3_ASAP7_75t_L g1594 ( 
.A(n_1438),
.Y(n_1594)
);

INVx2_ASAP7_75t_L g1595 ( 
.A(n_1441),
.Y(n_1595)
);

AO21x2_ASAP7_75t_L g1596 ( 
.A1(n_1430),
.A2(n_1541),
.B(n_1502),
.Y(n_1596)
);

INVx3_ASAP7_75t_L g1597 ( 
.A(n_1438),
.Y(n_1597)
);

INVxp33_ASAP7_75t_L g1598 ( 
.A(n_1534),
.Y(n_1598)
);

HB1xp67_ASAP7_75t_L g1599 ( 
.A(n_1448),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1485),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1433),
.Y(n_1601)
);

BUFx2_ASAP7_75t_L g1602 ( 
.A(n_1476),
.Y(n_1602)
);

BUFx3_ASAP7_75t_L g1603 ( 
.A(n_1529),
.Y(n_1603)
);

OAI21x1_ASAP7_75t_L g1604 ( 
.A1(n_1479),
.A2(n_1507),
.B(n_1466),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1430),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1468),
.Y(n_1606)
);

HB1xp67_ASAP7_75t_L g1607 ( 
.A(n_1509),
.Y(n_1607)
);

HB1xp67_ASAP7_75t_L g1608 ( 
.A(n_1474),
.Y(n_1608)
);

HB1xp67_ASAP7_75t_L g1609 ( 
.A(n_1426),
.Y(n_1609)
);

AND2x2_ASAP7_75t_L g1610 ( 
.A(n_1536),
.B(n_1450),
.Y(n_1610)
);

NAND2x1p5_ASAP7_75t_L g1611 ( 
.A(n_1505),
.B(n_1438),
.Y(n_1611)
);

AOI222xp33_ASAP7_75t_L g1612 ( 
.A1(n_1444),
.A2(n_1461),
.B1(n_1437),
.B2(n_1477),
.C1(n_1473),
.C2(n_1423),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1459),
.B(n_1487),
.Y(n_1613)
);

HB1xp67_ASAP7_75t_L g1614 ( 
.A(n_1503),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_L g1615 ( 
.A(n_1487),
.B(n_1467),
.Y(n_1615)
);

INVx2_ASAP7_75t_L g1616 ( 
.A(n_1492),
.Y(n_1616)
);

OR2x2_ASAP7_75t_L g1617 ( 
.A(n_1484),
.B(n_1432),
.Y(n_1617)
);

OA21x2_ASAP7_75t_L g1618 ( 
.A1(n_1490),
.A2(n_1496),
.B(n_1494),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1495),
.Y(n_1619)
);

INVx2_ASAP7_75t_L g1620 ( 
.A(n_1508),
.Y(n_1620)
);

CKINVDCx5p33_ASAP7_75t_R g1621 ( 
.A(n_1471),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1482),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1412),
.Y(n_1623)
);

OAI21x1_ASAP7_75t_L g1624 ( 
.A1(n_1419),
.A2(n_1493),
.B(n_1531),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1410),
.Y(n_1625)
);

HB1xp67_ASAP7_75t_L g1626 ( 
.A(n_1512),
.Y(n_1626)
);

AO21x2_ASAP7_75t_L g1627 ( 
.A1(n_1500),
.A2(n_1480),
.B(n_1410),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1512),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1521),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1521),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1539),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1539),
.Y(n_1632)
);

OAI21x1_ASAP7_75t_L g1633 ( 
.A1(n_1535),
.A2(n_1423),
.B(n_1434),
.Y(n_1633)
);

OR2x2_ASAP7_75t_L g1634 ( 
.A(n_1478),
.B(n_1499),
.Y(n_1634)
);

AND2x4_ASAP7_75t_L g1635 ( 
.A(n_1440),
.B(n_1447),
.Y(n_1635)
);

INVx2_ASAP7_75t_SL g1636 ( 
.A(n_1488),
.Y(n_1636)
);

AND2x2_ASAP7_75t_L g1637 ( 
.A(n_1561),
.B(n_1413),
.Y(n_1637)
);

AND2x2_ASAP7_75t_L g1638 ( 
.A(n_1561),
.B(n_1413),
.Y(n_1638)
);

AND2x4_ASAP7_75t_L g1639 ( 
.A(n_1559),
.B(n_1447),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_L g1640 ( 
.A(n_1554),
.B(n_1486),
.Y(n_1640)
);

NOR2xp33_ASAP7_75t_L g1641 ( 
.A(n_1556),
.B(n_1453),
.Y(n_1641)
);

AND2x2_ASAP7_75t_L g1642 ( 
.A(n_1570),
.B(n_1414),
.Y(n_1642)
);

INVx3_ASAP7_75t_L g1643 ( 
.A(n_1575),
.Y(n_1643)
);

AND2x2_ASAP7_75t_L g1644 ( 
.A(n_1578),
.B(n_1414),
.Y(n_1644)
);

AND2x2_ASAP7_75t_L g1645 ( 
.A(n_1590),
.B(n_1414),
.Y(n_1645)
);

INVxp67_ASAP7_75t_L g1646 ( 
.A(n_1618),
.Y(n_1646)
);

BUFx3_ASAP7_75t_L g1647 ( 
.A(n_1627),
.Y(n_1647)
);

BUFx2_ASAP7_75t_L g1648 ( 
.A(n_1627),
.Y(n_1648)
);

BUFx2_ASAP7_75t_L g1649 ( 
.A(n_1627),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_L g1650 ( 
.A(n_1584),
.B(n_1483),
.Y(n_1650)
);

BUFx8_ASAP7_75t_SL g1651 ( 
.A(n_1621),
.Y(n_1651)
);

AOI22xp33_ASAP7_75t_L g1652 ( 
.A1(n_1552),
.A2(n_1518),
.B1(n_1454),
.B2(n_1417),
.Y(n_1652)
);

OR2x2_ASAP7_75t_L g1653 ( 
.A(n_1593),
.B(n_1543),
.Y(n_1653)
);

OR2x2_ASAP7_75t_L g1654 ( 
.A(n_1593),
.B(n_1520),
.Y(n_1654)
);

NOR2xp33_ASAP7_75t_L g1655 ( 
.A(n_1598),
.B(n_1453),
.Y(n_1655)
);

OAI221xp5_ASAP7_75t_L g1656 ( 
.A1(n_1552),
.A2(n_1572),
.B1(n_1551),
.B2(n_1586),
.C(n_1560),
.Y(n_1656)
);

AND2x2_ASAP7_75t_L g1657 ( 
.A(n_1596),
.B(n_1504),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1596),
.B(n_1435),
.Y(n_1658)
);

AND2x4_ASAP7_75t_L g1659 ( 
.A(n_1559),
.B(n_1491),
.Y(n_1659)
);

AND2x2_ASAP7_75t_L g1660 ( 
.A(n_1596),
.B(n_1498),
.Y(n_1660)
);

AND2x2_ASAP7_75t_L g1661 ( 
.A(n_1579),
.B(n_1569),
.Y(n_1661)
);

AND2x2_ASAP7_75t_L g1662 ( 
.A(n_1579),
.B(n_1491),
.Y(n_1662)
);

OAI21x1_ASAP7_75t_L g1663 ( 
.A1(n_1545),
.A2(n_1473),
.B(n_1425),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_L g1664 ( 
.A(n_1550),
.B(n_1428),
.Y(n_1664)
);

OR2x2_ASAP7_75t_L g1665 ( 
.A(n_1577),
.B(n_1462),
.Y(n_1665)
);

INVx3_ASAP7_75t_SL g1666 ( 
.A(n_1621),
.Y(n_1666)
);

INVx3_ASAP7_75t_L g1667 ( 
.A(n_1559),
.Y(n_1667)
);

OR2x2_ASAP7_75t_L g1668 ( 
.A(n_1577),
.B(n_1576),
.Y(n_1668)
);

BUFx6f_ASAP7_75t_L g1669 ( 
.A(n_1633),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_L g1670 ( 
.A(n_1572),
.B(n_1473),
.Y(n_1670)
);

HB1xp67_ASAP7_75t_L g1671 ( 
.A(n_1577),
.Y(n_1671)
);

AND2x2_ASAP7_75t_L g1672 ( 
.A(n_1580),
.B(n_1471),
.Y(n_1672)
);

NOR2xp33_ASAP7_75t_L g1673 ( 
.A(n_1615),
.B(n_1537),
.Y(n_1673)
);

HB1xp67_ASAP7_75t_L g1674 ( 
.A(n_1577),
.Y(n_1674)
);

OR2x2_ASAP7_75t_L g1675 ( 
.A(n_1577),
.B(n_1514),
.Y(n_1675)
);

AND2x2_ASAP7_75t_L g1676 ( 
.A(n_1583),
.B(n_1514),
.Y(n_1676)
);

AND2x2_ASAP7_75t_L g1677 ( 
.A(n_1583),
.B(n_1537),
.Y(n_1677)
);

HB1xp67_ASAP7_75t_L g1678 ( 
.A(n_1588),
.Y(n_1678)
);

BUFx2_ASAP7_75t_L g1679 ( 
.A(n_1602),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_L g1680 ( 
.A(n_1567),
.B(n_1461),
.Y(n_1680)
);

BUFx2_ASAP7_75t_L g1681 ( 
.A(n_1602),
.Y(n_1681)
);

NAND2xp5_ASAP7_75t_L g1682 ( 
.A(n_1567),
.B(n_1606),
.Y(n_1682)
);

NAND2xp5_ASAP7_75t_SL g1683 ( 
.A(n_1665),
.B(n_1564),
.Y(n_1683)
);

AND2x2_ASAP7_75t_L g1684 ( 
.A(n_1637),
.B(n_1618),
.Y(n_1684)
);

OAI21xp5_ASAP7_75t_L g1685 ( 
.A1(n_1656),
.A2(n_1560),
.B(n_1544),
.Y(n_1685)
);

AND2x2_ASAP7_75t_L g1686 ( 
.A(n_1637),
.B(n_1618),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_SL g1687 ( 
.A(n_1665),
.B(n_1564),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_L g1688 ( 
.A(n_1678),
.B(n_1547),
.Y(n_1688)
);

AOI21xp33_ASAP7_75t_L g1689 ( 
.A1(n_1675),
.A2(n_1586),
.B(n_1613),
.Y(n_1689)
);

AND2x2_ASAP7_75t_L g1690 ( 
.A(n_1637),
.B(n_1638),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_L g1691 ( 
.A(n_1682),
.B(n_1557),
.Y(n_1691)
);

AOI22xp33_ASAP7_75t_L g1692 ( 
.A1(n_1656),
.A2(n_1544),
.B1(n_1565),
.B2(n_1581),
.Y(n_1692)
);

OAI221xp5_ASAP7_75t_L g1693 ( 
.A1(n_1670),
.A2(n_1612),
.B1(n_1549),
.B2(n_1566),
.C(n_1548),
.Y(n_1693)
);

NAND2xp5_ASAP7_75t_SL g1694 ( 
.A(n_1675),
.B(n_1581),
.Y(n_1694)
);

NOR2xp33_ASAP7_75t_L g1695 ( 
.A(n_1641),
.B(n_1574),
.Y(n_1695)
);

NAND2xp5_ASAP7_75t_L g1696 ( 
.A(n_1640),
.B(n_1571),
.Y(n_1696)
);

AOI221xp5_ASAP7_75t_L g1697 ( 
.A1(n_1670),
.A2(n_1587),
.B1(n_1607),
.B2(n_1599),
.C(n_1608),
.Y(n_1697)
);

AND2x2_ASAP7_75t_L g1698 ( 
.A(n_1672),
.B(n_1609),
.Y(n_1698)
);

AND2x2_ASAP7_75t_L g1699 ( 
.A(n_1642),
.B(n_1592),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_SL g1700 ( 
.A(n_1680),
.B(n_1548),
.Y(n_1700)
);

NAND3xp33_ASAP7_75t_L g1701 ( 
.A(n_1658),
.B(n_1585),
.C(n_1565),
.Y(n_1701)
);

OAI22xp33_ASAP7_75t_SL g1702 ( 
.A1(n_1680),
.A2(n_1585),
.B1(n_1611),
.B2(n_1617),
.Y(n_1702)
);

AND2x2_ASAP7_75t_L g1703 ( 
.A(n_1642),
.B(n_1592),
.Y(n_1703)
);

OAI21xp5_ASAP7_75t_SL g1704 ( 
.A1(n_1652),
.A2(n_1582),
.B(n_1573),
.Y(n_1704)
);

OAI22xp5_ASAP7_75t_L g1705 ( 
.A1(n_1650),
.A2(n_1565),
.B1(n_1611),
.B2(n_1587),
.Y(n_1705)
);

NOR3xp33_ASAP7_75t_SL g1706 ( 
.A(n_1664),
.B(n_1650),
.C(n_1673),
.Y(n_1706)
);

AOI221xp5_ASAP7_75t_L g1707 ( 
.A1(n_1658),
.A2(n_1582),
.B1(n_1610),
.B2(n_1614),
.C(n_1601),
.Y(n_1707)
);

OAI21xp33_ASAP7_75t_L g1708 ( 
.A1(n_1658),
.A2(n_1610),
.B(n_1604),
.Y(n_1708)
);

OAI211xp5_ASAP7_75t_L g1709 ( 
.A1(n_1671),
.A2(n_1565),
.B(n_1601),
.C(n_1546),
.Y(n_1709)
);

OAI21xp33_ASAP7_75t_L g1710 ( 
.A1(n_1657),
.A2(n_1604),
.B(n_1616),
.Y(n_1710)
);

NOR2xp33_ASAP7_75t_L g1711 ( 
.A(n_1672),
.B(n_1574),
.Y(n_1711)
);

NAND3xp33_ASAP7_75t_L g1712 ( 
.A(n_1653),
.B(n_1616),
.C(n_1623),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_L g1713 ( 
.A(n_1644),
.B(n_1589),
.Y(n_1713)
);

AND2x2_ASAP7_75t_L g1714 ( 
.A(n_1662),
.B(n_1605),
.Y(n_1714)
);

AND2x2_ASAP7_75t_L g1715 ( 
.A(n_1662),
.B(n_1600),
.Y(n_1715)
);

OAI221xp5_ASAP7_75t_L g1716 ( 
.A1(n_1655),
.A2(n_1611),
.B1(n_1617),
.B2(n_1636),
.C(n_1634),
.Y(n_1716)
);

AND2x2_ASAP7_75t_L g1717 ( 
.A(n_1662),
.B(n_1595),
.Y(n_1717)
);

NAND3xp33_ASAP7_75t_L g1718 ( 
.A(n_1653),
.B(n_1623),
.C(n_1628),
.Y(n_1718)
);

AND2x2_ASAP7_75t_L g1719 ( 
.A(n_1657),
.B(n_1558),
.Y(n_1719)
);

NAND3xp33_ASAP7_75t_L g1720 ( 
.A(n_1654),
.B(n_1628),
.C(n_1632),
.Y(n_1720)
);

NAND2xp5_ASAP7_75t_SL g1721 ( 
.A(n_1676),
.B(n_1563),
.Y(n_1721)
);

AOI22xp33_ASAP7_75t_L g1722 ( 
.A1(n_1676),
.A2(n_1635),
.B1(n_1594),
.B2(n_1597),
.Y(n_1722)
);

NAND3xp33_ASAP7_75t_L g1723 ( 
.A(n_1654),
.B(n_1629),
.C(n_1631),
.Y(n_1723)
);

NOR2xp33_ASAP7_75t_R g1724 ( 
.A(n_1666),
.B(n_1591),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_L g1725 ( 
.A(n_1645),
.B(n_1553),
.Y(n_1725)
);

NAND3xp33_ASAP7_75t_L g1726 ( 
.A(n_1671),
.B(n_1629),
.C(n_1632),
.Y(n_1726)
);

OAI22xp5_ASAP7_75t_L g1727 ( 
.A1(n_1664),
.A2(n_1635),
.B1(n_1622),
.B2(n_1591),
.Y(n_1727)
);

HB1xp67_ASAP7_75t_L g1728 ( 
.A(n_1679),
.Y(n_1728)
);

NOR2xp33_ASAP7_75t_L g1729 ( 
.A(n_1677),
.B(n_1603),
.Y(n_1729)
);

OAI22xp5_ASAP7_75t_L g1730 ( 
.A1(n_1666),
.A2(n_1635),
.B1(n_1622),
.B2(n_1603),
.Y(n_1730)
);

NOR3xp33_ASAP7_75t_L g1731 ( 
.A(n_1660),
.B(n_1624),
.C(n_1625),
.Y(n_1731)
);

NAND4xp25_ASAP7_75t_L g1732 ( 
.A(n_1668),
.B(n_1619),
.C(n_1620),
.D(n_1555),
.Y(n_1732)
);

AND2x2_ASAP7_75t_L g1733 ( 
.A(n_1684),
.B(n_1661),
.Y(n_1733)
);

AND2x2_ASAP7_75t_L g1734 ( 
.A(n_1684),
.B(n_1661),
.Y(n_1734)
);

NAND2xp5_ASAP7_75t_L g1735 ( 
.A(n_1686),
.B(n_1668),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1728),
.Y(n_1736)
);

AND2x4_ASAP7_75t_L g1737 ( 
.A(n_1719),
.B(n_1667),
.Y(n_1737)
);

HB1xp67_ASAP7_75t_L g1738 ( 
.A(n_1715),
.Y(n_1738)
);

OR2x6_ASAP7_75t_L g1739 ( 
.A(n_1701),
.B(n_1667),
.Y(n_1739)
);

INVx2_ASAP7_75t_L g1740 ( 
.A(n_1699),
.Y(n_1740)
);

AND2x4_ASAP7_75t_L g1741 ( 
.A(n_1731),
.B(n_1643),
.Y(n_1741)
);

AND2x2_ASAP7_75t_L g1742 ( 
.A(n_1703),
.B(n_1690),
.Y(n_1742)
);

AND2x2_ASAP7_75t_L g1743 ( 
.A(n_1690),
.B(n_1646),
.Y(n_1743)
);

INVx2_ASAP7_75t_L g1744 ( 
.A(n_1717),
.Y(n_1744)
);

AND2x2_ASAP7_75t_L g1745 ( 
.A(n_1715),
.B(n_1660),
.Y(n_1745)
);

OR2x2_ASAP7_75t_L g1746 ( 
.A(n_1688),
.B(n_1674),
.Y(n_1746)
);

OR2x2_ASAP7_75t_L g1747 ( 
.A(n_1683),
.B(n_1674),
.Y(n_1747)
);

AND2x2_ASAP7_75t_L g1748 ( 
.A(n_1714),
.B(n_1660),
.Y(n_1748)
);

INVx2_ASAP7_75t_L g1749 ( 
.A(n_1725),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_L g1750 ( 
.A(n_1691),
.B(n_1683),
.Y(n_1750)
);

HB1xp67_ASAP7_75t_L g1751 ( 
.A(n_1726),
.Y(n_1751)
);

INVxp67_ASAP7_75t_SL g1752 ( 
.A(n_1687),
.Y(n_1752)
);

AND2x2_ASAP7_75t_L g1753 ( 
.A(n_1708),
.B(n_1647),
.Y(n_1753)
);

HB1xp67_ASAP7_75t_L g1754 ( 
.A(n_1720),
.Y(n_1754)
);

AND2x4_ASAP7_75t_L g1755 ( 
.A(n_1712),
.B(n_1669),
.Y(n_1755)
);

INVxp67_ASAP7_75t_SL g1756 ( 
.A(n_1687),
.Y(n_1756)
);

BUFx2_ASAP7_75t_L g1757 ( 
.A(n_1732),
.Y(n_1757)
);

NOR2xp33_ASAP7_75t_L g1758 ( 
.A(n_1700),
.B(n_1677),
.Y(n_1758)
);

INVx3_ASAP7_75t_L g1759 ( 
.A(n_1713),
.Y(n_1759)
);

AND2x2_ASAP7_75t_L g1760 ( 
.A(n_1710),
.B(n_1648),
.Y(n_1760)
);

AND2x2_ASAP7_75t_L g1761 ( 
.A(n_1694),
.B(n_1649),
.Y(n_1761)
);

AND2x2_ASAP7_75t_L g1762 ( 
.A(n_1694),
.B(n_1649),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1723),
.Y(n_1763)
);

INVx2_ASAP7_75t_L g1764 ( 
.A(n_1740),
.Y(n_1764)
);

OR2x2_ASAP7_75t_L g1765 ( 
.A(n_1735),
.B(n_1696),
.Y(n_1765)
);

AND2x2_ASAP7_75t_L g1766 ( 
.A(n_1745),
.B(n_1698),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1738),
.Y(n_1767)
);

AND2x4_ASAP7_75t_L g1768 ( 
.A(n_1737),
.B(n_1659),
.Y(n_1768)
);

AND2x2_ASAP7_75t_L g1769 ( 
.A(n_1745),
.B(n_1639),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_L g1770 ( 
.A(n_1763),
.B(n_1700),
.Y(n_1770)
);

AND2x4_ASAP7_75t_L g1771 ( 
.A(n_1737),
.B(n_1659),
.Y(n_1771)
);

NOR2xp33_ASAP7_75t_L g1772 ( 
.A(n_1758),
.B(n_1666),
.Y(n_1772)
);

OR2x2_ASAP7_75t_L g1773 ( 
.A(n_1735),
.B(n_1681),
.Y(n_1773)
);

AOI22xp33_ASAP7_75t_L g1774 ( 
.A1(n_1758),
.A2(n_1692),
.B1(n_1705),
.B2(n_1689),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1738),
.Y(n_1775)
);

INVx3_ASAP7_75t_L g1776 ( 
.A(n_1737),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1744),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1744),
.Y(n_1778)
);

AND2x2_ASAP7_75t_L g1779 ( 
.A(n_1742),
.B(n_1659),
.Y(n_1779)
);

A2O1A1Ixp33_ASAP7_75t_L g1780 ( 
.A1(n_1757),
.A2(n_1706),
.B(n_1685),
.C(n_1697),
.Y(n_1780)
);

INVx2_ASAP7_75t_L g1781 ( 
.A(n_1740),
.Y(n_1781)
);

NAND2xp5_ASAP7_75t_L g1782 ( 
.A(n_1763),
.B(n_1707),
.Y(n_1782)
);

AOI221x1_ASAP7_75t_L g1783 ( 
.A1(n_1763),
.A2(n_1702),
.B1(n_1718),
.B2(n_1630),
.C(n_1631),
.Y(n_1783)
);

AOI211xp5_ASAP7_75t_L g1784 ( 
.A1(n_1754),
.A2(n_1693),
.B(n_1704),
.C(n_1716),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1743),
.Y(n_1785)
);

AND2x2_ASAP7_75t_L g1786 ( 
.A(n_1748),
.B(n_1659),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1743),
.Y(n_1787)
);

OR2x6_ASAP7_75t_L g1788 ( 
.A(n_1739),
.B(n_1663),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1743),
.Y(n_1789)
);

OR2x2_ASAP7_75t_L g1790 ( 
.A(n_1752),
.B(n_1709),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1749),
.Y(n_1791)
);

BUFx2_ASAP7_75t_L g1792 ( 
.A(n_1755),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1749),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1749),
.Y(n_1794)
);

INVxp33_ASAP7_75t_L g1795 ( 
.A(n_1750),
.Y(n_1795)
);

AND2x4_ASAP7_75t_L g1796 ( 
.A(n_1737),
.B(n_1755),
.Y(n_1796)
);

NOR2xp67_ASAP7_75t_SL g1797 ( 
.A(n_1754),
.B(n_1669),
.Y(n_1797)
);

NAND2xp5_ASAP7_75t_L g1798 ( 
.A(n_1782),
.B(n_1752),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1767),
.Y(n_1799)
);

AND2x4_ASAP7_75t_L g1800 ( 
.A(n_1768),
.B(n_1741),
.Y(n_1800)
);

OR2x2_ASAP7_75t_L g1801 ( 
.A(n_1770),
.B(n_1751),
.Y(n_1801)
);

OAI22xp33_ASAP7_75t_SL g1802 ( 
.A1(n_1782),
.A2(n_1739),
.B1(n_1751),
.B2(n_1757),
.Y(n_1802)
);

OA21x2_ASAP7_75t_L g1803 ( 
.A1(n_1783),
.A2(n_1756),
.B(n_1741),
.Y(n_1803)
);

AND2x2_ASAP7_75t_L g1804 ( 
.A(n_1768),
.B(n_1756),
.Y(n_1804)
);

OR2x2_ASAP7_75t_L g1805 ( 
.A(n_1770),
.B(n_1746),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1767),
.Y(n_1806)
);

NAND2xp5_ASAP7_75t_L g1807 ( 
.A(n_1784),
.B(n_1757),
.Y(n_1807)
);

AND2x2_ASAP7_75t_L g1808 ( 
.A(n_1768),
.B(n_1733),
.Y(n_1808)
);

NAND2xp5_ASAP7_75t_L g1809 ( 
.A(n_1784),
.B(n_1750),
.Y(n_1809)
);

NAND2xp5_ASAP7_75t_L g1810 ( 
.A(n_1795),
.B(n_1780),
.Y(n_1810)
);

AOI211xp5_ASAP7_75t_L g1811 ( 
.A1(n_1790),
.A2(n_1721),
.B(n_1727),
.C(n_1760),
.Y(n_1811)
);

NOR2xp33_ASAP7_75t_L g1812 ( 
.A(n_1772),
.B(n_1651),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1775),
.Y(n_1813)
);

AND2x2_ASAP7_75t_L g1814 ( 
.A(n_1768),
.B(n_1734),
.Y(n_1814)
);

AND2x2_ASAP7_75t_L g1815 ( 
.A(n_1771),
.B(n_1769),
.Y(n_1815)
);

INVx2_ASAP7_75t_L g1816 ( 
.A(n_1764),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1775),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1785),
.Y(n_1818)
);

NAND2x1p5_ASAP7_75t_L g1819 ( 
.A(n_1797),
.B(n_1755),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1785),
.Y(n_1820)
);

AND2x2_ASAP7_75t_L g1821 ( 
.A(n_1771),
.B(n_1734),
.Y(n_1821)
);

NOR2x1_ASAP7_75t_L g1822 ( 
.A(n_1790),
.B(n_1739),
.Y(n_1822)
);

NAND2xp5_ASAP7_75t_L g1823 ( 
.A(n_1774),
.B(n_1759),
.Y(n_1823)
);

AND2x2_ASAP7_75t_L g1824 ( 
.A(n_1771),
.B(n_1734),
.Y(n_1824)
);

INVx1_ASAP7_75t_SL g1825 ( 
.A(n_1765),
.Y(n_1825)
);

NAND2xp5_ASAP7_75t_L g1826 ( 
.A(n_1765),
.B(n_1759),
.Y(n_1826)
);

OR2x2_ASAP7_75t_L g1827 ( 
.A(n_1787),
.B(n_1746),
.Y(n_1827)
);

HB1xp67_ASAP7_75t_L g1828 ( 
.A(n_1787),
.Y(n_1828)
);

INVx5_ASAP7_75t_L g1829 ( 
.A(n_1788),
.Y(n_1829)
);

INVx2_ASAP7_75t_L g1830 ( 
.A(n_1764),
.Y(n_1830)
);

AND2x4_ASAP7_75t_L g1831 ( 
.A(n_1771),
.B(n_1741),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1789),
.Y(n_1832)
);

HB1xp67_ASAP7_75t_L g1833 ( 
.A(n_1789),
.Y(n_1833)
);

OAI21xp5_ASAP7_75t_L g1834 ( 
.A1(n_1783),
.A2(n_1739),
.B(n_1753),
.Y(n_1834)
);

INVx2_ASAP7_75t_L g1835 ( 
.A(n_1764),
.Y(n_1835)
);

OR2x2_ASAP7_75t_L g1836 ( 
.A(n_1773),
.B(n_1746),
.Y(n_1836)
);

BUFx2_ASAP7_75t_L g1837 ( 
.A(n_1792),
.Y(n_1837)
);

AND2x4_ASAP7_75t_L g1838 ( 
.A(n_1796),
.B(n_1741),
.Y(n_1838)
);

NAND2x1p5_ASAP7_75t_L g1839 ( 
.A(n_1797),
.B(n_1755),
.Y(n_1839)
);

INVx2_ASAP7_75t_L g1840 ( 
.A(n_1781),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1773),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1791),
.Y(n_1842)
);

OR2x2_ASAP7_75t_L g1843 ( 
.A(n_1777),
.B(n_1747),
.Y(n_1843)
);

INVx2_ASAP7_75t_L g1844 ( 
.A(n_1837),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1813),
.Y(n_1845)
);

AND2x2_ASAP7_75t_L g1846 ( 
.A(n_1815),
.B(n_1804),
.Y(n_1846)
);

INVx1_ASAP7_75t_SL g1847 ( 
.A(n_1837),
.Y(n_1847)
);

NOR2xp33_ASAP7_75t_L g1848 ( 
.A(n_1812),
.B(n_1711),
.Y(n_1848)
);

INVxp67_ASAP7_75t_L g1849 ( 
.A(n_1807),
.Y(n_1849)
);

INVx3_ASAP7_75t_L g1850 ( 
.A(n_1803),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1813),
.Y(n_1851)
);

INVx2_ASAP7_75t_L g1852 ( 
.A(n_1803),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1799),
.Y(n_1853)
);

OR2x2_ASAP7_75t_L g1854 ( 
.A(n_1801),
.B(n_1777),
.Y(n_1854)
);

INVx2_ASAP7_75t_L g1855 ( 
.A(n_1803),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1806),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1817),
.Y(n_1857)
);

AND2x2_ASAP7_75t_L g1858 ( 
.A(n_1815),
.B(n_1792),
.Y(n_1858)
);

AND2x2_ASAP7_75t_L g1859 ( 
.A(n_1804),
.B(n_1796),
.Y(n_1859)
);

NAND2xp5_ASAP7_75t_L g1860 ( 
.A(n_1809),
.B(n_1791),
.Y(n_1860)
);

INVx1_ASAP7_75t_SL g1861 ( 
.A(n_1801),
.Y(n_1861)
);

BUFx3_ASAP7_75t_L g1862 ( 
.A(n_1810),
.Y(n_1862)
);

INVx2_ASAP7_75t_SL g1863 ( 
.A(n_1838),
.Y(n_1863)
);

AND2x2_ASAP7_75t_L g1864 ( 
.A(n_1808),
.B(n_1796),
.Y(n_1864)
);

AND2x2_ASAP7_75t_L g1865 ( 
.A(n_1808),
.B(n_1796),
.Y(n_1865)
);

INVxp67_ASAP7_75t_L g1866 ( 
.A(n_1798),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1820),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1820),
.Y(n_1868)
);

AND2x2_ASAP7_75t_L g1869 ( 
.A(n_1814),
.B(n_1779),
.Y(n_1869)
);

AOI22xp33_ASAP7_75t_L g1870 ( 
.A1(n_1823),
.A2(n_1739),
.B1(n_1788),
.B2(n_1753),
.Y(n_1870)
);

INVx2_ASAP7_75t_SL g1871 ( 
.A(n_1838),
.Y(n_1871)
);

NAND2xp5_ASAP7_75t_L g1872 ( 
.A(n_1825),
.B(n_1793),
.Y(n_1872)
);

NAND2xp5_ASAP7_75t_L g1873 ( 
.A(n_1841),
.B(n_1766),
.Y(n_1873)
);

AND2x2_ASAP7_75t_L g1874 ( 
.A(n_1814),
.B(n_1779),
.Y(n_1874)
);

INVx1_ASAP7_75t_SL g1875 ( 
.A(n_1822),
.Y(n_1875)
);

OR2x2_ASAP7_75t_L g1876 ( 
.A(n_1805),
.B(n_1778),
.Y(n_1876)
);

AND2x2_ASAP7_75t_L g1877 ( 
.A(n_1821),
.B(n_1786),
.Y(n_1877)
);

INVx1_ASAP7_75t_SL g1878 ( 
.A(n_1805),
.Y(n_1878)
);

CKINVDCx16_ASAP7_75t_R g1879 ( 
.A(n_1834),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1828),
.Y(n_1880)
);

INVx1_ASAP7_75t_SL g1881 ( 
.A(n_1833),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1818),
.Y(n_1882)
);

INVx2_ASAP7_75t_L g1883 ( 
.A(n_1850),
.Y(n_1883)
);

INVx1_ASAP7_75t_SL g1884 ( 
.A(n_1847),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_1844),
.Y(n_1885)
);

OR2x2_ASAP7_75t_L g1886 ( 
.A(n_1873),
.B(n_1836),
.Y(n_1886)
);

INVx2_ASAP7_75t_SL g1887 ( 
.A(n_1844),
.Y(n_1887)
);

INVx2_ASAP7_75t_L g1888 ( 
.A(n_1850),
.Y(n_1888)
);

AOI22xp5_ASAP7_75t_L g1889 ( 
.A1(n_1879),
.A2(n_1811),
.B1(n_1802),
.B2(n_1739),
.Y(n_1889)
);

OAI332xp33_ASAP7_75t_L g1890 ( 
.A1(n_1879),
.A2(n_1836),
.A3(n_1832),
.B1(n_1827),
.B2(n_1826),
.B3(n_1747),
.C1(n_1843),
.C2(n_1840),
.Y(n_1890)
);

AOI21xp33_ASAP7_75t_SL g1891 ( 
.A1(n_1849),
.A2(n_1839),
.B(n_1819),
.Y(n_1891)
);

NAND2xp5_ASAP7_75t_SL g1892 ( 
.A(n_1862),
.B(n_1819),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1844),
.Y(n_1893)
);

AOI21xp33_ASAP7_75t_L g1894 ( 
.A1(n_1875),
.A2(n_1739),
.B(n_1788),
.Y(n_1894)
);

INVx1_ASAP7_75t_SL g1895 ( 
.A(n_1847),
.Y(n_1895)
);

OAI32xp33_ASAP7_75t_L g1896 ( 
.A1(n_1850),
.A2(n_1819),
.A3(n_1839),
.B1(n_1827),
.B2(n_1747),
.Y(n_1896)
);

NOR2xp33_ASAP7_75t_L g1897 ( 
.A(n_1862),
.B(n_1848),
.Y(n_1897)
);

OAI22xp5_ASAP7_75t_L g1898 ( 
.A1(n_1862),
.A2(n_1839),
.B1(n_1829),
.B2(n_1788),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1845),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1845),
.Y(n_1900)
);

OAI21xp5_ASAP7_75t_L g1901 ( 
.A1(n_1875),
.A2(n_1829),
.B(n_1788),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1851),
.Y(n_1902)
);

INVx1_ASAP7_75t_L g1903 ( 
.A(n_1851),
.Y(n_1903)
);

NOR2xp33_ASAP7_75t_L g1904 ( 
.A(n_1866),
.B(n_1729),
.Y(n_1904)
);

INVxp67_ASAP7_75t_SL g1905 ( 
.A(n_1850),
.Y(n_1905)
);

AOI33xp33_ASAP7_75t_L g1906 ( 
.A1(n_1861),
.A2(n_1760),
.A3(n_1761),
.B1(n_1762),
.B2(n_1753),
.B3(n_1842),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1867),
.Y(n_1907)
);

AOI221xp5_ASAP7_75t_SL g1908 ( 
.A1(n_1852),
.A2(n_1760),
.B1(n_1824),
.B2(n_1821),
.C(n_1761),
.Y(n_1908)
);

NAND2xp5_ASAP7_75t_L g1909 ( 
.A(n_1861),
.B(n_1766),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1867),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1868),
.Y(n_1911)
);

INVx2_ASAP7_75t_L g1912 ( 
.A(n_1887),
.Y(n_1912)
);

AND2x4_ASAP7_75t_L g1913 ( 
.A(n_1887),
.B(n_1863),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1905),
.Y(n_1914)
);

AND2x4_ASAP7_75t_L g1915 ( 
.A(n_1884),
.B(n_1863),
.Y(n_1915)
);

INVx2_ASAP7_75t_SL g1916 ( 
.A(n_1883),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1885),
.Y(n_1917)
);

INVxp67_ASAP7_75t_L g1918 ( 
.A(n_1897),
.Y(n_1918)
);

INVx1_ASAP7_75t_L g1919 ( 
.A(n_1893),
.Y(n_1919)
);

NAND2xp5_ASAP7_75t_L g1920 ( 
.A(n_1895),
.B(n_1878),
.Y(n_1920)
);

AND2x2_ASAP7_75t_L g1921 ( 
.A(n_1897),
.B(n_1846),
.Y(n_1921)
);

NAND2xp33_ASAP7_75t_L g1922 ( 
.A(n_1889),
.B(n_1852),
.Y(n_1922)
);

OAI22xp5_ASAP7_75t_L g1923 ( 
.A1(n_1892),
.A2(n_1870),
.B1(n_1852),
.B2(n_1855),
.Y(n_1923)
);

INVx1_ASAP7_75t_L g1924 ( 
.A(n_1883),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1888),
.Y(n_1925)
);

INVx2_ASAP7_75t_L g1926 ( 
.A(n_1888),
.Y(n_1926)
);

AND2x4_ASAP7_75t_L g1927 ( 
.A(n_1892),
.B(n_1871),
.Y(n_1927)
);

AND2x2_ASAP7_75t_L g1928 ( 
.A(n_1891),
.B(n_1846),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1899),
.Y(n_1929)
);

INVx1_ASAP7_75t_L g1930 ( 
.A(n_1900),
.Y(n_1930)
);

INVx1_ASAP7_75t_L g1931 ( 
.A(n_1902),
.Y(n_1931)
);

INVx1_ASAP7_75t_SL g1932 ( 
.A(n_1909),
.Y(n_1932)
);

AOI21xp5_ASAP7_75t_L g1933 ( 
.A1(n_1890),
.A2(n_1855),
.B(n_1860),
.Y(n_1933)
);

AND2x2_ASAP7_75t_L g1934 ( 
.A(n_1901),
.B(n_1871),
.Y(n_1934)
);

NAND2xp5_ASAP7_75t_SL g1935 ( 
.A(n_1915),
.B(n_1878),
.Y(n_1935)
);

AND2x2_ASAP7_75t_L g1936 ( 
.A(n_1921),
.B(n_1904),
.Y(n_1936)
);

NOR2xp33_ASAP7_75t_SL g1937 ( 
.A(n_1918),
.B(n_1881),
.Y(n_1937)
);

NAND2xp5_ASAP7_75t_L g1938 ( 
.A(n_1915),
.B(n_1904),
.Y(n_1938)
);

AOI211xp5_ASAP7_75t_L g1939 ( 
.A1(n_1933),
.A2(n_1896),
.B(n_1898),
.C(n_1855),
.Y(n_1939)
);

OAI221xp5_ASAP7_75t_L g1940 ( 
.A1(n_1922),
.A2(n_1908),
.B1(n_1894),
.B2(n_1886),
.C(n_1860),
.Y(n_1940)
);

OAI222xp33_ASAP7_75t_L g1941 ( 
.A1(n_1923),
.A2(n_1881),
.B1(n_1829),
.B2(n_1880),
.C1(n_1858),
.C2(n_1859),
.Y(n_1941)
);

AOI221x1_ASAP7_75t_L g1942 ( 
.A1(n_1914),
.A2(n_1911),
.B1(n_1910),
.B2(n_1907),
.C(n_1903),
.Y(n_1942)
);

NAND4xp25_ASAP7_75t_L g1943 ( 
.A(n_1920),
.B(n_1921),
.C(n_1932),
.D(n_1934),
.Y(n_1943)
);

AOI221xp5_ASAP7_75t_SL g1944 ( 
.A1(n_1922),
.A2(n_1880),
.B1(n_1858),
.B2(n_1856),
.C(n_1853),
.Y(n_1944)
);

NAND2xp5_ASAP7_75t_L g1945 ( 
.A(n_1912),
.B(n_1906),
.Y(n_1945)
);

AOI211xp5_ASAP7_75t_L g1946 ( 
.A1(n_1934),
.A2(n_1856),
.B(n_1857),
.C(n_1853),
.Y(n_1946)
);

NOR2x1_ASAP7_75t_SL g1947 ( 
.A(n_1928),
.B(n_1857),
.Y(n_1947)
);

AOI21xp33_ASAP7_75t_SL g1948 ( 
.A1(n_1915),
.A2(n_1872),
.B(n_1695),
.Y(n_1948)
);

NOR2x1_ASAP7_75t_L g1949 ( 
.A(n_1912),
.B(n_1868),
.Y(n_1949)
);

OAI21xp5_ASAP7_75t_L g1950 ( 
.A1(n_1941),
.A2(n_1927),
.B(n_1928),
.Y(n_1950)
);

NAND2xp5_ASAP7_75t_L g1951 ( 
.A(n_1936),
.B(n_1927),
.Y(n_1951)
);

NOR2x1p5_ASAP7_75t_L g1952 ( 
.A(n_1938),
.B(n_1927),
.Y(n_1952)
);

AO22x2_ASAP7_75t_L g1953 ( 
.A1(n_1942),
.A2(n_1916),
.B1(n_1930),
.B2(n_1929),
.Y(n_1953)
);

NOR2x1_ASAP7_75t_SL g1954 ( 
.A(n_1935),
.B(n_1916),
.Y(n_1954)
);

NOR2x1_ASAP7_75t_L g1955 ( 
.A(n_1943),
.B(n_1926),
.Y(n_1955)
);

INVx1_ASAP7_75t_L g1956 ( 
.A(n_1949),
.Y(n_1956)
);

NAND3xp33_ASAP7_75t_L g1957 ( 
.A(n_1939),
.B(n_1919),
.C(n_1917),
.Y(n_1957)
);

INVx1_ASAP7_75t_L g1958 ( 
.A(n_1947),
.Y(n_1958)
);

NAND2x1_ASAP7_75t_SL g1959 ( 
.A(n_1937),
.B(n_1913),
.Y(n_1959)
);

NAND4xp75_ASAP7_75t_L g1960 ( 
.A(n_1944),
.B(n_1925),
.C(n_1924),
.D(n_1926),
.Y(n_1960)
);

NAND3xp33_ASAP7_75t_L g1961 ( 
.A(n_1945),
.B(n_1913),
.C(n_1931),
.Y(n_1961)
);

NAND3xp33_ASAP7_75t_SL g1962 ( 
.A(n_1950),
.B(n_1945),
.C(n_1948),
.Y(n_1962)
);

NAND4xp25_ASAP7_75t_SL g1963 ( 
.A(n_1957),
.B(n_1940),
.C(n_1906),
.D(n_1946),
.Y(n_1963)
);

OAI211xp5_ASAP7_75t_SL g1964 ( 
.A1(n_1955),
.A2(n_1872),
.B(n_1882),
.C(n_1854),
.Y(n_1964)
);

AOI211x1_ASAP7_75t_SL g1965 ( 
.A1(n_1961),
.A2(n_1913),
.B(n_1830),
.C(n_1835),
.Y(n_1965)
);

A2O1A1Ixp33_ASAP7_75t_L g1966 ( 
.A1(n_1959),
.A2(n_1829),
.B(n_1882),
.C(n_1859),
.Y(n_1966)
);

OAI211xp5_ASAP7_75t_SL g1967 ( 
.A1(n_1951),
.A2(n_1854),
.B(n_1876),
.C(n_1721),
.Y(n_1967)
);

INVx2_ASAP7_75t_L g1968 ( 
.A(n_1954),
.Y(n_1968)
);

INVx1_ASAP7_75t_L g1969 ( 
.A(n_1953),
.Y(n_1969)
);

OAI211xp5_ASAP7_75t_L g1970 ( 
.A1(n_1969),
.A2(n_1956),
.B(n_1958),
.C(n_1953),
.Y(n_1970)
);

NAND2xp5_ASAP7_75t_SL g1971 ( 
.A(n_1968),
.B(n_1829),
.Y(n_1971)
);

INVx1_ASAP7_75t_L g1972 ( 
.A(n_1964),
.Y(n_1972)
);

INVx1_ASAP7_75t_L g1973 ( 
.A(n_1965),
.Y(n_1973)
);

AOI22xp5_ASAP7_75t_L g1974 ( 
.A1(n_1963),
.A2(n_1952),
.B1(n_1960),
.B2(n_1864),
.Y(n_1974)
);

AOI22xp5_ASAP7_75t_L g1975 ( 
.A1(n_1962),
.A2(n_1864),
.B1(n_1865),
.B2(n_1838),
.Y(n_1975)
);

NOR2xp33_ASAP7_75t_L g1976 ( 
.A(n_1966),
.B(n_1865),
.Y(n_1976)
);

AND2x4_ASAP7_75t_L g1977 ( 
.A(n_1971),
.B(n_1975),
.Y(n_1977)
);

OR2x2_ASAP7_75t_L g1978 ( 
.A(n_1972),
.B(n_1876),
.Y(n_1978)
);

NOR2xp33_ASAP7_75t_L g1979 ( 
.A(n_1974),
.B(n_1967),
.Y(n_1979)
);

AND2x2_ASAP7_75t_L g1980 ( 
.A(n_1976),
.B(n_1869),
.Y(n_1980)
);

NAND3xp33_ASAP7_75t_L g1981 ( 
.A(n_1970),
.B(n_1874),
.C(n_1869),
.Y(n_1981)
);

OAI221xp5_ASAP7_75t_SL g1982 ( 
.A1(n_1973),
.A2(n_1874),
.B1(n_1877),
.B2(n_1843),
.C(n_1636),
.Y(n_1982)
);

AOI21xp5_ASAP7_75t_L g1983 ( 
.A1(n_1977),
.A2(n_1830),
.B(n_1816),
.Y(n_1983)
);

INVx3_ASAP7_75t_SL g1984 ( 
.A(n_1978),
.Y(n_1984)
);

AND2x4_ASAP7_75t_L g1985 ( 
.A(n_1980),
.B(n_1877),
.Y(n_1985)
);

XOR2x1_ASAP7_75t_L g1986 ( 
.A(n_1981),
.B(n_1800),
.Y(n_1986)
);

INVx1_ASAP7_75t_L g1987 ( 
.A(n_1986),
.Y(n_1987)
);

NAND5xp2_ASAP7_75t_L g1988 ( 
.A(n_1987),
.B(n_1979),
.C(n_1982),
.D(n_1983),
.E(n_1984),
.Y(n_1988)
);

OAI22xp5_ASAP7_75t_L g1989 ( 
.A1(n_1988),
.A2(n_1985),
.B1(n_1840),
.B2(n_1835),
.Y(n_1989)
);

INVx1_ASAP7_75t_L g1990 ( 
.A(n_1988),
.Y(n_1990)
);

AOI21xp33_ASAP7_75t_L g1991 ( 
.A1(n_1990),
.A2(n_1816),
.B(n_1800),
.Y(n_1991)
);

OAI221xp5_ASAP7_75t_L g1992 ( 
.A1(n_1989),
.A2(n_1776),
.B1(n_1793),
.B2(n_1794),
.C(n_1736),
.Y(n_1992)
);

INVx1_ASAP7_75t_L g1993 ( 
.A(n_1991),
.Y(n_1993)
);

INVx1_ASAP7_75t_L g1994 ( 
.A(n_1992),
.Y(n_1994)
);

AOI21xp5_ASAP7_75t_L g1995 ( 
.A1(n_1993),
.A2(n_1994),
.B(n_1831),
.Y(n_1995)
);

AOI22xp5_ASAP7_75t_SL g1996 ( 
.A1(n_1995),
.A2(n_1831),
.B1(n_1800),
.B2(n_1824),
.Y(n_1996)
);

OAI221xp5_ASAP7_75t_R g1997 ( 
.A1(n_1996),
.A2(n_1724),
.B1(n_1831),
.B2(n_1722),
.C(n_1562),
.Y(n_1997)
);

AOI211xp5_ASAP7_75t_L g1998 ( 
.A1(n_1997),
.A2(n_1730),
.B(n_1626),
.C(n_1568),
.Y(n_1998)
);


endmodule