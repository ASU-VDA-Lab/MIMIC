module fake_jpeg_3687_n_36 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_36);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_36;

wire n_13;
wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_32;
wire n_15;

NOR2xp33_ASAP7_75t_L g13 ( 
.A(n_7),
.B(n_4),
.Y(n_13)
);

INVx4_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_SL g16 ( 
.A(n_1),
.B(n_3),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_18),
.Y(n_23)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_19),
.Y(n_21)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_20),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_19),
.B(n_16),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_22),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g26 ( 
.A1(n_24),
.A2(n_20),
.B1(n_15),
.B2(n_17),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_26),
.B(n_28),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_23),
.B(n_13),
.C(n_17),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g30 ( 
.A(n_27),
.B(n_25),
.C(n_21),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g28 ( 
.A1(n_21),
.A2(n_15),
.B1(n_16),
.B2(n_2),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g31 ( 
.A(n_30),
.B(n_0),
.C(n_1),
.Y(n_31)
);

XNOR2xp5_ASAP7_75t_SL g33 ( 
.A(n_31),
.B(n_32),
.Y(n_33)
);

XOR2xp5_ASAP7_75t_L g32 ( 
.A(n_29),
.B(n_5),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g34 ( 
.A(n_33),
.B(n_6),
.C(n_8),
.Y(n_34)
);

O2A1O1Ixp33_ASAP7_75t_SL g35 ( 
.A1(n_34),
.A2(n_9),
.B(n_10),
.C(n_12),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_35),
.Y(n_36)
);


endmodule