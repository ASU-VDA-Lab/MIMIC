module fake_jpeg_1026_n_120 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_8, n_15, n_7, n_120);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_8;
input n_15;
input n_7;

output n_120;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

BUFx8_ASAP7_75t_L g32 ( 
.A(n_27),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

CKINVDCx14_ASAP7_75t_R g36 ( 
.A(n_28),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_29),
.Y(n_39)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_14),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_43),
.B(n_47),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

INVx13_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_46),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_32),
.B(n_0),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_36),
.Y(n_48)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_48),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

CKINVDCx12_ASAP7_75t_R g54 ( 
.A(n_49),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_44),
.A2(n_40),
.B1(n_33),
.B2(n_41),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

AOI32xp33_ASAP7_75t_L g55 ( 
.A1(n_43),
.A2(n_40),
.A3(n_42),
.B1(n_37),
.B2(n_33),
.Y(n_55)
);

OR2x2_ASAP7_75t_L g71 ( 
.A(n_55),
.B(n_31),
.Y(n_71)
);

O2A1O1Ixp33_ASAP7_75t_L g56 ( 
.A1(n_44),
.A2(n_45),
.B(n_46),
.C(n_48),
.Y(n_56)
);

OAI21xp33_ASAP7_75t_L g68 ( 
.A1(n_56),
.A2(n_35),
.B(n_38),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_49),
.A2(n_41),
.B1(n_42),
.B2(n_37),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_57),
.A2(n_47),
.B1(n_49),
.B2(n_45),
.Y(n_61)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_50),
.Y(n_60)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_60),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_61),
.A2(n_65),
.B1(n_59),
.B2(n_71),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_53),
.B(n_39),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_62),
.B(n_63),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_53),
.B(n_1),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_52),
.B(n_1),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_64),
.B(n_66),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_58),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_56),
.B(n_49),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_67),
.B(n_69),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_68),
.B(n_70),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_58),
.B(n_2),
.Y(n_69)
);

XOR2xp5_ASAP7_75t_L g70 ( 
.A(n_54),
.B(n_35),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_71),
.B(n_30),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_70),
.B(n_15),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_72),
.B(n_73),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_68),
.B(n_16),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_74),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_93)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_61),
.Y(n_78)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_78),
.Y(n_87)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_65),
.Y(n_79)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_79),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_80),
.B(n_81),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_62),
.B(n_2),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_67),
.A2(n_59),
.B(n_4),
.Y(n_84)
);

NAND2x1_ASAP7_75t_L g86 ( 
.A(n_84),
.B(n_3),
.Y(n_86)
);

INVx1_ASAP7_75t_SL g102 ( 
.A(n_86),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_83),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_88),
.A2(n_90),
.B1(n_93),
.B2(n_84),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_82),
.B(n_5),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_89),
.B(n_92),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_83),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_72),
.B(n_19),
.C(n_23),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_91),
.B(n_96),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_75),
.B(n_76),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_77),
.B(n_9),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_95),
.B(n_74),
.C(n_73),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_97),
.B(n_100),
.C(n_104),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_98),
.Y(n_109)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_87),
.Y(n_99)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_99),
.Y(n_111)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_94),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_91),
.B(n_25),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_SL g107 ( 
.A(n_101),
.B(n_10),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_88),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_103),
.A2(n_11),
.B(n_13),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_93),
.A2(n_86),
.B1(n_90),
.B2(n_85),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_107),
.B(n_102),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_110),
.B(n_103),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_112),
.A2(n_113),
.B1(n_114),
.B2(n_102),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_111),
.B(n_105),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_115),
.B(n_116),
.C(n_107),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_114),
.B(n_108),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_117),
.B(n_116),
.C(n_106),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_118),
.B(n_101),
.C(n_109),
.Y(n_119)
);

AOI221xp5_ASAP7_75t_L g120 ( 
.A1(n_119),
.A2(n_22),
.B1(n_18),
.B2(n_20),
.C(n_21),
.Y(n_120)
);


endmodule