module fake_jpeg_23894_n_306 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_306);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_306;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_14;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_301;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_145;
wire n_18;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_303;
wire n_90;
wire n_304;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_300;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_302;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_305;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_270;
wire n_260;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_282;
wire n_258;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_7),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_3),
.Y(n_14)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_2),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_4),
.B(n_8),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx24_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_5),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_24),
.Y(n_28)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_24),
.Y(n_29)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_24),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

BUFx10_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_17),
.B(n_12),
.Y(n_32)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_25),
.B(n_0),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_33),
.B(n_15),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_27),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_34),
.B(n_35),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_27),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_36),
.B(n_22),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_43),
.B(n_44),
.Y(n_60)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

CKINVDCx16_ASAP7_75t_R g64 ( 
.A(n_45),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_32),
.B(n_17),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_47),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_33),
.A2(n_21),
.B1(n_15),
.B2(n_23),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_50),
.A2(n_31),
.B1(n_36),
.B2(n_21),
.Y(n_59)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_29),
.Y(n_51)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_52),
.B(n_33),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_28),
.Y(n_53)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_53),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_32),
.B(n_19),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_54),
.B(n_32),
.Y(n_71)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_55),
.Y(n_93)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_53),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_56),
.B(n_72),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_38),
.A2(n_15),
.B1(n_21),
.B2(n_19),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_57),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_SL g94 ( 
.A(n_59),
.B(n_74),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_52),
.A2(n_31),
.B1(n_23),
.B2(n_21),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_61),
.B(n_36),
.C(n_48),
.Y(n_87)
);

HB1xp67_ASAP7_75t_L g62 ( 
.A(n_53),
.Y(n_62)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_62),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_52),
.B(n_33),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_63),
.B(n_36),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_38),
.A2(n_21),
.B1(n_15),
.B2(n_23),
.Y(n_65)
);

OAI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_65),
.A2(n_66),
.B1(n_51),
.B2(n_46),
.Y(n_90)
);

OAI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_50),
.A2(n_31),
.B1(n_34),
.B2(n_35),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_67),
.Y(n_96)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_70),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_71),
.B(n_39),
.Y(n_76)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

CKINVDCx12_ASAP7_75t_R g73 ( 
.A(n_39),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_73),
.B(n_22),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_76),
.B(n_82),
.Y(n_107)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_70),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_77),
.B(n_79),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_55),
.A2(n_40),
.B1(n_44),
.B2(n_43),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_78),
.Y(n_101)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_58),
.Y(n_79)
);

XOR2xp5_ASAP7_75t_L g81 ( 
.A(n_63),
.B(n_74),
.Y(n_81)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_81),
.B(n_87),
.Y(n_113)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_58),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_84),
.B(n_85),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_68),
.B(n_35),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_74),
.B(n_48),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_88),
.B(n_97),
.Y(n_99)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_60),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_89),
.B(n_95),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_90),
.A2(n_69),
.B1(n_75),
.B2(n_70),
.Y(n_103)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_58),
.Y(n_91)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_91),
.Y(n_105)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_73),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_83),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_98),
.B(n_115),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_92),
.A2(n_61),
.B1(n_59),
.B2(n_68),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_100),
.A2(n_110),
.B1(n_96),
.B2(n_80),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_81),
.B(n_71),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_102),
.B(n_104),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_103),
.A2(n_119),
.B1(n_93),
.B2(n_69),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_82),
.B(n_64),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_SL g109 ( 
.A(n_94),
.B(n_70),
.C(n_64),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_109),
.A2(n_112),
.B(n_86),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_88),
.A2(n_75),
.B1(n_56),
.B2(n_72),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_85),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_111),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_92),
.A2(n_46),
.B(n_25),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_76),
.Y(n_115)
);

INVx13_ASAP7_75t_L g116 ( 
.A(n_77),
.Y(n_116)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_116),
.Y(n_139)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_80),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_117),
.B(n_118),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_87),
.Y(n_118)
);

OAI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_93),
.A2(n_69),
.B1(n_48),
.B2(n_35),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_109),
.A2(n_94),
.B(n_97),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_121),
.A2(n_141),
.B(n_144),
.Y(n_154)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_106),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_122),
.B(n_123),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_106),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_SL g124 ( 
.A(n_113),
.B(n_89),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_124),
.A2(n_126),
.B(n_137),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_125),
.A2(n_129),
.B1(n_136),
.B2(n_110),
.Y(n_148)
);

NOR2x1_ASAP7_75t_L g128 ( 
.A(n_115),
.B(n_34),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_128),
.B(n_135),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_103),
.A2(n_86),
.B1(n_91),
.B2(n_84),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_113),
.B(n_37),
.C(n_79),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_130),
.B(n_134),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_131),
.A2(n_133),
.B1(n_105),
.B2(n_117),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_116),
.B(n_96),
.Y(n_132)
);

CKINVDCx14_ASAP7_75t_R g151 ( 
.A(n_132),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_100),
.A2(n_34),
.B1(n_49),
.B2(n_41),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_102),
.B(n_37),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_111),
.B(n_13),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_101),
.A2(n_49),
.B1(n_41),
.B2(n_13),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_112),
.A2(n_37),
.B(n_28),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_99),
.B(n_37),
.C(n_49),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_138),
.B(n_105),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_104),
.B(n_20),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_140),
.B(n_114),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_99),
.A2(n_14),
.B(n_26),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_107),
.A2(n_37),
.B(n_28),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_145),
.B(n_146),
.Y(n_181)
);

CKINVDCx12_ASAP7_75t_R g146 ( 
.A(n_139),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_L g172 ( 
.A1(n_148),
.A2(n_141),
.B1(n_136),
.B2(n_116),
.Y(n_172)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_120),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_149),
.B(n_152),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_131),
.A2(n_107),
.B1(n_114),
.B2(n_98),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_150),
.A2(n_166),
.B1(n_30),
.B2(n_29),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_143),
.B(n_128),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_139),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_153),
.B(n_158),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_155),
.B(n_67),
.C(n_30),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_143),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_156),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_142),
.B(n_108),
.Y(n_157)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_157),
.Y(n_195)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_138),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_121),
.A2(n_108),
.B(n_119),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_159),
.A2(n_170),
.B(n_20),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_135),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_161),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_129),
.A2(n_127),
.B1(n_130),
.B2(n_133),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_162),
.A2(n_37),
.B1(n_67),
.B2(n_28),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_142),
.B(n_105),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_163),
.B(n_164),
.Y(n_190)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_144),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_123),
.B(n_122),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_165),
.Y(n_182)
);

NAND2x1_ASAP7_75t_SL g168 ( 
.A(n_137),
.B(n_126),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_168),
.A2(n_134),
.B(n_124),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_140),
.B(n_16),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_172),
.A2(n_177),
.B1(n_188),
.B2(n_191),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_173),
.A2(n_154),
.B(n_157),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_156),
.B(n_22),
.Y(n_174)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_174),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_153),
.B(n_150),
.Y(n_175)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_175),
.Y(n_212)
);

MAJx2_ASAP7_75t_L g178 ( 
.A(n_160),
.B(n_22),
.C(n_11),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_178),
.B(n_159),
.Y(n_199)
);

HB1xp67_ASAP7_75t_L g183 ( 
.A(n_146),
.Y(n_183)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_183),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_149),
.B(n_22),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_184),
.B(n_185),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_151),
.B(n_16),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_186),
.B(n_155),
.C(n_147),
.Y(n_198)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_166),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_187),
.B(n_189),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_164),
.A2(n_162),
.B1(n_160),
.B2(n_148),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_158),
.A2(n_14),
.B1(n_18),
.B2(n_26),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_167),
.B(n_18),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_192),
.B(n_170),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_193),
.A2(n_167),
.B1(n_163),
.B2(n_145),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_165),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_194),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_173),
.B(n_147),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_197),
.B(n_199),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_198),
.B(n_214),
.C(n_215),
.Y(n_232)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_200),
.Y(n_218)
);

BUFx12f_ASAP7_75t_L g202 ( 
.A(n_179),
.Y(n_202)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_202),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_188),
.B(n_154),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_203),
.B(n_204),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_207),
.A2(n_177),
.B1(n_187),
.B2(n_194),
.Y(n_217)
);

OR2x2_ASAP7_75t_L g208 ( 
.A(n_180),
.B(n_152),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_208),
.B(n_209),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_176),
.Y(n_209)
);

AO22x1_ASAP7_75t_SL g210 ( 
.A1(n_190),
.A2(n_168),
.B1(n_169),
.B2(n_161),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_210),
.A2(n_182),
.B1(n_195),
.B2(n_178),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_176),
.A2(n_169),
.B(n_168),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_211),
.A2(n_195),
.B1(n_186),
.B2(n_189),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_190),
.B(n_11),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_182),
.B(n_30),
.C(n_29),
.Y(n_215)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_217),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_212),
.A2(n_193),
.B1(n_180),
.B2(n_179),
.Y(n_220)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_220),
.Y(n_244)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_202),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_221),
.B(n_222),
.Y(n_245)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_202),
.Y(n_222)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_214),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_225),
.B(n_229),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_197),
.B(n_171),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_226),
.B(n_228),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_203),
.B(n_171),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_201),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_230),
.A2(n_234),
.B(n_210),
.Y(n_239)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_208),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_231),
.B(n_235),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_196),
.B(n_181),
.Y(n_233)
);

CKINVDCx14_ASAP7_75t_R g252 ( 
.A(n_233),
.Y(n_252)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_215),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_210),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_236),
.B(n_199),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_232),
.B(n_198),
.C(n_213),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_238),
.B(n_250),
.C(n_251),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_239),
.B(n_1),
.Y(n_268)
);

BUFx12_ASAP7_75t_L g241 ( 
.A(n_227),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_241),
.B(n_246),
.Y(n_262)
);

HB1xp67_ASAP7_75t_L g242 ( 
.A(n_228),
.Y(n_242)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_242),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_219),
.A2(n_209),
.B(n_216),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_SL g264 ( 
.A1(n_243),
.A2(n_0),
.B(n_1),
.Y(n_264)
);

INVx13_ASAP7_75t_L g246 ( 
.A(n_217),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_230),
.Y(n_247)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_247),
.Y(n_260)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_249),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_232),
.B(n_223),
.C(n_226),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_223),
.B(n_205),
.C(n_206),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_241),
.B(n_191),
.Y(n_254)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_254),
.Y(n_269)
);

OR2x2_ASAP7_75t_L g255 ( 
.A(n_246),
.B(n_224),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_255),
.B(n_259),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_247),
.A2(n_224),
.B1(n_218),
.B2(n_2),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_256),
.B(n_257),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_240),
.A2(n_239),
.B1(n_244),
.B2(n_237),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_241),
.B(n_11),
.Y(n_259)
);

HB1xp67_ASAP7_75t_L g263 ( 
.A(n_245),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_263),
.B(n_265),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_264),
.A2(n_243),
.B(n_249),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_253),
.B(n_10),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_237),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_266),
.B(n_268),
.C(n_1),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_270),
.B(n_268),
.Y(n_281)
);

AND2x2_ASAP7_75t_L g272 ( 
.A(n_261),
.B(n_250),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_272),
.B(n_277),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_260),
.A2(n_238),
.B(n_252),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_L g286 ( 
.A1(n_274),
.A2(n_275),
.B(n_256),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_262),
.A2(n_251),
.B(n_248),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_267),
.A2(n_10),
.B1(n_9),
.B2(n_4),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_276),
.B(n_279),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_266),
.B(n_9),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_278),
.B(n_3),
.Y(n_288)
);

HB1xp67_ASAP7_75t_L g279 ( 
.A(n_255),
.Y(n_279)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_281),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_280),
.B(n_269),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_282),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_SL g284 ( 
.A1(n_271),
.A2(n_258),
.B(n_261),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_284),
.B(n_288),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_273),
.B(n_257),
.Y(n_285)
);

AOI322xp5_ASAP7_75t_L g296 ( 
.A1(n_285),
.A2(n_286),
.A3(n_287),
.B1(n_290),
.B2(n_6),
.C1(n_30),
.C2(n_29),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_273),
.A2(n_10),
.B1(n_4),
.B2(n_5),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_SL g290 ( 
.A(n_275),
.B(n_3),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_289),
.B(n_4),
.C(n_5),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_293),
.B(n_294),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_289),
.B(n_5),
.C(n_6),
.Y(n_294)
);

O2A1O1Ixp33_ASAP7_75t_SL g299 ( 
.A1(n_296),
.A2(n_283),
.B(n_6),
.C(n_30),
.Y(n_299)
);

INVxp33_ASAP7_75t_L g298 ( 
.A(n_292),
.Y(n_298)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_298),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_299),
.B(n_292),
.Y(n_300)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_300),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_302),
.A2(n_301),
.B(n_295),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_303),
.B(n_297),
.C(n_291),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_304),
.A2(n_6),
.B1(n_30),
.B2(n_29),
.Y(n_305)
);

AO21x1_ASAP7_75t_L g306 ( 
.A1(n_305),
.A2(n_29),
.B(n_156),
.Y(n_306)
);


endmodule