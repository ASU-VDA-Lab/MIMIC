module fake_jpeg_14824_n_39 (n_3, n_2, n_1, n_0, n_4, n_5, n_39);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_39;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx4_ASAP7_75t_L g6 ( 
.A(n_4),
.Y(n_6)
);

NOR2xp33_ASAP7_75t_L g7 ( 
.A(n_4),
.B(n_3),
.Y(n_7)
);

INVx11_ASAP7_75t_L g8 ( 
.A(n_3),
.Y(n_8)
);

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_3),
.Y(n_9)
);

INVx8_ASAP7_75t_L g10 ( 
.A(n_2),
.Y(n_10)
);

AOI21xp33_ASAP7_75t_SL g11 ( 
.A1(n_2),
.A2(n_5),
.B(n_0),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_7),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_12),
.B(n_6),
.Y(n_18)
);

AOI22xp5_ASAP7_75t_L g13 ( 
.A1(n_11),
.A2(n_6),
.B1(n_10),
.B2(n_2),
.Y(n_13)
);

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_13),
.A2(n_15),
.B1(n_16),
.B2(n_1),
.Y(n_19)
);

AND2x4_ASAP7_75t_L g14 ( 
.A(n_11),
.B(n_0),
.Y(n_14)
);

AOI21xp5_ASAP7_75t_L g17 ( 
.A1(n_14),
.A2(n_1),
.B(n_7),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_SL g15 ( 
.A1(n_6),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_15)
);

AOI22xp33_ASAP7_75t_L g16 ( 
.A1(n_6),
.A2(n_4),
.B1(n_5),
.B2(n_0),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_SL g24 ( 
.A1(n_17),
.A2(n_18),
.B(n_19),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_12),
.B(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_20),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_22),
.B(n_14),
.Y(n_26)
);

OAI21xp5_ASAP7_75t_L g23 ( 
.A1(n_19),
.A2(n_14),
.B(n_13),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_23),
.B(n_25),
.C(n_14),
.Y(n_27)
);

OAI21xp5_ASAP7_75t_SL g25 ( 
.A1(n_17),
.A2(n_14),
.B(n_15),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g32 ( 
.A(n_26),
.B(n_27),
.C(n_28),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g28 ( 
.A(n_24),
.B(n_9),
.C(n_8),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_21),
.B(n_10),
.Y(n_29)
);

XOR2xp5_ASAP7_75t_L g30 ( 
.A(n_29),
.B(n_23),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_30),
.B(n_9),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_L g31 ( 
.A1(n_28),
.A2(n_10),
.B1(n_8),
.B2(n_9),
.Y(n_31)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_31),
.B(n_9),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_33),
.A2(n_8),
.B1(n_31),
.B2(n_1),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_34),
.B(n_35),
.Y(n_37)
);

XNOR2xp5_ASAP7_75t_L g35 ( 
.A(n_32),
.B(n_10),
.Y(n_35)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_36),
.Y(n_38)
);

AOI21xp5_ASAP7_75t_L g39 ( 
.A1(n_38),
.A2(n_37),
.B(n_35),
.Y(n_39)
);


endmodule