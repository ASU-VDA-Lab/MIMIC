module fake_ariane_1623_n_865 (n_83, n_8, n_56, n_60, n_160, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_158, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_865);

input n_83;
input n_8;
input n_56;
input n_60;
input n_160;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_158;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_865;

wire n_295;
wire n_356;
wire n_556;
wire n_170;
wire n_190;
wire n_698;
wire n_695;
wire n_180;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_581;
wire n_294;
wire n_646;
wire n_197;
wire n_640;
wire n_463;
wire n_830;
wire n_176;
wire n_691;
wire n_404;
wire n_172;
wire n_678;
wire n_651;
wire n_347;
wire n_423;
wire n_183;
wire n_469;
wire n_479;
wire n_726;
wire n_603;
wire n_373;
wire n_299;
wire n_836;
wire n_541;
wire n_499;
wire n_789;
wire n_788;
wire n_850;
wire n_771;
wire n_564;
wire n_610;
wire n_205;
wire n_752;
wire n_341;
wire n_421;
wire n_245;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_760;
wire n_690;
wire n_416;
wire n_283;
wire n_525;
wire n_187;
wire n_806;
wire n_367;
wire n_713;
wire n_649;
wire n_598;
wire n_374;
wire n_345;
wire n_318;
wire n_817;
wire n_244;
wire n_643;
wire n_679;
wire n_226;
wire n_781;
wire n_220;
wire n_261;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_189;
wire n_717;
wire n_819;
wire n_286;
wire n_443;
wire n_586;
wire n_864;
wire n_686;
wire n_605;
wire n_776;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_826;
wire n_524;
wire n_634;
wire n_391;
wire n_349;
wire n_756;
wire n_466;
wire n_346;
wire n_214;
wire n_764;
wire n_348;
wire n_552;
wire n_462;
wire n_607;
wire n_670;
wire n_410;
wire n_379;
wire n_445;
wire n_515;
wire n_807;
wire n_765;
wire n_264;
wire n_737;
wire n_198;
wire n_232;
wire n_441;
wire n_568;
wire n_385;
wire n_637;
wire n_327;
wire n_766;
wire n_372;
wire n_377;
wire n_396;
wire n_802;
wire n_631;
wire n_399;
wire n_554;
wire n_520;
wire n_714;
wire n_279;
wire n_702;
wire n_207;
wire n_790;
wire n_857;
wire n_363;
wire n_720;
wire n_354;
wire n_813;
wire n_725;
wire n_419;
wire n_230;
wire n_270;
wire n_194;
wire n_633;
wire n_338;
wire n_285;
wire n_473;
wire n_186;
wire n_801;
wire n_202;
wire n_193;
wire n_761;
wire n_733;
wire n_818;
wire n_500;
wire n_665;
wire n_336;
wire n_731;
wire n_754;
wire n_779;
wire n_315;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_829;
wire n_668;
wire n_339;
wire n_758;
wire n_738;
wire n_833;
wire n_672;
wire n_487;
wire n_740;
wire n_167;
wire n_422;
wire n_648;
wire n_784;
wire n_269;
wire n_597;
wire n_816;
wire n_855;
wire n_259;
wire n_835;
wire n_808;
wire n_446;
wire n_553;
wire n_753;
wire n_566;
wire n_814;
wire n_578;
wire n_701;
wire n_625;
wire n_405;
wire n_557;
wire n_169;
wire n_173;
wire n_858;
wire n_242;
wire n_645;
wire n_309;
wire n_320;
wire n_331;
wire n_559;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_822;
wire n_344;
wire n_381;
wire n_795;
wire n_426;
wire n_433;
wire n_481;
wire n_600;
wire n_721;
wire n_840;
wire n_398;
wire n_210;
wire n_200;
wire n_529;
wire n_502;
wire n_253;
wire n_561;
wire n_770;
wire n_218;
wire n_821;
wire n_839;
wire n_271;
wire n_507;
wire n_486;
wire n_465;
wire n_759;
wire n_247;
wire n_569;
wire n_567;
wire n_825;
wire n_732;
wire n_240;
wire n_369;
wire n_224;
wire n_787;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_222;
wire n_478;
wire n_703;
wire n_748;
wire n_786;
wire n_510;
wire n_831;
wire n_256;
wire n_326;
wire n_681;
wire n_778;
wire n_227;
wire n_188;
wire n_323;
wire n_550;
wire n_635;
wire n_707;
wire n_330;
wire n_400;
wire n_689;
wire n_694;
wire n_282;
wire n_328;
wire n_368;
wire n_590;
wire n_699;
wire n_727;
wire n_277;
wire n_248;
wire n_301;
wire n_467;
wire n_432;
wire n_545;
wire n_536;
wire n_644;
wire n_293;
wire n_823;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_859;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_693;
wire n_863;
wire n_303;
wire n_671;
wire n_442;
wire n_777;
wire n_168;
wire n_352;
wire n_538;
wire n_206;
wire n_576;
wire n_843;
wire n_511;
wire n_611;
wire n_238;
wire n_365;
wire n_455;
wire n_429;
wire n_654;
wire n_588;
wire n_638;
wire n_334;
wire n_192;
wire n_729;
wire n_661;
wire n_488;
wire n_775;
wire n_667;
wire n_300;
wire n_533;
wire n_505;
wire n_846;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_512;
wire n_715;
wire n_579;
wire n_844;
wire n_459;
wire n_685;
wire n_221;
wire n_321;
wire n_458;
wire n_361;
wire n_383;
wire n_623;
wire n_838;
wire n_237;
wire n_780;
wire n_861;
wire n_175;
wire n_711;
wire n_453;
wire n_734;
wire n_491;
wire n_810;
wire n_181;
wire n_723;
wire n_617;
wire n_616;
wire n_658;
wire n_630;
wire n_705;
wire n_570;
wire n_260;
wire n_362;
wire n_543;
wire n_310;
wire n_709;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_281;
wire n_628;
wire n_809;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_743;
wire n_225;
wire n_235;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_297;
wire n_662;
wire n_641;
wire n_503;
wire n_700;
wire n_290;
wire n_527;
wire n_741;
wire n_747;
wire n_772;
wire n_847;
wire n_371;
wire n_845;
wire n_199;
wire n_639;
wire n_217;
wire n_452;
wire n_673;
wire n_676;
wire n_178;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_201;
wire n_572;
wire n_343;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_582;
wire n_284;
wire n_448;
wire n_593;
wire n_755;
wire n_710;
wire n_860;
wire n_249;
wire n_534;
wire n_355;
wire n_212;
wire n_444;
wire n_609;
wire n_278;
wire n_851;
wire n_255;
wire n_560;
wire n_450;
wire n_257;
wire n_842;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_468;
wire n_853;
wire n_526;
wire n_742;
wire n_716;
wire n_182;
wire n_696;
wire n_674;
wire n_482;
wire n_316;
wire n_196;
wire n_798;
wire n_769;
wire n_820;
wire n_577;
wire n_407;
wire n_774;
wire n_254;
wire n_596;
wire n_476;
wire n_460;
wire n_219;
wire n_832;
wire n_535;
wire n_231;
wire n_366;
wire n_744;
wire n_762;
wire n_656;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_848;
wire n_804;
wire n_280;
wire n_215;
wire n_252;
wire n_629;
wire n_664;
wire n_454;
wire n_298;
wire n_532;
wire n_415;
wire n_794;
wire n_763;
wire n_655;
wire n_544;
wire n_540;
wire n_216;
wire n_692;
wire n_599;
wire n_768;
wire n_514;
wire n_418;
wire n_537;
wire n_223;
wire n_403;
wire n_750;
wire n_834;
wire n_389;
wire n_800;
wire n_657;
wire n_513;
wire n_837;
wire n_288;
wire n_179;
wire n_812;
wire n_395;
wire n_621;
wire n_195;
wire n_606;
wire n_213;
wire n_862;
wire n_304;
wire n_659;
wire n_583;
wire n_509;
wire n_724;
wire n_306;
wire n_666;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_203;
wire n_378;
wire n_436;
wire n_757;
wire n_375;
wire n_324;
wire n_585;
wire n_669;
wire n_785;
wire n_827;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_622;
wire n_697;
wire n_472;
wire n_296;
wire n_265;
wire n_746;
wire n_208;
wire n_456;
wire n_292;
wire n_793;
wire n_852;
wire n_174;
wire n_275;
wire n_704;
wire n_204;
wire n_751;
wire n_615;
wire n_521;
wire n_496;
wire n_739;
wire n_342;
wire n_246;
wire n_517;
wire n_530;
wire n_792;
wire n_824;
wire n_428;
wire n_358;
wire n_580;
wire n_608;
wire n_494;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_563;
wire n_229;
wire n_394;
wire n_250;
wire n_773;
wire n_317;
wire n_243;
wire n_803;
wire n_329;
wire n_718;
wire n_185;
wire n_340;
wire n_749;
wire n_289;
wire n_548;
wire n_542;
wire n_815;
wire n_523;
wire n_268;
wire n_266;
wire n_470;
wire n_457;
wire n_632;
wire n_184;
wire n_177;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_782;
wire n_856;
wire n_425;
wire n_431;
wire n_811;
wire n_508;
wire n_624;
wire n_791;
wire n_618;
wire n_411;
wire n_484;
wire n_712;
wire n_849;
wire n_353;
wire n_736;
wire n_767;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_382;
wire n_191;
wire n_797;
wire n_489;
wire n_480;
wire n_211;
wire n_642;
wire n_408;
wire n_828;
wire n_595;
wire n_322;
wire n_251;
wire n_506;
wire n_602;
wire n_799;
wire n_558;
wire n_592;
wire n_397;
wire n_841;
wire n_854;
wire n_471;
wire n_351;
wire n_393;
wire n_474;
wire n_653;
wire n_359;
wire n_573;
wire n_796;
wire n_805;
wire n_531;
wire n_783;
wire n_675;

INVx1_ASAP7_75t_L g167 ( 
.A(n_157),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_100),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_163),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_160),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_147),
.Y(n_171)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_46),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_91),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_155),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_15),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_133),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_146),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_165),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_152),
.Y(n_179)
);

BUFx10_ASAP7_75t_L g180 ( 
.A(n_88),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_42),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_162),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_80),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_39),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g185 ( 
.A(n_86),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_131),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_113),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_153),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_130),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_164),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_135),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_12),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_18),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_84),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_156),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_74),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_48),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_95),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_159),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_92),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_117),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_3),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_34),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_61),
.Y(n_204)
);

INVx1_ASAP7_75t_SL g205 ( 
.A(n_9),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_52),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_76),
.Y(n_207)
);

BUFx3_ASAP7_75t_L g208 ( 
.A(n_141),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_166),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_127),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_114),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_158),
.Y(n_212)
);

BUFx2_ASAP7_75t_L g213 ( 
.A(n_96),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_144),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_6),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_128),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_161),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_104),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_9),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_45),
.Y(n_220)
);

BUFx2_ASAP7_75t_L g221 ( 
.A(n_59),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_17),
.Y(n_222)
);

BUFx3_ASAP7_75t_L g223 ( 
.A(n_1),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_140),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_149),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_14),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_69),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_43),
.Y(n_228)
);

INVx1_ASAP7_75t_SL g229 ( 
.A(n_20),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_14),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_23),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_68),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_26),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_151),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_223),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_193),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_192),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_202),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_223),
.Y(n_239)
);

INVxp67_ASAP7_75t_SL g240 ( 
.A(n_219),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_222),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_226),
.Y(n_242)
);

INVxp33_ASAP7_75t_SL g243 ( 
.A(n_175),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_231),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_175),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_213),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_168),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_215),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_221),
.Y(n_249)
);

INVxp33_ASAP7_75t_SL g250 ( 
.A(n_233),
.Y(n_250)
);

INVx1_ASAP7_75t_SL g251 ( 
.A(n_231),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_233),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_194),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_180),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_180),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_194),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_180),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_167),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_173),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_230),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_212),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_208),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_212),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_176),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g265 ( 
.A(n_205),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_177),
.Y(n_266)
);

INVxp33_ASAP7_75t_SL g267 ( 
.A(n_229),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_185),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_208),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_169),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_178),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_181),
.Y(n_272)
);

HB1xp67_ASAP7_75t_L g273 ( 
.A(n_169),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_183),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_170),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_184),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_186),
.Y(n_277)
);

INVxp33_ASAP7_75t_SL g278 ( 
.A(n_170),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_247),
.Y(n_279)
);

INVx3_ASAP7_75t_L g280 ( 
.A(n_247),
.Y(n_280)
);

OAI21x1_ASAP7_75t_L g281 ( 
.A1(n_258),
.A2(n_188),
.B(n_172),
.Y(n_281)
);

INVx3_ASAP7_75t_L g282 ( 
.A(n_247),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_247),
.Y(n_283)
);

BUFx6f_ASAP7_75t_L g284 ( 
.A(n_262),
.Y(n_284)
);

HB1xp67_ASAP7_75t_L g285 ( 
.A(n_265),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_254),
.B(n_190),
.Y(n_286)
);

BUFx6f_ASAP7_75t_L g287 ( 
.A(n_262),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_259),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_266),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_272),
.B(n_195),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_274),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_276),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_277),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_241),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_242),
.Y(n_295)
);

BUFx6f_ASAP7_75t_L g296 ( 
.A(n_235),
.Y(n_296)
);

OAI21x1_ASAP7_75t_L g297 ( 
.A1(n_239),
.A2(n_188),
.B(n_172),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_240),
.Y(n_298)
);

AND2x4_ASAP7_75t_L g299 ( 
.A(n_255),
.B(n_204),
.Y(n_299)
);

BUFx3_ASAP7_75t_L g300 ( 
.A(n_257),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_237),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_238),
.Y(n_302)
);

INVx3_ASAP7_75t_L g303 ( 
.A(n_246),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_249),
.B(n_264),
.Y(n_304)
);

OA21x2_ASAP7_75t_L g305 ( 
.A1(n_245),
.A2(n_203),
.B(n_201),
.Y(n_305)
);

INVx3_ASAP7_75t_L g306 ( 
.A(n_271),
.Y(n_306)
);

INVx3_ASAP7_75t_L g307 ( 
.A(n_236),
.Y(n_307)
);

BUFx2_ASAP7_75t_L g308 ( 
.A(n_270),
.Y(n_308)
);

INVx4_ASAP7_75t_L g309 ( 
.A(n_248),
.Y(n_309)
);

INVx3_ASAP7_75t_L g310 ( 
.A(n_260),
.Y(n_310)
);

BUFx6f_ASAP7_75t_L g311 ( 
.A(n_278),
.Y(n_311)
);

BUFx6f_ASAP7_75t_L g312 ( 
.A(n_273),
.Y(n_312)
);

INVx3_ASAP7_75t_L g313 ( 
.A(n_251),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_252),
.Y(n_314)
);

AND2x2_ASAP7_75t_L g315 ( 
.A(n_269),
.B(n_171),
.Y(n_315)
);

BUFx8_ASAP7_75t_L g316 ( 
.A(n_269),
.Y(n_316)
);

NAND2xp33_ASAP7_75t_L g317 ( 
.A(n_270),
.B(n_171),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_275),
.Y(n_318)
);

AND2x4_ASAP7_75t_L g319 ( 
.A(n_275),
.B(n_204),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_243),
.Y(n_320)
);

BUFx6f_ASAP7_75t_L g321 ( 
.A(n_250),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_268),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_267),
.Y(n_323)
);

BUFx6f_ASAP7_75t_L g324 ( 
.A(n_253),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_263),
.B(n_207),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_256),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_256),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_294),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_294),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_308),
.B(n_244),
.Y(n_330)
);

INVx3_ASAP7_75t_L g331 ( 
.A(n_284),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_308),
.B(n_244),
.Y(n_332)
);

INVxp67_ASAP7_75t_L g333 ( 
.A(n_285),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_284),
.Y(n_334)
);

INVx3_ASAP7_75t_L g335 ( 
.A(n_284),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_294),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_319),
.A2(n_174),
.B1(n_209),
.B2(n_232),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_284),
.Y(n_338)
);

BUFx3_ASAP7_75t_L g339 ( 
.A(n_284),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_295),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_309),
.B(n_220),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_298),
.B(n_174),
.Y(n_342)
);

INVxp67_ASAP7_75t_L g343 ( 
.A(n_285),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_295),
.Y(n_344)
);

NAND2xp33_ASAP7_75t_SL g345 ( 
.A(n_309),
.B(n_261),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_295),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_319),
.A2(n_225),
.B1(n_227),
.B2(n_228),
.Y(n_347)
);

INVx3_ASAP7_75t_L g348 ( 
.A(n_284),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_284),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_281),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_288),
.Y(n_351)
);

AND2x2_ASAP7_75t_L g352 ( 
.A(n_291),
.B(n_292),
.Y(n_352)
);

OAI22xp33_ASAP7_75t_R g353 ( 
.A1(n_320),
.A2(n_314),
.B1(n_318),
.B2(n_286),
.Y(n_353)
);

INVx3_ASAP7_75t_L g354 ( 
.A(n_287),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_304),
.B(n_179),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_288),
.Y(n_356)
);

BUFx4f_ASAP7_75t_L g357 ( 
.A(n_305),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_289),
.Y(n_358)
);

HB1xp67_ASAP7_75t_L g359 ( 
.A(n_315),
.Y(n_359)
);

AND2x6_ASAP7_75t_L g360 ( 
.A(n_306),
.B(n_168),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_281),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_289),
.Y(n_362)
);

BUFx2_ASAP7_75t_L g363 ( 
.A(n_315),
.Y(n_363)
);

INVxp67_ASAP7_75t_L g364 ( 
.A(n_313),
.Y(n_364)
);

BUFx6f_ASAP7_75t_L g365 ( 
.A(n_287),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_287),
.Y(n_366)
);

BUFx6f_ASAP7_75t_L g367 ( 
.A(n_287),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_281),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_287),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_293),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_293),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_287),
.Y(n_372)
);

AND2x2_ASAP7_75t_L g373 ( 
.A(n_291),
.B(n_261),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_291),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_292),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_292),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_296),
.Y(n_377)
);

INVx1_ASAP7_75t_SL g378 ( 
.A(n_313),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_296),
.Y(n_379)
);

AND2x2_ASAP7_75t_L g380 ( 
.A(n_298),
.B(n_182),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_287),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_296),
.Y(n_382)
);

INVx3_ASAP7_75t_L g383 ( 
.A(n_280),
.Y(n_383)
);

HB1xp67_ASAP7_75t_L g384 ( 
.A(n_315),
.Y(n_384)
);

BUFx8_ASAP7_75t_L g385 ( 
.A(n_321),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_296),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_296),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_296),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_296),
.Y(n_389)
);

INVx3_ASAP7_75t_L g390 ( 
.A(n_280),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_298),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_L g392 ( 
.A1(n_319),
.A2(n_234),
.B1(n_224),
.B2(n_218),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_290),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_326),
.A2(n_217),
.B1(n_216),
.B2(n_214),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_SL g395 ( 
.A(n_357),
.B(n_311),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_352),
.Y(n_396)
);

INVxp67_ASAP7_75t_L g397 ( 
.A(n_330),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_328),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_378),
.B(n_307),
.Y(n_399)
);

INVx2_ASAP7_75t_SL g400 ( 
.A(n_373),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_355),
.B(n_306),
.Y(n_401)
);

NAND3xp33_ASAP7_75t_L g402 ( 
.A(n_333),
.B(n_304),
.C(n_320),
.Y(n_402)
);

INVxp33_ASAP7_75t_L g403 ( 
.A(n_330),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_393),
.B(n_380),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_380),
.B(n_306),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_364),
.B(n_306),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_391),
.B(n_307),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_342),
.B(n_307),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_352),
.B(n_307),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_351),
.Y(n_410)
);

NAND2xp33_ASAP7_75t_L g411 ( 
.A(n_341),
.B(n_311),
.Y(n_411)
);

XOR2xp5_ASAP7_75t_L g412 ( 
.A(n_332),
.B(n_324),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_392),
.B(n_310),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_356),
.B(n_310),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_SL g415 ( 
.A(n_385),
.B(n_316),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_358),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_329),
.Y(n_417)
);

OA21x2_ASAP7_75t_L g418 ( 
.A1(n_350),
.A2(n_297),
.B(n_290),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_SL g419 ( 
.A(n_357),
.B(n_311),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_353),
.A2(n_319),
.B1(n_312),
.B2(n_310),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_SL g421 ( 
.A(n_357),
.B(n_311),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_336),
.Y(n_422)
);

INVx8_ASAP7_75t_L g423 ( 
.A(n_360),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_362),
.B(n_310),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_SL g425 ( 
.A(n_385),
.B(n_311),
.Y(n_425)
);

BUFx6f_ASAP7_75t_SL g426 ( 
.A(n_360),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_370),
.B(n_309),
.Y(n_427)
);

BUFx3_ASAP7_75t_L g428 ( 
.A(n_385),
.Y(n_428)
);

NAND2xp33_ASAP7_75t_L g429 ( 
.A(n_341),
.B(n_311),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_340),
.Y(n_430)
);

AND2x2_ASAP7_75t_L g431 ( 
.A(n_343),
.B(n_313),
.Y(n_431)
);

INVxp67_ASAP7_75t_L g432 ( 
.A(n_332),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_371),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_347),
.B(n_312),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_344),
.B(n_309),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_346),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_374),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_375),
.B(n_309),
.Y(n_438)
);

NOR3xp33_ASAP7_75t_L g439 ( 
.A(n_363),
.B(n_317),
.C(n_318),
.Y(n_439)
);

BUFx6f_ASAP7_75t_SL g440 ( 
.A(n_360),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_376),
.B(n_312),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_386),
.Y(n_442)
);

AND2x2_ASAP7_75t_L g443 ( 
.A(n_373),
.B(n_313),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_SL g444 ( 
.A(n_365),
.B(n_311),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_337),
.B(n_312),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_383),
.B(n_312),
.Y(n_446)
);

BUFx6f_ASAP7_75t_L g447 ( 
.A(n_365),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_383),
.Y(n_448)
);

NAND2xp33_ASAP7_75t_L g449 ( 
.A(n_360),
.B(n_321),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_365),
.B(n_321),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_386),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_383),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_390),
.B(n_312),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_390),
.B(n_312),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_390),
.B(n_314),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_377),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_379),
.Y(n_457)
);

AND2x2_ASAP7_75t_L g458 ( 
.A(n_363),
.B(n_313),
.Y(n_458)
);

NOR3xp33_ASAP7_75t_L g459 ( 
.A(n_345),
.B(n_318),
.C(n_303),
.Y(n_459)
);

BUFx6f_ASAP7_75t_L g460 ( 
.A(n_365),
.Y(n_460)
);

NAND2xp33_ASAP7_75t_L g461 ( 
.A(n_360),
.B(n_321),
.Y(n_461)
);

OA21x2_ASAP7_75t_L g462 ( 
.A1(n_350),
.A2(n_297),
.B(n_283),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_331),
.B(n_323),
.Y(n_463)
);

AOI22xp5_ASAP7_75t_L g464 ( 
.A1(n_413),
.A2(n_353),
.B1(n_345),
.B2(n_359),
.Y(n_464)
);

AO22x2_ASAP7_75t_L g465 ( 
.A1(n_412),
.A2(n_327),
.B1(n_326),
.B2(n_319),
.Y(n_465)
);

AND2x4_ASAP7_75t_L g466 ( 
.A(n_443),
.B(n_324),
.Y(n_466)
);

AO22x2_ASAP7_75t_L g467 ( 
.A1(n_397),
.A2(n_327),
.B1(n_325),
.B2(n_322),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_413),
.B(n_321),
.Y(n_468)
);

AO22x2_ASAP7_75t_L g469 ( 
.A1(n_432),
.A2(n_327),
.B1(n_325),
.B2(n_322),
.Y(n_469)
);

AND2x2_ASAP7_75t_L g470 ( 
.A(n_458),
.B(n_384),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_410),
.Y(n_471)
);

A2O1A1Ixp33_ASAP7_75t_L g472 ( 
.A1(n_445),
.A2(n_286),
.B(n_300),
.C(n_321),
.Y(n_472)
);

HB1xp67_ASAP7_75t_L g473 ( 
.A(n_400),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_399),
.B(n_321),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_416),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_398),
.Y(n_476)
);

AO22x2_ASAP7_75t_L g477 ( 
.A1(n_439),
.A2(n_322),
.B1(n_323),
.B2(n_316),
.Y(n_477)
);

AO22x2_ASAP7_75t_L g478 ( 
.A1(n_404),
.A2(n_323),
.B1(n_316),
.B2(n_324),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_433),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_396),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_SL g481 ( 
.A(n_399),
.B(n_394),
.Y(n_481)
);

AO22x2_ASAP7_75t_L g482 ( 
.A1(n_420),
.A2(n_316),
.B1(n_324),
.B2(n_303),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_405),
.B(n_303),
.Y(n_483)
);

OAI221xp5_ASAP7_75t_L g484 ( 
.A1(n_402),
.A2(n_302),
.B1(n_301),
.B2(n_300),
.C(n_303),
.Y(n_484)
);

AO22x2_ASAP7_75t_L g485 ( 
.A1(n_459),
.A2(n_316),
.B1(n_324),
.B2(n_299),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_428),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_401),
.B(n_301),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_409),
.B(n_302),
.Y(n_488)
);

INVx3_ASAP7_75t_L g489 ( 
.A(n_428),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_417),
.Y(n_490)
);

NAND2xp33_ASAP7_75t_L g491 ( 
.A(n_427),
.B(n_360),
.Y(n_491)
);

AND2x4_ASAP7_75t_L g492 ( 
.A(n_431),
.B(n_324),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_422),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_437),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_398),
.Y(n_495)
);

AO22x2_ASAP7_75t_L g496 ( 
.A1(n_403),
.A2(n_324),
.B1(n_299),
.B2(n_368),
.Y(n_496)
);

AO22x2_ASAP7_75t_L g497 ( 
.A1(n_395),
.A2(n_299),
.B1(n_361),
.B2(n_368),
.Y(n_497)
);

AO22x2_ASAP7_75t_L g498 ( 
.A1(n_395),
.A2(n_299),
.B1(n_361),
.B2(n_300),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_426),
.Y(n_499)
);

AO22x2_ASAP7_75t_L g500 ( 
.A1(n_419),
.A2(n_299),
.B1(n_305),
.B2(n_387),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_430),
.Y(n_501)
);

OR2x2_ASAP7_75t_L g502 ( 
.A(n_455),
.B(n_305),
.Y(n_502)
);

AOI22xp5_ASAP7_75t_L g503 ( 
.A1(n_445),
.A2(n_305),
.B1(n_388),
.B2(n_382),
.Y(n_503)
);

CKINVDCx20_ASAP7_75t_R g504 ( 
.A(n_425),
.Y(n_504)
);

AND2x4_ASAP7_75t_L g505 ( 
.A(n_425),
.B(n_339),
.Y(n_505)
);

OR2x6_ASAP7_75t_L g506 ( 
.A(n_423),
.B(n_297),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_430),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_436),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_426),
.Y(n_509)
);

NAND2xp33_ASAP7_75t_L g510 ( 
.A(n_447),
.B(n_365),
.Y(n_510)
);

AO22x2_ASAP7_75t_L g511 ( 
.A1(n_419),
.A2(n_305),
.B1(n_389),
.B2(n_372),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_436),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_440),
.Y(n_513)
);

AO22x2_ASAP7_75t_L g514 ( 
.A1(n_421),
.A2(n_381),
.B1(n_372),
.B2(n_369),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_464),
.B(n_434),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_476),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_SL g517 ( 
.A(n_468),
.B(n_421),
.Y(n_517)
);

NOR2x1_ASAP7_75t_R g518 ( 
.A(n_486),
.B(n_415),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_470),
.B(n_434),
.Y(n_519)
);

BUFx6f_ASAP7_75t_L g520 ( 
.A(n_505),
.Y(n_520)
);

AOI21xp5_ASAP7_75t_L g521 ( 
.A1(n_474),
.A2(n_408),
.B(n_411),
.Y(n_521)
);

OR2x2_ASAP7_75t_L g522 ( 
.A(n_473),
.B(n_463),
.Y(n_522)
);

A2O1A1Ixp33_ASAP7_75t_L g523 ( 
.A1(n_481),
.A2(n_408),
.B(n_414),
.C(n_424),
.Y(n_523)
);

AO32x1_ASAP7_75t_L g524 ( 
.A1(n_495),
.A2(n_508),
.A3(n_507),
.B1(n_501),
.B2(n_512),
.Y(n_524)
);

AOI22x1_ASAP7_75t_L g525 ( 
.A1(n_497),
.A2(n_448),
.B1(n_452),
.B2(n_457),
.Y(n_525)
);

AOI22x1_ASAP7_75t_L g526 ( 
.A1(n_497),
.A2(n_456),
.B1(n_460),
.B2(n_447),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_487),
.B(n_406),
.Y(n_527)
);

AOI21xp5_ASAP7_75t_L g528 ( 
.A1(n_510),
.A2(n_429),
.B(n_407),
.Y(n_528)
);

A2O1A1Ixp33_ASAP7_75t_SL g529 ( 
.A1(n_483),
.A2(n_454),
.B(n_438),
.C(n_435),
.Y(n_529)
);

AOI21x1_ASAP7_75t_L g530 ( 
.A1(n_511),
.A2(n_441),
.B(n_444),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_490),
.Y(n_531)
);

BUFx3_ASAP7_75t_L g532 ( 
.A(n_489),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_471),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_493),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_475),
.Y(n_535)
);

BUFx12f_ASAP7_75t_L g536 ( 
.A(n_499),
.Y(n_536)
);

INVx5_ASAP7_75t_L g537 ( 
.A(n_506),
.Y(n_537)
);

OAI21xp5_ASAP7_75t_L g538 ( 
.A1(n_472),
.A2(n_454),
.B(n_453),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_494),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_480),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_SL g541 ( 
.A(n_502),
.B(n_447),
.Y(n_541)
);

AND2x2_ASAP7_75t_L g542 ( 
.A(n_492),
.B(n_446),
.Y(n_542)
);

INVx11_ASAP7_75t_L g543 ( 
.A(n_509),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_479),
.Y(n_544)
);

OAI22xp5_ASAP7_75t_L g545 ( 
.A1(n_488),
.A2(n_450),
.B1(n_444),
.B2(n_460),
.Y(n_545)
);

AOI22xp5_ASAP7_75t_L g546 ( 
.A1(n_482),
.A2(n_450),
.B1(n_461),
.B2(n_449),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_466),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_467),
.B(n_442),
.Y(n_548)
);

BUFx6f_ASAP7_75t_L g549 ( 
.A(n_506),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_496),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_467),
.B(n_451),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_SL g552 ( 
.A(n_503),
.B(n_447),
.Y(n_552)
);

AOI21xp5_ASAP7_75t_L g553 ( 
.A1(n_491),
.A2(n_460),
.B(n_418),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_469),
.B(n_460),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_469),
.B(n_418),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_465),
.B(n_418),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_533),
.Y(n_557)
);

OAI22xp5_ASAP7_75t_L g558 ( 
.A1(n_515),
.A2(n_482),
.B1(n_484),
.B2(n_504),
.Y(n_558)
);

OAI22xp5_ASAP7_75t_SL g559 ( 
.A1(n_536),
.A2(n_513),
.B1(n_477),
.B2(n_478),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_519),
.B(n_465),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_516),
.Y(n_561)
);

O2A1O1Ixp33_ASAP7_75t_L g562 ( 
.A1(n_523),
.A2(n_331),
.B(n_348),
.C(n_335),
.Y(n_562)
);

AND2x2_ASAP7_75t_L g563 ( 
.A(n_544),
.B(n_496),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_516),
.Y(n_564)
);

NOR2x1_ASAP7_75t_L g565 ( 
.A(n_532),
.B(n_331),
.Y(n_565)
);

OR2x2_ASAP7_75t_L g566 ( 
.A(n_550),
.B(n_556),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_531),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_544),
.B(n_477),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_535),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_SL g570 ( 
.A(n_527),
.B(n_367),
.Y(n_570)
);

AND2x2_ASAP7_75t_L g571 ( 
.A(n_531),
.B(n_498),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_540),
.Y(n_572)
);

BUFx12f_ASAP7_75t_L g573 ( 
.A(n_549),
.Y(n_573)
);

BUFx6f_ASAP7_75t_L g574 ( 
.A(n_549),
.Y(n_574)
);

AND2x4_ASAP7_75t_L g575 ( 
.A(n_537),
.B(n_339),
.Y(n_575)
);

AND2x2_ASAP7_75t_L g576 ( 
.A(n_534),
.B(n_498),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_522),
.B(n_478),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_534),
.B(n_485),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_539),
.B(n_485),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_539),
.Y(n_580)
);

AOI22xp33_ASAP7_75t_L g581 ( 
.A1(n_540),
.A2(n_500),
.B1(n_511),
.B2(n_514),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_548),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_SL g583 ( 
.A(n_520),
.B(n_367),
.Y(n_583)
);

AOI22xp33_ASAP7_75t_L g584 ( 
.A1(n_520),
.A2(n_500),
.B1(n_514),
.B2(n_440),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_543),
.Y(n_585)
);

HB1xp67_ASAP7_75t_L g586 ( 
.A(n_554),
.Y(n_586)
);

OAI21xp5_ASAP7_75t_L g587 ( 
.A1(n_523),
.A2(n_348),
.B(n_335),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_555),
.Y(n_588)
);

OAI22xp5_ASAP7_75t_L g589 ( 
.A1(n_521),
.A2(n_348),
.B1(n_354),
.B2(n_335),
.Y(n_589)
);

BUFx2_ASAP7_75t_L g590 ( 
.A(n_549),
.Y(n_590)
);

AOI22xp33_ASAP7_75t_SL g591 ( 
.A1(n_526),
.A2(n_520),
.B1(n_551),
.B2(n_547),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_532),
.B(n_354),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_524),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_SL g594 ( 
.A(n_520),
.B(n_367),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_585),
.Y(n_595)
);

NOR2xp33_ASAP7_75t_L g596 ( 
.A(n_585),
.B(n_518),
.Y(n_596)
);

AOI21xp5_ASAP7_75t_L g597 ( 
.A1(n_562),
.A2(n_553),
.B(n_517),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_557),
.Y(n_598)
);

OR2x6_ASAP7_75t_L g599 ( 
.A(n_573),
.B(n_549),
.Y(n_599)
);

AOI22xp33_ASAP7_75t_L g600 ( 
.A1(n_558),
.A2(n_542),
.B1(n_525),
.B2(n_552),
.Y(n_600)
);

AND2x4_ASAP7_75t_L g601 ( 
.A(n_590),
.B(n_574),
.Y(n_601)
);

A2O1A1Ixp33_ASAP7_75t_SL g602 ( 
.A1(n_587),
.A2(n_538),
.B(n_528),
.C(n_545),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_567),
.Y(n_603)
);

BUFx6f_ASAP7_75t_SL g604 ( 
.A(n_574),
.Y(n_604)
);

O2A1O1Ixp33_ASAP7_75t_L g605 ( 
.A1(n_570),
.A2(n_529),
.B(n_517),
.C(n_552),
.Y(n_605)
);

INVx3_ASAP7_75t_L g606 ( 
.A(n_575),
.Y(n_606)
);

AND2x4_ASAP7_75t_L g607 ( 
.A(n_590),
.B(n_537),
.Y(n_607)
);

INVx3_ASAP7_75t_L g608 ( 
.A(n_575),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_SL g609 ( 
.A(n_574),
.B(n_537),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_569),
.B(n_537),
.Y(n_610)
);

AOI21xp5_ASAP7_75t_L g611 ( 
.A1(n_589),
.A2(n_529),
.B(n_541),
.Y(n_611)
);

INVx3_ASAP7_75t_SL g612 ( 
.A(n_574),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_567),
.Y(n_613)
);

NAND2x1p5_ASAP7_75t_L g614 ( 
.A(n_575),
.B(n_574),
.Y(n_614)
);

INVx3_ASAP7_75t_L g615 ( 
.A(n_573),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_580),
.B(n_541),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_572),
.Y(n_617)
);

CKINVDCx20_ASAP7_75t_R g618 ( 
.A(n_559),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_580),
.Y(n_619)
);

AOI21xp5_ASAP7_75t_L g620 ( 
.A1(n_583),
.A2(n_546),
.B(n_524),
.Y(n_620)
);

CKINVDCx11_ASAP7_75t_R g621 ( 
.A(n_588),
.Y(n_621)
);

A2O1A1Ixp33_ASAP7_75t_L g622 ( 
.A1(n_591),
.A2(n_423),
.B(n_338),
.C(n_334),
.Y(n_622)
);

INVx1_ASAP7_75t_SL g623 ( 
.A(n_586),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_563),
.B(n_280),
.Y(n_624)
);

OAI22xp5_ASAP7_75t_L g625 ( 
.A1(n_592),
.A2(n_530),
.B1(n_354),
.B2(n_462),
.Y(n_625)
);

OR2x2_ASAP7_75t_SL g626 ( 
.A(n_577),
.B(n_168),
.Y(n_626)
);

AOI21xp5_ASAP7_75t_L g627 ( 
.A1(n_594),
.A2(n_524),
.B(n_423),
.Y(n_627)
);

BUFx2_ASAP7_75t_L g628 ( 
.A(n_565),
.Y(n_628)
);

AOI21xp5_ASAP7_75t_L g629 ( 
.A1(n_588),
.A2(n_462),
.B(n_367),
.Y(n_629)
);

OR2x6_ASAP7_75t_L g630 ( 
.A(n_563),
.B(n_334),
.Y(n_630)
);

AOI21xp5_ASAP7_75t_L g631 ( 
.A1(n_581),
.A2(n_462),
.B(n_367),
.Y(n_631)
);

NAND2x1p5_ASAP7_75t_L g632 ( 
.A(n_564),
.B(n_280),
.Y(n_632)
);

AOI21xp5_ASAP7_75t_L g633 ( 
.A1(n_584),
.A2(n_349),
.B(n_338),
.Y(n_633)
);

BUFx2_ASAP7_75t_L g634 ( 
.A(n_566),
.Y(n_634)
);

BUFx5_ASAP7_75t_L g635 ( 
.A(n_564),
.Y(n_635)
);

OR2x2_ASAP7_75t_L g636 ( 
.A(n_560),
.B(n_282),
.Y(n_636)
);

AOI22xp33_ASAP7_75t_L g637 ( 
.A1(n_568),
.A2(n_381),
.B1(n_369),
.B2(n_366),
.Y(n_637)
);

A2O1A1Ixp33_ASAP7_75t_SL g638 ( 
.A1(n_593),
.A2(n_282),
.B(n_283),
.C(n_279),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_634),
.B(n_566),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_598),
.B(n_571),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_623),
.B(n_571),
.Y(n_641)
);

OAI22xp5_ASAP7_75t_L g642 ( 
.A1(n_600),
.A2(n_579),
.B1(n_578),
.B2(n_576),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_619),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_621),
.B(n_576),
.Y(n_644)
);

AOI21xp5_ASAP7_75t_L g645 ( 
.A1(n_602),
.A2(n_593),
.B(n_582),
.Y(n_645)
);

OR2x2_ASAP7_75t_L g646 ( 
.A(n_630),
.B(n_561),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_595),
.Y(n_647)
);

INVx1_ASAP7_75t_SL g648 ( 
.A(n_612),
.Y(n_648)
);

BUFx2_ASAP7_75t_L g649 ( 
.A(n_615),
.Y(n_649)
);

OR2x2_ASAP7_75t_L g650 ( 
.A(n_630),
.B(n_561),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_617),
.B(n_0),
.Y(n_651)
);

AND2x2_ASAP7_75t_L g652 ( 
.A(n_606),
.B(n_0),
.Y(n_652)
);

NAND3xp33_ASAP7_75t_L g653 ( 
.A(n_610),
.B(n_279),
.C(n_168),
.Y(n_653)
);

A2O1A1Ixp33_ASAP7_75t_L g654 ( 
.A1(n_631),
.A2(n_199),
.B(n_189),
.C(n_191),
.Y(n_654)
);

BUFx6f_ASAP7_75t_L g655 ( 
.A(n_607),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_624),
.B(n_1),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_606),
.B(n_2),
.Y(n_657)
);

OAI22xp5_ASAP7_75t_L g658 ( 
.A1(n_626),
.A2(n_206),
.B1(n_196),
.B2(n_197),
.Y(n_658)
);

OAI22xp5_ASAP7_75t_L g659 ( 
.A1(n_622),
.A2(n_210),
.B1(n_198),
.B2(n_200),
.Y(n_659)
);

OAI22xp5_ASAP7_75t_L g660 ( 
.A1(n_618),
.A2(n_211),
.B1(n_187),
.B2(n_366),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_608),
.B(n_2),
.Y(n_661)
);

OAI22xp5_ASAP7_75t_L g662 ( 
.A1(n_615),
.A2(n_349),
.B1(n_282),
.B2(n_5),
.Y(n_662)
);

AND2x2_ASAP7_75t_L g663 ( 
.A(n_608),
.B(n_3),
.Y(n_663)
);

O2A1O1Ixp33_ASAP7_75t_L g664 ( 
.A1(n_605),
.A2(n_282),
.B(n_5),
.C(n_6),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_616),
.Y(n_665)
);

INVx1_ASAP7_75t_SL g666 ( 
.A(n_601),
.Y(n_666)
);

HB1xp67_ASAP7_75t_L g667 ( 
.A(n_625),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_601),
.B(n_4),
.Y(n_668)
);

NOR2xp33_ASAP7_75t_SL g669 ( 
.A(n_596),
.B(n_28),
.Y(n_669)
);

OR2x2_ASAP7_75t_L g670 ( 
.A(n_636),
.B(n_4),
.Y(n_670)
);

O2A1O1Ixp33_ASAP7_75t_L g671 ( 
.A1(n_638),
.A2(n_7),
.B(n_8),
.C(n_10),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_628),
.B(n_7),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_599),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_607),
.B(n_8),
.Y(n_674)
);

CKINVDCx6p67_ASAP7_75t_R g675 ( 
.A(n_599),
.Y(n_675)
);

AND2x2_ASAP7_75t_L g676 ( 
.A(n_614),
.B(n_635),
.Y(n_676)
);

AND2x2_ASAP7_75t_L g677 ( 
.A(n_635),
.B(n_10),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_SL g678 ( 
.A(n_635),
.B(n_11),
.Y(n_678)
);

OA222x2_ASAP7_75t_L g679 ( 
.A1(n_670),
.A2(n_613),
.B1(n_603),
.B2(n_620),
.C1(n_611),
.C2(n_597),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_665),
.Y(n_680)
);

AOI22xp33_ASAP7_75t_L g681 ( 
.A1(n_642),
.A2(n_658),
.B1(n_641),
.B2(n_650),
.Y(n_681)
);

AOI22xp33_ASAP7_75t_L g682 ( 
.A1(n_646),
.A2(n_637),
.B1(n_633),
.B2(n_635),
.Y(n_682)
);

AOI22xp33_ASAP7_75t_L g683 ( 
.A1(n_640),
.A2(n_644),
.B1(n_667),
.B2(n_643),
.Y(n_683)
);

AOI22xp33_ASAP7_75t_L g684 ( 
.A1(n_667),
.A2(n_635),
.B1(n_627),
.B2(n_609),
.Y(n_684)
);

BUFx2_ASAP7_75t_L g685 ( 
.A(n_676),
.Y(n_685)
);

OAI21xp33_ASAP7_75t_L g686 ( 
.A1(n_678),
.A2(n_629),
.B(n_632),
.Y(n_686)
);

AOI22xp33_ASAP7_75t_L g687 ( 
.A1(n_643),
.A2(n_604),
.B1(n_12),
.B2(n_13),
.Y(n_687)
);

HB1xp67_ASAP7_75t_L g688 ( 
.A(n_639),
.Y(n_688)
);

OAI21xp33_ASAP7_75t_L g689 ( 
.A1(n_678),
.A2(n_11),
.B(n_13),
.Y(n_689)
);

OAI22xp33_ASAP7_75t_L g690 ( 
.A1(n_669),
.A2(n_604),
.B1(n_16),
.B2(n_17),
.Y(n_690)
);

OAI22xp5_ASAP7_75t_L g691 ( 
.A1(n_664),
.A2(n_15),
.B1(n_16),
.B2(n_18),
.Y(n_691)
);

AOI22xp33_ASAP7_75t_L g692 ( 
.A1(n_659),
.A2(n_19),
.B1(n_20),
.B2(n_21),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_666),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_645),
.Y(n_694)
);

AOI22xp33_ASAP7_75t_L g695 ( 
.A1(n_662),
.A2(n_19),
.B1(n_21),
.B2(n_22),
.Y(n_695)
);

BUFx12f_ASAP7_75t_L g696 ( 
.A(n_647),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_651),
.Y(n_697)
);

AND2x2_ASAP7_75t_L g698 ( 
.A(n_677),
.B(n_22),
.Y(n_698)
);

AND2x2_ASAP7_75t_L g699 ( 
.A(n_652),
.B(n_23),
.Y(n_699)
);

OAI22xp5_ASAP7_75t_L g700 ( 
.A1(n_656),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_700)
);

AND2x2_ASAP7_75t_L g701 ( 
.A(n_663),
.B(n_24),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_649),
.B(n_25),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_655),
.Y(n_703)
);

OAI22xp33_ASAP7_75t_L g704 ( 
.A1(n_674),
.A2(n_27),
.B1(n_29),
.B2(n_30),
.Y(n_704)
);

BUFx3_ASAP7_75t_L g705 ( 
.A(n_655),
.Y(n_705)
);

OAI22xp5_ASAP7_75t_L g706 ( 
.A1(n_654),
.A2(n_27),
.B1(n_31),
.B2(n_32),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_648),
.B(n_33),
.Y(n_707)
);

OAI22xp5_ASAP7_75t_SL g708 ( 
.A1(n_673),
.A2(n_35),
.B1(n_36),
.B2(n_37),
.Y(n_708)
);

INVx3_ASAP7_75t_L g709 ( 
.A(n_705),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_680),
.Y(n_710)
);

AOI21xp5_ASAP7_75t_L g711 ( 
.A1(n_689),
.A2(n_654),
.B(n_671),
.Y(n_711)
);

AND2x2_ASAP7_75t_L g712 ( 
.A(n_685),
.B(n_655),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_680),
.Y(n_713)
);

OAI21xp5_ASAP7_75t_L g714 ( 
.A1(n_689),
.A2(n_672),
.B(n_668),
.Y(n_714)
);

O2A1O1Ixp33_ASAP7_75t_SL g715 ( 
.A1(n_702),
.A2(n_657),
.B(n_661),
.C(n_647),
.Y(n_715)
);

AOI211xp5_ASAP7_75t_L g716 ( 
.A1(n_700),
.A2(n_660),
.B(n_673),
.C(n_653),
.Y(n_716)
);

OR2x2_ASAP7_75t_L g717 ( 
.A(n_688),
.B(n_655),
.Y(n_717)
);

O2A1O1Ixp33_ASAP7_75t_SL g718 ( 
.A1(n_700),
.A2(n_675),
.B(n_40),
.C(n_41),
.Y(n_718)
);

AND2x2_ASAP7_75t_L g719 ( 
.A(n_685),
.B(n_675),
.Y(n_719)
);

OR2x2_ASAP7_75t_L g720 ( 
.A(n_693),
.B(n_38),
.Y(n_720)
);

AND2x2_ASAP7_75t_L g721 ( 
.A(n_679),
.B(n_44),
.Y(n_721)
);

AND2x2_ASAP7_75t_L g722 ( 
.A(n_679),
.B(n_47),
.Y(n_722)
);

A2O1A1Ixp33_ASAP7_75t_L g723 ( 
.A1(n_691),
.A2(n_49),
.B(n_50),
.C(n_51),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_694),
.Y(n_724)
);

NOR2x1_ASAP7_75t_SL g725 ( 
.A(n_705),
.B(n_53),
.Y(n_725)
);

NAND3xp33_ASAP7_75t_L g726 ( 
.A(n_694),
.B(n_54),
.C(n_55),
.Y(n_726)
);

AND2x2_ASAP7_75t_L g727 ( 
.A(n_703),
.B(n_56),
.Y(n_727)
);

HB1xp67_ASAP7_75t_L g728 ( 
.A(n_697),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_693),
.Y(n_729)
);

A2O1A1Ixp33_ASAP7_75t_L g730 ( 
.A1(n_697),
.A2(n_706),
.B(n_698),
.C(n_681),
.Y(n_730)
);

AOI22xp33_ASAP7_75t_L g731 ( 
.A1(n_721),
.A2(n_708),
.B1(n_683),
.B2(n_690),
.Y(n_731)
);

OR2x2_ASAP7_75t_L g732 ( 
.A(n_717),
.B(n_703),
.Y(n_732)
);

AND2x2_ASAP7_75t_L g733 ( 
.A(n_712),
.B(n_705),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_710),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_724),
.Y(n_735)
);

BUFx2_ASAP7_75t_L g736 ( 
.A(n_724),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_710),
.B(n_698),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_713),
.Y(n_738)
);

OR2x2_ASAP7_75t_L g739 ( 
.A(n_717),
.B(n_684),
.Y(n_739)
);

HB1xp67_ASAP7_75t_L g740 ( 
.A(n_713),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_728),
.B(n_699),
.Y(n_741)
);

AND2x2_ASAP7_75t_L g742 ( 
.A(n_712),
.B(n_699),
.Y(n_742)
);

NOR2x1_ASAP7_75t_SL g743 ( 
.A(n_719),
.B(n_696),
.Y(n_743)
);

INVx4_ASAP7_75t_L g744 ( 
.A(n_721),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_729),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_729),
.Y(n_746)
);

AOI21xp5_ASAP7_75t_L g747 ( 
.A1(n_731),
.A2(n_722),
.B(n_718),
.Y(n_747)
);

O2A1O1Ixp33_ASAP7_75t_L g748 ( 
.A1(n_741),
.A2(n_730),
.B(n_714),
.C(n_715),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_745),
.Y(n_749)
);

INVx1_ASAP7_75t_SL g750 ( 
.A(n_742),
.Y(n_750)
);

INVx1_ASAP7_75t_SL g751 ( 
.A(n_742),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_736),
.Y(n_752)
);

AOI21x1_ASAP7_75t_L g753 ( 
.A1(n_736),
.A2(n_722),
.B(n_719),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_740),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_746),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_746),
.Y(n_756)
);

HB1xp67_ASAP7_75t_L g757 ( 
.A(n_734),
.Y(n_757)
);

OR2x2_ASAP7_75t_L g758 ( 
.A(n_744),
.B(n_709),
.Y(n_758)
);

HB1xp67_ASAP7_75t_L g759 ( 
.A(n_757),
.Y(n_759)
);

AND2x4_ASAP7_75t_SL g760 ( 
.A(n_754),
.B(n_744),
.Y(n_760)
);

OR2x2_ASAP7_75t_L g761 ( 
.A(n_750),
.B(n_737),
.Y(n_761)
);

AND2x2_ASAP7_75t_L g762 ( 
.A(n_751),
.B(n_744),
.Y(n_762)
);

AND2x2_ASAP7_75t_L g763 ( 
.A(n_753),
.B(n_743),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_749),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_747),
.B(n_739),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_755),
.Y(n_766)
);

AND2x2_ASAP7_75t_L g767 ( 
.A(n_758),
.B(n_743),
.Y(n_767)
);

INVx2_ASAP7_75t_SL g768 ( 
.A(n_758),
.Y(n_768)
);

OA21x2_ASAP7_75t_L g769 ( 
.A1(n_765),
.A2(n_752),
.B(n_756),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_764),
.Y(n_770)
);

NAND4xp25_ASAP7_75t_L g771 ( 
.A(n_762),
.B(n_748),
.C(n_711),
.D(n_716),
.Y(n_771)
);

AND2x2_ASAP7_75t_L g772 ( 
.A(n_762),
.B(n_752),
.Y(n_772)
);

OR2x2_ASAP7_75t_L g773 ( 
.A(n_761),
.B(n_757),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_759),
.Y(n_774)
);

OAI22xp5_ASAP7_75t_L g775 ( 
.A1(n_760),
.A2(n_739),
.B1(n_709),
.B2(n_733),
.Y(n_775)
);

INVxp67_ASAP7_75t_SL g776 ( 
.A(n_769),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_774),
.Y(n_777)
);

OAI21xp33_ASAP7_75t_L g778 ( 
.A1(n_771),
.A2(n_768),
.B(n_760),
.Y(n_778)
);

AND2x2_ASAP7_75t_L g779 ( 
.A(n_772),
.B(n_767),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_769),
.B(n_759),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_770),
.Y(n_781)
);

NOR2xp67_ASAP7_75t_L g782 ( 
.A(n_779),
.B(n_773),
.Y(n_782)
);

INVx1_ASAP7_75t_SL g783 ( 
.A(n_780),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_776),
.Y(n_784)
);

INVx1_ASAP7_75t_SL g785 ( 
.A(n_777),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_776),
.Y(n_786)
);

HB1xp67_ASAP7_75t_L g787 ( 
.A(n_781),
.Y(n_787)
);

INVx1_ASAP7_75t_SL g788 ( 
.A(n_778),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_776),
.Y(n_789)
);

INVx2_ASAP7_75t_SL g790 ( 
.A(n_780),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_776),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_787),
.Y(n_792)
);

OAI22xp5_ASAP7_75t_L g793 ( 
.A1(n_782),
.A2(n_783),
.B1(n_788),
.B2(n_789),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_785),
.B(n_768),
.Y(n_794)
);

AOI332xp33_ASAP7_75t_L g795 ( 
.A1(n_784),
.A2(n_766),
.A3(n_763),
.B1(n_695),
.B2(n_692),
.B3(n_701),
.C1(n_687),
.C2(n_775),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_787),
.Y(n_796)
);

OAI22xp5_ASAP7_75t_L g797 ( 
.A1(n_791),
.A2(n_696),
.B1(n_733),
.B2(n_723),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_792),
.Y(n_798)
);

INVxp67_ASAP7_75t_L g799 ( 
.A(n_793),
.Y(n_799)
);

NOR2xp33_ASAP7_75t_L g800 ( 
.A(n_794),
.B(n_790),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_796),
.Y(n_801)
);

NOR2xp33_ASAP7_75t_L g802 ( 
.A(n_799),
.B(n_790),
.Y(n_802)
);

NOR3xp33_ASAP7_75t_L g803 ( 
.A(n_800),
.B(n_786),
.C(n_797),
.Y(n_803)
);

NAND2xp33_ASAP7_75t_SL g804 ( 
.A(n_802),
.B(n_798),
.Y(n_804)
);

AND2x2_ASAP7_75t_L g805 ( 
.A(n_803),
.B(n_801),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_802),
.Y(n_806)
);

AOI211x1_ASAP7_75t_L g807 ( 
.A1(n_805),
.A2(n_795),
.B(n_701),
.C(n_707),
.Y(n_807)
);

AOI221xp5_ASAP7_75t_L g808 ( 
.A1(n_804),
.A2(n_704),
.B1(n_726),
.B2(n_708),
.C(n_735),
.Y(n_808)
);

BUFx2_ASAP7_75t_L g809 ( 
.A(n_806),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_809),
.B(n_738),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_807),
.Y(n_811)
);

NAND3xp33_ASAP7_75t_SL g812 ( 
.A(n_808),
.B(n_720),
.C(n_727),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_810),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_SL g814 ( 
.A(n_811),
.B(n_727),
.Y(n_814)
);

NOR3xp33_ASAP7_75t_L g815 ( 
.A(n_812),
.B(n_720),
.C(n_735),
.Y(n_815)
);

NOR2x1_ASAP7_75t_L g816 ( 
.A(n_811),
.B(n_709),
.Y(n_816)
);

NOR2x1p5_ASAP7_75t_L g817 ( 
.A(n_810),
.B(n_732),
.Y(n_817)
);

NAND4xp75_ASAP7_75t_L g818 ( 
.A(n_811),
.B(n_725),
.C(n_738),
.D(n_60),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_810),
.Y(n_819)
);

OR2x2_ASAP7_75t_L g820 ( 
.A(n_819),
.B(n_732),
.Y(n_820)
);

AOI221xp5_ASAP7_75t_L g821 ( 
.A1(n_814),
.A2(n_686),
.B1(n_725),
.B2(n_682),
.C(n_63),
.Y(n_821)
);

AOI22xp33_ASAP7_75t_L g822 ( 
.A1(n_813),
.A2(n_686),
.B1(n_58),
.B2(n_62),
.Y(n_822)
);

INVx1_ASAP7_75t_SL g823 ( 
.A(n_816),
.Y(n_823)
);

OAI22xp33_ASAP7_75t_L g824 ( 
.A1(n_818),
.A2(n_57),
.B1(n_64),
.B2(n_65),
.Y(n_824)
);

NAND3x1_ASAP7_75t_L g825 ( 
.A(n_815),
.B(n_66),
.C(n_67),
.Y(n_825)
);

AOI22xp5_ASAP7_75t_L g826 ( 
.A1(n_817),
.A2(n_70),
.B1(n_71),
.B2(n_72),
.Y(n_826)
);

OAI221xp5_ASAP7_75t_L g827 ( 
.A1(n_816),
.A2(n_73),
.B1(n_75),
.B2(n_77),
.C(n_78),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_820),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_823),
.Y(n_829)
);

HB1xp67_ASAP7_75t_L g830 ( 
.A(n_825),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_826),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_824),
.Y(n_832)
);

INVx4_ASAP7_75t_L g833 ( 
.A(n_827),
.Y(n_833)
);

BUFx6f_ASAP7_75t_L g834 ( 
.A(n_822),
.Y(n_834)
);

AOI22xp5_ASAP7_75t_L g835 ( 
.A1(n_821),
.A2(n_79),
.B1(n_81),
.B2(n_82),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_820),
.Y(n_836)
);

INVx2_ASAP7_75t_L g837 ( 
.A(n_825),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_820),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_825),
.Y(n_839)
);

OR2x6_ASAP7_75t_L g840 ( 
.A(n_829),
.B(n_83),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_830),
.B(n_85),
.Y(n_841)
);

NAND3xp33_ASAP7_75t_SL g842 ( 
.A(n_837),
.B(n_87),
.C(n_89),
.Y(n_842)
);

NAND5xp2_ASAP7_75t_L g843 ( 
.A(n_828),
.B(n_90),
.C(n_93),
.D(n_94),
.E(n_97),
.Y(n_843)
);

OA22x2_ASAP7_75t_L g844 ( 
.A1(n_833),
.A2(n_98),
.B1(n_99),
.B2(n_101),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_839),
.Y(n_845)
);

NAND3x1_ASAP7_75t_L g846 ( 
.A(n_836),
.B(n_102),
.C(n_103),
.Y(n_846)
);

NAND4xp75_ASAP7_75t_L g847 ( 
.A(n_838),
.B(n_105),
.C(n_106),
.D(n_107),
.Y(n_847)
);

XNOR2xp5_ASAP7_75t_L g848 ( 
.A(n_846),
.B(n_832),
.Y(n_848)
);

NAND4xp25_ASAP7_75t_SL g849 ( 
.A(n_845),
.B(n_835),
.C(n_831),
.D(n_834),
.Y(n_849)
);

NOR4xp25_ASAP7_75t_L g850 ( 
.A(n_841),
.B(n_834),
.C(n_109),
.D(n_110),
.Y(n_850)
);

OAI211xp5_ASAP7_75t_L g851 ( 
.A1(n_842),
.A2(n_108),
.B(n_111),
.C(n_112),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_844),
.Y(n_852)
);

XNOR2xp5_ASAP7_75t_L g853 ( 
.A(n_840),
.B(n_115),
.Y(n_853)
);

OAI22xp5_ASAP7_75t_L g854 ( 
.A1(n_852),
.A2(n_847),
.B1(n_843),
.B2(n_119),
.Y(n_854)
);

OAI22xp5_ASAP7_75t_L g855 ( 
.A1(n_848),
.A2(n_116),
.B1(n_118),
.B2(n_120),
.Y(n_855)
);

AOI221xp5_ASAP7_75t_L g856 ( 
.A1(n_849),
.A2(n_121),
.B1(n_122),
.B2(n_123),
.C(n_124),
.Y(n_856)
);

AOI22xp5_ASAP7_75t_L g857 ( 
.A1(n_854),
.A2(n_853),
.B1(n_851),
.B2(n_850),
.Y(n_857)
);

NAND4xp25_ASAP7_75t_SL g858 ( 
.A(n_857),
.B(n_856),
.C(n_855),
.D(n_129),
.Y(n_858)
);

AOI31xp67_ASAP7_75t_L g859 ( 
.A1(n_858),
.A2(n_125),
.A3(n_126),
.B(n_132),
.Y(n_859)
);

NAND3xp33_ASAP7_75t_L g860 ( 
.A(n_858),
.B(n_134),
.C(n_136),
.Y(n_860)
);

NAND2xp33_ASAP7_75t_L g861 ( 
.A(n_860),
.B(n_137),
.Y(n_861)
);

NOR2xp33_ASAP7_75t_L g862 ( 
.A(n_859),
.B(n_138),
.Y(n_862)
);

OR2x6_ASAP7_75t_L g863 ( 
.A(n_862),
.B(n_139),
.Y(n_863)
);

AOI221xp5_ASAP7_75t_L g864 ( 
.A1(n_863),
.A2(n_861),
.B1(n_143),
.B2(n_145),
.C(n_148),
.Y(n_864)
);

AOI211xp5_ASAP7_75t_L g865 ( 
.A1(n_864),
.A2(n_142),
.B(n_150),
.C(n_154),
.Y(n_865)
);


endmodule