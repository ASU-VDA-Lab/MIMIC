module fake_jpeg_1099_n_144 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_144);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_144;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_L g12 ( 
.A(n_0),
.B(n_6),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_9),
.Y(n_13)
);

INVx3_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_2),
.B(n_8),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_8),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_24),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_29),
.Y(n_59)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_30),
.Y(n_51)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_31),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_25),
.B(n_5),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_32),
.B(n_45),
.Y(n_64)
);

INVx6_ASAP7_75t_SL g33 ( 
.A(n_27),
.Y(n_33)
);

CKINVDCx6p67_ASAP7_75t_R g53 ( 
.A(n_33),
.Y(n_53)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

INVx2_ASAP7_75t_SL g57 ( 
.A(n_34),
.Y(n_57)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

BUFx10_ASAP7_75t_L g70 ( 
.A(n_35),
.Y(n_70)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

INVx3_ASAP7_75t_SL g62 ( 
.A(n_36),
.Y(n_62)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

AOI21xp5_ASAP7_75t_L g38 ( 
.A1(n_12),
.A2(n_1),
.B(n_2),
.Y(n_38)
);

OR2x2_ASAP7_75t_L g52 ( 
.A(n_38),
.B(n_41),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_14),
.A2(n_1),
.B1(n_5),
.B2(n_7),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_39),
.A2(n_13),
.B1(n_21),
.B2(n_23),
.Y(n_60)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_16),
.A2(n_14),
.B1(n_20),
.B2(n_11),
.Y(n_41)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_42),
.Y(n_71)
);

HB1xp67_ASAP7_75t_L g43 ( 
.A(n_11),
.Y(n_43)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_15),
.B(n_16),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_20),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_46),
.B(n_49),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_22),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_47),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_28),
.B(n_22),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_48),
.B(n_15),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_28),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_23),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_50),
.B(n_21),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_49),
.B(n_13),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_56),
.B(n_61),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_60),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_47),
.B(n_34),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_63),
.B(n_65),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_42),
.B(n_44),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_35),
.A2(n_36),
.B1(n_37),
.B2(n_40),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_67),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_39),
.B(n_29),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_68),
.B(n_69),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_36),
.A2(n_29),
.B1(n_35),
.B2(n_40),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_72),
.Y(n_78)
);

OAI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_41),
.A2(n_36),
.B1(n_40),
.B2(n_37),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_74),
.A2(n_72),
.B(n_67),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_45),
.B(n_50),
.Y(n_76)
);

CKINVDCx14_ASAP7_75t_R g88 ( 
.A(n_76),
.Y(n_88)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_58),
.Y(n_77)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_77),
.Y(n_102)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_62),
.Y(n_79)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_79),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_54),
.B(n_51),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_80),
.B(n_91),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_81),
.B(n_73),
.Y(n_95)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_66),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_85),
.B(n_87),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_57),
.B(n_55),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_86),
.Y(n_97)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_57),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_53),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_89),
.B(n_93),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_52),
.B(n_64),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_53),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_52),
.B(n_74),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_94),
.B(n_60),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_95),
.A2(n_90),
.B1(n_83),
.B2(n_81),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_96),
.B(n_108),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_91),
.B(n_71),
.C(n_75),
.Y(n_99)
);

XOR2x2_ASAP7_75t_L g112 ( 
.A(n_99),
.B(n_100),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_92),
.B(n_84),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_86),
.Y(n_101)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_101),
.Y(n_111)
);

FAx1_ASAP7_75t_SL g105 ( 
.A(n_94),
.B(n_53),
.CI(n_70),
.CON(n_105),
.SN(n_105)
);

OAI32xp33_ASAP7_75t_L g113 ( 
.A1(n_105),
.A2(n_106),
.A3(n_83),
.B1(n_90),
.B2(n_86),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_SL g106 ( 
.A(n_88),
.B(n_75),
.C(n_70),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_80),
.B(n_59),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_109),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_113),
.A2(n_105),
.B(n_95),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_96),
.A2(n_78),
.B1(n_82),
.B2(n_59),
.Y(n_114)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_114),
.Y(n_120)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_102),
.Y(n_115)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_115),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_99),
.B(n_108),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_116),
.B(n_117),
.Y(n_122)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_98),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_104),
.Y(n_118)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_118),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_112),
.B(n_100),
.C(n_103),
.Y(n_121)
);

BUFx2_ASAP7_75t_L g128 ( 
.A(n_121),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_111),
.B(n_107),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_125),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_126),
.A2(n_110),
.B(n_116),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_127),
.A2(n_126),
.B(n_124),
.Y(n_135)
);

INVxp67_ASAP7_75t_SL g129 ( 
.A(n_119),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_129),
.B(n_123),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_120),
.A2(n_95),
.B1(n_110),
.B2(n_105),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_131),
.A2(n_122),
.B1(n_124),
.B2(n_97),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_132),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_128),
.B(n_112),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_133),
.B(n_134),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_135),
.B(n_113),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_138),
.A2(n_130),
.B(n_109),
.Y(n_140)
);

BUFx24_ASAP7_75t_SL g139 ( 
.A(n_136),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_139),
.B(n_140),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_141),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_142),
.B(n_137),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_143),
.B(n_133),
.Y(n_144)
);


endmodule