module fake_aes_8591_n_46 (n_11, n_1, n_2, n_13, n_12, n_6, n_4, n_3, n_9, n_5, n_14, n_7, n_10, n_8, n_0, n_46);
input n_11;
input n_1;
input n_2;
input n_13;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_14;
input n_7;
input n_10;
input n_8;
input n_0;
output n_46;
wire n_45;
wire n_20;
wire n_38;
wire n_44;
wire n_36;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_41;
wire n_35;
wire n_17;
wire n_15;
wire n_42;
wire n_24;
wire n_19;
wire n_27;
wire n_21;
wire n_43;
wire n_40;
wire n_29;
wire n_39;
INVx2_ASAP7_75t_L g15 ( .A(n_14), .Y(n_15) );
CKINVDCx6p67_ASAP7_75t_R g16 ( .A(n_13), .Y(n_16) );
NOR2xp33_ASAP7_75t_L g17 ( .A(n_0), .B(n_5), .Y(n_17) );
INVx1_ASAP7_75t_L g18 ( .A(n_11), .Y(n_18) );
INVx5_ASAP7_75t_L g19 ( .A(n_6), .Y(n_19) );
INVx2_ASAP7_75t_L g20 ( .A(n_8), .Y(n_20) );
XNOR2x1_ASAP7_75t_L g21 ( .A(n_7), .B(n_10), .Y(n_21) );
INVx2_ASAP7_75t_L g22 ( .A(n_2), .Y(n_22) );
AND2x2_ASAP7_75t_L g23 ( .A(n_22), .B(n_0), .Y(n_23) );
NAND2xp5_ASAP7_75t_L g24 ( .A(n_15), .B(n_1), .Y(n_24) );
NOR2xp33_ASAP7_75t_R g25 ( .A(n_16), .B(n_9), .Y(n_25) );
INVx2_ASAP7_75t_L g26 ( .A(n_20), .Y(n_26) );
INVx2_ASAP7_75t_L g27 ( .A(n_26), .Y(n_27) );
OR2x6_ASAP7_75t_L g28 ( .A(n_23), .B(n_18), .Y(n_28) );
INVx1_ASAP7_75t_L g29 ( .A(n_24), .Y(n_29) );
AOI22xp33_ASAP7_75t_SL g30 ( .A1(n_29), .A2(n_21), .B1(n_25), .B2(n_24), .Y(n_30) );
INVx1_ASAP7_75t_L g31 ( .A(n_27), .Y(n_31) );
OR2x4_ASAP7_75t_L g32 ( .A(n_30), .B(n_28), .Y(n_32) );
OR2x2_ASAP7_75t_L g33 ( .A(n_31), .B(n_28), .Y(n_33) );
AOI22xp5_ASAP7_75t_L g34 ( .A1(n_32), .A2(n_18), .B1(n_17), .B2(n_19), .Y(n_34) );
AOI21xp5_ASAP7_75t_L g35 ( .A1(n_33), .A2(n_19), .B(n_12), .Y(n_35) );
CKINVDCx20_ASAP7_75t_R g36 ( .A(n_34), .Y(n_36) );
INVx2_ASAP7_75t_L g37 ( .A(n_35), .Y(n_37) );
INVx1_ASAP7_75t_L g38 ( .A(n_34), .Y(n_38) );
NAND3xp33_ASAP7_75t_L g39 ( .A(n_38), .B(n_19), .C(n_2), .Y(n_39) );
INVx1_ASAP7_75t_L g40 ( .A(n_36), .Y(n_40) );
NAND3xp33_ASAP7_75t_L g41 ( .A(n_37), .B(n_1), .C(n_3), .Y(n_41) );
OAI22xp5_ASAP7_75t_L g42 ( .A1(n_39), .A2(n_37), .B1(n_4), .B2(n_3), .Y(n_42) );
INVx1_ASAP7_75t_L g43 ( .A(n_41), .Y(n_43) );
INVx1_ASAP7_75t_L g44 ( .A(n_40), .Y(n_44) );
INVx1_ASAP7_75t_SL g45 ( .A(n_44), .Y(n_45) );
AOI22xp5_ASAP7_75t_L g46 ( .A1(n_45), .A2(n_43), .B1(n_42), .B2(n_4), .Y(n_46) );
endmodule