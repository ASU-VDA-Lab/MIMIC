module fake_jpeg_7375_n_319 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_319);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_319;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_6),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx4f_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_SL g24 ( 
.A(n_3),
.B(n_11),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_15),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_5),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_18),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_34),
.B(n_36),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_29),
.B(n_0),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_35),
.B(n_42),
.Y(n_45)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx2_ASAP7_75t_R g39 ( 
.A(n_18),
.Y(n_39)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_39),
.Y(n_56)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_29),
.B(n_0),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_43),
.B(n_20),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_35),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_48),
.B(n_55),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_35),
.B(n_24),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_51),
.B(n_57),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_35),
.B(n_32),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_52),
.B(n_54),
.Y(n_65)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_53),
.B(n_43),
.Y(n_80)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_42),
.B(n_24),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_42),
.B(n_22),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_60),
.Y(n_74)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_61),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_34),
.B(n_22),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_62),
.B(n_28),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_63),
.Y(n_76)
);

HB1xp67_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_64),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_47),
.A2(n_32),
.B1(n_19),
.B2(n_33),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_66),
.Y(n_110)
);

BUFx2_ASAP7_75t_L g69 ( 
.A(n_59),
.Y(n_69)
);

HB1xp67_ASAP7_75t_L g90 ( 
.A(n_69),
.Y(n_90)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_50),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_70),
.B(n_87),
.Y(n_94)
);

INVx1_ASAP7_75t_SL g73 ( 
.A(n_49),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_73),
.B(n_78),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_45),
.A2(n_40),
.B1(n_34),
.B2(n_43),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_75),
.A2(n_79),
.B1(n_20),
.B2(n_19),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_61),
.Y(n_77)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_77),
.Y(n_98)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_46),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_48),
.A2(n_40),
.B1(n_32),
.B2(n_33),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_80),
.B(n_86),
.Y(n_95)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_46),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_81),
.B(n_83),
.Y(n_116)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_62),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_58),
.Y(n_84)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_84),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_45),
.B(n_36),
.C(n_43),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_85),
.B(n_56),
.C(n_41),
.Y(n_106)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_57),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_55),
.B(n_28),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_88),
.B(n_89),
.Y(n_112)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_52),
.Y(n_89)
);

OA22x2_ASAP7_75t_L g91 ( 
.A1(n_74),
.A2(n_63),
.B1(n_60),
.B2(n_44),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_91),
.A2(n_100),
.B1(n_50),
.B2(n_38),
.Y(n_144)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_84),
.Y(n_92)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_92),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_86),
.A2(n_40),
.B1(n_83),
.B2(n_36),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_93),
.A2(n_104),
.B1(n_108),
.B2(n_113),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_77),
.A2(n_56),
.B(n_54),
.Y(n_96)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_96),
.B(n_71),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_65),
.B(n_51),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_97),
.B(n_103),
.Y(n_117)
);

O2A1O1Ixp33_ASAP7_75t_L g100 ( 
.A1(n_75),
.A2(n_63),
.B(n_60),
.C(n_44),
.Y(n_100)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_87),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_102),
.B(n_97),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_65),
.B(n_53),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_67),
.A2(n_33),
.B1(n_30),
.B2(n_19),
.Y(n_104)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_73),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_105),
.B(n_115),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_106),
.B(n_41),
.Y(n_140)
);

OR2x2_ASAP7_75t_L g107 ( 
.A(n_72),
.B(n_50),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_107),
.B(n_114),
.Y(n_138)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_70),
.Y(n_111)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_111),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_67),
.A2(n_30),
.B1(n_20),
.B2(n_59),
.Y(n_113)
);

AND2x2_ASAP7_75t_SL g114 ( 
.A(n_89),
.B(n_41),
.Y(n_114)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_70),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_110),
.A2(n_85),
.B1(n_76),
.B2(n_74),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_118),
.A2(n_139),
.B1(n_144),
.B2(n_95),
.Y(n_164)
);

AND2x2_ASAP7_75t_SL g119 ( 
.A(n_103),
.B(n_82),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_119),
.B(n_126),
.C(n_140),
.Y(n_152)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_101),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_120),
.B(n_124),
.Y(n_165)
);

OAI22x1_ASAP7_75t_L g121 ( 
.A1(n_110),
.A2(n_68),
.B1(n_76),
.B2(n_82),
.Y(n_121)
);

AOI22x1_ASAP7_75t_L g163 ( 
.A1(n_121),
.A2(n_91),
.B1(n_90),
.B2(n_100),
.Y(n_163)
);

NOR2x1_ASAP7_75t_L g122 ( 
.A(n_107),
.B(n_71),
.Y(n_122)
);

OAI21x1_ASAP7_75t_L g153 ( 
.A1(n_122),
.A2(n_126),
.B(n_121),
.Y(n_153)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_101),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_123),
.B(n_125),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_94),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_116),
.Y(n_125)
);

AND2x2_ASAP7_75t_SL g126 ( 
.A(n_98),
.B(n_71),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_114),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_127),
.B(n_135),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_115),
.B(n_68),
.Y(n_130)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_130),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g131 ( 
.A(n_92),
.Y(n_131)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_131),
.Y(n_160)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_109),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_132),
.B(n_109),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_116),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_114),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_136),
.B(n_142),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_99),
.B(n_58),
.Y(n_137)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_137),
.Y(n_162)
);

OAI22xp33_ASAP7_75t_L g139 ( 
.A1(n_98),
.A2(n_59),
.B1(n_69),
.B2(n_30),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_141),
.B(n_96),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_106),
.B(n_41),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_143),
.A2(n_91),
.B(n_108),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_129),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_145),
.B(n_150),
.Y(n_179)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_146),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_147),
.B(n_161),
.C(n_167),
.Y(n_188)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_131),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_148),
.B(n_156),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_128),
.B(n_105),
.Y(n_149)
);

CKINVDCx14_ASAP7_75t_R g187 ( 
.A(n_149),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_139),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_128),
.B(n_134),
.Y(n_151)
);

CKINVDCx14_ASAP7_75t_R g190 ( 
.A(n_151),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_153),
.A2(n_154),
.B(n_152),
.Y(n_205)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_132),
.Y(n_156)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_134),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_157),
.B(n_158),
.Y(n_180)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_144),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_119),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_159),
.B(n_166),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_140),
.B(n_95),
.C(n_102),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_163),
.A2(n_99),
.B1(n_26),
.B2(n_25),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_164),
.A2(n_171),
.B1(n_126),
.B2(n_133),
.Y(n_185)
);

INVx2_ASAP7_75t_SL g166 ( 
.A(n_123),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_SL g167 ( 
.A(n_122),
.B(n_107),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_119),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_169),
.B(n_170),
.Y(n_189)
);

HB1xp67_ASAP7_75t_L g170 ( 
.A(n_118),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_127),
.A2(n_91),
.B1(n_112),
.B2(n_111),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_138),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_172),
.B(n_175),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_138),
.Y(n_175)
);

FAx1_ASAP7_75t_SL g176 ( 
.A(n_117),
.B(n_38),
.CI(n_37),
.CON(n_176),
.SN(n_176)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_176),
.B(n_0),
.Y(n_201)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_156),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_182),
.B(n_200),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_167),
.A2(n_136),
.B(n_143),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_183),
.A2(n_205),
.B(n_154),
.Y(n_206)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_168),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_184),
.B(n_197),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_185),
.A2(n_186),
.B1(n_199),
.B2(n_152),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_158),
.A2(n_143),
.B1(n_141),
.B2(n_117),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_192),
.A2(n_184),
.B1(n_193),
.B2(n_31),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_173),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_193),
.B(n_194),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_165),
.Y(n_194)
);

BUFx4f_ASAP7_75t_SL g195 ( 
.A(n_157),
.Y(n_195)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_195),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_174),
.B(n_29),
.Y(n_196)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_196),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_176),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g198 ( 
.A(n_163),
.B(n_0),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_198),
.A2(n_26),
.B(n_17),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_164),
.A2(n_171),
.B1(n_163),
.B2(n_176),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_166),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_201),
.B(n_202),
.Y(n_228)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_145),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_161),
.B(n_27),
.Y(n_203)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_203),
.Y(n_221)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_155),
.Y(n_204)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_204),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_SL g242 ( 
.A(n_206),
.B(n_198),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_204),
.B(n_162),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_207),
.B(n_219),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_209),
.A2(n_212),
.B1(n_213),
.B2(n_225),
.Y(n_235)
);

NAND3xp33_ASAP7_75t_L g211 ( 
.A(n_186),
.B(n_147),
.C(n_2),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_211),
.B(n_220),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_199),
.A2(n_185),
.B1(n_189),
.B2(n_180),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_205),
.A2(n_160),
.B1(n_148),
.B2(n_16),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_195),
.Y(n_214)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_214),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_216),
.A2(n_217),
.B1(n_230),
.B2(n_16),
.Y(n_232)
);

FAx1_ASAP7_75t_SL g219 ( 
.A(n_188),
.B(n_38),
.CI(n_37),
.CON(n_219),
.SN(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_178),
.Y(n_220)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_181),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_223),
.B(n_226),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_188),
.B(n_160),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_224),
.B(n_229),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_179),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_225),
.B(n_228),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_191),
.B(n_25),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_196),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_227),
.B(n_182),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_183),
.B(n_38),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_198),
.A2(n_31),
.B(n_17),
.Y(n_230)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_232),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_235),
.A2(n_27),
.B1(n_23),
.B2(n_21),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_224),
.B(n_203),
.C(n_202),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_236),
.B(n_238),
.Y(n_267)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_208),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_SL g239 ( 
.A(n_206),
.B(n_197),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_SL g258 ( 
.A(n_239),
.B(n_242),
.Y(n_258)
);

INVxp33_ASAP7_75t_L g240 ( 
.A(n_210),
.Y(n_240)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_240),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_215),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_241),
.B(n_243),
.Y(n_254)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_215),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_212),
.A2(n_200),
.B1(n_190),
.B2(n_187),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_244),
.A2(n_222),
.B1(n_231),
.B2(n_214),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_209),
.B(n_229),
.C(n_221),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_245),
.B(n_247),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_213),
.B(n_177),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_219),
.B(n_177),
.C(n_195),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_248),
.B(n_219),
.Y(n_256)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_249),
.Y(n_260)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_217),
.Y(n_251)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_251),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_252),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_235),
.A2(n_230),
.B1(n_216),
.B2(n_218),
.Y(n_253)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_253),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_256),
.B(n_237),
.C(n_245),
.Y(n_277)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_261),
.Y(n_273)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_249),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_264),
.B(n_266),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_265),
.A2(n_257),
.B1(n_244),
.B2(n_260),
.Y(n_271)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_233),
.Y(n_266)
);

HB1xp67_ASAP7_75t_L g268 ( 
.A(n_239),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_268),
.B(n_247),
.Y(n_275)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_271),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_267),
.B(n_236),
.C(n_248),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_272),
.B(n_280),
.C(n_281),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_SL g274 ( 
.A(n_258),
.B(n_242),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_SL g288 ( 
.A(n_274),
.B(n_21),
.Y(n_288)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_275),
.Y(n_286)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_254),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_276),
.B(n_279),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_277),
.B(n_37),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_262),
.A2(n_246),
.B(n_240),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_278),
.A2(n_9),
.B(n_2),
.Y(n_294)
);

CKINVDCx14_ASAP7_75t_R g279 ( 
.A(n_261),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_259),
.B(n_237),
.C(n_234),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_259),
.B(n_250),
.C(n_37),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_263),
.B(n_255),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_282),
.B(n_27),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_273),
.A2(n_256),
.B1(n_258),
.B2(n_265),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_283),
.A2(n_288),
.B1(n_289),
.B2(n_274),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_SL g287 ( 
.A(n_272),
.B(n_12),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_287),
.B(n_292),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_270),
.A2(n_27),
.B1(n_23),
.B2(n_1),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_290),
.B(n_278),
.C(n_1),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_280),
.B(n_21),
.C(n_23),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_293),
.B(n_1),
.C(n_4),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_294),
.B(n_7),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_L g295 ( 
.A1(n_284),
.A2(n_281),
.B(n_269),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_295),
.B(n_297),
.C(n_298),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_296),
.A2(n_291),
.B1(n_285),
.B2(n_286),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_L g298 ( 
.A1(n_284),
.A2(n_9),
.B(n_3),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_299),
.B(n_300),
.C(n_302),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_290),
.B(n_4),
.C(n_7),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_293),
.B(n_4),
.C(n_7),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_303),
.B(n_301),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_304),
.B(n_305),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_299),
.B(n_289),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_308),
.A2(n_309),
.B(n_8),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_301),
.B(n_283),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_306),
.B(n_288),
.C(n_11),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g313 ( 
.A1(n_310),
.A2(n_312),
.B(n_308),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_SL g314 ( 
.A1(n_313),
.A2(n_311),
.B(n_307),
.Y(n_314)
);

NOR3xp33_ASAP7_75t_L g315 ( 
.A(n_314),
.B(n_8),
.C(n_11),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_L g316 ( 
.A1(n_315),
.A2(n_12),
.B(n_13),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_316),
.B(n_13),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_317),
.B(n_14),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_318),
.A2(n_14),
.B1(n_15),
.B2(n_257),
.Y(n_319)
);


endmodule