module real_jpeg_21536_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_201;
wire n_49;
wire n_114;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_194;
wire n_153;
wire n_104;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_281;
wire n_163;
wire n_276;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_238;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_262;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_195;
wire n_205;
wire n_110;
wire n_258;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_150;
wire n_74;
wire n_32;
wire n_20;
wire n_80;
wire n_228;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_225;
wire n_103;
wire n_259;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_279;
wire n_59;
wire n_169;
wire n_167;
wire n_128;
wire n_216;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_210;
wire n_53;
wire n_127;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_283;
wire n_101;
wire n_274;
wire n_256;
wire n_182;
wire n_273;
wire n_96;
wire n_253;
wire n_269;
wire n_89;

OAI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_0),
.A2(n_27),
.B1(n_31),
.B2(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

OAI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_0),
.A2(n_39),
.B1(n_77),
.B2(n_82),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_0),
.A2(n_34),
.B1(n_35),
.B2(n_39),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_0),
.A2(n_39),
.B1(n_47),
.B2(n_48),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_1),
.A2(n_47),
.B1(n_48),
.B2(n_55),
.Y(n_54)
);

CKINVDCx14_ASAP7_75t_R g55 ( 
.A(n_1),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_1),
.A2(n_27),
.B1(n_31),
.B2(n_55),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_1),
.A2(n_34),
.B1(n_35),
.B2(n_55),
.Y(n_121)
);

BUFx16f_ASAP7_75t_L g77 ( 
.A(n_2),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_3),
.A2(n_77),
.B1(n_82),
.B2(n_153),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_3),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_3),
.A2(n_47),
.B1(n_48),
.B2(n_153),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_3),
.A2(n_27),
.B1(n_31),
.B2(n_153),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_3),
.A2(n_34),
.B1(n_35),
.B2(n_153),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_4),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_4),
.B(n_79),
.Y(n_179)
);

AOI21xp33_ASAP7_75t_L g201 ( 
.A1(n_4),
.A2(n_14),
.B(n_35),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_4),
.A2(n_27),
.B1(n_31),
.B2(n_151),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_4),
.A2(n_61),
.B1(n_65),
.B2(n_210),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_4),
.B(n_183),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_4),
.B(n_47),
.Y(n_234)
);

AOI21xp33_ASAP7_75t_L g238 ( 
.A1(n_4),
.A2(n_47),
.B(n_234),
.Y(n_238)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_5),
.Y(n_64)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_5),
.Y(n_65)
);

BUFx8_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_7),
.A2(n_27),
.B1(n_30),
.B2(n_31),
.Y(n_26)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_7),
.A2(n_30),
.B1(n_34),
.B2(n_35),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_7),
.A2(n_30),
.B1(n_77),
.B2(n_82),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_7),
.A2(n_30),
.B1(n_47),
.B2(n_48),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_8),
.A2(n_77),
.B1(n_82),
.B2(n_99),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_8),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_8),
.A2(n_47),
.B1(n_48),
.B2(n_99),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_8),
.A2(n_34),
.B1(n_35),
.B2(n_99),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_8),
.A2(n_27),
.B1(n_31),
.B2(n_99),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_9),
.A2(n_77),
.B1(n_82),
.B2(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_9),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g147 ( 
.A1(n_9),
.A2(n_47),
.B1(n_48),
.B2(n_131),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_9),
.A2(n_34),
.B1(n_35),
.B2(n_131),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_9),
.A2(n_27),
.B1(n_31),
.B2(n_131),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_10),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_11),
.A2(n_47),
.B1(n_48),
.B2(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_11),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_11),
.A2(n_27),
.B1(n_31),
.B2(n_53),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_11),
.A2(n_34),
.B1(n_35),
.B2(n_53),
.Y(n_159)
);

INVx13_ASAP7_75t_L g46 ( 
.A(n_12),
.Y(n_46)
);

INVx13_ASAP7_75t_L g76 ( 
.A(n_13),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_13),
.A2(n_47),
.B1(n_48),
.B2(n_76),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_14),
.A2(n_34),
.B1(n_35),
.B2(n_36),
.Y(n_33)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

A2O1A1Ixp33_ASAP7_75t_L g41 ( 
.A1(n_14),
.A2(n_31),
.B(n_33),
.C(n_42),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_14),
.B(n_31),
.Y(n_42)
);

INVx11_ASAP7_75t_SL g29 ( 
.A(n_15),
.Y(n_29)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_134),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_133),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_108),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_20),
.B(n_108),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_87),
.B2(n_107),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_57),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_43),
.B(n_56),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_24),
.B(n_43),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_37),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_25),
.A2(n_41),
.B(n_241),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_32),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_26),
.Y(n_144)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_27),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_27),
.A2(n_31),
.B1(n_45),
.B2(n_51),
.Y(n_50)
);

A2O1A1Ixp33_ASAP7_75t_L g200 ( 
.A1(n_27),
.A2(n_36),
.B(n_151),
.C(n_201),
.Y(n_200)
);

NAND2xp33_ASAP7_75t_SL g235 ( 
.A(n_27),
.B(n_45),
.Y(n_235)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

AOI32xp33_ASAP7_75t_L g233 ( 
.A1(n_31),
.A2(n_48),
.A3(n_51),
.B1(n_234),
.B2(n_235),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_32),
.B(n_38),
.Y(n_70)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_33),
.A2(n_41),
.B1(n_69),
.B2(n_95),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_33),
.A2(n_37),
.B(n_95),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_33),
.A2(n_41),
.B1(n_204),
.B2(n_205),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_33),
.B(n_151),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_33),
.A2(n_41),
.B1(n_205),
.B2(n_225),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_33),
.A2(n_41),
.B1(n_225),
.B2(n_241),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_34),
.B(n_63),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_34),
.B(n_214),
.Y(n_213)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_40),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_SL g68 ( 
.A1(n_41),
.A2(n_69),
.B(n_70),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_41),
.A2(n_70),
.B(n_144),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_44),
.A2(n_50),
.B1(n_52),
.B2(n_54),
.Y(n_43)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_44),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_44),
.A2(n_50),
.B1(n_147),
.B2(n_148),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_44),
.A2(n_50),
.B1(n_182),
.B2(n_238),
.Y(n_237)
);

A2O1A1Ixp33_ASAP7_75t_L g44 ( 
.A1(n_45),
.A2(n_47),
.B(n_49),
.C(n_50),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_45),
.B(n_47),
.Y(n_49)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_45),
.Y(n_51)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_47),
.B(n_76),
.Y(n_157)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_48),
.A2(n_78),
.B1(n_150),
.B2(n_157),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_50),
.A2(n_52),
.B(n_103),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_50),
.B(n_106),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_50),
.B(n_126),
.Y(n_168)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_50),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_59),
.B1(n_71),
.B2(n_72),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_68),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_60),
.A2(n_73),
.B1(n_85),
.B2(n_86),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_60),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_60),
.A2(n_68),
.B1(n_86),
.B2(n_113),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_65),
.B(n_66),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_61),
.A2(n_121),
.B(n_122),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_61),
.A2(n_121),
.B1(n_159),
.B2(n_160),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_61),
.A2(n_64),
.B1(n_194),
.B2(n_210),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_61),
.A2(n_93),
.B(n_197),
.Y(n_226)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_62),
.B(n_91),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_62),
.A2(n_193),
.B1(n_195),
.B2(n_196),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_62),
.A2(n_67),
.B(n_123),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_63),
.B(n_67),
.Y(n_93)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_63),
.Y(n_160)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_64),
.B(n_92),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_65),
.A2(n_90),
.B(n_159),
.Y(n_178)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_65),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_65),
.B(n_151),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_67),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_68),
.Y(n_113)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_73),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_SL g73 ( 
.A1(n_74),
.A2(n_80),
.B(n_83),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_74),
.A2(n_98),
.B(n_100),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_74),
.A2(n_98),
.B1(n_130),
.B2(n_132),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_74),
.A2(n_130),
.B1(n_132),
.B2(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_75),
.A2(n_79),
.B1(n_150),
.B2(n_152),
.Y(n_149)
);

O2A1O1Ixp33_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_77),
.B(n_78),
.C(n_79),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_76),
.B(n_77),
.Y(n_78)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_77),
.Y(n_82)
);

HAxp5_ASAP7_75t_SL g150 ( 
.A(n_77),
.B(n_151),
.CON(n_150),
.SN(n_150)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_79),
.B(n_84),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_79),
.B(n_81),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_79),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_81),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_87),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_96),
.C(n_101),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_88),
.B(n_111),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_94),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_89),
.B(n_94),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_93),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_96),
.A2(n_97),
.B1(n_101),
.B2(n_102),
.Y(n_111)
);

CKINVDCx14_ASAP7_75t_R g96 ( 
.A(n_97),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_102),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_104),
.B(n_105),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_104),
.A2(n_125),
.B(n_127),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_104),
.A2(n_167),
.B(n_168),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_104),
.A2(n_181),
.B1(n_183),
.B2(n_184),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_112),
.C(n_114),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_109),
.A2(n_110),
.B1(n_112),
.B2(n_283),
.Y(n_282)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

CKINVDCx14_ASAP7_75t_R g283 ( 
.A(n_112),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_114),
.B(n_282),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_124),
.C(n_128),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_115),
.A2(n_116),
.B1(n_273),
.B2(n_274),
.Y(n_272)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_117),
.B(n_119),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_117),
.A2(n_118),
.B1(n_119),
.B2(n_120),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_118),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_120),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_124),
.A2(n_128),
.B1(n_129),
.B2(n_275),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_124),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_135),
.A2(n_279),
.B(n_284),
.Y(n_134)
);

O2A1O1Ixp33_ASAP7_75t_SL g135 ( 
.A1(n_136),
.A2(n_185),
.B(n_264),
.C(n_278),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_170),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_137),
.B(n_170),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_138),
.A2(n_139),
.B1(n_154),
.B2(n_169),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_SL g139 ( 
.A(n_140),
.B(n_141),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_140),
.B(n_141),
.C(n_169),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_145),
.C(n_149),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_142),
.A2(n_143),
.B1(n_145),
.B2(n_146),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_143),
.Y(n_142)
);

CKINVDCx14_ASAP7_75t_R g145 ( 
.A(n_146),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_147),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_148),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_SL g171 ( 
.A(n_149),
.B(n_172),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_152),
.Y(n_164)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_154),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_161),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_155),
.B(n_162),
.C(n_166),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_158),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_156),
.B(n_158),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_162),
.A2(n_163),
.B1(n_165),
.B2(n_166),
.Y(n_161)
);

CKINVDCx14_ASAP7_75t_R g162 ( 
.A(n_163),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_166),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_173),
.C(n_175),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_171),
.B(n_261),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_173),
.A2(n_174),
.B1(n_175),
.B2(n_176),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_174),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_176),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_179),
.C(n_180),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_177),
.A2(n_178),
.B1(n_179),
.B2(n_252),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_179),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_SL g250 ( 
.A(n_180),
.B(n_251),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_182),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_186),
.B(n_263),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_187),
.A2(n_258),
.B(n_262),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_188),
.A2(n_246),
.B(n_257),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_189),
.A2(n_228),
.B(n_245),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_190),
.A2(n_217),
.B(n_227),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_191),
.A2(n_206),
.B(n_216),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_198),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_192),
.B(n_198),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_194),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_197),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_199),
.A2(n_200),
.B1(n_202),
.B2(n_203),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_200),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_200),
.B(n_202),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_203),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_207),
.A2(n_211),
.B(n_215),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_209),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_208),
.B(n_209),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_212),
.B(n_213),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_219),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_218),
.B(n_219),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_226),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_221),
.A2(n_222),
.B1(n_223),
.B2(n_224),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_221),
.B(n_224),
.C(n_226),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_222),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_224),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_230),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_229),
.B(n_230),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_231),
.A2(n_236),
.B1(n_243),
.B2(n_244),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_231),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_233),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_232),
.B(n_233),
.Y(n_255)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_236),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_237),
.A2(n_239),
.B1(n_240),
.B2(n_242),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_237),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_239),
.B(n_242),
.C(n_243),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_240),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_248),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_247),
.B(n_248),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_249),
.A2(n_250),
.B1(n_253),
.B2(n_254),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_249),
.B(n_255),
.C(n_256),
.Y(n_259)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_254),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_256),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_260),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_259),
.B(n_260),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_266),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_SL g278 ( 
.A(n_265),
.B(n_266),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_267),
.A2(n_268),
.B1(n_276),
.B2(n_277),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_269),
.A2(n_270),
.B1(n_271),
.B2(n_272),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_269),
.B(n_272),
.C(n_277),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_276),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_281),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_280),
.B(n_281),
.Y(n_284)
);


endmodule