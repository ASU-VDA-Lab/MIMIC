module fake_jpeg_9020_n_225 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_225);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_225;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_127;
wire n_154;
wire n_76;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx3_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_15),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_2),
.B(n_14),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_9),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_11),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_9),
.B(n_8),
.Y(n_34)
);

INVx3_ASAP7_75t_SL g35 ( 
.A(n_23),
.Y(n_35)
);

BUFx10_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

NAND2xp33_ASAP7_75t_SL g60 ( 
.A(n_37),
.B(n_17),
.Y(n_60)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

OAI22xp33_ASAP7_75t_L g40 ( 
.A1(n_20),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_40),
.A2(n_18),
.B1(n_28),
.B2(n_22),
.Y(n_56)
);

INVx4_ASAP7_75t_SL g41 ( 
.A(n_26),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_41),
.A2(n_20),
.B1(n_31),
.B2(n_29),
.Y(n_47)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_42),
.B(n_23),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_0),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_44),
.B(n_45),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_0),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_46),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_47),
.A2(n_41),
.B1(n_37),
.B2(n_36),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_49),
.Y(n_77)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_50),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_38),
.A2(n_20),
.B1(n_29),
.B2(n_28),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_52),
.A2(n_56),
.B1(n_63),
.B2(n_19),
.Y(n_87)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

OR2x2_ASAP7_75t_SL g73 ( 
.A(n_54),
.B(n_55),
.Y(n_73)
);

OAI21xp33_ASAP7_75t_L g55 ( 
.A1(n_44),
.A2(n_1),
.B(n_3),
.Y(n_55)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

OR2x2_ASAP7_75t_SL g89 ( 
.A(n_58),
.B(n_41),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_44),
.B(n_24),
.Y(n_59)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_59),
.Y(n_72)
);

O2A1O1Ixp33_ASAP7_75t_L g67 ( 
.A1(n_60),
.A2(n_41),
.B(n_38),
.C(n_26),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_45),
.B(n_18),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_61),
.B(n_33),
.Y(n_79)
);

OAI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_38),
.A2(n_32),
.B1(n_30),
.B2(n_27),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_40),
.B(n_23),
.Y(n_64)
);

XNOR2xp5_ASAP7_75t_SL g83 ( 
.A(n_64),
.B(n_41),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_50),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_66),
.B(n_75),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_67),
.A2(n_87),
.B1(n_90),
.B2(n_33),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_61),
.B(n_42),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_69),
.B(n_53),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_49),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_70),
.Y(n_117)
);

INVx13_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_71),
.B(n_80),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_64),
.A2(n_37),
.B1(n_42),
.B2(n_36),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_74),
.A2(n_95),
.B1(n_51),
.B2(n_58),
.Y(n_101)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_56),
.Y(n_75)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_78),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_79),
.B(n_81),
.Y(n_115)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_46),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_57),
.B(n_21),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_46),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_82),
.B(n_84),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_83),
.B(n_48),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_57),
.B(n_21),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_59),
.B(n_25),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_85),
.B(n_88),
.Y(n_113)
);

NAND2x1_ASAP7_75t_SL g86 ( 
.A(n_60),
.B(n_43),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_86),
.A2(n_89),
.B(n_91),
.Y(n_114)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_62),
.Y(n_88)
);

AND2x2_ASAP7_75t_SL g91 ( 
.A(n_54),
.B(n_43),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_62),
.Y(n_92)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_92),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_46),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_93),
.B(n_22),
.Y(n_116)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_65),
.Y(n_94)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_94),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_65),
.A2(n_37),
.B1(n_36),
.B2(n_19),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_53),
.B(n_25),
.Y(n_96)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_96),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_97),
.B(n_102),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_101),
.A2(n_110),
.B1(n_67),
.B2(n_78),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_69),
.B(n_43),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_103),
.A2(n_91),
.B1(n_80),
.B2(n_17),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_66),
.B(n_39),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_104),
.B(n_108),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_106),
.B(n_83),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_68),
.B(n_72),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_75),
.A2(n_51),
.B1(n_43),
.B2(n_39),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_68),
.B(n_39),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_112),
.B(n_118),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_116),
.B(n_32),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_72),
.B(n_39),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_79),
.B(n_27),
.Y(n_119)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_119),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_79),
.B(n_30),
.Y(n_120)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_120),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_121),
.B(n_125),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_103),
.A2(n_107),
.B1(n_104),
.B2(n_102),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_122),
.A2(n_141),
.B1(n_115),
.B2(n_116),
.Y(n_146)
);

NAND3xp33_ASAP7_75t_L g123 ( 
.A(n_119),
.B(n_73),
.C(n_86),
.Y(n_123)
);

OAI211xp5_ASAP7_75t_L g163 ( 
.A1(n_123),
.A2(n_136),
.B(n_48),
.C(n_5),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_109),
.B(n_77),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_127),
.B(n_128),
.C(n_137),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_114),
.B(n_91),
.C(n_93),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_109),
.B(n_77),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_130),
.B(n_131),
.Y(n_155)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_118),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_114),
.A2(n_107),
.B(n_106),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_133),
.A2(n_113),
.B(n_111),
.Y(n_149)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_108),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_135),
.B(n_143),
.Y(n_152)
);

NOR3xp33_ASAP7_75t_SL g136 ( 
.A(n_120),
.B(n_73),
.C(n_89),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_106),
.B(n_74),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_138),
.A2(n_48),
.B1(n_5),
.B2(n_6),
.Y(n_164)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_113),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_139),
.B(n_100),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_110),
.Y(n_140)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_140),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_97),
.A2(n_95),
.B1(n_94),
.B2(n_71),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_142),
.A2(n_144),
.B1(n_117),
.B2(n_105),
.Y(n_153)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_112),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_101),
.A2(n_92),
.B1(n_88),
.B2(n_70),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_138),
.A2(n_143),
.B1(n_131),
.B2(n_144),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_145),
.A2(n_160),
.B1(n_154),
.B2(n_146),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_146),
.A2(n_149),
.B(n_153),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_132),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_147),
.B(n_151),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_135),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_150),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_132),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_124),
.B(n_111),
.Y(n_156)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_156),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_124),
.B(n_115),
.Y(n_157)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_157),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_127),
.B(n_76),
.C(n_105),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_159),
.B(n_4),
.C(n_7),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_122),
.A2(n_100),
.B1(n_98),
.B2(n_99),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_161),
.B(n_134),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_128),
.A2(n_98),
.B(n_24),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_162),
.B(n_133),
.C(n_137),
.Y(n_166)
);

AOI322xp5_ASAP7_75t_L g171 ( 
.A1(n_163),
.A2(n_129),
.A3(n_126),
.B1(n_136),
.B2(n_14),
.C1(n_16),
.C2(n_13),
.Y(n_171)
);

OAI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_164),
.A2(n_126),
.B1(n_157),
.B2(n_156),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_166),
.B(n_179),
.Y(n_187)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_154),
.B(n_134),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_167),
.A2(n_170),
.B(n_160),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_148),
.B(n_129),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_168),
.B(n_172),
.Y(n_183)
);

NOR3xp33_ASAP7_75t_SL g181 ( 
.A(n_171),
.B(n_149),
.C(n_16),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_155),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_174),
.B(n_178),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_176),
.A2(n_152),
.B1(n_162),
.B2(n_153),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_158),
.B(n_141),
.C(n_48),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_177),
.B(n_158),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_145),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_181),
.B(n_182),
.Y(n_194)
);

NOR3xp33_ASAP7_75t_SL g182 ( 
.A(n_173),
.B(n_151),
.C(n_147),
.Y(n_182)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_184),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_185),
.A2(n_190),
.B1(n_172),
.B2(n_179),
.Y(n_200)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_165),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_186),
.B(n_189),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_188),
.B(n_177),
.C(n_187),
.Y(n_199)
);

BUFx12_ASAP7_75t_L g189 ( 
.A(n_175),
.Y(n_189)
);

INVx13_ASAP7_75t_L g190 ( 
.A(n_175),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_178),
.A2(n_152),
.B1(n_159),
.B2(n_164),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_192),
.A2(n_167),
.B1(n_150),
.B2(n_9),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_191),
.A2(n_173),
.B(n_180),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_193),
.B(n_198),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_186),
.A2(n_169),
.B1(n_170),
.B2(n_167),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_195),
.A2(n_202),
.B1(n_150),
.B2(n_189),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_188),
.B(n_166),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_199),
.B(n_187),
.Y(n_208)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_200),
.Y(n_204)
);

NOR3xp33_ASAP7_75t_L g201 ( 
.A(n_182),
.B(n_161),
.C(n_181),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_201),
.B(n_183),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_203),
.B(n_205),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_197),
.A2(n_190),
.B1(n_184),
.B2(n_192),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_206),
.B(n_209),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_208),
.B(n_199),
.C(n_198),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_196),
.B(n_189),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_210),
.B(n_214),
.Y(n_216)
);

MAJx2_ASAP7_75t_L g213 ( 
.A(n_208),
.B(n_193),
.C(n_195),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_213),
.A2(n_204),
.B(n_207),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_207),
.B(n_194),
.C(n_202),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_212),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_215),
.A2(n_217),
.B1(n_218),
.B2(n_10),
.Y(n_221)
);

OAI321xp33_ASAP7_75t_L g218 ( 
.A1(n_212),
.A2(n_206),
.A3(n_13),
.B1(n_10),
.B2(n_11),
.C(n_12),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_216),
.B(n_211),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_219),
.B(n_220),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_216),
.B(n_4),
.C(n_7),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_221),
.A2(n_10),
.B(n_4),
.Y(n_223)
);

BUFx24_ASAP7_75t_SL g224 ( 
.A(n_223),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_224),
.B(n_222),
.Y(n_225)
);


endmodule