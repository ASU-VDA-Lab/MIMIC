module fake_aes_8951_n_1292 (n_117, n_219, n_44, n_133, n_149, n_220, n_81, n_69, n_214, n_267, n_204, n_221, n_249, n_185, n_22, n_203, n_57, n_88, n_52, n_244, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_107, n_158, n_278, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_240, n_254, n_9, n_161, n_262, n_10, n_177, n_130, n_189, n_103, n_239, n_19, n_87, n_137, n_180, n_104, n_277, n_160, n_98, n_74, n_206, n_276, n_154, n_272, n_7, n_29, n_195, n_165, n_146, n_45, n_85, n_250, n_237, n_181, n_101, n_62, n_255, n_36, n_47, n_215, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_217, n_139, n_229, n_230, n_274, n_16, n_13, n_198, n_169, n_193, n_273, n_252, n_152, n_113, n_241, n_95, n_124, n_156, n_238, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_247, n_197, n_201, n_242, n_260, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_202, n_210, n_38, n_64, n_142, n_184, n_245, n_265, n_191, n_264, n_232, n_200, n_46, n_31, n_208, n_211, n_58, n_122, n_187, n_138, n_126, n_275, n_178, n_118, n_258, n_253, n_32, n_0, n_179, n_84, n_131, n_112, n_266, n_55, n_205, n_12, n_86, n_143, n_213, n_235, n_243, n_182, n_263, n_166, n_162, n_186, n_75, n_163, n_226, n_105, n_159, n_174, n_227, n_248, n_268, n_231, n_72, n_136, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_256, n_67, n_77, n_216, n_20, n_2, n_147, n_199, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_212, n_228, n_92, n_11, n_223, n_251, n_25, n_30, n_59, n_236, n_150, n_218, n_168, n_194, n_3, n_18, n_110, n_261, n_66, n_134, n_222, n_234, n_1, n_164, n_233, n_271, n_82, n_106, n_175, n_15, n_173, n_190, n_145, n_270, n_246, n_153, n_61, n_259, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_207, n_257, n_224, n_96, n_269, n_225, n_39, n_1292);
input n_117;
input n_219;
input n_44;
input n_133;
input n_149;
input n_220;
input n_81;
input n_69;
input n_214;
input n_267;
input n_204;
input n_221;
input n_249;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_244;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_107;
input n_158;
input n_278;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_240;
input n_254;
input n_9;
input n_161;
input n_262;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_239;
input n_19;
input n_87;
input n_137;
input n_180;
input n_104;
input n_277;
input n_160;
input n_98;
input n_74;
input n_206;
input n_276;
input n_154;
input n_272;
input n_7;
input n_29;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_250;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_47;
input n_215;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_217;
input n_139;
input n_229;
input n_230;
input n_274;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_273;
input n_252;
input n_152;
input n_113;
input n_241;
input n_95;
input n_124;
input n_156;
input n_238;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_247;
input n_197;
input n_201;
input n_242;
input n_260;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_202;
input n_210;
input n_38;
input n_64;
input n_142;
input n_184;
input n_245;
input n_265;
input n_191;
input n_264;
input n_232;
input n_200;
input n_46;
input n_31;
input n_208;
input n_211;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_275;
input n_178;
input n_118;
input n_258;
input n_253;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_266;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_213;
input n_235;
input n_243;
input n_182;
input n_263;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_226;
input n_105;
input n_159;
input n_174;
input n_227;
input n_248;
input n_268;
input n_231;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_256;
input n_67;
input n_77;
input n_216;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_212;
input n_228;
input n_92;
input n_11;
input n_223;
input n_251;
input n_25;
input n_30;
input n_59;
input n_236;
input n_150;
input n_218;
input n_168;
input n_194;
input n_3;
input n_18;
input n_110;
input n_261;
input n_66;
input n_134;
input n_222;
input n_234;
input n_1;
input n_164;
input n_233;
input n_271;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_145;
input n_270;
input n_246;
input n_153;
input n_61;
input n_259;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_207;
input n_257;
input n_224;
input n_96;
input n_269;
input n_225;
input n_39;
output n_1292;
wire n_963;
wire n_1034;
wire n_949;
wire n_1277;
wire n_858;
wire n_646;
wire n_829;
wire n_1198;
wire n_667;
wire n_988;
wire n_311;
wire n_655;
wire n_903;
wire n_965;
wire n_918;
wire n_770;
wire n_1211;
wire n_878;
wire n_637;
wire n_564;
wire n_779;
wire n_528;
wire n_1128;
wire n_850;
wire n_672;
wire n_627;
wire n_1118;
wire n_1161;
wire n_1030;
wire n_807;
wire n_877;
wire n_545;
wire n_896;
wire n_334;
wire n_588;
wire n_1019;
wire n_940;
wire n_789;
wire n_1197;
wire n_1163;
wire n_387;
wire n_452;
wire n_518;
wire n_298;
wire n_411;
wire n_860;
wire n_1208;
wire n_305;
wire n_1201;
wire n_340;
wire n_373;
wire n_1194;
wire n_922;
wire n_465;
wire n_636;
wire n_914;
wire n_1005;
wire n_1097;
wire n_1125;
wire n_1017;
wire n_324;
wire n_773;
wire n_847;
wire n_668;
wire n_437;
wire n_680;
wire n_642;
wire n_1267;
wire n_830;
wire n_1112;
wire n_517;
wire n_502;
wire n_543;
wire n_312;
wire n_1159;
wire n_1250;
wire n_1002;
wire n_915;
wire n_367;
wire n_314;
wire n_999;
wire n_769;
wire n_624;
wire n_725;
wire n_1018;
wire n_979;
wire n_319;
wire n_499;
wire n_1033;
wire n_1063;
wire n_1010;
wire n_533;
wire n_490;
wire n_648;
wire n_613;
wire n_304;
wire n_892;
wire n_571;
wire n_610;
wire n_771;
wire n_474;
wire n_402;
wire n_413;
wire n_676;
wire n_950;
wire n_995;
wire n_938;
wire n_331;
wire n_746;
wire n_619;
wire n_501;
wire n_299;
wire n_699;
wire n_338;
wire n_551;
wire n_404;
wire n_1061;
wire n_509;
wire n_849;
wire n_864;
wire n_961;
wire n_1140;
wire n_611;
wire n_990;
wire n_800;
wire n_626;
wire n_1209;
wire n_926;
wire n_1274;
wire n_537;
wire n_660;
wire n_839;
wire n_1210;
wire n_1001;
wire n_1129;
wire n_450;
wire n_1099;
wire n_556;
wire n_1214;
wire n_379;
wire n_641;
wire n_966;
wire n_527;
wire n_797;
wire n_666;
wire n_954;
wire n_574;
wire n_823;
wire n_706;
wire n_822;
wire n_1181;
wire n_390;
wire n_514;
wire n_486;
wire n_568;
wire n_716;
wire n_899;
wire n_1066;
wire n_1251;
wire n_1199;
wire n_883;
wire n_573;
wire n_673;
wire n_1071;
wire n_1079;
wire n_315;
wire n_409;
wire n_295;
wire n_677;
wire n_1242;
wire n_283;
wire n_756;
wire n_1240;
wire n_1139;
wire n_577;
wire n_870;
wire n_790;
wire n_761;
wire n_1287;
wire n_472;
wire n_1100;
wire n_419;
wire n_1193;
wire n_1119;
wire n_825;
wire n_477;
wire n_815;
wire n_908;
wire n_429;
wire n_488;
wire n_821;
wire n_745;
wire n_684;
wire n_1281;
wire n_327;
wire n_1102;
wire n_723;
wire n_972;
wire n_997;
wire n_1244;
wire n_1184;
wire n_947;
wire n_620;
wire n_1141;
wire n_1213;
wire n_359;
wire n_1189;
wire n_923;
wire n_1205;
wire n_1172;
wire n_741;
wire n_1142;
wire n_1228;
wire n_831;
wire n_859;
wire n_1165;
wire n_930;
wire n_994;
wire n_410;
wire n_774;
wire n_1207;
wire n_377;
wire n_510;
wire n_1075;
wire n_1282;
wire n_493;
wire n_855;
wire n_722;
wire n_1083;
wire n_690;
wire n_1164;
wire n_281;
wire n_451;
wire n_487;
wire n_748;
wire n_824;
wire n_793;
wire n_753;
wire n_355;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_1226;
wire n_1233;
wire n_1067;
wire n_866;
wire n_1108;
wire n_350;
wire n_433;
wire n_483;
wire n_280;
wire n_395;
wire n_992;
wire n_361;
wire n_1077;
wire n_838;
wire n_705;
wire n_964;
wire n_590;
wire n_407;
wire n_1229;
wire n_792;
wire n_925;
wire n_1289;
wire n_957;
wire n_808;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_958;
wire n_468;
wire n_917;
wire n_523;
wire n_920;
wire n_1202;
wire n_911;
wire n_980;
wire n_817;
wire n_1056;
wire n_856;
wire n_661;
wire n_890;
wire n_787;
wire n_1015;
wire n_548;
wire n_1048;
wire n_973;
wire n_587;
wire n_476;
wire n_434;
wire n_489;
wire n_752;
wire n_1098;
wire n_1012;
wire n_461;
wire n_857;
wire n_1090;
wire n_786;
wire n_1121;
wire n_576;
wire n_1179;
wire n_796;
wire n_1216;
wire n_927;
wire n_840;
wire n_846;
wire n_968;
wire n_512;
wire n_586;
wire n_1246;
wire n_1276;
wire n_560;
wire n_697;
wire n_780;
wire n_447;
wire n_897;
wire n_1188;
wire n_580;
wire n_1009;
wire n_921;
wire n_854;
wire n_1011;
wire n_1155;
wire n_511;
wire n_467;
wire n_692;
wire n_644;
wire n_1116;
wire n_818;
wire n_738;
wire n_1225;
wire n_575;
wire n_711;
wire n_977;
wire n_884;
wire n_767;
wire n_293;
wire n_393;
wire n_550;
wire n_826;
wire n_399;
wire n_1235;
wire n_1171;
wire n_294;
wire n_459;
wire n_907;
wire n_310;
wire n_1062;
wire n_708;
wire n_1271;
wire n_307;
wire n_634;
wire n_696;
wire n_1203;
wire n_1013;
wire n_1000;
wire n_939;
wire n_953;
wire n_391;
wire n_478;
wire n_482;
wire n_394;
wire n_442;
wire n_485;
wire n_1248;
wire n_519;
wire n_329;
wire n_1020;
wire n_1106;
wire n_635;
wire n_731;
wire n_986;
wire n_507;
wire n_605;
wire n_704;
wire n_633;
wire n_873;
wire n_751;
wire n_1147;
wire n_466;
wire n_900;
wire n_952;
wire n_685;
wire n_308;
wire n_565;
wire n_1035;
wire n_475;
wire n_578;
wire n_542;
wire n_430;
wire n_943;
wire n_557;
wire n_842;
wire n_1269;
wire n_439;
wire n_614;
wire n_1107;
wire n_446;
wire n_423;
wire n_342;
wire n_799;
wire n_1050;
wire n_643;
wire n_874;
wire n_1049;
wire n_454;
wire n_687;
wire n_970;
wire n_984;
wire n_720;
wire n_1157;
wire n_806;
wire n_539;
wire n_1153;
wire n_317;
wire n_816;
wire n_522;
wire n_898;
wire n_1135;
wire n_669;
wire n_541;
wire n_363;
wire n_733;
wire n_894;
wire n_376;
wire n_744;
wire n_520;
wire n_681;
wire n_942;
wire n_1029;
wire n_508;
wire n_721;
wire n_1060;
wire n_438;
wire n_640;
wire n_1037;
wire n_686;
wire n_944;
wire n_1110;
wire n_498;
wire n_1069;
wire n_1123;
wire n_811;
wire n_530;
wire n_737;
wire n_1266;
wire n_795;
wire n_1232;
wire n_449;
wire n_734;
wire n_919;
wire n_763;
wire n_1174;
wire n_657;
wire n_583;
wire n_841;
wire n_582;
wire n_836;
wire n_561;
wire n_1096;
wire n_594;
wire n_531;
wire n_1136;
wire n_306;
wire n_1007;
wire n_1117;
wire n_424;
wire n_714;
wire n_932;
wire n_837;
wire n_867;
wire n_1070;
wire n_1270;
wire n_675;
wire n_504;
wire n_581;
wire n_698;
wire n_555;
wire n_901;
wire n_834;
wire n_727;
wire n_1038;
wire n_1162;
wire n_1103;
wire n_785;
wire n_375;
wire n_688;
wire n_323;
wire n_347;
wire n_515;
wire n_1290;
wire n_1234;
wire n_592;
wire n_1045;
wire n_1115;
wire n_521;
wire n_625;
wire n_585;
wire n_1190;
wire n_1237;
wire n_713;
wire n_457;
wire n_736;
wire n_287;
wire n_606;
wire n_332;
wire n_421;
wire n_1148;
wire n_739;
wire n_1166;
wire n_987;
wire n_1086;
wire n_406;
wire n_1236;
wire n_791;
wire n_707;
wire n_603;
wire n_1261;
wire n_885;
wire n_284;
wire n_500;
wire n_607;
wire n_496;
wire n_801;
wire n_1059;
wire n_309;
wire n_701;
wire n_612;
wire n_1032;
wire n_1284;
wire n_336;
wire n_464;
wire n_1243;
wire n_1196;
wire n_814;
wire n_985;
wire n_1191;
wire n_971;
wire n_904;
wire n_532;
wire n_400;
wire n_386;
wire n_432;
wire n_659;
wire n_316;
wire n_1185;
wire n_389;
wire n_436;
wire n_1217;
wire n_715;
wire n_330;
wire n_1087;
wire n_662;
wire n_617;
wire n_598;
wire n_732;
wire n_724;
wire n_599;
wire n_301;
wire n_609;
wire n_909;
wire n_1273;
wire n_366;
wire n_596;
wire n_1215;
wire n_286;
wire n_951;
wire n_321;
wire n_1024;
wire n_1016;
wire n_652;
wire n_333;
wire n_638;
wire n_563;
wire n_479;
wire n_623;
wire n_1222;
wire n_593;
wire n_872;
wire n_809;
wire n_1101;
wire n_1072;
wire n_865;
wire n_1064;
wire n_1254;
wire n_764;
wire n_426;
wire n_282;
wire n_969;
wire n_417;
wire n_1253;
wire n_632;
wire n_1182;
wire n_828;
wire n_1138;
wire n_506;
wire n_381;
wire n_1255;
wire n_313;
wire n_322;
wire n_427;
wire n_703;
wire n_415;
wire n_1272;
wire n_928;
wire n_352;
wire n_882;
wire n_871;
wire n_803;
wire n_805;
wire n_729;
wire n_693;
wire n_1036;
wire n_1145;
wire n_651;
wire n_747;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_959;
wire n_719;
wire n_1206;
wire n_1257;
wire n_710;
wire n_1178;
wire n_546;
wire n_412;
wire n_664;
wire n_1249;
wire n_788;
wire n_403;
wire n_516;
wire n_549;
wire n_832;
wire n_996;
wire n_285;
wire n_420;
wire n_1089;
wire n_1058;
wire n_388;
wire n_1082;
wire n_1052;
wire n_1055;
wire n_974;
wire n_591;
wire n_933;
wire n_1252;
wire n_416;
wire n_536;
wire n_1256;
wire n_1259;
wire n_956;
wire n_989;
wire n_754;
wire n_775;
wire n_616;
wire n_1227;
wire n_365;
wire n_495;
wire n_364;
wire n_566;
wire n_1144;
wire n_344;
wire n_503;
wire n_1279;
wire n_1152;
wire n_1068;
wire n_1149;
wire n_615;
wire n_1170;
wire n_804;
wire n_570;
wire n_1133;
wire n_440;
wire n_422;
wire n_679;
wire n_1131;
wire n_597;
wire n_1039;
wire n_835;
wire n_778;
wire n_1156;
wire n_1288;
wire n_300;
wire n_1042;
wire n_1130;
wire n_584;
wire n_912;
wire n_1043;
wire n_1283;
wire n_346;
wire n_397;
wire n_1008;
wire n_1109;
wire n_1026;
wire n_1027;
wire n_1040;
wire n_569;
wire n_946;
wire n_960;
wire n_1168;
wire n_343;
wire n_458;
wire n_1084;
wire n_618;
wire n_341;
wire n_470;
wire n_1085;
wire n_1073;
wire n_868;
wire n_473;
wire n_991;
wire n_843;
wire n_1263;
wire n_538;
wire n_492;
wire n_1150;
wire n_368;
wire n_650;
wire n_469;
wire n_1187;
wire n_742;
wire n_913;
wire n_845;
wire n_891;
wire n_1134;
wire n_494;
wire n_372;
wire n_631;
wire n_934;
wire n_425;
wire n_562;
wire n_1192;
wire n_983;
wire n_781;
wire n_709;
wire n_1105;
wire n_408;
wire n_290;
wire n_385;
wire n_1127;
wire n_1173;
wire n_663;
wire n_513;
wire n_1092;
wire n_1124;
wire n_1278;
wire n_998;
wire n_604;
wire n_1260;
wire n_755;
wire n_848;
wire n_1031;
wire n_1280;
wire n_292;
wire n_1158;
wire n_328;
wire n_743;
wire n_757;
wire n_750;
wire n_448;
wire n_645;
wire n_348;
wire n_1022;
wire n_802;
wire n_353;
wire n_993;
wire n_1122;
wire n_1224;
wire n_288;
wire n_383;
wire n_762;
wire n_981;
wire n_1095;
wire n_758;
wire n_544;
wire n_1175;
wire n_853;
wire n_296;
wire n_765;
wire n_1177;
wire n_462;
wire n_783;
wire n_1074;
wire n_463;
wire n_1003;
wire n_678;
wire n_1200;
wire n_384;
wire n_978;
wire n_547;
wire n_1247;
wire n_628;
wire n_812;
wire n_777;
wire n_351;
wire n_401;
wire n_345;
wire n_360;
wire n_481;
wire n_443;
wire n_694;
wire n_1262;
wire n_1078;
wire n_702;
wire n_572;
wire n_1094;
wire n_1204;
wire n_392;
wire n_1169;
wire n_975;
wire n_279;
wire n_303;
wire n_326;
wire n_289;
wire n_1081;
wire n_671;
wire n_540;
wire n_937;
wire n_1093;
wire n_955;
wire n_1275;
wire n_945;
wire n_554;
wire n_726;
wire n_712;
wire n_608;
wire n_567;
wire n_888;
wire n_455;
wire n_529;
wire n_1025;
wire n_1132;
wire n_630;
wire n_1180;
wire n_647;
wire n_844;
wire n_1160;
wire n_1245;
wire n_1195;
wire n_1241;
wire n_895;
wire n_798;
wire n_318;
wire n_887;
wire n_471;
wire n_1014;
wire n_665;
wire n_1154;
wire n_863;
wire n_1265;
wire n_730;
wire n_1212;
wire n_735;
wire n_1091;
wire n_784;
wire n_354;
wire n_1220;
wire n_893;
wire n_1028;
wire n_910;
wire n_935;
wire n_1046;
wire n_1183;
wire n_460;
wire n_813;
wire n_1076;
wire n_369;
wire n_1186;
wire n_1167;
wire n_674;
wire n_810;
wire n_982;
wire n_889;
wire n_689;
wire n_902;
wire n_1113;
wire n_1264;
wire n_760;
wire n_941;
wire n_302;
wire n_362;
wire n_931;
wire n_827;
wire n_1218;
wire n_1041;
wire n_1080;
wire n_1126;
wire n_1151;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_1065;
wire n_622;
wire n_601;
wire n_1176;
wire n_649;
wire n_526;
wire n_1047;
wire n_320;
wire n_768;
wire n_869;
wire n_880;
wire n_621;
wire n_370;
wire n_589;
wire n_505;
wire n_682;
wire n_906;
wire n_357;
wire n_653;
wire n_881;
wire n_374;
wire n_718;
wire n_1238;
wire n_1114;
wire n_1286;
wire n_948;
wire n_717;
wire n_861;
wire n_654;
wire n_1221;
wire n_428;
wire n_794;
wire n_1268;
wire n_639;
wire n_552;
wire n_1023;
wire n_1057;
wire n_435;
wire n_1051;
wire n_1088;
wire n_851;
wire n_396;
wire n_398;
wire n_445;
wire n_656;
wire n_1230;
wire n_553;
wire n_325;
wire n_349;
wire n_1021;
wire n_749;
wire n_535;
wire n_1006;
wire n_1054;
wire n_1231;
wire n_358;
wire n_456;
wire n_962;
wire n_782;
wire n_524;
wire n_1044;
wire n_875;
wire n_497;
wire n_728;
wire n_339;
wire n_1239;
wire n_924;
wire n_378;
wire n_441;
wire n_1285;
wire n_335;
wire n_700;
wire n_534;
wire n_766;
wire n_602;
wire n_1143;
wire n_629;
wire n_297;
wire n_1053;
wire n_1223;
wire n_967;
wire n_1258;
wire n_291;
wire n_418;
wire n_380;
wire n_356;
wire n_600;
wire n_371;
wire n_820;
wire n_558;
wire n_670;
wire n_1004;
wire n_683;
wire n_929;
wire n_1111;
wire n_976;
wire n_695;
wire n_1104;
wire n_1120;
wire n_1219;
wire n_595;
wire n_759;
wire n_559;
wire n_480;
wire n_453;
wire n_833;
wire n_1146;
wire n_414;
wire n_1137;
wire n_916;
wire n_740;
wire n_772;
wire n_819;
wire n_405;
wire n_491;
wire n_1291;
INVxp67_ASAP7_75t_SL g279 ( .A(n_183), .Y(n_279) );
INVxp33_ASAP7_75t_L g280 ( .A(n_212), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_23), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_12), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_184), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_229), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_112), .Y(n_285) );
BUFx3_ASAP7_75t_L g286 ( .A(n_131), .Y(n_286) );
INVx2_ASAP7_75t_L g287 ( .A(n_210), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_3), .Y(n_288) );
INVxp33_ASAP7_75t_L g289 ( .A(n_63), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_178), .Y(n_290) );
INVx2_ASAP7_75t_L g291 ( .A(n_250), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_197), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_171), .Y(n_293) );
CKINVDCx5p33_ASAP7_75t_R g294 ( .A(n_67), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_218), .Y(n_295) );
INVxp33_ASAP7_75t_L g296 ( .A(n_222), .Y(n_296) );
CKINVDCx16_ASAP7_75t_R g297 ( .A(n_1), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_126), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_273), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_148), .Y(n_300) );
INVx2_ASAP7_75t_L g301 ( .A(n_76), .Y(n_301) );
CKINVDCx16_ASAP7_75t_R g302 ( .A(n_54), .Y(n_302) );
CKINVDCx5p33_ASAP7_75t_R g303 ( .A(n_252), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_246), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_76), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_193), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_234), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_249), .Y(n_308) );
CKINVDCx5p33_ASAP7_75t_R g309 ( .A(n_138), .Y(n_309) );
CKINVDCx16_ASAP7_75t_R g310 ( .A(n_68), .Y(n_310) );
CKINVDCx5p33_ASAP7_75t_R g311 ( .A(n_27), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_144), .Y(n_312) );
INVxp33_ASAP7_75t_SL g313 ( .A(n_73), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_267), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_62), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_214), .Y(n_316) );
CKINVDCx20_ASAP7_75t_R g317 ( .A(n_245), .Y(n_317) );
INVxp33_ASAP7_75t_SL g318 ( .A(n_86), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_262), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_256), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_206), .Y(n_321) );
NOR2xp33_ASAP7_75t_L g322 ( .A(n_34), .B(n_53), .Y(n_322) );
INVxp33_ASAP7_75t_SL g323 ( .A(n_142), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_196), .Y(n_324) );
INVxp33_ASAP7_75t_SL g325 ( .A(n_26), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_276), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_264), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_150), .Y(n_328) );
CKINVDCx5p33_ASAP7_75t_R g329 ( .A(n_274), .Y(n_329) );
INVxp67_ASAP7_75t_SL g330 ( .A(n_96), .Y(n_330) );
INVxp33_ASAP7_75t_SL g331 ( .A(n_106), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_176), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_241), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_58), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_31), .Y(n_335) );
INVxp33_ASAP7_75t_SL g336 ( .A(n_81), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_141), .Y(n_337) );
INVxp67_ASAP7_75t_SL g338 ( .A(n_185), .Y(n_338) );
CKINVDCx20_ASAP7_75t_R g339 ( .A(n_101), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_59), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_104), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_87), .Y(n_342) );
HB1xp67_ASAP7_75t_L g343 ( .A(n_260), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_58), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_61), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_162), .Y(n_346) );
INVxp67_ASAP7_75t_SL g347 ( .A(n_103), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_158), .Y(n_348) );
CKINVDCx20_ASAP7_75t_R g349 ( .A(n_82), .Y(n_349) );
BUFx8_ASAP7_75t_SL g350 ( .A(n_186), .Y(n_350) );
CKINVDCx5p33_ASAP7_75t_R g351 ( .A(n_24), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_34), .Y(n_352) );
INVxp67_ASAP7_75t_SL g353 ( .A(n_27), .Y(n_353) );
INVxp33_ASAP7_75t_L g354 ( .A(n_59), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_110), .Y(n_355) );
CKINVDCx16_ASAP7_75t_R g356 ( .A(n_88), .Y(n_356) );
INVxp33_ASAP7_75t_L g357 ( .A(n_136), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_275), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_23), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_181), .Y(n_360) );
INVxp67_ASAP7_75t_SL g361 ( .A(n_205), .Y(n_361) );
CKINVDCx20_ASAP7_75t_R g362 ( .A(n_147), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_157), .Y(n_363) );
CKINVDCx20_ASAP7_75t_R g364 ( .A(n_172), .Y(n_364) );
CKINVDCx5p33_ASAP7_75t_R g365 ( .A(n_92), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_240), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_91), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_35), .Y(n_368) );
CKINVDCx5p33_ASAP7_75t_R g369 ( .A(n_44), .Y(n_369) );
BUFx6f_ASAP7_75t_SL g370 ( .A(n_5), .Y(n_370) );
INVxp33_ASAP7_75t_SL g371 ( .A(n_224), .Y(n_371) );
CKINVDCx5p33_ASAP7_75t_R g372 ( .A(n_191), .Y(n_372) );
CKINVDCx14_ASAP7_75t_R g373 ( .A(n_160), .Y(n_373) );
INVxp67_ASAP7_75t_SL g374 ( .A(n_152), .Y(n_374) );
INVxp33_ASAP7_75t_SL g375 ( .A(n_89), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_177), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_57), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_237), .Y(n_378) );
BUFx3_ASAP7_75t_L g379 ( .A(n_161), .Y(n_379) );
CKINVDCx5p33_ASAP7_75t_R g380 ( .A(n_90), .Y(n_380) );
INVxp67_ASAP7_75t_SL g381 ( .A(n_146), .Y(n_381) );
INVxp33_ASAP7_75t_SL g382 ( .A(n_188), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_65), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_140), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_208), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_85), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_44), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_31), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_107), .Y(n_389) );
CKINVDCx5p33_ASAP7_75t_R g390 ( .A(n_228), .Y(n_390) );
INVxp67_ASAP7_75t_L g391 ( .A(n_149), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_1), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_251), .Y(n_393) );
BUFx3_ASAP7_75t_L g394 ( .A(n_182), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_128), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_113), .Y(n_396) );
CKINVDCx5p33_ASAP7_75t_R g397 ( .A(n_0), .Y(n_397) );
CKINVDCx16_ASAP7_75t_R g398 ( .A(n_215), .Y(n_398) );
NOR2xp33_ASAP7_75t_L g399 ( .A(n_62), .B(n_239), .Y(n_399) );
BUFx3_ASAP7_75t_L g400 ( .A(n_187), .Y(n_400) );
INVxp33_ASAP7_75t_L g401 ( .A(n_15), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_221), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_121), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_100), .Y(n_404) );
INVxp67_ASAP7_75t_SL g405 ( .A(n_248), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_83), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_20), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_156), .Y(n_408) );
CKINVDCx16_ASAP7_75t_R g409 ( .A(n_166), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_7), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_81), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_139), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_93), .Y(n_413) );
HB1xp67_ASAP7_75t_L g414 ( .A(n_118), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_10), .Y(n_415) );
CKINVDCx20_ASAP7_75t_R g416 ( .A(n_61), .Y(n_416) );
AND2x4_ASAP7_75t_L g417 ( .A(n_301), .B(n_0), .Y(n_417) );
NAND2xp5_ASAP7_75t_SL g418 ( .A(n_280), .B(n_2), .Y(n_418) );
AND2x4_ASAP7_75t_L g419 ( .A(n_301), .B(n_2), .Y(n_419) );
INVx3_ASAP7_75t_L g420 ( .A(n_292), .Y(n_420) );
CKINVDCx5p33_ASAP7_75t_R g421 ( .A(n_370), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_292), .Y(n_422) );
INVx2_ASAP7_75t_L g423 ( .A(n_287), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_343), .B(n_3), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_414), .B(n_4), .Y(n_425) );
INVx6_ASAP7_75t_L g426 ( .A(n_286), .Y(n_426) );
INVx2_ASAP7_75t_L g427 ( .A(n_287), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_305), .B(n_4), .Y(n_428) );
INVx3_ASAP7_75t_L g429 ( .A(n_293), .Y(n_429) );
HB1xp67_ASAP7_75t_L g430 ( .A(n_370), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_305), .B(n_5), .Y(n_431) );
BUFx6f_ASAP7_75t_L g432 ( .A(n_286), .Y(n_432) );
INVx3_ASAP7_75t_L g433 ( .A(n_293), .Y(n_433) );
NAND2xp5_ASAP7_75t_SL g434 ( .A(n_296), .B(n_6), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_315), .B(n_6), .Y(n_435) );
INVx2_ASAP7_75t_L g436 ( .A(n_291), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_295), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_295), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_298), .Y(n_439) );
INVx2_ASAP7_75t_L g440 ( .A(n_291), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_298), .Y(n_441) );
BUFx6f_ASAP7_75t_L g442 ( .A(n_379), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_299), .Y(n_443) );
BUFx2_ASAP7_75t_L g444 ( .A(n_356), .Y(n_444) );
NAND2xp5_ASAP7_75t_SL g445 ( .A(n_357), .B(n_7), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_299), .Y(n_446) );
AND2x4_ASAP7_75t_L g447 ( .A(n_379), .B(n_8), .Y(n_447) );
BUFx6f_ASAP7_75t_L g448 ( .A(n_394), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_423), .Y(n_449) );
AND2x2_ASAP7_75t_L g450 ( .A(n_430), .B(n_398), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_423), .Y(n_451) );
OAI21xp33_ASAP7_75t_L g452 ( .A1(n_422), .A2(n_400), .B(n_394), .Y(n_452) );
BUFx6f_ASAP7_75t_L g453 ( .A(n_432), .Y(n_453) );
AND2x2_ASAP7_75t_SL g454 ( .A(n_447), .B(n_409), .Y(n_454) );
INVx3_ASAP7_75t_L g455 ( .A(n_417), .Y(n_455) );
OR2x6_ASAP7_75t_L g456 ( .A(n_430), .B(n_315), .Y(n_456) );
INVx4_ASAP7_75t_SL g457 ( .A(n_426), .Y(n_457) );
BUFx3_ASAP7_75t_L g458 ( .A(n_426), .Y(n_458) );
OAI22xp33_ASAP7_75t_SL g459 ( .A1(n_418), .A2(n_325), .B1(n_336), .B2(n_313), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_422), .B(n_283), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_423), .Y(n_461) );
AND2x2_ASAP7_75t_L g462 ( .A(n_444), .B(n_289), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_422), .B(n_284), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_423), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_427), .Y(n_465) );
AND2x6_ASAP7_75t_L g466 ( .A(n_447), .B(n_300), .Y(n_466) );
AOI22xp5_ASAP7_75t_L g467 ( .A1(n_417), .A2(n_325), .B1(n_336), .B2(n_313), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_444), .B(n_354), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_427), .Y(n_469) );
OR2x2_ASAP7_75t_L g470 ( .A(n_444), .B(n_297), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_427), .Y(n_471) );
BUFx6f_ASAP7_75t_L g472 ( .A(n_432), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_427), .Y(n_473) );
NAND2x1p5_ASAP7_75t_L g474 ( .A(n_417), .B(n_300), .Y(n_474) );
AND2x2_ASAP7_75t_L g475 ( .A(n_421), .B(n_373), .Y(n_475) );
BUFx3_ASAP7_75t_L g476 ( .A(n_426), .Y(n_476) );
OR2x2_ASAP7_75t_L g477 ( .A(n_424), .B(n_302), .Y(n_477) );
NAND2xp33_ASAP7_75t_L g478 ( .A(n_421), .B(n_303), .Y(n_478) );
BUFx2_ASAP7_75t_L g479 ( .A(n_447), .Y(n_479) );
OAI22xp5_ASAP7_75t_L g480 ( .A1(n_417), .A2(n_310), .B1(n_416), .B2(n_349), .Y(n_480) );
OR2x2_ASAP7_75t_L g481 ( .A(n_424), .B(n_401), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_436), .Y(n_482) );
BUFx3_ASAP7_75t_L g483 ( .A(n_426), .Y(n_483) );
AND2x4_ASAP7_75t_L g484 ( .A(n_447), .B(n_345), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_436), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_436), .Y(n_486) );
INVx2_ASAP7_75t_L g487 ( .A(n_432), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_436), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_438), .B(n_285), .Y(n_489) );
INVx3_ASAP7_75t_L g490 ( .A(n_417), .Y(n_490) );
INVx2_ASAP7_75t_L g491 ( .A(n_432), .Y(n_491) );
INVx2_ASAP7_75t_L g492 ( .A(n_432), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_474), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_481), .B(n_437), .Y(n_494) );
BUFx3_ASAP7_75t_L g495 ( .A(n_466), .Y(n_495) );
INVx2_ASAP7_75t_L g496 ( .A(n_449), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_474), .Y(n_497) );
INVx4_ASAP7_75t_L g498 ( .A(n_456), .Y(n_498) );
INVx3_ASAP7_75t_SL g499 ( .A(n_456), .Y(n_499) );
INVx3_ASAP7_75t_L g500 ( .A(n_455), .Y(n_500) );
BUFx6f_ASAP7_75t_L g501 ( .A(n_466), .Y(n_501) );
BUFx8_ASAP7_75t_L g502 ( .A(n_450), .Y(n_502) );
INVx5_ASAP7_75t_L g503 ( .A(n_466), .Y(n_503) );
AND2x4_ASAP7_75t_L g504 ( .A(n_456), .B(n_417), .Y(n_504) );
AND2x4_ASAP7_75t_L g505 ( .A(n_456), .B(n_419), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_481), .B(n_437), .Y(n_506) );
AND3x1_ASAP7_75t_L g507 ( .A(n_467), .B(n_425), .C(n_428), .Y(n_507) );
AOI22xp5_ASAP7_75t_L g508 ( .A1(n_454), .A2(n_418), .B1(n_445), .B2(n_434), .Y(n_508) );
INVx3_ASAP7_75t_L g509 ( .A(n_455), .Y(n_509) );
AOI21xp5_ASAP7_75t_L g510 ( .A1(n_479), .A2(n_439), .B(n_438), .Y(n_510) );
AOI22xp5_ASAP7_75t_L g511 ( .A1(n_454), .A2(n_445), .B1(n_434), .B2(n_447), .Y(n_511) );
AOI21xp5_ASAP7_75t_L g512 ( .A1(n_479), .A2(n_439), .B(n_438), .Y(n_512) );
NOR2xp33_ASAP7_75t_L g513 ( .A(n_455), .B(n_425), .Y(n_513) );
AND2x6_ASAP7_75t_L g514 ( .A(n_455), .B(n_447), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_454), .B(n_443), .Y(n_515) );
AOI22xp5_ASAP7_75t_L g516 ( .A1(n_467), .A2(n_370), .B1(n_419), .B2(n_311), .Y(n_516) );
AND2x4_ASAP7_75t_L g517 ( .A(n_456), .B(n_419), .Y(n_517) );
BUFx3_ASAP7_75t_L g518 ( .A(n_466), .Y(n_518) );
INVx3_ASAP7_75t_L g519 ( .A(n_490), .Y(n_519) );
NOR2xp33_ASAP7_75t_L g520 ( .A(n_490), .B(n_443), .Y(n_520) );
BUFx6f_ASAP7_75t_L g521 ( .A(n_466), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_474), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_474), .Y(n_523) );
NAND3xp33_ASAP7_75t_L g524 ( .A(n_477), .B(n_311), .C(n_294), .Y(n_524) );
INVx2_ASAP7_75t_L g525 ( .A(n_449), .Y(n_525) );
NAND2x1_ASAP7_75t_L g526 ( .A(n_466), .B(n_426), .Y(n_526) );
INVx2_ASAP7_75t_L g527 ( .A(n_451), .Y(n_527) );
BUFx2_ASAP7_75t_L g528 ( .A(n_456), .Y(n_528) );
OR2x6_ASAP7_75t_L g529 ( .A(n_480), .B(n_419), .Y(n_529) );
INVx2_ASAP7_75t_L g530 ( .A(n_451), .Y(n_530) );
AND2x2_ASAP7_75t_L g531 ( .A(n_462), .B(n_294), .Y(n_531) );
BUFx3_ASAP7_75t_L g532 ( .A(n_466), .Y(n_532) );
CKINVDCx5p33_ASAP7_75t_R g533 ( .A(n_480), .Y(n_533) );
NOR2xp33_ASAP7_75t_L g534 ( .A(n_490), .B(n_446), .Y(n_534) );
NOR2xp67_ASAP7_75t_L g535 ( .A(n_470), .B(n_420), .Y(n_535) );
INVx3_ASAP7_75t_L g536 ( .A(n_490), .Y(n_536) );
INVx2_ASAP7_75t_L g537 ( .A(n_461), .Y(n_537) );
CKINVDCx5p33_ASAP7_75t_R g538 ( .A(n_450), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_477), .B(n_446), .Y(n_539) );
BUFx2_ASAP7_75t_L g540 ( .A(n_450), .Y(n_540) );
NAND2xp5_ASAP7_75t_SL g541 ( .A(n_484), .B(n_419), .Y(n_541) );
CKINVDCx5p33_ASAP7_75t_R g542 ( .A(n_470), .Y(n_542) );
BUFx2_ASAP7_75t_L g543 ( .A(n_462), .Y(n_543) );
BUFx6f_ASAP7_75t_L g544 ( .A(n_466), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_484), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_484), .Y(n_546) );
INVx3_ASAP7_75t_SL g547 ( .A(n_466), .Y(n_547) );
BUFx3_ASAP7_75t_L g548 ( .A(n_458), .Y(n_548) );
INVx3_ASAP7_75t_L g549 ( .A(n_484), .Y(n_549) );
AND2x4_ASAP7_75t_L g550 ( .A(n_475), .B(n_419), .Y(n_550) );
INVx3_ASAP7_75t_L g551 ( .A(n_461), .Y(n_551) );
INVx4_ASAP7_75t_L g552 ( .A(n_457), .Y(n_552) );
CKINVDCx8_ASAP7_75t_R g553 ( .A(n_457), .Y(n_553) );
HB1xp67_ASAP7_75t_L g554 ( .A(n_468), .Y(n_554) );
NAND2xp5_ASAP7_75t_SL g555 ( .A(n_459), .B(n_439), .Y(n_555) );
OR2x6_ASAP7_75t_L g556 ( .A(n_468), .B(n_428), .Y(n_556) );
AOI22xp33_ASAP7_75t_L g557 ( .A1(n_464), .A2(n_441), .B1(n_429), .B2(n_433), .Y(n_557) );
AOI22xp33_ASAP7_75t_L g558 ( .A1(n_464), .A2(n_441), .B1(n_429), .B2(n_433), .Y(n_558) );
AOI22xp5_ASAP7_75t_L g559 ( .A1(n_459), .A2(n_369), .B1(n_397), .B2(n_351), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_465), .Y(n_560) );
AOI22xp5_ASAP7_75t_L g561 ( .A1(n_475), .A2(n_369), .B1(n_397), .B2(n_351), .Y(n_561) );
AOI22xp5_ASAP7_75t_L g562 ( .A1(n_475), .A2(n_339), .B1(n_362), .B2(n_317), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_460), .B(n_441), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_465), .Y(n_564) );
CKINVDCx5p33_ASAP7_75t_R g565 ( .A(n_460), .Y(n_565) );
INVx2_ASAP7_75t_L g566 ( .A(n_469), .Y(n_566) );
OR2x2_ASAP7_75t_L g567 ( .A(n_463), .B(n_431), .Y(n_567) );
CKINVDCx8_ASAP7_75t_R g568 ( .A(n_478), .Y(n_568) );
AND2x4_ASAP7_75t_L g569 ( .A(n_463), .B(n_431), .Y(n_569) );
INVx2_ASAP7_75t_L g570 ( .A(n_469), .Y(n_570) );
AOI21x1_ASAP7_75t_L g571 ( .A1(n_489), .A2(n_440), .B(n_435), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_471), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_489), .B(n_420), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_551), .Y(n_574) );
INVx2_ASAP7_75t_SL g575 ( .A(n_499), .Y(n_575) );
INVx2_ASAP7_75t_SL g576 ( .A(n_499), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_551), .Y(n_577) );
BUFx3_ASAP7_75t_L g578 ( .A(n_547), .Y(n_578) );
BUFx10_ASAP7_75t_L g579 ( .A(n_504), .Y(n_579) );
NOR2xp33_ASAP7_75t_L g580 ( .A(n_554), .B(n_318), .Y(n_580) );
AND2x2_ASAP7_75t_L g581 ( .A(n_569), .B(n_471), .Y(n_581) );
AOI22xp33_ASAP7_75t_L g582 ( .A1(n_529), .A2(n_452), .B1(n_482), .B2(n_473), .Y(n_582) );
NOR2xp33_ASAP7_75t_L g583 ( .A(n_554), .B(n_318), .Y(n_583) );
BUFx2_ASAP7_75t_L g584 ( .A(n_498), .Y(n_584) );
AND2x4_ASAP7_75t_L g585 ( .A(n_498), .B(n_435), .Y(n_585) );
INVx4_ASAP7_75t_L g586 ( .A(n_498), .Y(n_586) );
INVx3_ASAP7_75t_L g587 ( .A(n_501), .Y(n_587) );
AOI22xp33_ASAP7_75t_L g588 ( .A1(n_529), .A2(n_452), .B1(n_482), .B2(n_473), .Y(n_588) );
BUFx6f_ASAP7_75t_L g589 ( .A(n_501), .Y(n_589) );
AO21x2_ASAP7_75t_L g590 ( .A1(n_555), .A2(n_306), .B(n_304), .Y(n_590) );
AO21x2_ASAP7_75t_L g591 ( .A1(n_555), .A2(n_306), .B(n_304), .Y(n_591) );
OR2x2_ASAP7_75t_L g592 ( .A(n_542), .B(n_485), .Y(n_592) );
INVx2_ASAP7_75t_L g593 ( .A(n_496), .Y(n_593) );
BUFx6f_ASAP7_75t_L g594 ( .A(n_501), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_545), .Y(n_595) );
HB1xp67_ASAP7_75t_L g596 ( .A(n_504), .Y(n_596) );
INVx2_ASAP7_75t_L g597 ( .A(n_496), .Y(n_597) );
INVx2_ASAP7_75t_L g598 ( .A(n_525), .Y(n_598) );
BUFx8_ASAP7_75t_SL g599 ( .A(n_529), .Y(n_599) );
INVx5_ASAP7_75t_L g600 ( .A(n_501), .Y(n_600) );
INVx4_ASAP7_75t_L g601 ( .A(n_547), .Y(n_601) );
AOI21xp5_ASAP7_75t_L g602 ( .A1(n_541), .A2(n_476), .B(n_458), .Y(n_602) );
HB1xp67_ASAP7_75t_L g603 ( .A(n_504), .Y(n_603) );
AND2x2_ASAP7_75t_L g604 ( .A(n_569), .B(n_485), .Y(n_604) );
INVxp67_ASAP7_75t_SL g605 ( .A(n_528), .Y(n_605) );
BUFx12f_ASAP7_75t_L g606 ( .A(n_502), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_525), .Y(n_607) );
INVx3_ASAP7_75t_L g608 ( .A(n_521), .Y(n_608) );
AOI22xp33_ASAP7_75t_L g609 ( .A1(n_505), .A2(n_488), .B1(n_486), .B2(n_331), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_565), .B(n_486), .Y(n_610) );
AOI21xp5_ASAP7_75t_L g611 ( .A1(n_541), .A2(n_476), .B(n_458), .Y(n_611) );
CKINVDCx20_ASAP7_75t_R g612 ( .A(n_502), .Y(n_612) );
INVx2_ASAP7_75t_L g613 ( .A(n_527), .Y(n_613) );
BUFx3_ASAP7_75t_L g614 ( .A(n_521), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_527), .Y(n_615) );
AOI221xp5_ASAP7_75t_L g616 ( .A1(n_507), .A2(n_353), .B1(n_282), .B2(n_334), .C(n_288), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_546), .Y(n_617) );
INVx2_ASAP7_75t_L g618 ( .A(n_530), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_549), .Y(n_619) );
AND2x2_ASAP7_75t_L g620 ( .A(n_569), .B(n_488), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_530), .Y(n_621) );
CKINVDCx20_ASAP7_75t_R g622 ( .A(n_502), .Y(n_622) );
NAND2xp5_ASAP7_75t_SL g623 ( .A(n_565), .B(n_303), .Y(n_623) );
OR2x6_ASAP7_75t_SL g624 ( .A(n_542), .B(n_309), .Y(n_624) );
BUFx6f_ASAP7_75t_L g625 ( .A(n_521), .Y(n_625) );
BUFx12f_ASAP7_75t_L g626 ( .A(n_533), .Y(n_626) );
INVx3_ASAP7_75t_L g627 ( .A(n_521), .Y(n_627) );
BUFx2_ASAP7_75t_L g628 ( .A(n_505), .Y(n_628) );
AOI21xp5_ASAP7_75t_L g629 ( .A1(n_510), .A2(n_483), .B(n_476), .Y(n_629) );
INVxp67_ASAP7_75t_SL g630 ( .A(n_493), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_537), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_537), .Y(n_632) );
A2O1A1Ixp33_ASAP7_75t_SL g633 ( .A1(n_513), .A2(n_492), .B(n_491), .C(n_487), .Y(n_633) );
AND2x2_ASAP7_75t_L g634 ( .A(n_567), .B(n_420), .Y(n_634) );
AOI22xp33_ASAP7_75t_L g635 ( .A1(n_505), .A2(n_331), .B1(n_371), .B2(n_323), .Y(n_635) );
NOR2xp33_ASAP7_75t_L g636 ( .A(n_556), .B(n_323), .Y(n_636) );
CKINVDCx20_ASAP7_75t_R g637 ( .A(n_538), .Y(n_637) );
HB1xp67_ASAP7_75t_L g638 ( .A(n_517), .Y(n_638) );
INVx2_ASAP7_75t_L g639 ( .A(n_566), .Y(n_639) );
OAI22xp5_ASAP7_75t_L g640 ( .A1(n_497), .A2(n_364), .B1(n_375), .B2(n_371), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_566), .Y(n_641) );
INVx2_ASAP7_75t_SL g642 ( .A(n_522), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_570), .Y(n_643) );
OR2x6_ASAP7_75t_L g644 ( .A(n_517), .B(n_345), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_549), .Y(n_645) );
INVx5_ASAP7_75t_L g646 ( .A(n_544), .Y(n_646) );
INVx2_ASAP7_75t_L g647 ( .A(n_570), .Y(n_647) );
BUFx3_ASAP7_75t_L g648 ( .A(n_544), .Y(n_648) );
INVx6_ASAP7_75t_L g649 ( .A(n_503), .Y(n_649) );
AOI22xp33_ASAP7_75t_L g650 ( .A1(n_517), .A2(n_382), .B1(n_375), .B2(n_420), .Y(n_650) );
AOI21xp5_ASAP7_75t_L g651 ( .A1(n_512), .A2(n_483), .B(n_487), .Y(n_651) );
BUFx2_ASAP7_75t_L g652 ( .A(n_523), .Y(n_652) );
BUFx12f_ASAP7_75t_L g653 ( .A(n_533), .Y(n_653) );
INVx1_ASAP7_75t_L g654 ( .A(n_560), .Y(n_654) );
INVx1_ASAP7_75t_L g655 ( .A(n_564), .Y(n_655) );
INVx2_ASAP7_75t_L g656 ( .A(n_500), .Y(n_656) );
AOI21xp5_ASAP7_75t_L g657 ( .A1(n_515), .A2(n_483), .B(n_487), .Y(n_657) );
BUFx2_ASAP7_75t_L g658 ( .A(n_495), .Y(n_658) );
BUFx6f_ASAP7_75t_L g659 ( .A(n_544), .Y(n_659) );
INVx2_ASAP7_75t_SL g660 ( .A(n_544), .Y(n_660) );
BUFx2_ASAP7_75t_L g661 ( .A(n_495), .Y(n_661) );
NOR2x1_ASAP7_75t_L g662 ( .A(n_524), .B(n_420), .Y(n_662) );
INVx1_ASAP7_75t_L g663 ( .A(n_572), .Y(n_663) );
INVx4_ASAP7_75t_L g664 ( .A(n_503), .Y(n_664) );
NOR2xp33_ASAP7_75t_L g665 ( .A(n_556), .B(n_382), .Y(n_665) );
INVx3_ASAP7_75t_L g666 ( .A(n_518), .Y(n_666) );
A2O1A1Ixp33_ASAP7_75t_L g667 ( .A1(n_513), .A2(n_433), .B(n_429), .C(n_440), .Y(n_667) );
AND2x4_ASAP7_75t_L g668 ( .A(n_550), .B(n_457), .Y(n_668) );
INVx1_ASAP7_75t_L g669 ( .A(n_500), .Y(n_669) );
BUFx3_ASAP7_75t_L g670 ( .A(n_518), .Y(n_670) );
BUFx12f_ASAP7_75t_L g671 ( .A(n_538), .Y(n_671) );
INVx1_ASAP7_75t_L g672 ( .A(n_509), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_539), .B(n_494), .Y(n_673) );
HB1xp67_ASAP7_75t_L g674 ( .A(n_540), .Y(n_674) );
AND2x4_ASAP7_75t_L g675 ( .A(n_550), .B(n_457), .Y(n_675) );
AOI22xp33_ASAP7_75t_L g676 ( .A1(n_556), .A2(n_429), .B1(n_433), .B2(n_426), .Y(n_676) );
AND2x2_ASAP7_75t_L g677 ( .A(n_506), .B(n_429), .Y(n_677) );
BUFx2_ASAP7_75t_L g678 ( .A(n_532), .Y(n_678) );
AND2x4_ASAP7_75t_L g679 ( .A(n_550), .B(n_457), .Y(n_679) );
BUFx2_ASAP7_75t_L g680 ( .A(n_532), .Y(n_680) );
CKINVDCx5p33_ASAP7_75t_R g681 ( .A(n_562), .Y(n_681) );
INVx1_ASAP7_75t_L g682 ( .A(n_509), .Y(n_682) );
AND2x2_ASAP7_75t_L g683 ( .A(n_531), .B(n_433), .Y(n_683) );
HB1xp67_ASAP7_75t_L g684 ( .A(n_535), .Y(n_684) );
BUFx3_ASAP7_75t_L g685 ( .A(n_503), .Y(n_685) );
INVx2_ASAP7_75t_L g686 ( .A(n_581), .Y(n_686) );
OAI221xp5_ASAP7_75t_L g687 ( .A1(n_616), .A2(n_559), .B1(n_516), .B2(n_543), .C(n_508), .Y(n_687) );
AOI221xp5_ASAP7_75t_L g688 ( .A1(n_673), .A2(n_561), .B1(n_534), .B2(n_520), .C(n_563), .Y(n_688) );
AND2x4_ASAP7_75t_L g689 ( .A(n_581), .B(n_503), .Y(n_689) );
INVxp67_ASAP7_75t_SL g690 ( .A(n_652), .Y(n_690) );
AOI22xp33_ASAP7_75t_L g691 ( .A1(n_683), .A2(n_514), .B1(n_511), .B2(n_520), .Y(n_691) );
INVx6_ASAP7_75t_L g692 ( .A(n_606), .Y(n_692) );
OR2x6_ASAP7_75t_L g693 ( .A(n_606), .B(n_526), .Y(n_693) );
AOI22xp33_ASAP7_75t_SL g694 ( .A1(n_637), .A2(n_387), .B1(n_411), .B2(n_410), .Y(n_694) );
AND2x4_ASAP7_75t_L g695 ( .A(n_604), .B(n_519), .Y(n_695) );
INVx1_ASAP7_75t_L g696 ( .A(n_592), .Y(n_696) );
AND2x4_ASAP7_75t_L g697 ( .A(n_604), .B(n_519), .Y(n_697) );
INVx2_ASAP7_75t_L g698 ( .A(n_620), .Y(n_698) );
NAND2x1p5_ASAP7_75t_L g699 ( .A(n_586), .B(n_552), .Y(n_699) );
CKINVDCx14_ASAP7_75t_R g700 ( .A(n_612), .Y(n_700) );
INVx1_ASAP7_75t_L g701 ( .A(n_592), .Y(n_701) );
O2A1O1Ixp33_ASAP7_75t_SL g702 ( .A1(n_633), .A2(n_308), .B(n_312), .C(n_307), .Y(n_702) );
OAI22xp5_ASAP7_75t_L g703 ( .A1(n_610), .A2(n_573), .B1(n_534), .B2(n_558), .Y(n_703) );
OAI21x1_ASAP7_75t_L g704 ( .A1(n_657), .A2(n_571), .B(n_492), .Y(n_704) );
AOI22xp33_ASAP7_75t_L g705 ( .A1(n_683), .A2(n_514), .B1(n_536), .B2(n_557), .Y(n_705) );
INVx2_ASAP7_75t_L g706 ( .A(n_620), .Y(n_706) );
AOI221xp5_ASAP7_75t_L g707 ( .A1(n_580), .A2(n_558), .B1(n_557), .B2(n_335), .C(n_344), .Y(n_707) );
INVx1_ASAP7_75t_SL g708 ( .A(n_637), .Y(n_708) );
INVx5_ASAP7_75t_L g709 ( .A(n_579), .Y(n_709) );
AOI22xp33_ASAP7_75t_L g710 ( .A1(n_644), .A2(n_514), .B1(n_536), .B2(n_281), .Y(n_710) );
AOI221xp5_ASAP7_75t_L g711 ( .A1(n_583), .A2(n_383), .B1(n_392), .B2(n_388), .C(n_359), .Y(n_711) );
AOI22xp33_ASAP7_75t_L g712 ( .A1(n_644), .A2(n_514), .B1(n_340), .B2(n_368), .Y(n_712) );
INVx2_ASAP7_75t_L g713 ( .A(n_593), .Y(n_713) );
INVx3_ASAP7_75t_L g714 ( .A(n_586), .Y(n_714) );
NAND3x1_ASAP7_75t_L g715 ( .A(n_624), .B(n_322), .C(n_387), .Y(n_715) );
HB1xp67_ASAP7_75t_L g716 ( .A(n_652), .Y(n_716) );
OR2x6_ASAP7_75t_L g717 ( .A(n_644), .B(n_552), .Y(n_717) );
OAI22xp5_ASAP7_75t_L g718 ( .A1(n_644), .A2(n_630), .B1(n_642), .B2(n_588), .Y(n_718) );
AO31x2_ASAP7_75t_L g719 ( .A1(n_667), .A2(n_440), .A3(n_492), .B(n_491), .Y(n_719) );
AOI22xp33_ASAP7_75t_L g720 ( .A1(n_654), .A2(n_514), .B1(n_377), .B2(n_407), .Y(n_720) );
INVx1_ASAP7_75t_L g721 ( .A(n_634), .Y(n_721) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_634), .B(n_568), .Y(n_722) );
CKINVDCx5p33_ASAP7_75t_R g723 ( .A(n_612), .Y(n_723) );
OAI22xp33_ASAP7_75t_L g724 ( .A1(n_624), .A2(n_410), .B1(n_411), .B2(n_352), .Y(n_724) );
INVx3_ASAP7_75t_L g725 ( .A(n_586), .Y(n_725) );
BUFx2_ASAP7_75t_L g726 ( .A(n_671), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_585), .B(n_548), .Y(n_727) );
CKINVDCx5p33_ASAP7_75t_R g728 ( .A(n_622), .Y(n_728) );
AOI22xp33_ASAP7_75t_L g729 ( .A1(n_654), .A2(n_415), .B1(n_440), .B2(n_548), .Y(n_729) );
INVx1_ASAP7_75t_L g730 ( .A(n_655), .Y(n_730) );
AOI22xp33_ASAP7_75t_SL g731 ( .A1(n_622), .A2(n_400), .B1(n_307), .B2(n_312), .Y(n_731) );
INVx2_ASAP7_75t_L g732 ( .A(n_593), .Y(n_732) );
INVx2_ASAP7_75t_L g733 ( .A(n_597), .Y(n_733) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_585), .B(n_309), .Y(n_734) );
INVx3_ASAP7_75t_L g735 ( .A(n_579), .Y(n_735) );
OA21x2_ASAP7_75t_L g736 ( .A1(n_651), .A2(n_491), .B(n_314), .Y(n_736) );
OAI221xp5_ASAP7_75t_L g737 ( .A1(n_636), .A2(n_279), .B1(n_381), .B2(n_374), .C(n_361), .Y(n_737) );
INVx1_ASAP7_75t_L g738 ( .A(n_655), .Y(n_738) );
AOI221xp5_ASAP7_75t_L g739 ( .A1(n_674), .A2(n_391), .B1(n_399), .B2(n_314), .C(n_316), .Y(n_739) );
INVx1_ASAP7_75t_L g740 ( .A(n_663), .Y(n_740) );
INVx2_ASAP7_75t_L g741 ( .A(n_597), .Y(n_741) );
AOI22xp33_ASAP7_75t_L g742 ( .A1(n_663), .A2(n_308), .B1(n_319), .B2(n_316), .Y(n_742) );
INVx8_ASAP7_75t_L g743 ( .A(n_599), .Y(n_743) );
AOI22xp33_ASAP7_75t_L g744 ( .A1(n_677), .A2(n_319), .B1(n_321), .B2(n_320), .Y(n_744) );
BUFx4f_ASAP7_75t_SL g745 ( .A(n_671), .Y(n_745) );
INVx3_ASAP7_75t_L g746 ( .A(n_579), .Y(n_746) );
NAND2xp5_ASAP7_75t_L g747 ( .A(n_585), .B(n_329), .Y(n_747) );
OAI22xp5_ASAP7_75t_L g748 ( .A1(n_642), .A2(n_553), .B1(n_365), .B2(n_372), .Y(n_748) );
INVx2_ASAP7_75t_L g749 ( .A(n_598), .Y(n_749) );
INVx1_ASAP7_75t_L g750 ( .A(n_595), .Y(n_750) );
INVx1_ASAP7_75t_L g751 ( .A(n_617), .Y(n_751) );
BUFx2_ASAP7_75t_R g752 ( .A(n_681), .Y(n_752) );
INVxp67_ASAP7_75t_SL g753 ( .A(n_607), .Y(n_753) );
AOI22xp5_ASAP7_75t_L g754 ( .A1(n_640), .A2(n_329), .B1(n_372), .B2(n_365), .Y(n_754) );
INVx2_ASAP7_75t_L g755 ( .A(n_598), .Y(n_755) );
OAI22xp5_ASAP7_75t_L g756 ( .A1(n_582), .A2(n_553), .B1(n_390), .B2(n_380), .Y(n_756) );
INVx1_ASAP7_75t_L g757 ( .A(n_677), .Y(n_757) );
INVx1_ASAP7_75t_L g758 ( .A(n_607), .Y(n_758) );
HB1xp67_ASAP7_75t_L g759 ( .A(n_584), .Y(n_759) );
INVx1_ASAP7_75t_L g760 ( .A(n_615), .Y(n_760) );
AND2x2_ASAP7_75t_L g761 ( .A(n_665), .B(n_380), .Y(n_761) );
INVx1_ASAP7_75t_L g762 ( .A(n_615), .Y(n_762) );
AOI22xp33_ASAP7_75t_L g763 ( .A1(n_621), .A2(n_320), .B1(n_324), .B2(n_321), .Y(n_763) );
INVxp67_ASAP7_75t_SL g764 ( .A(n_621), .Y(n_764) );
AOI22xp33_ASAP7_75t_L g765 ( .A1(n_631), .A2(n_324), .B1(n_327), .B2(n_326), .Y(n_765) );
INVx3_ASAP7_75t_L g766 ( .A(n_601), .Y(n_766) );
AND2x2_ASAP7_75t_L g767 ( .A(n_681), .B(n_390), .Y(n_767) );
NAND2xp5_ASAP7_75t_L g768 ( .A(n_628), .B(n_552), .Y(n_768) );
AND2x4_ASAP7_75t_L g769 ( .A(n_584), .B(n_330), .Y(n_769) );
INVx1_ASAP7_75t_L g770 ( .A(n_631), .Y(n_770) );
AND2x2_ASAP7_75t_L g771 ( .A(n_635), .B(n_8), .Y(n_771) );
OAI221xp5_ASAP7_75t_L g772 ( .A1(n_650), .A2(n_347), .B1(n_405), .B2(n_338), .C(n_328), .Y(n_772) );
AOI22xp5_ASAP7_75t_L g773 ( .A1(n_605), .A2(n_628), .B1(n_576), .B2(n_575), .Y(n_773) );
BUFx6f_ASAP7_75t_L g774 ( .A(n_589), .Y(n_774) );
OAI22x1_ASAP7_75t_L g775 ( .A1(n_623), .A2(n_326), .B1(n_328), .B2(n_327), .Y(n_775) );
AOI22xp33_ASAP7_75t_L g776 ( .A1(n_632), .A2(n_386), .B1(n_412), .B2(n_385), .Y(n_776) );
INVx1_ASAP7_75t_SL g777 ( .A(n_575), .Y(n_777) );
AOI22xp33_ASAP7_75t_L g778 ( .A1(n_632), .A2(n_386), .B1(n_412), .B2(n_385), .Y(n_778) );
A2O1A1Ixp33_ASAP7_75t_L g779 ( .A1(n_641), .A2(n_332), .B(n_333), .C(n_290), .Y(n_779) );
AOI22xp33_ASAP7_75t_L g780 ( .A1(n_641), .A2(n_426), .B1(n_442), .B2(n_432), .Y(n_780) );
AOI22xp33_ASAP7_75t_L g781 ( .A1(n_643), .A2(n_442), .B1(n_448), .B2(n_432), .Y(n_781) );
INVx2_ASAP7_75t_L g782 ( .A(n_613), .Y(n_782) );
AOI22xp33_ASAP7_75t_L g783 ( .A1(n_643), .A2(n_442), .B1(n_448), .B2(n_432), .Y(n_783) );
NAND2x1p5_ASAP7_75t_L g784 ( .A(n_576), .B(n_337), .Y(n_784) );
OR2x2_ASAP7_75t_L g785 ( .A(n_613), .B(n_618), .Y(n_785) );
BUFx2_ASAP7_75t_SL g786 ( .A(n_601), .Y(n_786) );
INVx1_ASAP7_75t_L g787 ( .A(n_684), .Y(n_787) );
NAND3xp33_ASAP7_75t_SL g788 ( .A(n_609), .B(n_342), .C(n_341), .Y(n_788) );
OAI21xp5_ASAP7_75t_L g789 ( .A1(n_618), .A2(n_348), .B(n_346), .Y(n_789) );
AOI22xp33_ASAP7_75t_L g790 ( .A1(n_639), .A2(n_442), .B1(n_448), .B2(n_355), .Y(n_790) );
AND2x4_ASAP7_75t_L g791 ( .A(n_601), .B(n_358), .Y(n_791) );
CKINVDCx11_ASAP7_75t_R g792 ( .A(n_626), .Y(n_792) );
OAI21x1_ASAP7_75t_L g793 ( .A1(n_639), .A2(n_363), .B(n_360), .Y(n_793) );
INVx1_ASAP7_75t_L g794 ( .A(n_647), .Y(n_794) );
OAI22xp5_ASAP7_75t_L g795 ( .A1(n_647), .A2(n_396), .B1(n_366), .B2(n_376), .Y(n_795) );
AOI21xp5_ASAP7_75t_L g796 ( .A1(n_629), .A2(n_472), .B(n_453), .Y(n_796) );
AND2x2_ASAP7_75t_L g797 ( .A(n_626), .B(n_9), .Y(n_797) );
INVx4_ASAP7_75t_L g798 ( .A(n_600), .Y(n_798) );
INVx2_ASAP7_75t_L g799 ( .A(n_619), .Y(n_799) );
OAI22xp5_ASAP7_75t_L g800 ( .A1(n_596), .A2(n_403), .B1(n_367), .B2(n_384), .Y(n_800) );
CKINVDCx5p33_ASAP7_75t_R g801 ( .A(n_653), .Y(n_801) );
OR2x2_ASAP7_75t_L g802 ( .A(n_603), .B(n_9), .Y(n_802) );
INVx1_ASAP7_75t_L g803 ( .A(n_645), .Y(n_803) );
INVx3_ASAP7_75t_L g804 ( .A(n_664), .Y(n_804) );
OAI22xp5_ASAP7_75t_L g805 ( .A1(n_638), .A2(n_404), .B1(n_378), .B2(n_393), .Y(n_805) );
OAI22xp33_ASAP7_75t_L g806 ( .A1(n_653), .A2(n_406), .B1(n_389), .B2(n_395), .Y(n_806) );
OR2x2_ASAP7_75t_L g807 ( .A(n_676), .B(n_10), .Y(n_807) );
BUFx12f_ASAP7_75t_L g808 ( .A(n_792), .Y(n_808) );
AOI221xp5_ASAP7_75t_L g809 ( .A1(n_724), .A2(n_682), .B1(n_669), .B2(n_672), .C(n_574), .Y(n_809) );
NAND3xp33_ASAP7_75t_L g810 ( .A(n_731), .B(n_662), .C(n_448), .Y(n_810) );
AOI21xp5_ASAP7_75t_L g811 ( .A1(n_796), .A2(n_577), .B(n_574), .Y(n_811) );
AOI22xp33_ASAP7_75t_L g812 ( .A1(n_724), .A2(n_590), .B1(n_591), .B2(n_577), .Y(n_812) );
BUFx6f_ASAP7_75t_L g813 ( .A(n_774), .Y(n_813) );
OR2x6_ASAP7_75t_L g814 ( .A(n_717), .B(n_578), .Y(n_814) );
OAI22xp5_ASAP7_75t_L g815 ( .A1(n_753), .A2(n_658), .B1(n_678), .B2(n_661), .Y(n_815) );
INVx2_ASAP7_75t_L g816 ( .A(n_785), .Y(n_816) );
NAND2xp5_ASAP7_75t_L g817 ( .A(n_696), .B(n_669), .Y(n_817) );
AOI22xp33_ASAP7_75t_L g818 ( .A1(n_771), .A2(n_591), .B1(n_590), .B2(n_672), .Y(n_818) );
NAND2xp5_ASAP7_75t_L g819 ( .A(n_701), .B(n_682), .Y(n_819) );
NOR2xp67_ASAP7_75t_L g820 ( .A(n_723), .B(n_600), .Y(n_820) );
NAND3xp33_ASAP7_75t_L g821 ( .A(n_731), .B(n_448), .C(n_442), .Y(n_821) );
INVxp67_ASAP7_75t_L g822 ( .A(n_690), .Y(n_822) );
NOR2xp33_ASAP7_75t_L g823 ( .A(n_687), .B(n_656), .Y(n_823) );
INVx3_ASAP7_75t_L g824 ( .A(n_709), .Y(n_824) );
OAI22xp33_ASAP7_75t_L g825 ( .A1(n_753), .A2(n_578), .B1(n_661), .B2(n_658), .Y(n_825) );
INVx1_ASAP7_75t_L g826 ( .A(n_750), .Y(n_826) );
AND2x2_ASAP7_75t_L g827 ( .A(n_767), .B(n_590), .Y(n_827) );
AOI22xp33_ASAP7_75t_L g828 ( .A1(n_694), .A2(n_591), .B1(n_656), .B2(n_678), .Y(n_828) );
OAI22xp5_ASAP7_75t_SL g829 ( .A1(n_700), .A2(n_680), .B1(n_600), .B2(n_646), .Y(n_829) );
A2O1A1Ixp33_ASAP7_75t_L g830 ( .A1(n_764), .A2(n_602), .B(n_611), .C(n_666), .Y(n_830) );
AOI221xp5_ASAP7_75t_L g831 ( .A1(n_711), .A2(n_408), .B1(n_402), .B2(n_413), .C(n_442), .Y(n_831) );
AOI22xp33_ASAP7_75t_SL g832 ( .A1(n_690), .A2(n_680), .B1(n_646), .B2(n_600), .Y(n_832) );
OAI221xp5_ASAP7_75t_L g833 ( .A1(n_694), .A2(n_666), .B1(n_670), .B2(n_660), .C(n_614), .Y(n_833) );
AOI22xp33_ASAP7_75t_SL g834 ( .A1(n_764), .A2(n_646), .B1(n_600), .B2(n_670), .Y(n_834) );
BUFx4f_ASAP7_75t_SL g835 ( .A(n_726), .Y(n_835) );
OR2x2_ASAP7_75t_L g836 ( .A(n_708), .B(n_660), .Y(n_836) );
AOI221xp5_ASAP7_75t_L g837 ( .A1(n_806), .A2(n_448), .B1(n_442), .B2(n_675), .C(n_668), .Y(n_837) );
INVx1_ASAP7_75t_SL g838 ( .A(n_745), .Y(n_838) );
AOI22xp33_ASAP7_75t_SL g839 ( .A1(n_716), .A2(n_646), .B1(n_666), .B2(n_648), .Y(n_839) );
INVx2_ASAP7_75t_L g840 ( .A(n_713), .Y(n_840) );
INVx1_ASAP7_75t_L g841 ( .A(n_751), .Y(n_841) );
INVx1_ASAP7_75t_L g842 ( .A(n_730), .Y(n_842) );
INVx2_ASAP7_75t_L g843 ( .A(n_732), .Y(n_843) );
INVx2_ASAP7_75t_SL g844 ( .A(n_692), .Y(n_844) );
AND2x2_ASAP7_75t_L g845 ( .A(n_686), .B(n_668), .Y(n_845) );
OR2x2_ASAP7_75t_L g846 ( .A(n_698), .B(n_614), .Y(n_846) );
OAI211xp5_ASAP7_75t_L g847 ( .A1(n_737), .A2(n_442), .B(n_448), .C(n_664), .Y(n_847) );
INVxp67_ASAP7_75t_SL g848 ( .A(n_716), .Y(n_848) );
OAI22xp5_ASAP7_75t_L g849 ( .A1(n_712), .A2(n_589), .B1(n_594), .B2(n_625), .Y(n_849) );
NAND3xp33_ASAP7_75t_L g850 ( .A(n_779), .B(n_448), .C(n_453), .Y(n_850) );
AOI22xp33_ASAP7_75t_L g851 ( .A1(n_788), .A2(n_648), .B1(n_350), .B2(n_675), .Y(n_851) );
INVx1_ASAP7_75t_L g852 ( .A(n_738), .Y(n_852) );
INVx1_ASAP7_75t_L g853 ( .A(n_740), .Y(n_853) );
AOI221xp5_ASAP7_75t_L g854 ( .A1(n_806), .A2(n_679), .B1(n_675), .B2(n_668), .C(n_627), .Y(n_854) );
OAI211xp5_ASAP7_75t_L g855 ( .A1(n_739), .A2(n_664), .B(n_608), .C(n_587), .Y(n_855) );
AOI22xp33_ASAP7_75t_L g856 ( .A1(n_757), .A2(n_679), .B1(n_625), .B2(n_659), .Y(n_856) );
BUFx3_ASAP7_75t_L g857 ( .A(n_692), .Y(n_857) );
AOI22xp33_ASAP7_75t_L g858 ( .A1(n_688), .A2(n_679), .B1(n_685), .B2(n_587), .Y(n_858) );
AOI221xp5_ASAP7_75t_L g859 ( .A1(n_772), .A2(n_608), .B1(n_587), .B2(n_627), .C(n_685), .Y(n_859) );
AOI221xp5_ASAP7_75t_L g860 ( .A1(n_721), .A2(n_608), .B1(n_627), .B2(n_453), .C(n_472), .Y(n_860) );
AOI22xp33_ASAP7_75t_L g861 ( .A1(n_712), .A2(n_649), .B1(n_646), .B2(n_659), .Y(n_861) );
BUFx2_ASAP7_75t_L g862 ( .A(n_728), .Y(n_862) );
AOI22xp33_ASAP7_75t_L g863 ( .A1(n_722), .A2(n_649), .B1(n_659), .B2(n_625), .Y(n_863) );
OAI221xp5_ASAP7_75t_L g864 ( .A1(n_691), .A2(n_649), .B1(n_659), .B2(n_625), .C(n_594), .Y(n_864) );
AO21x2_ASAP7_75t_L g865 ( .A1(n_702), .A2(n_472), .B(n_453), .Y(n_865) );
OA21x2_ASAP7_75t_L g866 ( .A1(n_704), .A2(n_472), .B(n_453), .Y(n_866) );
AOI22xp33_ASAP7_75t_L g867 ( .A1(n_691), .A2(n_659), .B1(n_625), .B2(n_594), .Y(n_867) );
INVx1_ASAP7_75t_L g868 ( .A(n_758), .Y(n_868) );
AND2x2_ASAP7_75t_L g869 ( .A(n_706), .B(n_11), .Y(n_869) );
NAND2xp5_ASAP7_75t_L g870 ( .A(n_695), .B(n_589), .Y(n_870) );
HB1xp67_ASAP7_75t_L g871 ( .A(n_759), .Y(n_871) );
OAI211xp5_ASAP7_75t_L g872 ( .A1(n_754), .A2(n_453), .B(n_472), .C(n_589), .Y(n_872) );
AOI22xp33_ASAP7_75t_L g873 ( .A1(n_807), .A2(n_703), .B1(n_762), .B2(n_760), .Y(n_873) );
A2O1A1Ixp33_ASAP7_75t_L g874 ( .A1(n_710), .A2(n_594), .B(n_589), .C(n_472), .Y(n_874) );
AOI22xp33_ASAP7_75t_L g875 ( .A1(n_770), .A2(n_594), .B1(n_649), .B2(n_472), .Y(n_875) );
BUFx2_ASAP7_75t_L g876 ( .A(n_700), .Y(n_876) );
INVx1_ASAP7_75t_L g877 ( .A(n_802), .Y(n_877) );
AOI22xp33_ASAP7_75t_SL g878 ( .A1(n_743), .A2(n_11), .B1(n_12), .B2(n_13), .Y(n_878) );
OA21x2_ASAP7_75t_L g879 ( .A1(n_793), .A2(n_453), .B(n_94), .Y(n_879) );
AND2x4_ASAP7_75t_L g880 ( .A(n_709), .B(n_13), .Y(n_880) );
OAI21xp5_ASAP7_75t_SL g881 ( .A1(n_784), .A2(n_14), .B(n_15), .Y(n_881) );
BUFx6f_ASAP7_75t_L g882 ( .A(n_774), .Y(n_882) );
OAI22xp5_ASAP7_75t_L g883 ( .A1(n_717), .A2(n_14), .B1(n_16), .B2(n_17), .Y(n_883) );
CKINVDCx20_ASAP7_75t_R g884 ( .A(n_745), .Y(n_884) );
OAI21x1_ASAP7_75t_L g885 ( .A1(n_736), .A2(n_95), .B(n_84), .Y(n_885) );
AOI22xp33_ASAP7_75t_SL g886 ( .A1(n_743), .A2(n_16), .B1(n_17), .B2(n_18), .Y(n_886) );
OAI21xp5_ASAP7_75t_L g887 ( .A1(n_720), .A2(n_18), .B(n_19), .Y(n_887) );
NAND2xp5_ASAP7_75t_L g888 ( .A(n_695), .B(n_19), .Y(n_888) );
AOI221xp5_ASAP7_75t_L g889 ( .A1(n_707), .A2(n_20), .B1(n_21), .B2(n_22), .C(n_24), .Y(n_889) );
AND2x2_ASAP7_75t_L g890 ( .A(n_761), .B(n_797), .Y(n_890) );
NOR2xp33_ASAP7_75t_L g891 ( .A(n_697), .B(n_21), .Y(n_891) );
AOI221xp5_ASAP7_75t_L g892 ( .A1(n_744), .A2(n_22), .B1(n_25), .B2(n_26), .C(n_28), .Y(n_892) );
AOI21xp5_ASAP7_75t_L g893 ( .A1(n_702), .A2(n_98), .B(n_97), .Y(n_893) );
AND2x2_ASAP7_75t_L g894 ( .A(n_697), .B(n_25), .Y(n_894) );
AOI221xp5_ASAP7_75t_L g895 ( .A1(n_744), .A2(n_28), .B1(n_29), .B2(n_30), .C(n_32), .Y(n_895) );
CKINVDCx5p33_ASAP7_75t_R g896 ( .A(n_743), .Y(n_896) );
A2O1A1Ixp33_ASAP7_75t_L g897 ( .A1(n_710), .A2(n_29), .B(n_30), .C(n_32), .Y(n_897) );
INVx4_ASAP7_75t_L g898 ( .A(n_709), .Y(n_898) );
AOI22xp33_ASAP7_75t_SL g899 ( .A1(n_718), .A2(n_33), .B1(n_35), .B2(n_36), .Y(n_899) );
INVx4_ASAP7_75t_L g900 ( .A(n_709), .Y(n_900) );
INVx2_ASAP7_75t_L g901 ( .A(n_733), .Y(n_901) );
OAI22xp5_ASAP7_75t_L g902 ( .A1(n_717), .A2(n_33), .B1(n_36), .B2(n_37), .Y(n_902) );
INVx1_ASAP7_75t_L g903 ( .A(n_803), .Y(n_903) );
AOI22xp5_ASAP7_75t_L g904 ( .A1(n_715), .A2(n_37), .B1(n_38), .B2(n_39), .Y(n_904) );
INVx2_ASAP7_75t_L g905 ( .A(n_741), .Y(n_905) );
AND2x2_ASAP7_75t_L g906 ( .A(n_784), .B(n_38), .Y(n_906) );
AOI221xp5_ASAP7_75t_L g907 ( .A1(n_779), .A2(n_39), .B1(n_40), .B2(n_41), .C(n_42), .Y(n_907) );
AND2x4_ASAP7_75t_L g908 ( .A(n_689), .B(n_40), .Y(n_908) );
AOI22xp33_ASAP7_75t_L g909 ( .A1(n_789), .A2(n_41), .B1(n_42), .B2(n_43), .Y(n_909) );
INVx3_ASAP7_75t_L g910 ( .A(n_798), .Y(n_910) );
AOI22xp33_ASAP7_75t_L g911 ( .A1(n_705), .A2(n_43), .B1(n_45), .B2(n_46), .Y(n_911) );
BUFx6f_ASAP7_75t_L g912 ( .A(n_774), .Y(n_912) );
AND2x2_ASAP7_75t_L g913 ( .A(n_777), .B(n_45), .Y(n_913) );
OAI211xp5_ASAP7_75t_L g914 ( .A1(n_742), .A2(n_46), .B(n_47), .C(n_48), .Y(n_914) );
INVx3_ASAP7_75t_SL g915 ( .A(n_692), .Y(n_915) );
OAI33xp33_ASAP7_75t_L g916 ( .A1(n_795), .A2(n_47), .A3(n_48), .B1(n_49), .B2(n_50), .B3(n_51), .Y(n_916) );
CKINVDCx11_ASAP7_75t_R g917 ( .A(n_693), .Y(n_917) );
AOI221xp5_ASAP7_75t_L g918 ( .A1(n_800), .A2(n_49), .B1(n_50), .B2(n_51), .C(n_52), .Y(n_918) );
AOI22xp33_ASAP7_75t_L g919 ( .A1(n_705), .A2(n_52), .B1(n_53), .B2(n_54), .Y(n_919) );
AOI22xp33_ASAP7_75t_L g920 ( .A1(n_775), .A2(n_55), .B1(n_56), .B2(n_57), .Y(n_920) );
INVx1_ASAP7_75t_L g921 ( .A(n_799), .Y(n_921) );
OAI22xp5_ASAP7_75t_L g922 ( .A1(n_720), .A2(n_55), .B1(n_56), .B2(n_60), .Y(n_922) );
BUFx3_ASAP7_75t_L g923 ( .A(n_801), .Y(n_923) );
NAND3xp33_ASAP7_75t_L g924 ( .A(n_904), .B(n_765), .C(n_763), .Y(n_924) );
INVx1_ASAP7_75t_L g925 ( .A(n_826), .Y(n_925) );
AOI22xp33_ASAP7_75t_L g926 ( .A1(n_899), .A2(n_759), .B1(n_791), .B2(n_742), .Y(n_926) );
AND2x2_ASAP7_75t_L g927 ( .A(n_890), .B(n_769), .Y(n_927) );
AND2x2_ASAP7_75t_L g928 ( .A(n_906), .B(n_769), .Y(n_928) );
NAND2xp33_ASAP7_75t_L g929 ( .A(n_851), .B(n_748), .Y(n_929) );
INVx2_ASAP7_75t_L g930 ( .A(n_866), .Y(n_930) );
AOI222xp33_ASAP7_75t_L g931 ( .A1(n_887), .A2(n_805), .B1(n_787), .B2(n_765), .C1(n_763), .C2(n_776), .Y(n_931) );
INVx2_ASAP7_75t_L g932 ( .A(n_866), .Y(n_932) );
AND2x4_ASAP7_75t_SL g933 ( .A(n_884), .B(n_693), .Y(n_933) );
AOI221xp5_ASAP7_75t_L g934 ( .A1(n_877), .A2(n_778), .B1(n_776), .B2(n_729), .C(n_747), .Y(n_934) );
OAI211xp5_ASAP7_75t_SL g935 ( .A1(n_878), .A2(n_778), .B(n_773), .C(n_734), .Y(n_935) );
OAI22xp33_ASAP7_75t_L g936 ( .A1(n_881), .A2(n_693), .B1(n_725), .B2(n_714), .Y(n_936) );
INVx1_ASAP7_75t_L g937 ( .A(n_841), .Y(n_937) );
OAI21xp33_ASAP7_75t_L g938 ( .A1(n_899), .A2(n_752), .B(n_791), .Y(n_938) );
INVx2_ASAP7_75t_L g939 ( .A(n_840), .Y(n_939) );
AOI22xp5_ASAP7_75t_L g940 ( .A1(n_854), .A2(n_786), .B1(n_689), .B2(n_756), .Y(n_940) );
INVx2_ASAP7_75t_SL g941 ( .A(n_835), .Y(n_941) );
AOI22xp33_ASAP7_75t_L g942 ( .A1(n_823), .A2(n_729), .B1(n_714), .B2(n_725), .Y(n_942) );
INVxp67_ASAP7_75t_SL g943 ( .A(n_816), .Y(n_943) );
AOI33xp33_ASAP7_75t_L g944 ( .A1(n_878), .A2(n_790), .A3(n_781), .B1(n_783), .B2(n_780), .B3(n_794), .Y(n_944) );
AOI21xp5_ASAP7_75t_SL g945 ( .A1(n_880), .A2(n_798), .B(n_699), .Y(n_945) );
OAI22xp5_ASAP7_75t_L g946 ( .A1(n_873), .A2(n_727), .B1(n_782), .B2(n_749), .Y(n_946) );
OAI22xp5_ASAP7_75t_L g947 ( .A1(n_873), .A2(n_755), .B1(n_766), .B2(n_746), .Y(n_947) );
AOI22xp5_ASAP7_75t_L g948 ( .A1(n_827), .A2(n_735), .B1(n_746), .B2(n_766), .Y(n_948) );
OAI33xp33_ASAP7_75t_L g949 ( .A1(n_883), .A2(n_768), .A3(n_63), .B1(n_64), .B2(n_65), .B3(n_66), .Y(n_949) );
AND2x2_ASAP7_75t_L g950 ( .A(n_894), .B(n_735), .Y(n_950) );
OAI211xp5_ASAP7_75t_L g951 ( .A1(n_886), .A2(n_790), .B(n_783), .C(n_781), .Y(n_951) );
INVx4_ASAP7_75t_R g952 ( .A(n_838), .Y(n_952) );
INVx1_ASAP7_75t_L g953 ( .A(n_903), .Y(n_953) );
OAI33xp33_ASAP7_75t_L g954 ( .A1(n_902), .A2(n_60), .A3(n_64), .B1(n_66), .B2(n_67), .B3(n_68), .Y(n_954) );
AOI22xp33_ASAP7_75t_L g955 ( .A1(n_916), .A2(n_736), .B1(n_804), .B2(n_780), .Y(n_955) );
NAND2xp5_ASAP7_75t_L g956 ( .A(n_842), .B(n_719), .Y(n_956) );
AOI221xp5_ASAP7_75t_L g957 ( .A1(n_922), .A2(n_804), .B1(n_699), .B2(n_719), .C(n_774), .Y(n_957) );
AND2x2_ASAP7_75t_L g958 ( .A(n_908), .B(n_69), .Y(n_958) );
AOI22xp33_ASAP7_75t_L g959 ( .A1(n_809), .A2(n_736), .B1(n_719), .B2(n_71), .Y(n_959) );
OAI211xp5_ASAP7_75t_L g960 ( .A1(n_886), .A2(n_719), .B(n_70), .C(n_71), .Y(n_960) );
AOI22xp5_ASAP7_75t_L g961 ( .A1(n_908), .A2(n_69), .B1(n_70), .B2(n_72), .Y(n_961) );
INVx5_ASAP7_75t_SL g962 ( .A(n_814), .Y(n_962) );
INVx2_ASAP7_75t_L g963 ( .A(n_843), .Y(n_963) );
AOI21xp5_ASAP7_75t_L g964 ( .A1(n_874), .A2(n_189), .B(n_277), .Y(n_964) );
OAI21xp5_ASAP7_75t_L g965 ( .A1(n_821), .A2(n_72), .B(n_73), .Y(n_965) );
OAI33xp33_ASAP7_75t_L g966 ( .A1(n_888), .A2(n_74), .A3(n_75), .B1(n_77), .B2(n_78), .B3(n_79), .Y(n_966) );
CKINVDCx5p33_ASAP7_75t_R g967 ( .A(n_808), .Y(n_967) );
AOI22xp33_ASAP7_75t_L g968 ( .A1(n_911), .A2(n_74), .B1(n_75), .B2(n_77), .Y(n_968) );
OAI321xp33_ASAP7_75t_L g969 ( .A1(n_911), .A2(n_78), .A3(n_79), .B1(n_80), .B2(n_82), .C(n_99), .Y(n_969) );
BUFx2_ASAP7_75t_L g970 ( .A(n_835), .Y(n_970) );
AOI22xp33_ASAP7_75t_L g971 ( .A1(n_907), .A2(n_80), .B1(n_102), .B2(n_105), .Y(n_971) );
OAI221xp5_ASAP7_75t_L g972 ( .A1(n_920), .A2(n_108), .B1(n_109), .B2(n_111), .C(n_114), .Y(n_972) );
AND2x2_ASAP7_75t_L g973 ( .A(n_913), .B(n_115), .Y(n_973) );
INVx2_ASAP7_75t_L g974 ( .A(n_901), .Y(n_974) );
OAI21x1_ASAP7_75t_L g975 ( .A1(n_811), .A2(n_116), .B(n_117), .Y(n_975) );
AOI21xp33_ASAP7_75t_SL g976 ( .A1(n_915), .A2(n_119), .B(n_120), .Y(n_976) );
AOI21xp33_ASAP7_75t_L g977 ( .A1(n_847), .A2(n_122), .B(n_123), .Y(n_977) );
AND2x6_ASAP7_75t_L g978 ( .A(n_880), .B(n_124), .Y(n_978) );
INVx2_ASAP7_75t_L g979 ( .A(n_905), .Y(n_979) );
AOI221xp5_ASAP7_75t_L g980 ( .A1(n_889), .A2(n_125), .B1(n_127), .B2(n_129), .C(n_130), .Y(n_980) );
NOR2xp33_ASAP7_75t_L g981 ( .A(n_845), .B(n_132), .Y(n_981) );
BUFx2_ASAP7_75t_L g982 ( .A(n_898), .Y(n_982) );
AOI221xp5_ASAP7_75t_L g983 ( .A1(n_831), .A2(n_133), .B1(n_134), .B2(n_135), .C(n_137), .Y(n_983) );
OAI31xp33_ASAP7_75t_L g984 ( .A1(n_914), .A2(n_143), .A3(n_145), .B(n_151), .Y(n_984) );
INVx1_ASAP7_75t_L g985 ( .A(n_852), .Y(n_985) );
OAI22xp5_ASAP7_75t_L g986 ( .A1(n_920), .A2(n_153), .B1(n_154), .B2(n_155), .Y(n_986) );
OAI33xp33_ASAP7_75t_L g987 ( .A1(n_853), .A2(n_159), .A3(n_163), .B1(n_164), .B2(n_165), .B3(n_167), .Y(n_987) );
NAND2xp5_ASAP7_75t_L g988 ( .A(n_868), .B(n_168), .Y(n_988) );
AO21x2_ASAP7_75t_L g989 ( .A1(n_865), .A2(n_169), .B(n_170), .Y(n_989) );
OA21x2_ASAP7_75t_L g990 ( .A1(n_885), .A2(n_173), .B(n_174), .Y(n_990) );
OAI21x1_ASAP7_75t_L g991 ( .A1(n_849), .A2(n_175), .B(n_179), .Y(n_991) );
AOI221xp5_ASAP7_75t_L g992 ( .A1(n_918), .A2(n_180), .B1(n_190), .B2(n_192), .C(n_194), .Y(n_992) );
INVx2_ASAP7_75t_L g993 ( .A(n_813), .Y(n_993) );
AOI22xp5_ASAP7_75t_L g994 ( .A1(n_891), .A2(n_195), .B1(n_198), .B2(n_199), .Y(n_994) );
OAI211xp5_ASAP7_75t_L g995 ( .A1(n_851), .A2(n_200), .B(n_201), .C(n_202), .Y(n_995) );
OAI22xp5_ASAP7_75t_L g996 ( .A1(n_822), .A2(n_203), .B1(n_204), .B2(n_207), .Y(n_996) );
BUFx3_ASAP7_75t_L g997 ( .A(n_915), .Y(n_997) );
AOI222xp33_ASAP7_75t_L g998 ( .A1(n_917), .A2(n_209), .B1(n_211), .B2(n_213), .C1(n_216), .C2(n_217), .Y(n_998) );
OAI221xp5_ASAP7_75t_L g999 ( .A1(n_858), .A2(n_219), .B1(n_220), .B2(n_223), .C(n_225), .Y(n_999) );
NAND2xp5_ASAP7_75t_L g1000 ( .A(n_848), .B(n_278), .Y(n_1000) );
OAI211xp5_ASAP7_75t_L g1001 ( .A1(n_909), .A2(n_226), .B(n_227), .C(n_230), .Y(n_1001) );
OAI221xp5_ASAP7_75t_L g1002 ( .A1(n_909), .A2(n_231), .B1(n_232), .B2(n_233), .C(n_235), .Y(n_1002) );
AND2x2_ASAP7_75t_L g1003 ( .A(n_848), .B(n_236), .Y(n_1003) );
OAI211xp5_ASAP7_75t_L g1004 ( .A1(n_892), .A2(n_238), .B(n_242), .C(n_243), .Y(n_1004) );
AOI221xp5_ASAP7_75t_L g1005 ( .A1(n_895), .A2(n_244), .B1(n_247), .B2(n_253), .C(n_254), .Y(n_1005) );
NOR2xp33_ASAP7_75t_SL g1006 ( .A(n_896), .B(n_272), .Y(n_1006) );
OAI221xp5_ASAP7_75t_L g1007 ( .A1(n_837), .A2(n_255), .B1(n_257), .B2(n_258), .C(n_259), .Y(n_1007) );
NAND3xp33_ASAP7_75t_L g1008 ( .A(n_897), .B(n_261), .C(n_263), .Y(n_1008) );
INVx1_ASAP7_75t_L g1009 ( .A(n_921), .Y(n_1009) );
OAI22xp5_ASAP7_75t_L g1010 ( .A1(n_822), .A2(n_828), .B1(n_814), .B2(n_810), .Y(n_1010) );
NAND2xp5_ASAP7_75t_L g1011 ( .A(n_869), .B(n_265), .Y(n_1011) );
AOI21xp5_ASAP7_75t_L g1012 ( .A1(n_864), .A2(n_266), .B(n_268), .Y(n_1012) );
BUFx3_ASAP7_75t_L g1013 ( .A(n_857), .Y(n_1013) );
OAI31xp33_ASAP7_75t_L g1014 ( .A1(n_825), .A2(n_269), .A3(n_270), .B(n_271), .Y(n_1014) );
OAI21xp5_ASAP7_75t_SL g1015 ( .A1(n_876), .A2(n_828), .B(n_919), .Y(n_1015) );
AND2x2_ASAP7_75t_L g1016 ( .A(n_871), .B(n_820), .Y(n_1016) );
AOI22xp33_ASAP7_75t_L g1017 ( .A1(n_871), .A2(n_862), .B1(n_850), .B2(n_814), .Y(n_1017) );
OAI321xp33_ASAP7_75t_L g1018 ( .A1(n_812), .A2(n_825), .A3(n_833), .B1(n_855), .B2(n_818), .C(n_829), .Y(n_1018) );
INVx1_ASAP7_75t_L g1019 ( .A(n_817), .Y(n_1019) );
INVx2_ASAP7_75t_L g1020 ( .A(n_813), .Y(n_1020) );
NAND2xp5_ASAP7_75t_L g1021 ( .A(n_819), .B(n_836), .Y(n_1021) );
OAI211xp5_ASAP7_75t_SL g1022 ( .A1(n_844), .A2(n_812), .B(n_824), .C(n_818), .Y(n_1022) );
INVx2_ASAP7_75t_L g1023 ( .A(n_813), .Y(n_1023) );
AOI22xp33_ASAP7_75t_L g1024 ( .A1(n_898), .A2(n_900), .B1(n_824), .B2(n_815), .Y(n_1024) );
HB1xp67_ASAP7_75t_L g1025 ( .A(n_943), .Y(n_1025) );
AOI221xp5_ASAP7_75t_L g1026 ( .A1(n_938), .A2(n_923), .B1(n_830), .B2(n_910), .C(n_900), .Y(n_1026) );
AND2x2_ASAP7_75t_L g1027 ( .A(n_939), .B(n_910), .Y(n_1027) );
AND2x2_ASAP7_75t_L g1028 ( .A(n_939), .B(n_867), .Y(n_1028) );
INVx1_ASAP7_75t_L g1029 ( .A(n_956), .Y(n_1029) );
INVx1_ASAP7_75t_L g1030 ( .A(n_930), .Y(n_1030) );
INVx2_ASAP7_75t_L g1031 ( .A(n_930), .Y(n_1031) );
INVx5_ASAP7_75t_L g1032 ( .A(n_978), .Y(n_1032) );
AND2x2_ASAP7_75t_L g1033 ( .A(n_963), .B(n_867), .Y(n_1033) );
NAND2xp33_ASAP7_75t_L g1034 ( .A(n_978), .B(n_861), .Y(n_1034) );
INVx2_ASAP7_75t_L g1035 ( .A(n_932), .Y(n_1035) );
INVx2_ASAP7_75t_SL g1036 ( .A(n_982), .Y(n_1036) );
HB1xp67_ASAP7_75t_L g1037 ( .A(n_963), .Y(n_1037) );
AND2x2_ASAP7_75t_L g1038 ( .A(n_974), .B(n_813), .Y(n_1038) );
INVx1_ASAP7_75t_L g1039 ( .A(n_932), .Y(n_1039) );
AOI21xp5_ASAP7_75t_L g1040 ( .A1(n_936), .A2(n_872), .B(n_865), .Y(n_1040) );
INVx2_ASAP7_75t_L g1041 ( .A(n_974), .Y(n_1041) );
INVx1_ASAP7_75t_L g1042 ( .A(n_979), .Y(n_1042) );
NAND3xp33_ASAP7_75t_L g1043 ( .A(n_929), .B(n_1015), .C(n_961), .Y(n_1043) );
INVx1_ASAP7_75t_L g1044 ( .A(n_979), .Y(n_1044) );
OR2x2_ASAP7_75t_L g1045 ( .A(n_1021), .B(n_870), .Y(n_1045) );
NOR3xp33_ASAP7_75t_L g1046 ( .A(n_935), .B(n_832), .C(n_839), .Y(n_1046) );
HB1xp67_ASAP7_75t_L g1047 ( .A(n_1016), .Y(n_1047) );
OR2x2_ASAP7_75t_L g1048 ( .A(n_985), .B(n_846), .Y(n_1048) );
INVx1_ASAP7_75t_L g1049 ( .A(n_925), .Y(n_1049) );
NAND2xp5_ASAP7_75t_L g1050 ( .A(n_1019), .B(n_832), .Y(n_1050) );
AND2x2_ASAP7_75t_L g1051 ( .A(n_937), .B(n_882), .Y(n_1051) );
INVx1_ASAP7_75t_L g1052 ( .A(n_953), .Y(n_1052) );
INVx1_ASAP7_75t_L g1053 ( .A(n_1009), .Y(n_1053) );
AND2x4_ASAP7_75t_L g1054 ( .A(n_993), .B(n_912), .Y(n_1054) );
OA21x2_ASAP7_75t_L g1055 ( .A1(n_957), .A2(n_893), .B(n_875), .Y(n_1055) );
AOI221xp5_ASAP7_75t_L g1056 ( .A1(n_949), .A2(n_859), .B1(n_860), .B2(n_856), .C(n_863), .Y(n_1056) );
OR2x2_ASAP7_75t_L g1057 ( .A(n_962), .B(n_856), .Y(n_1057) );
INVx4_ASAP7_75t_L g1058 ( .A(n_978), .Y(n_1058) );
BUFx3_ASAP7_75t_L g1059 ( .A(n_997), .Y(n_1059) );
OAI211xp5_ASAP7_75t_L g1060 ( .A1(n_926), .A2(n_834), .B(n_839), .C(n_875), .Y(n_1060) );
OAI33xp33_ASAP7_75t_L g1061 ( .A1(n_936), .A2(n_834), .A3(n_879), .B1(n_882), .B2(n_912), .B3(n_1010), .Y(n_1061) );
INVx1_ASAP7_75t_L g1062 ( .A(n_993), .Y(n_1062) );
OAI221xp5_ASAP7_75t_L g1063 ( .A1(n_926), .A2(n_879), .B1(n_882), .B2(n_912), .C(n_968), .Y(n_1063) );
BUFx3_ASAP7_75t_L g1064 ( .A(n_997), .Y(n_1064) );
NAND3xp33_ASAP7_75t_L g1065 ( .A(n_1017), .B(n_882), .C(n_912), .Y(n_1065) );
INVx1_ASAP7_75t_L g1066 ( .A(n_1020), .Y(n_1066) );
INVx4_ASAP7_75t_L g1067 ( .A(n_978), .Y(n_1067) );
NAND2xp5_ASAP7_75t_L g1068 ( .A(n_928), .B(n_927), .Y(n_1068) );
BUFx2_ASAP7_75t_L g1069 ( .A(n_978), .Y(n_1069) );
AND2x2_ASAP7_75t_L g1070 ( .A(n_1020), .B(n_1023), .Y(n_1070) );
AOI222xp33_ASAP7_75t_L g1071 ( .A1(n_954), .A2(n_924), .B1(n_958), .B2(n_966), .C1(n_934), .C2(n_933), .Y(n_1071) );
AOI33xp33_ASAP7_75t_L g1072 ( .A1(n_968), .A2(n_933), .A3(n_959), .B1(n_950), .B2(n_941), .B3(n_1017), .Y(n_1072) );
BUFx3_ASAP7_75t_L g1073 ( .A(n_970), .Y(n_1073) );
INVx2_ASAP7_75t_L g1074 ( .A(n_1023), .Y(n_1074) );
AND2x2_ASAP7_75t_L g1075 ( .A(n_959), .B(n_1003), .Y(n_1075) );
AND2x2_ASAP7_75t_L g1076 ( .A(n_1024), .B(n_948), .Y(n_1076) );
NAND2xp5_ASAP7_75t_L g1077 ( .A(n_931), .B(n_962), .Y(n_1077) );
AND2x2_ASAP7_75t_L g1078 ( .A(n_1024), .B(n_955), .Y(n_1078) );
INVx1_ASAP7_75t_L g1079 ( .A(n_1022), .Y(n_1079) );
INVx2_ASAP7_75t_L g1080 ( .A(n_989), .Y(n_1080) );
INVxp67_ASAP7_75t_SL g1081 ( .A(n_946), .Y(n_1081) );
NAND2xp5_ASAP7_75t_L g1082 ( .A(n_962), .B(n_1013), .Y(n_1082) );
AND2x2_ASAP7_75t_L g1083 ( .A(n_955), .B(n_973), .Y(n_1083) );
OR2x2_ASAP7_75t_L g1084 ( .A(n_1000), .B(n_947), .Y(n_1084) );
INVx1_ASAP7_75t_L g1085 ( .A(n_988), .Y(n_1085) );
AOI22xp33_ASAP7_75t_L g1086 ( .A1(n_998), .A2(n_942), .B1(n_972), .B2(n_971), .Y(n_1086) );
INVx2_ASAP7_75t_L g1087 ( .A(n_990), .Y(n_1087) );
INVx1_ASAP7_75t_L g1088 ( .A(n_990), .Y(n_1088) );
AND2x2_ASAP7_75t_L g1089 ( .A(n_942), .B(n_944), .Y(n_1089) );
OAI21x1_ASAP7_75t_L g1090 ( .A1(n_991), .A2(n_964), .B(n_975), .Y(n_1090) );
OAI21x1_ASAP7_75t_L g1091 ( .A1(n_1012), .A2(n_990), .B(n_965), .Y(n_1091) );
AND2x4_ASAP7_75t_L g1092 ( .A(n_1008), .B(n_994), .Y(n_1092) );
AND2x2_ASAP7_75t_L g1093 ( .A(n_944), .B(n_981), .Y(n_1093) );
OR2x2_ASAP7_75t_L g1094 ( .A(n_1013), .B(n_945), .Y(n_1094) );
BUFx2_ASAP7_75t_L g1095 ( .A(n_940), .Y(n_1095) );
AOI21xp5_ASAP7_75t_L g1096 ( .A1(n_1018), .A2(n_987), .B(n_977), .Y(n_1096) );
NAND2xp33_ASAP7_75t_L g1097 ( .A(n_971), .B(n_986), .Y(n_1097) );
OAI221xp5_ASAP7_75t_L g1098 ( .A1(n_960), .A2(n_1014), .B1(n_984), .B2(n_995), .C(n_981), .Y(n_1098) );
HB1xp67_ASAP7_75t_L g1099 ( .A(n_1011), .Y(n_1099) );
INVx1_ASAP7_75t_L g1100 ( .A(n_996), .Y(n_1100) );
AOI33xp33_ASAP7_75t_L g1101 ( .A1(n_992), .A2(n_980), .A3(n_1005), .B1(n_952), .B2(n_983), .B3(n_969), .Y(n_1101) );
OAI31xp33_ASAP7_75t_L g1102 ( .A1(n_951), .A2(n_1001), .A3(n_1002), .B(n_1004), .Y(n_1102) );
INVx1_ASAP7_75t_L g1103 ( .A(n_976), .Y(n_1103) );
INVx1_ASAP7_75t_L g1104 ( .A(n_999), .Y(n_1104) );
AO21x2_ASAP7_75t_L g1105 ( .A1(n_1007), .A2(n_1006), .B(n_967), .Y(n_1105) );
HB1xp67_ASAP7_75t_L g1106 ( .A(n_943), .Y(n_1106) );
AND2x4_ASAP7_75t_L g1107 ( .A(n_930), .B(n_932), .Y(n_1107) );
INVx1_ASAP7_75t_L g1108 ( .A(n_956), .Y(n_1108) );
BUFx2_ASAP7_75t_SL g1109 ( .A(n_978), .Y(n_1109) );
HB1xp67_ASAP7_75t_L g1110 ( .A(n_943), .Y(n_1110) );
AND2x2_ASAP7_75t_L g1111 ( .A(n_939), .B(n_963), .Y(n_1111) );
INVx1_ASAP7_75t_L g1112 ( .A(n_1049), .Y(n_1112) );
INVx2_ASAP7_75t_L g1113 ( .A(n_1031), .Y(n_1113) );
INVx1_ASAP7_75t_L g1114 ( .A(n_1049), .Y(n_1114) );
NAND2xp5_ASAP7_75t_L g1115 ( .A(n_1025), .B(n_1106), .Y(n_1115) );
AND2x2_ASAP7_75t_L g1116 ( .A(n_1029), .B(n_1108), .Y(n_1116) );
OR2x2_ASAP7_75t_L g1117 ( .A(n_1110), .B(n_1047), .Y(n_1117) );
INVx2_ASAP7_75t_L g1118 ( .A(n_1031), .Y(n_1118) );
INVx2_ASAP7_75t_SL g1119 ( .A(n_1036), .Y(n_1119) );
INVx1_ASAP7_75t_L g1120 ( .A(n_1052), .Y(n_1120) );
OR2x2_ASAP7_75t_L g1121 ( .A(n_1036), .B(n_1037), .Y(n_1121) );
INVx2_ASAP7_75t_SL g1122 ( .A(n_1032), .Y(n_1122) );
AND2x2_ASAP7_75t_L g1123 ( .A(n_1029), .B(n_1108), .Y(n_1123) );
AOI31xp33_ASAP7_75t_L g1124 ( .A1(n_1043), .A2(n_1094), .A3(n_1026), .B(n_1071), .Y(n_1124) );
INVx2_ASAP7_75t_L g1125 ( .A(n_1035), .Y(n_1125) );
BUFx2_ASAP7_75t_L g1126 ( .A(n_1059), .Y(n_1126) );
OR2x2_ASAP7_75t_L g1127 ( .A(n_1030), .B(n_1039), .Y(n_1127) );
INVx1_ASAP7_75t_SL g1128 ( .A(n_1059), .Y(n_1128) );
NAND2xp5_ASAP7_75t_L g1129 ( .A(n_1053), .B(n_1052), .Y(n_1129) );
OR2x2_ASAP7_75t_L g1130 ( .A(n_1053), .B(n_1045), .Y(n_1130) );
OAI322xp33_ASAP7_75t_L g1131 ( .A1(n_1079), .A2(n_1077), .A3(n_1048), .B1(n_1045), .B2(n_1050), .C1(n_1089), .C2(n_1081), .Y(n_1131) );
INVx1_ASAP7_75t_L g1132 ( .A(n_1048), .Y(n_1132) );
AND2x2_ASAP7_75t_L g1133 ( .A(n_1107), .B(n_1039), .Y(n_1133) );
AND2x2_ASAP7_75t_L g1134 ( .A(n_1107), .B(n_1111), .Y(n_1134) );
INVx1_ASAP7_75t_L g1135 ( .A(n_1042), .Y(n_1135) );
NAND2xp5_ASAP7_75t_L g1136 ( .A(n_1089), .B(n_1093), .Y(n_1136) );
NOR2xp33_ASAP7_75t_SL g1137 ( .A(n_1058), .B(n_1067), .Y(n_1137) );
INVx1_ASAP7_75t_L g1138 ( .A(n_1042), .Y(n_1138) );
NAND2xp5_ASAP7_75t_L g1139 ( .A(n_1093), .B(n_1111), .Y(n_1139) );
OAI221xp5_ASAP7_75t_L g1140 ( .A1(n_1086), .A2(n_1099), .B1(n_1046), .B2(n_1079), .C(n_1102), .Y(n_1140) );
AOI22xp5_ASAP7_75t_L g1141 ( .A1(n_1095), .A2(n_1097), .B1(n_1076), .B2(n_1060), .Y(n_1141) );
NOR4xp25_ASAP7_75t_L g1142 ( .A(n_1072), .B(n_1068), .C(n_1063), .D(n_1098), .Y(n_1142) );
BUFx3_ASAP7_75t_L g1143 ( .A(n_1064), .Y(n_1143) );
NAND3xp33_ASAP7_75t_L g1144 ( .A(n_1103), .B(n_1096), .C(n_1056), .Y(n_1144) );
OR2x2_ASAP7_75t_L g1145 ( .A(n_1044), .B(n_1041), .Y(n_1145) );
CKINVDCx16_ASAP7_75t_R g1146 ( .A(n_1073), .Y(n_1146) );
NOR2xp33_ASAP7_75t_L g1147 ( .A(n_1095), .B(n_1085), .Y(n_1147) );
NOR2xp33_ASAP7_75t_L g1148 ( .A(n_1085), .B(n_1076), .Y(n_1148) );
NOR2xp33_ASAP7_75t_L g1149 ( .A(n_1073), .B(n_1094), .Y(n_1149) );
INVx1_ASAP7_75t_L g1150 ( .A(n_1051), .Y(n_1150) );
INVx1_ASAP7_75t_L g1151 ( .A(n_1051), .Y(n_1151) );
OR2x2_ASAP7_75t_L g1152 ( .A(n_1041), .B(n_1064), .Y(n_1152) );
INVx1_ASAP7_75t_L g1153 ( .A(n_1027), .Y(n_1153) );
AND2x4_ASAP7_75t_L g1154 ( .A(n_1058), .B(n_1067), .Y(n_1154) );
NAND2xp5_ASAP7_75t_L g1155 ( .A(n_1027), .B(n_1075), .Y(n_1155) );
INVx2_ASAP7_75t_L g1156 ( .A(n_1035), .Y(n_1156) );
OR2x2_ASAP7_75t_L g1157 ( .A(n_1069), .B(n_1066), .Y(n_1157) );
OAI221xp5_ASAP7_75t_L g1158 ( .A1(n_1103), .A2(n_1100), .B1(n_1034), .B2(n_1104), .C(n_1082), .Y(n_1158) );
INVx1_ASAP7_75t_L g1159 ( .A(n_1062), .Y(n_1159) );
AOI22xp33_ASAP7_75t_L g1160 ( .A1(n_1075), .A2(n_1104), .B1(n_1109), .B2(n_1100), .Y(n_1160) );
OR2x2_ASAP7_75t_L g1161 ( .A(n_1062), .B(n_1066), .Y(n_1161) );
NAND2xp5_ASAP7_75t_SL g1162 ( .A(n_1032), .B(n_1065), .Y(n_1162) );
AND2x2_ASAP7_75t_L g1163 ( .A(n_1028), .B(n_1033), .Y(n_1163) );
INVx1_ASAP7_75t_L g1164 ( .A(n_1070), .Y(n_1164) );
INVx2_ASAP7_75t_L g1165 ( .A(n_1074), .Y(n_1165) );
OAI31xp33_ASAP7_75t_L g1166 ( .A1(n_1078), .A2(n_1092), .A3(n_1083), .B(n_1057), .Y(n_1166) );
AND2x2_ASAP7_75t_L g1167 ( .A(n_1033), .B(n_1070), .Y(n_1167) );
NAND2xp5_ASAP7_75t_L g1168 ( .A(n_1078), .B(n_1083), .Y(n_1168) );
AND2x2_ASAP7_75t_L g1169 ( .A(n_1074), .B(n_1038), .Y(n_1169) );
NAND2xp5_ASAP7_75t_L g1170 ( .A(n_1038), .B(n_1084), .Y(n_1170) );
INVx1_ASAP7_75t_L g1171 ( .A(n_1057), .Y(n_1171) );
OR2x2_ASAP7_75t_L g1172 ( .A(n_1109), .B(n_1084), .Y(n_1172) );
NOR2xp33_ASAP7_75t_L g1173 ( .A(n_1061), .B(n_1105), .Y(n_1173) );
BUFx2_ASAP7_75t_L g1174 ( .A(n_1143), .Y(n_1174) );
AND2x2_ASAP7_75t_L g1175 ( .A(n_1134), .B(n_1088), .Y(n_1175) );
INVx1_ASAP7_75t_L g1176 ( .A(n_1112), .Y(n_1176) );
NAND2xp5_ASAP7_75t_L g1177 ( .A(n_1136), .B(n_1032), .Y(n_1177) );
AND2x2_ASAP7_75t_L g1178 ( .A(n_1134), .B(n_1088), .Y(n_1178) );
AND2x2_ASAP7_75t_L g1179 ( .A(n_1163), .B(n_1167), .Y(n_1179) );
NAND2xp5_ASAP7_75t_L g1180 ( .A(n_1148), .B(n_1032), .Y(n_1180) );
INVx1_ASAP7_75t_L g1181 ( .A(n_1129), .Y(n_1181) );
AND2x2_ASAP7_75t_L g1182 ( .A(n_1163), .B(n_1032), .Y(n_1182) );
AND2x2_ASAP7_75t_L g1183 ( .A(n_1167), .B(n_1032), .Y(n_1183) );
INVx1_ASAP7_75t_L g1184 ( .A(n_1114), .Y(n_1184) );
OR2x2_ASAP7_75t_L g1185 ( .A(n_1117), .B(n_1080), .Y(n_1185) );
INVx1_ASAP7_75t_L g1186 ( .A(n_1120), .Y(n_1186) );
INVx1_ASAP7_75t_L g1187 ( .A(n_1127), .Y(n_1187) );
OAI22xp5_ASAP7_75t_L g1188 ( .A1(n_1146), .A2(n_1040), .B1(n_1092), .B2(n_1054), .Y(n_1188) );
NAND2xp5_ASAP7_75t_L g1189 ( .A(n_1148), .B(n_1054), .Y(n_1189) );
NOR2xp33_ASAP7_75t_L g1190 ( .A(n_1140), .B(n_1105), .Y(n_1190) );
INVx1_ASAP7_75t_L g1191 ( .A(n_1127), .Y(n_1191) );
INVx1_ASAP7_75t_L g1192 ( .A(n_1161), .Y(n_1192) );
INVx1_ASAP7_75t_SL g1193 ( .A(n_1128), .Y(n_1193) );
INVx1_ASAP7_75t_L g1194 ( .A(n_1161), .Y(n_1194) );
NAND2xp5_ASAP7_75t_L g1195 ( .A(n_1116), .B(n_1054), .Y(n_1195) );
AND2x4_ASAP7_75t_L g1196 ( .A(n_1154), .B(n_1054), .Y(n_1196) );
AND2x2_ASAP7_75t_SL g1197 ( .A(n_1154), .B(n_1137), .Y(n_1197) );
NAND2xp5_ASAP7_75t_L g1198 ( .A(n_1116), .B(n_1092), .Y(n_1198) );
NOR3xp33_ASAP7_75t_L g1199 ( .A(n_1144), .B(n_1101), .C(n_1092), .Y(n_1199) );
INVx1_ASAP7_75t_L g1200 ( .A(n_1115), .Y(n_1200) );
NAND2xp5_ASAP7_75t_L g1201 ( .A(n_1123), .B(n_1105), .Y(n_1201) );
OR2x2_ASAP7_75t_L g1202 ( .A(n_1139), .B(n_1087), .Y(n_1202) );
NAND2xp5_ASAP7_75t_L g1203 ( .A(n_1123), .B(n_1055), .Y(n_1203) );
XNOR2x1_ASAP7_75t_L g1204 ( .A(n_1141), .B(n_1091), .Y(n_1204) );
INVx1_ASAP7_75t_L g1205 ( .A(n_1159), .Y(n_1205) );
AND2x2_ASAP7_75t_L g1206 ( .A(n_1133), .B(n_1055), .Y(n_1206) );
CKINVDCx16_ASAP7_75t_R g1207 ( .A(n_1143), .Y(n_1207) );
NAND3xp33_ASAP7_75t_L g1208 ( .A(n_1173), .B(n_1055), .C(n_1091), .Y(n_1208) );
NAND2xp5_ASAP7_75t_L g1209 ( .A(n_1147), .B(n_1055), .Y(n_1209) );
INVx1_ASAP7_75t_L g1210 ( .A(n_1130), .Y(n_1210) );
INVx1_ASAP7_75t_L g1211 ( .A(n_1135), .Y(n_1211) );
INVx2_ASAP7_75t_L g1212 ( .A(n_1113), .Y(n_1212) );
OAI33xp33_ASAP7_75t_L g1213 ( .A1(n_1132), .A2(n_1090), .A3(n_1168), .B1(n_1155), .B2(n_1171), .B3(n_1170), .Y(n_1213) );
NAND2x1_ASAP7_75t_L g1214 ( .A(n_1154), .B(n_1090), .Y(n_1214) );
NAND2x1p5_ASAP7_75t_L g1215 ( .A(n_1122), .B(n_1162), .Y(n_1215) );
OAI21xp33_ASAP7_75t_L g1216 ( .A1(n_1190), .A2(n_1124), .B(n_1173), .Y(n_1216) );
NAND2xp5_ASAP7_75t_L g1217 ( .A(n_1179), .B(n_1147), .Y(n_1217) );
NAND2xp5_ASAP7_75t_L g1218 ( .A(n_1179), .B(n_1164), .Y(n_1218) );
INVx2_ASAP7_75t_L g1219 ( .A(n_1212), .Y(n_1219) );
NOR2xp33_ASAP7_75t_L g1220 ( .A(n_1207), .B(n_1158), .Y(n_1220) );
INVx1_ASAP7_75t_SL g1221 ( .A(n_1193), .Y(n_1221) );
NOR3xp33_ASAP7_75t_L g1222 ( .A(n_1199), .B(n_1131), .C(n_1149), .Y(n_1222) );
INVx1_ASAP7_75t_L g1223 ( .A(n_1176), .Y(n_1223) );
NAND2xp5_ASAP7_75t_L g1224 ( .A(n_1200), .B(n_1153), .Y(n_1224) );
XNOR2x2_ASAP7_75t_L g1225 ( .A(n_1188), .B(n_1149), .Y(n_1225) );
INVx1_ASAP7_75t_L g1226 ( .A(n_1187), .Y(n_1226) );
NAND2xp5_ASAP7_75t_L g1227 ( .A(n_1187), .B(n_1150), .Y(n_1227) );
AND2x2_ASAP7_75t_L g1228 ( .A(n_1206), .B(n_1133), .Y(n_1228) );
NAND2xp5_ASAP7_75t_L g1229 ( .A(n_1191), .B(n_1151), .Y(n_1229) );
AOI21xp33_ASAP7_75t_SL g1230 ( .A1(n_1197), .A2(n_1142), .B(n_1119), .Y(n_1230) );
INVx1_ASAP7_75t_L g1231 ( .A(n_1191), .Y(n_1231) );
INVx1_ASAP7_75t_L g1232 ( .A(n_1192), .Y(n_1232) );
INVx1_ASAP7_75t_L g1233 ( .A(n_1176), .Y(n_1233) );
NOR2xp33_ASAP7_75t_L g1234 ( .A(n_1210), .B(n_1126), .Y(n_1234) );
INVx1_ASAP7_75t_SL g1235 ( .A(n_1174), .Y(n_1235) );
OR2x2_ASAP7_75t_L g1236 ( .A(n_1202), .B(n_1121), .Y(n_1236) );
INVx1_ASAP7_75t_L g1237 ( .A(n_1184), .Y(n_1237) );
INVx1_ASAP7_75t_L g1238 ( .A(n_1184), .Y(n_1238) );
AND2x2_ASAP7_75t_L g1239 ( .A(n_1206), .B(n_1169), .Y(n_1239) );
INVx1_ASAP7_75t_L g1240 ( .A(n_1192), .Y(n_1240) );
OAI221xp5_ASAP7_75t_L g1241 ( .A1(n_1204), .A2(n_1166), .B1(n_1160), .B2(n_1119), .C(n_1172), .Y(n_1241) );
CKINVDCx20_ASAP7_75t_R g1242 ( .A(n_1195), .Y(n_1242) );
NAND2xp5_ASAP7_75t_L g1243 ( .A(n_1194), .B(n_1160), .Y(n_1243) );
OR2x2_ASAP7_75t_L g1244 ( .A(n_1202), .B(n_1152), .Y(n_1244) );
INVx1_ASAP7_75t_SL g1245 ( .A(n_1196), .Y(n_1245) );
XNOR2x1_ASAP7_75t_L g1246 ( .A(n_1182), .B(n_1157), .Y(n_1246) );
OAI22xp5_ASAP7_75t_L g1247 ( .A1(n_1180), .A2(n_1145), .B1(n_1138), .B2(n_1125), .Y(n_1247) );
INVxp67_ASAP7_75t_L g1248 ( .A(n_1201), .Y(n_1248) );
NOR2x1_ASAP7_75t_L g1249 ( .A(n_1214), .B(n_1113), .Y(n_1249) );
NAND3xp33_ASAP7_75t_L g1250 ( .A(n_1208), .B(n_1165), .C(n_1125), .Y(n_1250) );
INVx8_ASAP7_75t_L g1251 ( .A(n_1196), .Y(n_1251) );
AND2x2_ASAP7_75t_L g1252 ( .A(n_1182), .B(n_1183), .Y(n_1252) );
AND2x2_ASAP7_75t_L g1253 ( .A(n_1175), .B(n_1165), .Y(n_1253) );
INVxp67_ASAP7_75t_SL g1254 ( .A(n_1215), .Y(n_1254) );
INVx1_ASAP7_75t_L g1255 ( .A(n_1186), .Y(n_1255) );
BUFx2_ASAP7_75t_L g1256 ( .A(n_1196), .Y(n_1256) );
OAI22xp5_ASAP7_75t_L g1257 ( .A1(n_1215), .A2(n_1118), .B1(n_1156), .B2(n_1198), .Y(n_1257) );
INVxp67_ASAP7_75t_L g1258 ( .A(n_1185), .Y(n_1258) );
INVx2_ASAP7_75t_L g1259 ( .A(n_1212), .Y(n_1259) );
INVx1_ASAP7_75t_L g1260 ( .A(n_1236), .Y(n_1260) );
OAI211xp5_ASAP7_75t_L g1261 ( .A1(n_1230), .A2(n_1216), .B(n_1222), .C(n_1220), .Y(n_1261) );
AOI21xp33_ASAP7_75t_L g1262 ( .A1(n_1241), .A2(n_1221), .B(n_1254), .Y(n_1262) );
INVx1_ASAP7_75t_L g1263 ( .A(n_1236), .Y(n_1263) );
NAND2xp5_ASAP7_75t_L g1264 ( .A(n_1248), .B(n_1243), .Y(n_1264) );
OAI211xp5_ASAP7_75t_L g1265 ( .A1(n_1251), .A2(n_1225), .B(n_1214), .C(n_1235), .Y(n_1265) );
AOI22xp33_ASAP7_75t_L g1266 ( .A1(n_1225), .A2(n_1213), .B1(n_1177), .B2(n_1234), .Y(n_1266) );
NOR3xp33_ASAP7_75t_L g1267 ( .A(n_1257), .B(n_1250), .C(n_1247), .Y(n_1267) );
NAND4xp25_ASAP7_75t_L g1268 ( .A(n_1209), .B(n_1256), .C(n_1249), .D(n_1245), .Y(n_1268) );
INVx1_ASAP7_75t_SL g1269 ( .A(n_1244), .Y(n_1269) );
AOI221xp5_ASAP7_75t_L g1270 ( .A1(n_1261), .A2(n_1258), .B1(n_1224), .B2(n_1240), .C(n_1231), .Y(n_1270) );
OAI221xp5_ASAP7_75t_L g1271 ( .A1(n_1265), .A2(n_1258), .B1(n_1246), .B2(n_1215), .C(n_1217), .Y(n_1271) );
AOI22x1_ASAP7_75t_L g1272 ( .A1(n_1269), .A2(n_1252), .B1(n_1239), .B2(n_1228), .Y(n_1272) );
NAND3x1_ASAP7_75t_L g1273 ( .A(n_1267), .B(n_1218), .C(n_1251), .Y(n_1273) );
AND2x2_ASAP7_75t_L g1274 ( .A(n_1260), .B(n_1228), .Y(n_1274) );
AOI22xp5_ASAP7_75t_L g1275 ( .A1(n_1262), .A2(n_1242), .B1(n_1226), .B2(n_1232), .Y(n_1275) );
NAND4xp25_ASAP7_75t_L g1276 ( .A(n_1266), .B(n_1203), .C(n_1189), .D(n_1227), .Y(n_1276) );
AOI22xp33_ASAP7_75t_L g1277 ( .A1(n_1271), .A2(n_1268), .B1(n_1266), .B2(n_1264), .Y(n_1277) );
INVxp67_ASAP7_75t_SL g1278 ( .A(n_1272), .Y(n_1278) );
INVx1_ASAP7_75t_L g1279 ( .A(n_1274), .Y(n_1279) );
NAND3xp33_ASAP7_75t_SL g1280 ( .A(n_1270), .B(n_1242), .C(n_1263), .Y(n_1280) );
INVx1_ASAP7_75t_L g1281 ( .A(n_1275), .Y(n_1281) );
AOI322xp5_ASAP7_75t_L g1282 ( .A1(n_1278), .A2(n_1276), .A3(n_1273), .B1(n_1239), .B2(n_1253), .C1(n_1229), .C2(n_1175), .Y(n_1282) );
AOI22xp5_ASAP7_75t_L g1283 ( .A1(n_1280), .A2(n_1255), .B1(n_1181), .B2(n_1233), .Y(n_1283) );
OR3x1_ASAP7_75t_L g1284 ( .A(n_1281), .B(n_1223), .C(n_1238), .Y(n_1284) );
INVx2_ASAP7_75t_SL g1285 ( .A(n_1283), .Y(n_1285) );
INVx1_ASAP7_75t_L g1286 ( .A(n_1284), .Y(n_1286) );
AOI22xp5_ASAP7_75t_L g1287 ( .A1(n_1286), .A2(n_1277), .B1(n_1279), .B2(n_1282), .Y(n_1287) );
AOI221xp5_ASAP7_75t_L g1288 ( .A1(n_1285), .A2(n_1237), .B1(n_1233), .B2(n_1205), .C(n_1211), .Y(n_1288) );
BUFx2_ASAP7_75t_L g1289 ( .A(n_1287), .Y(n_1289) );
OR2x2_ASAP7_75t_L g1290 ( .A(n_1288), .B(n_1237), .Y(n_1290) );
AOI221xp5_ASAP7_75t_L g1291 ( .A1(n_1289), .A2(n_1205), .B1(n_1211), .B2(n_1259), .C(n_1219), .Y(n_1291) );
AOI21xp5_ASAP7_75t_L g1292 ( .A1(n_1291), .A2(n_1290), .B(n_1178), .Y(n_1292) );
endmodule