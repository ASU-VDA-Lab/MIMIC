module real_aes_6184_n_100 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_100);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_100;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_693;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_649;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_725;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_552;
wire n_602;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_749;
wire n_358;
wire n_275;
wire n_214;
wire n_385;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_637;
wire n_526;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_101;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_741;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_717;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_639;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g555 ( .A1(n_0), .A2(n_162), .B(n_556), .C(n_559), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_1), .B(n_500), .Y(n_560) );
INVx1_ASAP7_75t_L g109 ( .A(n_2), .Y(n_109) );
INVx1_ASAP7_75t_L g196 ( .A(n_3), .Y(n_196) );
NAND2xp5_ASAP7_75t_SL g534 ( .A(n_4), .B(n_154), .Y(n_534) );
AOI21xp5_ASAP7_75t_L g493 ( .A1(n_5), .A2(n_469), .B(n_494), .Y(n_493) );
AO21x2_ASAP7_75t_L g484 ( .A1(n_6), .A2(n_139), .B(n_485), .Y(n_484) );
AOI22xp33_ASAP7_75t_L g225 ( .A1(n_7), .A2(n_35), .B1(n_148), .B2(n_226), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_8), .B(n_139), .Y(n_165) );
AND2x6_ASAP7_75t_L g163 ( .A(n_9), .B(n_164), .Y(n_163) );
A2O1A1Ixp33_ASAP7_75t_L g458 ( .A1(n_10), .A2(n_163), .B(n_459), .C(n_461), .Y(n_458) );
INVx1_ASAP7_75t_L g106 ( .A(n_11), .Y(n_106) );
NOR2xp33_ASAP7_75t_L g125 ( .A(n_11), .B(n_36), .Y(n_125) );
INVx1_ASAP7_75t_L g144 ( .A(n_12), .Y(n_144) );
INVx1_ASAP7_75t_L g189 ( .A(n_13), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_14), .B(n_152), .Y(n_232) );
NAND2xp5_ASAP7_75t_SL g490 ( .A(n_15), .B(n_154), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_16), .B(n_140), .Y(n_201) );
AO32x2_ASAP7_75t_L g223 ( .A1(n_17), .A2(n_139), .A3(n_169), .B1(n_180), .B2(n_224), .Y(n_223) );
NAND2xp5_ASAP7_75t_SL g236 ( .A(n_18), .B(n_148), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_19), .B(n_140), .Y(n_198) );
AOI22xp33_ASAP7_75t_L g227 ( .A1(n_20), .A2(n_52), .B1(n_148), .B2(n_226), .Y(n_227) );
AOI22xp33_ASAP7_75t_SL g248 ( .A1(n_21), .A2(n_80), .B1(n_148), .B2(n_152), .Y(n_248) );
NAND2xp5_ASAP7_75t_SL g218 ( .A(n_22), .B(n_148), .Y(n_218) );
A2O1A1Ixp33_ASAP7_75t_L g519 ( .A1(n_23), .A2(n_180), .B(n_459), .C(n_520), .Y(n_519) );
A2O1A1Ixp33_ASAP7_75t_L g487 ( .A1(n_24), .A2(n_180), .B(n_459), .C(n_488), .Y(n_487) );
BUFx6f_ASAP7_75t_L g156 ( .A(n_25), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_26), .B(n_182), .Y(n_181) );
CKINVDCx20_ASAP7_75t_R g126 ( .A(n_27), .Y(n_126) );
AOI21xp5_ASAP7_75t_L g552 ( .A1(n_28), .A2(n_469), .B(n_553), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_29), .B(n_182), .Y(n_220) );
INVx2_ASAP7_75t_L g150 ( .A(n_30), .Y(n_150) );
A2O1A1Ixp33_ASAP7_75t_L g507 ( .A1(n_31), .A2(n_471), .B(n_479), .C(n_508), .Y(n_507) );
NAND2xp5_ASAP7_75t_SL g172 ( .A(n_32), .B(n_148), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_33), .B(n_182), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_34), .B(n_234), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g105 ( .A(n_36), .B(n_106), .Y(n_105) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_37), .B(n_518), .Y(n_517) );
CKINVDCx20_ASAP7_75t_R g465 ( .A(n_38), .Y(n_465) );
AOI222xp33_ASAP7_75t_SL g127 ( .A1(n_39), .A2(n_78), .B1(n_128), .B2(n_733), .C1(n_734), .C2(n_738), .Y(n_127) );
CKINVDCx16_ASAP7_75t_R g733 ( .A(n_39), .Y(n_733) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_40), .B(n_154), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_41), .B(n_469), .Y(n_486) );
OAI22xp5_ASAP7_75t_SL g748 ( .A1(n_42), .A2(n_77), .B1(n_442), .B2(n_749), .Y(n_748) );
CKINVDCx20_ASAP7_75t_R g749 ( .A(n_42), .Y(n_749) );
A2O1A1Ixp33_ASAP7_75t_L g470 ( .A1(n_43), .A2(n_471), .B(n_473), .C(n_479), .Y(n_470) );
NAND2xp5_ASAP7_75t_SL g147 ( .A(n_44), .B(n_148), .Y(n_147) );
INVx1_ASAP7_75t_L g557 ( .A(n_45), .Y(n_557) );
AOI22xp33_ASAP7_75t_L g246 ( .A1(n_46), .A2(n_89), .B1(n_226), .B2(n_247), .Y(n_246) );
INVx1_ASAP7_75t_L g474 ( .A(n_47), .Y(n_474) );
NAND2xp5_ASAP7_75t_SL g158 ( .A(n_48), .B(n_148), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_49), .B(n_148), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_50), .B(n_469), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_51), .B(n_160), .Y(n_159) );
AOI22xp33_ASAP7_75t_SL g205 ( .A1(n_53), .A2(n_58), .B1(n_148), .B2(n_152), .Y(n_205) );
CKINVDCx20_ASAP7_75t_R g525 ( .A(n_54), .Y(n_525) );
NAND2xp5_ASAP7_75t_SL g177 ( .A(n_55), .B(n_148), .Y(n_177) );
NAND2xp5_ASAP7_75t_SL g231 ( .A(n_56), .B(n_148), .Y(n_231) );
AOI22xp33_ASAP7_75t_L g100 ( .A1(n_57), .A2(n_101), .B1(n_114), .B2(n_752), .Y(n_100) );
INVx1_ASAP7_75t_L g164 ( .A(n_59), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_60), .B(n_469), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_61), .B(n_500), .Y(n_499) );
A2O1A1Ixp33_ASAP7_75t_L g496 ( .A1(n_62), .A2(n_160), .B(n_192), .C(n_497), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_63), .B(n_148), .Y(n_197) );
INVx1_ASAP7_75t_L g143 ( .A(n_64), .Y(n_143) );
CKINVDCx20_ASAP7_75t_R g119 ( .A(n_65), .Y(n_119) );
NAND2xp5_ASAP7_75t_SL g510 ( .A(n_66), .B(n_154), .Y(n_510) );
AO32x2_ASAP7_75t_L g244 ( .A1(n_67), .A2(n_139), .A3(n_180), .B1(n_245), .B2(n_249), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_68), .B(n_155), .Y(n_462) );
INVx1_ASAP7_75t_L g175 ( .A(n_69), .Y(n_175) );
INVx1_ASAP7_75t_L g215 ( .A(n_70), .Y(n_215) );
CKINVDCx16_ASAP7_75t_R g554 ( .A(n_71), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_72), .B(n_476), .Y(n_521) );
A2O1A1Ixp33_ASAP7_75t_L g531 ( .A1(n_73), .A2(n_459), .B(n_479), .C(n_532), .Y(n_531) );
NAND2xp5_ASAP7_75t_SL g216 ( .A(n_74), .B(n_152), .Y(n_216) );
CKINVDCx16_ASAP7_75t_R g495 ( .A(n_75), .Y(n_495) );
INVx1_ASAP7_75t_L g113 ( .A(n_76), .Y(n_113) );
OAI22xp5_ASAP7_75t_SL g130 ( .A1(n_77), .A2(n_131), .B1(n_441), .B2(n_442), .Y(n_130) );
CKINVDCx20_ASAP7_75t_R g442 ( .A(n_77), .Y(n_442) );
NAND2xp5_ASAP7_75t_SL g522 ( .A(n_79), .B(n_475), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_81), .B(n_226), .Y(n_237) );
CKINVDCx20_ASAP7_75t_R g512 ( .A(n_82), .Y(n_512) );
NAND2xp5_ASAP7_75t_SL g219 ( .A(n_83), .B(n_152), .Y(n_219) );
INVx2_ASAP7_75t_L g141 ( .A(n_84), .Y(n_141) );
CKINVDCx20_ASAP7_75t_R g538 ( .A(n_85), .Y(n_538) );
NAND2xp5_ASAP7_75t_SL g463 ( .A(n_86), .B(n_179), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_87), .B(n_152), .Y(n_151) );
INVx2_ASAP7_75t_L g110 ( .A(n_88), .Y(n_110) );
OR2x2_ASAP7_75t_L g122 ( .A(n_88), .B(n_123), .Y(n_122) );
OR2x2_ASAP7_75t_L g445 ( .A(n_88), .B(n_124), .Y(n_445) );
AOI22xp33_ASAP7_75t_L g204 ( .A1(n_90), .A2(n_99), .B1(n_152), .B2(n_153), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_91), .B(n_469), .Y(n_506) );
INVx1_ASAP7_75t_L g509 ( .A(n_92), .Y(n_509) );
INVxp67_ASAP7_75t_L g498 ( .A(n_93), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_94), .B(n_152), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_95), .B(n_113), .Y(n_112) );
INVx1_ASAP7_75t_L g455 ( .A(n_96), .Y(n_455) );
INVx1_ASAP7_75t_L g533 ( .A(n_97), .Y(n_533) );
AND2x2_ASAP7_75t_L g481 ( .A(n_98), .B(n_182), .Y(n_481) );
INVx1_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
INVx2_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
INVx3_ASAP7_75t_SL g752 ( .A(n_103), .Y(n_752) );
AND2x2_ASAP7_75t_L g103 ( .A(n_104), .B(n_107), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
CKINVDCx14_ASAP7_75t_R g107 ( .A(n_108), .Y(n_107) );
NAND3xp33_ASAP7_75t_SL g108 ( .A(n_109), .B(n_110), .C(n_111), .Y(n_108) );
AND2x2_ASAP7_75t_L g124 ( .A(n_109), .B(n_125), .Y(n_124) );
OR2x2_ASAP7_75t_L g732 ( .A(n_110), .B(n_124), .Y(n_732) );
NOR2x2_ASAP7_75t_L g740 ( .A(n_110), .B(n_123), .Y(n_740) );
INVx1_ASAP7_75t_SL g111 ( .A(n_112), .Y(n_111) );
AOI22x1_ASAP7_75t_L g114 ( .A1(n_115), .A2(n_127), .B1(n_741), .B2(n_742), .Y(n_114) );
NOR2xp33_ASAP7_75t_L g115 ( .A(n_116), .B(n_120), .Y(n_115) );
INVx1_ASAP7_75t_SL g116 ( .A(n_117), .Y(n_116) );
BUFx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
INVx2_ASAP7_75t_SL g741 ( .A(n_118), .Y(n_741) );
INVx2_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
AOI21xp5_ASAP7_75t_L g742 ( .A1(n_120), .A2(n_743), .B(n_750), .Y(n_742) );
NOR2xp33_ASAP7_75t_SL g120 ( .A(n_121), .B(n_126), .Y(n_120) );
HB1xp67_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
INVx1_ASAP7_75t_SL g751 ( .A(n_122), .Y(n_751) );
INVx2_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
OAI22xp5_ASAP7_75t_SL g128 ( .A1(n_129), .A2(n_443), .B1(n_446), .B2(n_730), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
OAI22xp5_ASAP7_75t_SL g734 ( .A1(n_130), .A2(n_735), .B1(n_736), .B2(n_737), .Y(n_734) );
INVx2_ASAP7_75t_L g441 ( .A(n_131), .Y(n_441) );
OAI22xp5_ASAP7_75t_L g746 ( .A1(n_131), .A2(n_441), .B1(n_747), .B2(n_748), .Y(n_746) );
NAND2x1p5_ASAP7_75t_L g131 ( .A(n_132), .B(n_365), .Y(n_131) );
AND2x2_ASAP7_75t_SL g132 ( .A(n_133), .B(n_323), .Y(n_132) );
NOR4xp25_ASAP7_75t_L g133 ( .A(n_134), .B(n_263), .C(n_299), .D(n_313), .Y(n_133) );
OAI221xp5_ASAP7_75t_SL g134 ( .A1(n_135), .A2(n_207), .B1(n_239), .B2(n_250), .C(n_254), .Y(n_134) );
NAND2xp5_ASAP7_75t_SL g397 ( .A(n_135), .B(n_398), .Y(n_397) );
OR2x2_ASAP7_75t_L g135 ( .A(n_136), .B(n_183), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
AND2x2_ASAP7_75t_L g137 ( .A(n_138), .B(n_166), .Y(n_137) );
AND2x2_ASAP7_75t_L g260 ( .A(n_138), .B(n_167), .Y(n_260) );
INVx3_ASAP7_75t_L g268 ( .A(n_138), .Y(n_268) );
AND2x2_ASAP7_75t_L g322 ( .A(n_138), .B(n_186), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_138), .B(n_185), .Y(n_358) );
AND2x2_ASAP7_75t_L g416 ( .A(n_138), .B(n_278), .Y(n_416) );
OA21x2_ASAP7_75t_L g138 ( .A1(n_139), .A2(n_145), .B(n_165), .Y(n_138) );
INVx4_ASAP7_75t_L g206 ( .A(n_139), .Y(n_206) );
AOI21xp5_ASAP7_75t_L g485 ( .A1(n_139), .A2(n_486), .B(n_487), .Y(n_485) );
HB1xp67_ASAP7_75t_L g492 ( .A(n_139), .Y(n_492) );
BUFx6f_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
INVx1_ASAP7_75t_L g169 ( .A(n_140), .Y(n_169) );
AND2x2_ASAP7_75t_L g140 ( .A(n_141), .B(n_142), .Y(n_140) );
AND2x2_ASAP7_75t_SL g182 ( .A(n_141), .B(n_142), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_143), .B(n_144), .Y(n_142) );
OAI21xp5_ASAP7_75t_L g145 ( .A1(n_146), .A2(n_157), .B(n_163), .Y(n_145) );
AOI21xp5_ASAP7_75t_L g146 ( .A1(n_147), .A2(n_151), .B(n_154), .Y(n_146) );
INVx3_ASAP7_75t_L g214 ( .A(n_148), .Y(n_214) );
HB1xp67_ASAP7_75t_L g535 ( .A(n_148), .Y(n_535) );
BUFx6f_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx1_ASAP7_75t_L g226 ( .A(n_149), .Y(n_226) );
BUFx3_ASAP7_75t_L g247 ( .A(n_149), .Y(n_247) );
AND2x6_ASAP7_75t_L g459 ( .A(n_149), .B(n_460), .Y(n_459) );
INVx2_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx1_ASAP7_75t_L g153 ( .A(n_150), .Y(n_153) );
INVx1_ASAP7_75t_L g161 ( .A(n_150), .Y(n_161) );
INVx2_ASAP7_75t_L g190 ( .A(n_152), .Y(n_190) );
INVx3_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx2_ASAP7_75t_L g162 ( .A(n_154), .Y(n_162) );
AOI21xp5_ASAP7_75t_L g171 ( .A1(n_154), .A2(n_172), .B(n_173), .Y(n_171) );
O2A1O1Ixp5_ASAP7_75t_SL g213 ( .A1(n_154), .A2(n_214), .B(n_215), .C(n_216), .Y(n_213) );
NOR2xp33_ASAP7_75t_L g497 ( .A(n_154), .B(n_498), .Y(n_497) );
INVx5_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
OAI22xp5_ASAP7_75t_SL g245 ( .A1(n_155), .A2(n_179), .B1(n_246), .B2(n_248), .Y(n_245) );
INVx3_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
BUFx6f_ASAP7_75t_L g179 ( .A(n_156), .Y(n_179) );
BUFx6f_ASAP7_75t_L g194 ( .A(n_156), .Y(n_194) );
INVx1_ASAP7_75t_L g234 ( .A(n_156), .Y(n_234) );
AND2x2_ASAP7_75t_L g457 ( .A(n_156), .B(n_161), .Y(n_457) );
INVx1_ASAP7_75t_L g460 ( .A(n_156), .Y(n_460) );
AOI21xp5_ASAP7_75t_L g157 ( .A1(n_158), .A2(n_159), .B(n_162), .Y(n_157) );
INVx2_ASAP7_75t_L g176 ( .A(n_160), .Y(n_176) );
INVx1_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
O2A1O1Ixp33_ASAP7_75t_L g195 ( .A1(n_162), .A2(n_176), .B(n_196), .C(n_197), .Y(n_195) );
OAI22xp5_ASAP7_75t_L g203 ( .A1(n_162), .A2(n_179), .B1(n_204), .B2(n_205), .Y(n_203) );
OAI22xp5_ASAP7_75t_L g224 ( .A1(n_162), .A2(n_179), .B1(n_225), .B2(n_227), .Y(n_224) );
BUFx3_ASAP7_75t_L g180 ( .A(n_163), .Y(n_180) );
OAI21xp5_ASAP7_75t_L g187 ( .A1(n_163), .A2(n_188), .B(n_195), .Y(n_187) );
OAI21xp5_ASAP7_75t_L g212 ( .A1(n_163), .A2(n_213), .B(n_217), .Y(n_212) );
OAI21xp5_ASAP7_75t_L g229 ( .A1(n_163), .A2(n_230), .B(n_235), .Y(n_229) );
NAND2x1p5_ASAP7_75t_L g456 ( .A(n_163), .B(n_457), .Y(n_456) );
AND2x4_ASAP7_75t_L g469 ( .A(n_163), .B(n_457), .Y(n_469) );
INVx4_ASAP7_75t_SL g480 ( .A(n_163), .Y(n_480) );
AND2x2_ASAP7_75t_L g251 ( .A(n_166), .B(n_252), .Y(n_251) );
AND2x2_ASAP7_75t_L g265 ( .A(n_166), .B(n_186), .Y(n_265) );
INVx2_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_167), .B(n_186), .Y(n_280) );
AND2x2_ASAP7_75t_L g292 ( .A(n_167), .B(n_268), .Y(n_292) );
OR2x2_ASAP7_75t_L g294 ( .A(n_167), .B(n_252), .Y(n_294) );
AND2x2_ASAP7_75t_L g329 ( .A(n_167), .B(n_252), .Y(n_329) );
HB1xp67_ASAP7_75t_L g374 ( .A(n_167), .Y(n_374) );
INVx1_ASAP7_75t_L g382 ( .A(n_167), .Y(n_382) );
OA21x2_ASAP7_75t_L g167 ( .A1(n_168), .A2(n_170), .B(n_181), .Y(n_167) );
OA21x2_ASAP7_75t_L g186 ( .A1(n_168), .A2(n_187), .B(n_198), .Y(n_186) );
INVx2_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
NOR2xp33_ASAP7_75t_L g464 ( .A(n_169), .B(n_465), .Y(n_464) );
OAI21xp5_ASAP7_75t_L g170 ( .A1(n_171), .A2(n_174), .B(n_180), .Y(n_170) );
O2A1O1Ixp5_ASAP7_75t_L g174 ( .A1(n_175), .A2(n_176), .B(n_177), .C(n_178), .Y(n_174) );
AOI21xp5_ASAP7_75t_L g520 ( .A1(n_176), .A2(n_521), .B(n_522), .Y(n_520) );
AOI21xp5_ASAP7_75t_L g235 ( .A1(n_178), .A2(n_236), .B(n_237), .Y(n_235) );
INVx2_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
INVx4_ASAP7_75t_L g558 ( .A(n_179), .Y(n_558) );
NAND3xp33_ASAP7_75t_L g202 ( .A(n_180), .B(n_203), .C(n_206), .Y(n_202) );
OA21x2_ASAP7_75t_L g211 ( .A1(n_182), .A2(n_212), .B(n_220), .Y(n_211) );
OA21x2_ASAP7_75t_L g228 ( .A1(n_182), .A2(n_229), .B(n_238), .Y(n_228) );
INVx2_ASAP7_75t_L g249 ( .A(n_182), .Y(n_249) );
AOI21xp5_ASAP7_75t_L g467 ( .A1(n_182), .A2(n_468), .B(n_470), .Y(n_467) );
AOI21xp5_ASAP7_75t_L g505 ( .A1(n_182), .A2(n_506), .B(n_507), .Y(n_505) );
INVx1_ASAP7_75t_L g526 ( .A(n_182), .Y(n_526) );
OAI221xp5_ASAP7_75t_L g299 ( .A1(n_183), .A2(n_300), .B1(n_304), .B2(n_308), .C(n_309), .Y(n_299) );
INVx1_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
AND2x2_ASAP7_75t_L g259 ( .A(n_184), .B(n_260), .Y(n_259) );
AND2x2_ASAP7_75t_L g184 ( .A(n_185), .B(n_199), .Y(n_184) );
INVx2_ASAP7_75t_L g258 ( .A(n_185), .Y(n_258) );
AND2x2_ASAP7_75t_L g311 ( .A(n_185), .B(n_312), .Y(n_311) );
AND2x2_ASAP7_75t_L g330 ( .A(n_185), .B(n_268), .Y(n_330) );
INVx2_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
AND2x2_ASAP7_75t_L g393 ( .A(n_186), .B(n_268), .Y(n_393) );
O2A1O1Ixp33_ASAP7_75t_L g188 ( .A1(n_189), .A2(n_190), .B(n_191), .C(n_192), .Y(n_188) );
AOI21xp5_ASAP7_75t_L g461 ( .A1(n_190), .A2(n_462), .B(n_463), .Y(n_461) );
AOI21xp5_ASAP7_75t_L g488 ( .A1(n_190), .A2(n_489), .B(n_490), .Y(n_488) );
O2A1O1Ixp33_ASAP7_75t_L g532 ( .A1(n_192), .A2(n_533), .B(n_534), .C(n_535), .Y(n_532) );
INVx1_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
AOI21xp5_ASAP7_75t_L g217 ( .A1(n_193), .A2(n_218), .B(n_219), .Y(n_217) );
INVx4_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
INVx2_ASAP7_75t_L g476 ( .A(n_194), .Y(n_476) );
AND2x2_ASAP7_75t_L g315 ( .A(n_199), .B(n_260), .Y(n_315) );
OAI322xp33_ASAP7_75t_L g383 ( .A1(n_199), .A2(n_339), .A3(n_384), .B1(n_386), .B2(n_389), .C1(n_391), .C2(n_395), .Y(n_383) );
INVx3_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
NOR2x1_ASAP7_75t_L g266 ( .A(n_200), .B(n_267), .Y(n_266) );
INVx2_ASAP7_75t_L g279 ( .A(n_200), .Y(n_279) );
AND2x2_ASAP7_75t_L g388 ( .A(n_200), .B(n_268), .Y(n_388) );
AND2x2_ASAP7_75t_L g420 ( .A(n_200), .B(n_292), .Y(n_420) );
OR2x2_ASAP7_75t_L g423 ( .A(n_200), .B(n_424), .Y(n_423) );
AND2x4_ASAP7_75t_L g200 ( .A(n_201), .B(n_202), .Y(n_200) );
INVx1_ASAP7_75t_L g253 ( .A(n_201), .Y(n_253) );
AO21x1_ASAP7_75t_L g252 ( .A1(n_203), .A2(n_206), .B(n_253), .Y(n_252) );
AO21x2_ASAP7_75t_L g453 ( .A1(n_206), .A2(n_454), .B(n_464), .Y(n_453) );
INVx3_ASAP7_75t_L g500 ( .A(n_206), .Y(n_500) );
NOR2xp33_ASAP7_75t_L g511 ( .A(n_206), .B(n_512), .Y(n_511) );
AO21x2_ASAP7_75t_L g529 ( .A1(n_206), .A2(n_530), .B(n_537), .Y(n_529) );
NOR2xp33_ASAP7_75t_L g537 ( .A(n_206), .B(n_538), .Y(n_537) );
INVx1_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
AND2x2_ASAP7_75t_L g208 ( .A(n_209), .B(n_221), .Y(n_208) );
INVx1_ASAP7_75t_L g436 ( .A(n_209), .Y(n_436) );
INVx1_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
OR2x2_ASAP7_75t_L g241 ( .A(n_210), .B(n_228), .Y(n_241) );
INVx2_ASAP7_75t_L g276 ( .A(n_210), .Y(n_276) );
INVx2_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
INVx2_ASAP7_75t_L g298 ( .A(n_211), .Y(n_298) );
HB1xp67_ASAP7_75t_L g306 ( .A(n_211), .Y(n_306) );
OR2x2_ASAP7_75t_L g430 ( .A(n_211), .B(n_431), .Y(n_430) );
AND2x2_ASAP7_75t_L g255 ( .A(n_221), .B(n_256), .Y(n_255) );
AND2x2_ASAP7_75t_L g295 ( .A(n_221), .B(n_296), .Y(n_295) );
AND2x2_ASAP7_75t_L g347 ( .A(n_221), .B(n_348), .Y(n_347) );
AND2x2_ASAP7_75t_L g221 ( .A(n_222), .B(n_228), .Y(n_221) );
AND2x2_ASAP7_75t_L g242 ( .A(n_222), .B(n_243), .Y(n_242) );
NOR2xp67_ASAP7_75t_L g302 ( .A(n_222), .B(n_303), .Y(n_302) );
AND2x2_ASAP7_75t_L g356 ( .A(n_222), .B(n_244), .Y(n_356) );
OR2x2_ASAP7_75t_L g364 ( .A(n_222), .B(n_298), .Y(n_364) );
INVx2_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
BUFx2_ASAP7_75t_L g273 ( .A(n_223), .Y(n_273) );
AND2x2_ASAP7_75t_L g283 ( .A(n_223), .B(n_284), .Y(n_283) );
AND2x2_ASAP7_75t_L g307 ( .A(n_223), .B(n_228), .Y(n_307) );
AND2x2_ASAP7_75t_L g371 ( .A(n_223), .B(n_244), .Y(n_371) );
NOR2xp33_ASAP7_75t_L g261 ( .A(n_228), .B(n_262), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_228), .B(n_276), .Y(n_275) );
INVx2_ASAP7_75t_L g284 ( .A(n_228), .Y(n_284) );
INVx1_ASAP7_75t_L g289 ( .A(n_228), .Y(n_289) );
AND2x2_ASAP7_75t_L g301 ( .A(n_228), .B(n_302), .Y(n_301) );
HB1xp67_ASAP7_75t_L g379 ( .A(n_228), .Y(n_379) );
INVx1_ASAP7_75t_L g431 ( .A(n_228), .Y(n_431) );
AOI21xp5_ASAP7_75t_L g230 ( .A1(n_231), .A2(n_232), .B(n_233), .Y(n_230) );
INVx1_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_240), .B(n_242), .Y(n_239) );
AND2x2_ASAP7_75t_L g408 ( .A(n_240), .B(n_317), .Y(n_408) );
INVx2_ASAP7_75t_SL g240 ( .A(n_241), .Y(n_240) );
AND2x2_ASAP7_75t_L g335 ( .A(n_242), .B(n_336), .Y(n_335) );
AND2x2_ASAP7_75t_L g434 ( .A(n_242), .B(n_369), .Y(n_434) );
INVx1_ASAP7_75t_L g256 ( .A(n_243), .Y(n_256) );
AND2x2_ASAP7_75t_L g282 ( .A(n_243), .B(n_276), .Y(n_282) );
BUFx2_ASAP7_75t_L g341 ( .A(n_243), .Y(n_341) );
INVx1_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
BUFx6f_ASAP7_75t_L g262 ( .A(n_244), .Y(n_262) );
INVx1_ASAP7_75t_L g272 ( .A(n_244), .Y(n_272) );
HB1xp67_ASAP7_75t_L g478 ( .A(n_247), .Y(n_478) );
INVx2_ASAP7_75t_L g559 ( .A(n_247), .Y(n_559) );
INVx1_ASAP7_75t_L g523 ( .A(n_249), .Y(n_523) );
NOR2xp67_ASAP7_75t_L g410 ( .A(n_250), .B(n_257), .Y(n_410) );
INVx2_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
AOI32xp33_ASAP7_75t_L g254 ( .A1(n_251), .A2(n_255), .A3(n_257), .B1(n_259), .B2(n_261), .Y(n_254) );
AND2x2_ASAP7_75t_L g394 ( .A(n_251), .B(n_267), .Y(n_394) );
AND2x2_ASAP7_75t_L g432 ( .A(n_251), .B(n_330), .Y(n_432) );
INVx1_ASAP7_75t_L g312 ( .A(n_252), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_256), .B(n_318), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_257), .B(n_292), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_257), .B(n_260), .Y(n_308) );
NAND2xp5_ASAP7_75t_SL g411 ( .A(n_257), .B(n_329), .Y(n_411) );
OR2x2_ASAP7_75t_L g425 ( .A(n_257), .B(n_294), .Y(n_425) );
INVx3_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
AND2x2_ASAP7_75t_L g352 ( .A(n_258), .B(n_260), .Y(n_352) );
OR2x2_ASAP7_75t_L g361 ( .A(n_258), .B(n_348), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_260), .B(n_311), .Y(n_333) );
INVx2_ASAP7_75t_L g348 ( .A(n_262), .Y(n_348) );
OR2x2_ASAP7_75t_L g363 ( .A(n_262), .B(n_364), .Y(n_363) );
AND2x2_ASAP7_75t_L g378 ( .A(n_262), .B(n_379), .Y(n_378) );
A2O1A1Ixp33_ASAP7_75t_L g435 ( .A1(n_262), .A2(n_355), .B(n_436), .C(n_437), .Y(n_435) );
OAI321xp33_ASAP7_75t_L g263 ( .A1(n_264), .A2(n_269), .A3(n_274), .B1(n_277), .B2(n_281), .C(n_285), .Y(n_263) );
INVx1_ASAP7_75t_L g376 ( .A(n_264), .Y(n_376) );
NAND2x1p5_ASAP7_75t_L g264 ( .A(n_265), .B(n_266), .Y(n_264) );
AND2x2_ASAP7_75t_L g387 ( .A(n_265), .B(n_388), .Y(n_387) );
INVx1_ASAP7_75t_L g339 ( .A(n_267), .Y(n_339) );
INVx2_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_268), .B(n_382), .Y(n_399) );
OAI221xp5_ASAP7_75t_L g406 ( .A1(n_269), .A2(n_407), .B1(n_409), .B2(n_411), .C(n_412), .Y(n_406) );
INVx1_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
AND2x2_ASAP7_75t_L g270 ( .A(n_271), .B(n_273), .Y(n_270) );
AND2x2_ASAP7_75t_L g344 ( .A(n_271), .B(n_318), .Y(n_344) );
HB1xp67_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_272), .B(n_298), .Y(n_297) );
INVx2_ASAP7_75t_L g317 ( .A(n_273), .Y(n_317) );
A2O1A1Ixp33_ASAP7_75t_L g359 ( .A1(n_274), .A2(n_315), .B(n_360), .C(n_362), .Y(n_359) );
INVx1_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
AND2x2_ASAP7_75t_L g326 ( .A(n_276), .B(n_283), .Y(n_326) );
BUFx2_ASAP7_75t_L g336 ( .A(n_276), .Y(n_336) );
INVx1_ASAP7_75t_L g351 ( .A(n_276), .Y(n_351) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
NOR2xp33_ASAP7_75t_L g278 ( .A(n_279), .B(n_280), .Y(n_278) );
OR2x2_ASAP7_75t_L g357 ( .A(n_279), .B(n_358), .Y(n_357) );
INVx1_ASAP7_75t_L g440 ( .A(n_279), .Y(n_440) );
INVx1_ASAP7_75t_L g433 ( .A(n_280), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_282), .B(n_283), .Y(n_281) );
AND2x2_ASAP7_75t_L g286 ( .A(n_282), .B(n_287), .Y(n_286) );
AND2x2_ASAP7_75t_L g390 ( .A(n_282), .B(n_307), .Y(n_390) );
INVx1_ASAP7_75t_L g319 ( .A(n_283), .Y(n_319) );
AOI22xp5_ASAP7_75t_L g285 ( .A1(n_286), .A2(n_290), .B1(n_293), .B2(n_295), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_287), .B(n_403), .Y(n_402) );
INVxp67_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
AND2x4_ASAP7_75t_L g355 ( .A(n_288), .B(n_356), .Y(n_355) );
BUFx3_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
AND2x2_ASAP7_75t_SL g318 ( .A(n_289), .B(n_298), .Y(n_318) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
AND2x2_ASAP7_75t_L g310 ( .A(n_292), .B(n_311), .Y(n_310) );
INVx1_ASAP7_75t_SL g293 ( .A(n_294), .Y(n_293) );
OR2x2_ASAP7_75t_L g320 ( .A(n_294), .B(n_321), .Y(n_320) );
INVx1_ASAP7_75t_SL g296 ( .A(n_297), .Y(n_296) );
OAI221xp5_ASAP7_75t_L g414 ( .A1(n_297), .A2(n_415), .B1(n_417), .B2(n_418), .C(n_419), .Y(n_414) );
INVx1_ASAP7_75t_L g303 ( .A(n_298), .Y(n_303) );
HB1xp67_ASAP7_75t_L g369 ( .A(n_298), .Y(n_369) );
INVx1_ASAP7_75t_SL g300 ( .A(n_301), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_301), .B(n_420), .Y(n_419) );
OAI21xp5_ASAP7_75t_L g309 ( .A1(n_302), .A2(n_307), .B(n_310), .Y(n_309) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_305), .B(n_315), .Y(n_412) );
AND2x2_ASAP7_75t_L g305 ( .A(n_306), .B(n_307), .Y(n_305) );
INVx1_ASAP7_75t_L g381 ( .A(n_306), .Y(n_381) );
AND2x2_ASAP7_75t_L g340 ( .A(n_307), .B(n_341), .Y(n_340) );
INVx2_ASAP7_75t_L g429 ( .A(n_307), .Y(n_429) );
INVx1_ASAP7_75t_L g345 ( .A(n_310), .Y(n_345) );
INVx1_ASAP7_75t_L g400 ( .A(n_311), .Y(n_400) );
OAI22xp5_ASAP7_75t_L g313 ( .A1(n_314), .A2(n_316), .B1(n_319), .B2(n_320), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_317), .B(n_318), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_317), .B(n_351), .Y(n_350) );
INVx2_ASAP7_75t_L g385 ( .A(n_318), .Y(n_385) );
NAND2xp5_ASAP7_75t_SL g422 ( .A(n_318), .B(n_356), .Y(n_422) );
OR2x2_ASAP7_75t_L g395 ( .A(n_319), .B(n_348), .Y(n_395) );
INVx1_ASAP7_75t_L g334 ( .A(n_320), .Y(n_334) );
INVx1_ASAP7_75t_SL g321 ( .A(n_322), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_322), .B(n_373), .Y(n_372) );
NOR3xp33_ASAP7_75t_L g323 ( .A(n_324), .B(n_342), .C(n_353), .Y(n_323) );
OAI211xp5_ASAP7_75t_L g324 ( .A1(n_325), .A2(n_327), .B(n_331), .C(n_337), .Y(n_324) );
INVxp67_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
AOI221xp5_ASAP7_75t_L g396 ( .A1(n_326), .A2(n_397), .B1(n_401), .B2(n_404), .C(n_406), .Y(n_396) );
INVx1_ASAP7_75t_SL g327 ( .A(n_328), .Y(n_327) );
AND2x2_ASAP7_75t_L g328 ( .A(n_329), .B(n_330), .Y(n_328) );
AND2x2_ASAP7_75t_L g338 ( .A(n_329), .B(n_339), .Y(n_338) );
AND2x2_ASAP7_75t_L g392 ( .A(n_329), .B(n_393), .Y(n_392) );
OAI211xp5_ASAP7_75t_L g377 ( .A1(n_330), .A2(n_378), .B(n_380), .C(n_382), .Y(n_377) );
INVx2_ASAP7_75t_L g424 ( .A(n_330), .Y(n_424) );
OAI21xp5_ASAP7_75t_SL g331 ( .A1(n_332), .A2(n_334), .B(n_335), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
AND2x2_ASAP7_75t_L g403 ( .A(n_336), .B(n_356), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_338), .B(n_340), .Y(n_337) );
OAI21xp5_ASAP7_75t_SL g342 ( .A1(n_343), .A2(n_345), .B(n_346), .Y(n_342) );
INVxp67_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
OAI21xp5_ASAP7_75t_SL g346 ( .A1(n_347), .A2(n_349), .B(n_352), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_347), .B(n_376), .Y(n_375) );
INVxp67_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_352), .B(n_439), .Y(n_438) );
OAI21xp33_ASAP7_75t_L g353 ( .A1(n_354), .A2(n_357), .B(n_359), .Y(n_353) );
INVx1_ASAP7_75t_SL g354 ( .A(n_355), .Y(n_354) );
AND2x2_ASAP7_75t_L g380 ( .A(n_356), .B(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
AND4x1_ASAP7_75t_L g365 ( .A(n_366), .B(n_396), .C(n_413), .D(n_435), .Y(n_365) );
NOR2xp33_ASAP7_75t_L g366 ( .A(n_367), .B(n_383), .Y(n_366) );
OAI211xp5_ASAP7_75t_SL g367 ( .A1(n_368), .A2(n_372), .B(n_375), .C(n_377), .Y(n_367) );
OR2x2_ASAP7_75t_L g368 ( .A(n_369), .B(n_370), .Y(n_368) );
INVx1_ASAP7_75t_SL g370 ( .A(n_371), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_371), .B(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
NOR2xp33_ASAP7_75t_L g404 ( .A(n_382), .B(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
NOR2xp33_ASAP7_75t_L g391 ( .A(n_392), .B(n_394), .Y(n_391) );
INVx1_ASAP7_75t_L g417 ( .A(n_392), .Y(n_417) );
INVx2_ASAP7_75t_SL g405 ( .A(n_393), .Y(n_405) );
OR2x2_ASAP7_75t_L g398 ( .A(n_399), .B(n_400), .Y(n_398) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g418 ( .A(n_403), .Y(n_418) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
NOR2xp33_ASAP7_75t_SL g413 ( .A(n_414), .B(n_421), .Y(n_413) );
INVx1_ASAP7_75t_SL g415 ( .A(n_416), .Y(n_415) );
OAI221xp5_ASAP7_75t_SL g421 ( .A1(n_422), .A2(n_423), .B1(n_425), .B2(n_426), .C(n_427), .Y(n_421) );
AOI22xp5_ASAP7_75t_L g427 ( .A1(n_428), .A2(n_432), .B1(n_433), .B2(n_434), .Y(n_427) );
NAND2xp5_ASAP7_75t_SL g428 ( .A(n_429), .B(n_430), .Y(n_428) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx2_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx2_ASAP7_75t_L g735 ( .A(n_444), .Y(n_735) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx2_ASAP7_75t_L g736 ( .A(n_446), .Y(n_736) );
OR3x1_ASAP7_75t_L g446 ( .A(n_447), .B(n_628), .C(n_693), .Y(n_446) );
NAND4xp25_ASAP7_75t_SL g447 ( .A(n_448), .B(n_569), .C(n_595), .D(n_618), .Y(n_447) );
AOI221xp5_ASAP7_75t_L g448 ( .A1(n_449), .A2(n_501), .B1(n_539), .B2(n_546), .C(n_561), .Y(n_448) );
CKINVDCx14_ASAP7_75t_R g449 ( .A(n_450), .Y(n_449) );
OAI22xp5_ASAP7_75t_L g716 ( .A1(n_450), .A2(n_562), .B1(n_586), .B2(n_717), .Y(n_716) );
OR2x2_ASAP7_75t_L g450 ( .A(n_451), .B(n_482), .Y(n_450) );
INVx1_ASAP7_75t_SL g622 ( .A(n_451), .Y(n_622) );
OR2x2_ASAP7_75t_L g451 ( .A(n_452), .B(n_466), .Y(n_451) );
OR2x2_ASAP7_75t_L g544 ( .A(n_452), .B(n_545), .Y(n_544) );
AND2x2_ASAP7_75t_L g564 ( .A(n_452), .B(n_483), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_452), .B(n_491), .Y(n_577) );
AND2x2_ASAP7_75t_L g594 ( .A(n_452), .B(n_466), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_452), .B(n_542), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_452), .B(n_593), .Y(n_705) );
NOR2xp33_ASAP7_75t_L g715 ( .A(n_452), .B(n_482), .Y(n_715) );
AOI211xp5_ASAP7_75t_SL g726 ( .A1(n_452), .A2(n_632), .B(n_727), .C(n_728), .Y(n_726) );
INVx5_ASAP7_75t_SL g452 ( .A(n_453), .Y(n_452) );
NAND2xp5_ASAP7_75t_SL g598 ( .A(n_453), .B(n_483), .Y(n_598) );
AND2x2_ASAP7_75t_L g601 ( .A(n_453), .B(n_484), .Y(n_601) );
OR2x2_ASAP7_75t_L g646 ( .A(n_453), .B(n_483), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_453), .B(n_491), .Y(n_655) );
OAI21xp5_ASAP7_75t_L g454 ( .A1(n_455), .A2(n_456), .B(n_458), .Y(n_454) );
INVx5_ASAP7_75t_L g472 ( .A(n_459), .Y(n_472) );
INVx5_ASAP7_75t_SL g545 ( .A(n_466), .Y(n_545) );
AND2x2_ASAP7_75t_L g563 ( .A(n_466), .B(n_564), .Y(n_563) );
NOR2xp33_ASAP7_75t_L g645 ( .A(n_466), .B(n_646), .Y(n_645) );
AND2x2_ASAP7_75t_L g649 ( .A(n_466), .B(n_650), .Y(n_649) );
AND2x2_ASAP7_75t_L g681 ( .A(n_466), .B(n_491), .Y(n_681) );
OR2x2_ASAP7_75t_L g687 ( .A(n_466), .B(n_577), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_466), .B(n_637), .Y(n_696) );
OR2x6_ASAP7_75t_L g466 ( .A(n_467), .B(n_481), .Y(n_466) );
BUFx2_ASAP7_75t_L g518 ( .A(n_469), .Y(n_518) );
INVx2_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
O2A1O1Ixp33_ASAP7_75t_L g494 ( .A1(n_472), .A2(n_480), .B(n_495), .C(n_496), .Y(n_494) );
O2A1O1Ixp33_ASAP7_75t_SL g553 ( .A1(n_472), .A2(n_480), .B(n_554), .C(n_555), .Y(n_553) );
O2A1O1Ixp33_ASAP7_75t_L g473 ( .A1(n_474), .A2(n_475), .B(n_477), .C(n_478), .Y(n_473) );
O2A1O1Ixp33_ASAP7_75t_L g508 ( .A1(n_475), .A2(n_478), .B(n_509), .C(n_510), .Y(n_508) );
INVx2_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_483), .B(n_491), .Y(n_482) );
AND2x2_ASAP7_75t_L g578 ( .A(n_483), .B(n_545), .Y(n_578) );
INVx1_ASAP7_75t_SL g591 ( .A(n_483), .Y(n_591) );
OR2x2_ASAP7_75t_L g626 ( .A(n_483), .B(n_627), .Y(n_626) );
OR2x2_ASAP7_75t_L g632 ( .A(n_483), .B(n_491), .Y(n_632) );
AND2x2_ASAP7_75t_L g690 ( .A(n_483), .B(n_542), .Y(n_690) );
INVx2_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_484), .B(n_545), .Y(n_617) );
INVx3_ASAP7_75t_L g542 ( .A(n_491), .Y(n_542) );
OR2x2_ASAP7_75t_L g583 ( .A(n_491), .B(n_545), .Y(n_583) );
AND2x2_ASAP7_75t_L g593 ( .A(n_491), .B(n_591), .Y(n_593) );
HB1xp67_ASAP7_75t_L g641 ( .A(n_491), .Y(n_641) );
AND2x2_ASAP7_75t_L g650 ( .A(n_491), .B(n_564), .Y(n_650) );
OA21x2_ASAP7_75t_L g491 ( .A1(n_492), .A2(n_493), .B(n_499), .Y(n_491) );
OA21x2_ASAP7_75t_L g551 ( .A1(n_500), .A2(n_552), .B(n_560), .Y(n_551) );
AOI221xp5_ASAP7_75t_L g666 ( .A1(n_501), .A2(n_667), .B1(n_669), .B2(n_671), .C(n_674), .Y(n_666) );
INVx2_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
OR2x2_ASAP7_75t_L g502 ( .A(n_503), .B(n_513), .Y(n_502) );
AND2x2_ASAP7_75t_L g640 ( .A(n_503), .B(n_621), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_503), .B(n_699), .Y(n_703) );
OR2x2_ASAP7_75t_L g724 ( .A(n_503), .B(n_725), .Y(n_724) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_503), .B(n_729), .Y(n_728) );
BUFx2_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
INVx5_ASAP7_75t_L g571 ( .A(n_504), .Y(n_571) );
AND2x2_ASAP7_75t_L g648 ( .A(n_504), .B(n_515), .Y(n_648) );
AND2x2_ASAP7_75t_L g709 ( .A(n_504), .B(n_588), .Y(n_709) );
AND2x2_ASAP7_75t_L g722 ( .A(n_504), .B(n_542), .Y(n_722) );
OR2x6_ASAP7_75t_L g504 ( .A(n_505), .B(n_511), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_514), .B(n_527), .Y(n_513) );
AND2x4_ASAP7_75t_L g549 ( .A(n_514), .B(n_550), .Y(n_549) );
AND2x2_ASAP7_75t_L g567 ( .A(n_514), .B(n_568), .Y(n_567) );
INVx2_ASAP7_75t_L g574 ( .A(n_514), .Y(n_574) );
AND2x2_ASAP7_75t_L g643 ( .A(n_514), .B(n_621), .Y(n_643) );
AND2x2_ASAP7_75t_L g653 ( .A(n_514), .B(n_571), .Y(n_653) );
HB1xp67_ASAP7_75t_L g661 ( .A(n_514), .Y(n_661) );
AND2x2_ASAP7_75t_L g673 ( .A(n_514), .B(n_551), .Y(n_673) );
NOR2xp33_ASAP7_75t_L g677 ( .A(n_514), .B(n_605), .Y(n_677) );
AND2x2_ASAP7_75t_L g714 ( .A(n_514), .B(n_709), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_514), .B(n_588), .Y(n_725) );
OR2x2_ASAP7_75t_L g727 ( .A(n_514), .B(n_663), .Y(n_727) );
INVx5_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
AND2x2_ASAP7_75t_L g613 ( .A(n_515), .B(n_614), .Y(n_613) );
AND2x2_ASAP7_75t_L g623 ( .A(n_515), .B(n_568), .Y(n_623) );
AND2x2_ASAP7_75t_L g635 ( .A(n_515), .B(n_551), .Y(n_635) );
HB1xp67_ASAP7_75t_L g665 ( .A(n_515), .Y(n_665) );
AND2x4_ASAP7_75t_L g699 ( .A(n_515), .B(n_550), .Y(n_699) );
OR2x6_ASAP7_75t_L g515 ( .A(n_516), .B(n_524), .Y(n_515) );
AOI21xp5_ASAP7_75t_SL g516 ( .A1(n_517), .A2(n_519), .B(n_523), .Y(n_516) );
NOR2xp33_ASAP7_75t_L g524 ( .A(n_525), .B(n_526), .Y(n_524) );
BUFx2_ASAP7_75t_L g548 ( .A(n_527), .Y(n_548) );
HB1xp67_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
INVx2_ASAP7_75t_L g588 ( .A(n_528), .Y(n_588) );
AND2x2_ASAP7_75t_L g621 ( .A(n_528), .B(n_551), .Y(n_621) );
INVx2_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
AND2x2_ASAP7_75t_L g568 ( .A(n_529), .B(n_551), .Y(n_568) );
BUFx2_ASAP7_75t_L g614 ( .A(n_529), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_531), .B(n_536), .Y(n_530) );
INVx1_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_541), .B(n_543), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_541), .B(n_622), .Y(n_701) );
INVx1_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_542), .B(n_564), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_542), .B(n_545), .Y(n_603) );
AND2x2_ASAP7_75t_L g658 ( .A(n_542), .B(n_594), .Y(n_658) );
AOI221xp5_ASAP7_75t_SL g595 ( .A1(n_543), .A2(n_596), .B1(n_604), .B2(n_606), .C(n_610), .Y(n_595) );
INVx2_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
OR2x2_ASAP7_75t_L g590 ( .A(n_544), .B(n_591), .Y(n_590) );
OR2x2_ASAP7_75t_L g631 ( .A(n_544), .B(n_632), .Y(n_631) );
OAI321xp33_ASAP7_75t_L g638 ( .A1(n_544), .A2(n_597), .A3(n_639), .B1(n_641), .B2(n_642), .C(n_644), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_545), .B(n_690), .Y(n_689) );
INVx1_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_548), .B(n_549), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_548), .B(n_699), .Y(n_717) );
AND2x2_ASAP7_75t_L g604 ( .A(n_549), .B(n_605), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_549), .B(n_608), .Y(n_607) );
HB1xp67_ASAP7_75t_L g580 ( .A(n_550), .Y(n_580) );
AND2x2_ASAP7_75t_L g587 ( .A(n_550), .B(n_588), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_550), .B(n_662), .Y(n_692) );
INVx1_ASAP7_75t_L g729 ( .A(n_550), .Y(n_729) );
INVx2_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
NOR2xp33_ASAP7_75t_L g556 ( .A(n_557), .B(n_558), .Y(n_556) );
AOI21xp5_ASAP7_75t_L g561 ( .A1(n_562), .A2(n_565), .B(n_566), .Y(n_561) );
INVx1_ASAP7_75t_SL g562 ( .A(n_563), .Y(n_562) );
A2O1A1Ixp33_ASAP7_75t_L g721 ( .A1(n_563), .A2(n_673), .B(n_722), .C(n_723), .Y(n_721) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_564), .B(n_582), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_564), .B(n_602), .Y(n_668) );
INVx1_ASAP7_75t_SL g566 ( .A(n_567), .Y(n_566) );
INVx1_ASAP7_75t_L g611 ( .A(n_568), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_568), .B(n_571), .Y(n_625) );
NOR2xp33_ASAP7_75t_L g634 ( .A(n_568), .B(n_635), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_568), .B(n_653), .Y(n_652) );
AOI22xp33_ASAP7_75t_L g569 ( .A1(n_570), .A2(n_572), .B1(n_584), .B2(n_589), .Y(n_569) );
HB1xp67_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
OR2x2_ASAP7_75t_L g585 ( .A(n_571), .B(n_586), .Y(n_585) );
AND2x2_ASAP7_75t_L g608 ( .A(n_571), .B(n_609), .Y(n_608) );
AND2x2_ASAP7_75t_L g620 ( .A(n_571), .B(n_621), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_571), .B(n_614), .Y(n_656) );
OR2x2_ASAP7_75t_L g663 ( .A(n_571), .B(n_588), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_571), .B(n_673), .Y(n_672) );
AND2x2_ASAP7_75t_L g713 ( .A(n_571), .B(n_699), .Y(n_713) );
OAI22xp33_ASAP7_75t_L g572 ( .A1(n_573), .A2(n_575), .B1(n_579), .B2(n_581), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
AND2x2_ASAP7_75t_L g619 ( .A(n_574), .B(n_620), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_576), .B(n_578), .Y(n_575) );
INVx1_ASAP7_75t_SL g576 ( .A(n_577), .Y(n_576) );
OAI22xp33_ASAP7_75t_L g659 ( .A1(n_577), .A2(n_592), .B1(n_660), .B2(n_664), .Y(n_659) );
INVx1_ASAP7_75t_L g707 ( .A(n_578), .Y(n_707) );
INVx1_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
AOI221xp5_ASAP7_75t_L g618 ( .A1(n_582), .A2(n_619), .B1(n_622), .B2(n_623), .C(n_624), .Y(n_618) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
OR2x2_ASAP7_75t_L g597 ( .A(n_583), .B(n_598), .Y(n_597) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_587), .B(n_653), .Y(n_685) );
HB1xp67_ASAP7_75t_L g605 ( .A(n_588), .Y(n_605) );
INVx1_ASAP7_75t_L g609 ( .A(n_588), .Y(n_609) );
NAND2xp33_ASAP7_75t_L g589 ( .A(n_590), .B(n_592), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_593), .B(n_594), .Y(n_592) );
INVx1_ASAP7_75t_L g627 ( .A(n_594), .Y(n_627) );
AND2x2_ASAP7_75t_L g636 ( .A(n_594), .B(n_637), .Y(n_636) );
NAND2xp33_ASAP7_75t_L g596 ( .A(n_597), .B(n_599), .Y(n_596) );
INVx2_ASAP7_75t_SL g599 ( .A(n_600), .Y(n_599) );
AND2x4_ASAP7_75t_L g600 ( .A(n_601), .B(n_602), .Y(n_600) );
AND2x2_ASAP7_75t_L g680 ( .A(n_601), .B(n_681), .Y(n_680) );
INVx2_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
AOI221xp5_ASAP7_75t_L g629 ( .A1(n_604), .A2(n_630), .B1(n_633), .B2(n_636), .C(n_638), .Y(n_629) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_608), .B(n_665), .Y(n_664) );
AOI21xp33_ASAP7_75t_SL g610 ( .A1(n_611), .A2(n_612), .B(n_615), .Y(n_610) );
INVx2_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
CKINVDCx16_ASAP7_75t_R g712 ( .A(n_615), .Y(n_712) );
OR2x2_ASAP7_75t_L g615 ( .A(n_616), .B(n_617), .Y(n_615) );
OR2x2_ASAP7_75t_L g654 ( .A(n_617), .B(n_655), .Y(n_654) );
INVx1_ASAP7_75t_SL g675 ( .A(n_620), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_620), .B(n_680), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_623), .B(n_645), .Y(n_644) );
NOR2xp33_ASAP7_75t_L g624 ( .A(n_625), .B(n_626), .Y(n_624) );
NAND4xp25_ASAP7_75t_L g628 ( .A(n_629), .B(n_647), .C(n_666), .D(n_679), .Y(n_628) );
INVx1_ASAP7_75t_SL g630 ( .A(n_631), .Y(n_630) );
INVx1_ASAP7_75t_SL g637 ( .A(n_632), .Y(n_637) );
INVxp67_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
OR2x2_ASAP7_75t_L g670 ( .A(n_641), .B(n_646), .Y(n_670) );
INVxp67_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
AOI211xp5_ASAP7_75t_L g647 ( .A1(n_648), .A2(n_649), .B(n_651), .C(n_659), .Y(n_647) );
AOI211xp5_ASAP7_75t_L g718 ( .A1(n_649), .A2(n_691), .B(n_719), .C(n_726), .Y(n_718) );
INVx1_ASAP7_75t_SL g678 ( .A(n_650), .Y(n_678) );
OAI22xp5_ASAP7_75t_L g651 ( .A1(n_652), .A2(n_654), .B1(n_656), .B2(n_657), .Y(n_651) );
INVx1_ASAP7_75t_L g682 ( .A(n_656), .Y(n_682) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_661), .B(n_662), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_662), .B(n_699), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_662), .B(n_673), .Y(n_706) );
INVx2_ASAP7_75t_SL g662 ( .A(n_663), .Y(n_662) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
INVx1_ASAP7_75t_SL g669 ( .A(n_670), .Y(n_669) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
INVx1_ASAP7_75t_L g683 ( .A(n_673), .Y(n_683) );
AOI21xp33_ASAP7_75t_L g674 ( .A1(n_675), .A2(n_676), .B(n_678), .Y(n_674) );
INVxp33_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
AOI322xp5_ASAP7_75t_L g679 ( .A1(n_680), .A2(n_682), .A3(n_683), .B1(n_684), .B2(n_686), .C1(n_688), .C2(n_691), .Y(n_679) );
INVxp67_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
NAND3xp33_ASAP7_75t_SL g693 ( .A(n_694), .B(n_711), .C(n_718), .Y(n_693) );
AOI221xp5_ASAP7_75t_L g694 ( .A1(n_695), .A2(n_697), .B1(n_700), .B2(n_702), .C(n_704), .Y(n_694) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
INVx1_ASAP7_75t_SL g710 ( .A(n_699), .Y(n_710) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVxp67_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
OAI22xp33_ASAP7_75t_L g704 ( .A1(n_705), .A2(n_706), .B1(n_707), .B2(n_708), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_709), .B(n_710), .Y(n_708) );
AOI221xp5_ASAP7_75t_L g711 ( .A1(n_712), .A2(n_713), .B1(n_714), .B2(n_715), .C(n_716), .Y(n_711) );
NAND2xp33_ASAP7_75t_L g719 ( .A(n_720), .B(n_721), .Y(n_719) );
INVxp67_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx2_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
INVx2_ASAP7_75t_L g737 ( .A(n_731), .Y(n_737) );
INVx1_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
INVx1_ASAP7_75t_SL g738 ( .A(n_739), .Y(n_738) );
INVx3_ASAP7_75t_SL g739 ( .A(n_740), .Y(n_739) );
INVxp67_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
HB1xp67_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
INVx1_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
INVx1_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
INVx1_ASAP7_75t_SL g750 ( .A(n_751), .Y(n_750) );
endmodule