module fake_jpeg_3873_n_46 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_46);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_46;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_43;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx5_ASAP7_75t_L g7 ( 
.A(n_1),
.Y(n_7)
);

BUFx3_ASAP7_75t_L g8 ( 
.A(n_2),
.Y(n_8)
);

INVxp67_ASAP7_75t_L g9 ( 
.A(n_4),
.Y(n_9)
);

INVx2_ASAP7_75t_L g10 ( 
.A(n_2),
.Y(n_10)
);

NOR2xp33_ASAP7_75t_L g11 ( 
.A(n_2),
.B(n_0),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_4),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g13 ( 
.A(n_0),
.B(n_5),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_12),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_14),
.B(n_15),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_12),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_11),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_16),
.B(n_17),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g17 ( 
.A(n_7),
.B(n_0),
.C(n_1),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_18),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_11),
.B(n_1),
.Y(n_19)
);

CKINVDCx14_ASAP7_75t_R g22 ( 
.A(n_19),
.Y(n_22)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g24 ( 
.A(n_20),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_16),
.A2(n_10),
.B1(n_7),
.B2(n_13),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_21),
.A2(n_25),
.B1(n_17),
.B2(n_20),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_18),
.A2(n_10),
.B1(n_13),
.B2(n_9),
.Y(n_25)
);

CKINVDCx16_ASAP7_75t_R g28 ( 
.A(n_27),
.Y(n_28)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_25),
.Y(n_29)
);

INVxp33_ASAP7_75t_SL g36 ( 
.A(n_29),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_30),
.A2(n_31),
.B1(n_3),
.B2(n_29),
.Y(n_38)
);

CKINVDCx14_ASAP7_75t_R g31 ( 
.A(n_21),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_26),
.A2(n_8),
.B1(n_3),
.B2(n_6),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g35 ( 
.A1(n_32),
.A2(n_24),
.B1(n_5),
.B2(n_6),
.Y(n_35)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_33),
.A2(n_24),
.B1(n_22),
.B2(n_26),
.Y(n_34)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

AOI21xp5_ASAP7_75t_L g41 ( 
.A1(n_35),
.A2(n_38),
.B(n_33),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_36),
.B(n_30),
.C(n_32),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_39),
.B(n_35),
.Y(n_43)
);

CKINVDCx14_ASAP7_75t_R g42 ( 
.A(n_41),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_43),
.A2(n_40),
.B1(n_36),
.B2(n_37),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_44),
.B(n_42),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_45),
.B(n_3),
.Y(n_46)
);


endmodule