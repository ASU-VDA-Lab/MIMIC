module real_jpeg_25492_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_201;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_200;
wire n_56;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_242;
wire n_141;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_238;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_239;
wire n_162;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_211;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_150;
wire n_32;
wire n_20;
wire n_80;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_213;
wire n_179;
wire n_202;
wire n_216;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

INVx3_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g92 ( 
.A(n_1),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_2),
.B(n_46),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_2),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_2),
.B(n_74),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_2),
.B(n_55),
.C(n_57),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_2),
.A2(n_38),
.B1(n_39),
.B2(n_108),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_2),
.B(n_66),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_2),
.A2(n_54),
.B1(n_55),
.B2(n_108),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_2),
.B(n_27),
.C(n_92),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_2),
.A2(n_26),
.B(n_200),
.Y(n_225)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

INVx8_ASAP7_75t_SL g44 ( 
.A(n_4),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_5),
.A2(n_38),
.B1(n_39),
.B2(n_62),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g62 ( 
.A(n_5),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_5),
.A2(n_42),
.B1(n_62),
.B2(n_72),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_5),
.A2(n_54),
.B1(n_55),
.B2(n_62),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_5),
.A2(n_27),
.B1(n_31),
.B2(n_62),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_6),
.A2(n_27),
.B1(n_31),
.B2(n_32),
.Y(n_30)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_6),
.A2(n_32),
.B1(n_54),
.B2(n_55),
.Y(n_97)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_7),
.Y(n_57)
);

OAI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_8),
.A2(n_38),
.B1(n_39),
.B2(n_65),
.Y(n_64)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_8),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_8),
.A2(n_47),
.B1(n_65),
.B2(n_78),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_8),
.A2(n_54),
.B1(n_55),
.B2(n_65),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_8),
.A2(n_27),
.B1(n_31),
.B2(n_65),
.Y(n_170)
);

INVx13_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_10),
.A2(n_27),
.B1(n_31),
.B2(n_36),
.Y(n_35)
);

CKINVDCx14_ASAP7_75t_R g36 ( 
.A(n_10),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_10),
.A2(n_36),
.B1(n_54),
.B2(n_55),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_11),
.A2(n_27),
.B1(n_31),
.B2(n_85),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_11),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_12),
.A2(n_54),
.B1(n_55),
.B2(n_96),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_12),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_12),
.A2(n_38),
.B1(n_39),
.B2(n_96),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_L g154 ( 
.A1(n_12),
.A2(n_27),
.B1(n_31),
.B2(n_96),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_13),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_14),
.A2(n_47),
.B1(n_70),
.B2(n_71),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_14),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_14),
.A2(n_38),
.B1(n_39),
.B2(n_70),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g173 ( 
.A1(n_14),
.A2(n_54),
.B1(n_55),
.B2(n_70),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_14),
.A2(n_27),
.B1(n_31),
.B2(n_70),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_15),
.A2(n_27),
.B1(n_31),
.B2(n_118),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_15),
.Y(n_118)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_16),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_138),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_137),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_111),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_21),
.B(n_111),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_81),
.C(n_98),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_22),
.B(n_156),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_50),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_23),
.B(n_51),
.C(n_67),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_37),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_24),
.B(n_37),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_29),
.B1(n_33),
.B2(n_35),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_25),
.A2(n_211),
.B1(n_213),
.B2(n_214),
.Y(n_210)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_26),
.A2(n_83),
.B1(n_84),
.B2(n_86),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_26),
.A2(n_84),
.B1(n_117),
.B2(n_119),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_26),
.A2(n_28),
.B1(n_30),
.B2(n_154),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_26),
.B(n_170),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_26),
.A2(n_199),
.B(n_200),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_28),
.Y(n_26)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_27),
.Y(n_31)
);

OA22x2_ASAP7_75t_L g94 ( 
.A1(n_27),
.A2(n_31),
.B1(n_92),
.B2(n_93),
.Y(n_94)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_28),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_30),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_31),
.B(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_33),
.Y(n_119)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_34),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_34),
.B(n_108),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_35),
.Y(n_83)
);

AOI32xp33_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_41),
.A3(n_43),
.B1(n_45),
.B2(n_48),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_38),
.A2(n_39),
.B1(n_57),
.B2(n_58),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_38),
.A2(n_39),
.B1(n_43),
.B2(n_49),
.Y(n_74)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

NAND2xp33_ASAP7_75t_SL g48 ( 
.A(n_39),
.B(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_39),
.B(n_163),
.Y(n_162)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx11_ASAP7_75t_L g78 ( 
.A(n_41),
.Y(n_78)
);

OAI22xp33_ASAP7_75t_L g80 ( 
.A1(n_41),
.A2(n_42),
.B1(n_43),
.B2(n_49),
.Y(n_80)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVxp33_ASAP7_75t_L g109 ( 
.A(n_45),
.Y(n_109)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

OAI21xp33_ASAP7_75t_L g107 ( 
.A1(n_47),
.A2(n_108),
.B(n_109),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_67),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_SL g51 ( 
.A1(n_52),
.A2(n_60),
.B(n_63),
.Y(n_51)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_52),
.Y(n_105)
);

OAI21xp33_ASAP7_75t_L g176 ( 
.A1(n_52),
.A2(n_63),
.B(n_177),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_59),
.Y(n_52)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_53),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_53),
.A2(n_134),
.B(n_135),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_53),
.A2(n_135),
.B(n_150),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_54),
.A2(n_55),
.B1(n_57),
.B2(n_58),
.Y(n_53)
);

OAI22xp33_ASAP7_75t_L g91 ( 
.A1(n_54),
.A2(n_55),
.B1(n_92),
.B2(n_93),
.Y(n_91)
);

INVx4_ASAP7_75t_SL g54 ( 
.A(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_55),
.B(n_207),
.Y(n_206)
);

BUFx4f_ASAP7_75t_SL g55 ( 
.A(n_56),
.Y(n_55)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_57),
.Y(n_58)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_61),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_61),
.A2(n_66),
.B1(n_104),
.B2(n_105),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_64),
.B(n_66),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_64),
.B(n_105),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g67 ( 
.A1(n_68),
.A2(n_73),
.B(n_75),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_69),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_69),
.A2(n_74),
.B1(n_79),
.B2(n_131),
.Y(n_130)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_73),
.B(n_80),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_73),
.B(n_77),
.Y(n_110)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_79),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_79),
.A2(n_107),
.B(n_110),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_81),
.B(n_98),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_88),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_82),
.B(n_88),
.Y(n_136)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_87),
.B(n_201),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_89),
.A2(n_94),
.B1(n_95),
.B2(n_97),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_89),
.A2(n_187),
.B(n_188),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_89),
.A2(n_188),
.B(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_90),
.B(n_102),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_90),
.A2(n_121),
.B1(n_122),
.B2(n_123),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_90),
.A2(n_123),
.B1(n_172),
.B2(n_174),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_94),
.Y(n_90)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_92),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_94),
.A2(n_95),
.B(n_101),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_94),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_94),
.A2(n_101),
.B(n_173),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_94),
.B(n_108),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_97),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_103),
.C(n_106),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_99),
.A2(n_100),
.B1(n_103),
.B2(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_102),
.B(n_123),
.Y(n_188)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_103),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_104),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_106),
.B(n_145),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_113),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_114),
.A2(n_115),
.B1(n_126),
.B2(n_127),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_116),
.A2(n_120),
.B1(n_124),
.B2(n_125),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_116),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_120),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_136),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_130),
.B1(n_132),
.B2(n_133),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_139),
.B(n_242),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_157),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_155),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g243 ( 
.A(n_142),
.B(n_155),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_147),
.C(n_148),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_143),
.A2(n_144),
.B1(n_238),
.B2(n_239),
.Y(n_237)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_SL g239 ( 
.A(n_147),
.B(n_148),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_151),
.C(n_153),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_149),
.B(n_181),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_151),
.A2(n_152),
.B1(n_153),
.B2(n_182),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_153),
.Y(n_182)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_154),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_158),
.A2(n_236),
.B(n_241),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_189),
.B(n_235),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_178),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_160),
.B(n_178),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_171),
.C(n_175),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_161),
.B(n_231),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_SL g161 ( 
.A(n_162),
.B(n_164),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_162),
.B(n_164),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_165),
.A2(n_166),
.B(n_169),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_167),
.Y(n_166)
);

BUFx2_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_168),
.A2(n_212),
.B(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_169),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_170),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_171),
.A2(n_175),
.B1(n_176),
.B2(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_171),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_174),
.Y(n_187)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_179),
.A2(n_180),
.B1(n_183),
.B2(n_184),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_179),
.B(n_185),
.C(n_186),
.Y(n_240)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_186),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_190),
.A2(n_229),
.B(n_234),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_191),
.A2(n_208),
.B(n_228),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_192),
.B(n_202),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_192),
.B(n_202),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_198),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_194),
.A2(n_195),
.B1(n_196),
.B2(n_197),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_194),
.B(n_197),
.C(n_198),
.Y(n_233)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g214 ( 
.A(n_199),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_203),
.B(n_206),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_203),
.A2(n_204),
.B1(n_206),
.B2(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_206),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_209),
.A2(n_217),
.B(n_227),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_215),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_210),
.B(n_215),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g211 ( 
.A(n_212),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_218),
.A2(n_222),
.B(n_226),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_220),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_219),
.B(n_220),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_225),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_230),
.B(n_233),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_230),
.B(n_233),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_237),
.B(n_240),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_237),
.B(n_240),
.Y(n_241)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);


endmodule