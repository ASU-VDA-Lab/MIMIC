module fake_jpeg_28588_n_192 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_192);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_192;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_96;

BUFx24_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_13),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

CKINVDCx16_ASAP7_75t_R g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_30),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_34),
.B(n_36),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_31),
.B(n_0),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_37),
.B(n_45),
.Y(n_46)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_30),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_39),
.B(n_24),
.Y(n_62)
);

BUFx10_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

BUFx4f_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_28),
.B(n_29),
.Y(n_45)
);

OA22x2_ASAP7_75t_L g47 ( 
.A1(n_38),
.A2(n_18),
.B1(n_17),
.B2(n_29),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_47),
.B(n_42),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_36),
.A2(n_29),
.B1(n_33),
.B2(n_32),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_49),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_37),
.A2(n_32),
.B1(n_28),
.B2(n_19),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_54),
.A2(n_65),
.B1(n_26),
.B2(n_23),
.Y(n_69)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_56),
.Y(n_87)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_57),
.B(n_59),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_35),
.A2(n_29),
.B1(n_19),
.B2(n_22),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_58),
.A2(n_36),
.B1(n_44),
.B2(n_39),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_45),
.B(n_22),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_43),
.B(n_27),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_60),
.B(n_1),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_62),
.B(n_20),
.Y(n_76)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

INVx5_ASAP7_75t_SL g84 ( 
.A(n_64),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_42),
.A2(n_33),
.B1(n_27),
.B2(n_26),
.Y(n_65)
);

O2A1O1Ixp33_ASAP7_75t_L g67 ( 
.A1(n_47),
.A2(n_60),
.B(n_46),
.C(n_53),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_67),
.Y(n_94)
);

OR2x2_ASAP7_75t_L g105 ( 
.A(n_68),
.B(n_70),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_69),
.A2(n_80),
.B1(n_89),
.B2(n_79),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_50),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_71),
.B(n_72),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_63),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_SL g73 ( 
.A1(n_46),
.A2(n_40),
.B(n_36),
.Y(n_73)
);

XOR2xp5_ASAP7_75t_L g98 ( 
.A(n_73),
.B(n_86),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_74),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_48),
.B(n_20),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_75),
.B(n_83),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_76),
.B(n_77),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_65),
.B(n_23),
.Y(n_77)
);

A2O1A1Ixp33_ASAP7_75t_L g78 ( 
.A1(n_47),
.A2(n_40),
.B(n_9),
.C(n_10),
.Y(n_78)
);

NOR2xp67_ASAP7_75t_L g93 ( 
.A(n_78),
.B(n_1),
.Y(n_93)
);

OAI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_47),
.A2(n_34),
.B1(n_40),
.B2(n_25),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_61),
.Y(n_81)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_81),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_48),
.B(n_25),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_82),
.B(n_91),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_64),
.B(n_7),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_63),
.Y(n_85)
);

CKINVDCx6p67_ASAP7_75t_R g111 ( 
.A(n_85),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_61),
.A2(n_63),
.B(n_25),
.Y(n_86)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_55),
.Y(n_88)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_88),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_51),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_51),
.B(n_0),
.Y(n_90)
);

MAJx2_ASAP7_75t_L g113 ( 
.A(n_90),
.B(n_5),
.C(n_13),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_56),
.B(n_7),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_92),
.B(n_2),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_SL g130 ( 
.A(n_93),
.B(n_90),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_95),
.B(n_112),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_102),
.A2(n_109),
.B1(n_84),
.B2(n_72),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_71),
.B(n_11),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_103),
.B(n_107),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_92),
.B(n_52),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_104),
.B(n_108),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_66),
.B(n_6),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_67),
.B(n_52),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_69),
.A2(n_3),
.B1(n_5),
.B2(n_15),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_83),
.B(n_9),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_SL g131 ( 
.A(n_113),
.B(n_79),
.Y(n_131)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_110),
.Y(n_114)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_114),
.Y(n_134)
);

INVx13_ASAP7_75t_L g115 ( 
.A(n_111),
.Y(n_115)
);

CKINVDCx14_ASAP7_75t_R g136 ( 
.A(n_115),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_98),
.B(n_73),
.C(n_86),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_116),
.B(n_128),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_96),
.B(n_97),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_117),
.B(n_119),
.Y(n_148)
);

INVx1_ASAP7_75t_SL g118 ( 
.A(n_111),
.Y(n_118)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_118),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_106),
.B(n_81),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_108),
.B(n_68),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_120),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_106),
.B(n_90),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_121),
.B(n_122),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_111),
.Y(n_122)
);

AND2x6_ASAP7_75t_L g123 ( 
.A(n_98),
.B(n_78),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_123),
.B(n_126),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_95),
.B(n_104),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_111),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_127),
.B(n_130),
.Y(n_133)
);

XNOR2x1_ASAP7_75t_L g128 ( 
.A(n_94),
.B(n_68),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_131),
.B(n_113),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_132),
.A2(n_105),
.B1(n_125),
.B2(n_102),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_116),
.A2(n_94),
.B(n_105),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_135),
.Y(n_150)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_114),
.Y(n_138)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_138),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_140),
.B(n_120),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_120),
.A2(n_109),
.B1(n_93),
.B2(n_99),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_141),
.A2(n_132),
.B1(n_130),
.B2(n_123),
.Y(n_152)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_118),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_142),
.B(n_146),
.Y(n_149)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_125),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_147),
.B(n_131),
.C(n_128),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_152),
.A2(n_140),
.B1(n_143),
.B2(n_147),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_153),
.B(n_141),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_148),
.B(n_124),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_154),
.B(n_156),
.Y(n_167)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_144),
.Y(n_155)
);

BUFx2_ASAP7_75t_L g166 ( 
.A(n_155),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_139),
.B(n_129),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_145),
.B(n_122),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_157),
.A2(n_159),
.B(n_144),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_158),
.A2(n_143),
.B1(n_134),
.B2(n_100),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_136),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_137),
.B(n_100),
.C(n_101),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_160),
.B(n_137),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_161),
.B(n_165),
.C(n_168),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_150),
.A2(n_135),
.B(n_133),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_162),
.A2(n_150),
.B(n_152),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_163),
.A2(n_160),
.B(n_168),
.Y(n_176)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_164),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_153),
.B(n_133),
.Y(n_165)
);

OR2x2_ASAP7_75t_L g172 ( 
.A(n_169),
.B(n_151),
.Y(n_172)
);

AOI21x1_ASAP7_75t_L g170 ( 
.A1(n_162),
.A2(n_149),
.B(n_158),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_170),
.B(n_176),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_172),
.B(n_175),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_173),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_166),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_174),
.A2(n_167),
.B(n_155),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_178),
.B(n_101),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_172),
.B(n_163),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_179),
.B(n_165),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_182),
.B(n_183),
.Y(n_186)
);

OR2x2_ASAP7_75t_L g183 ( 
.A(n_177),
.B(n_115),
.Y(n_183)
);

NAND5xp2_ASAP7_75t_L g184 ( 
.A(n_180),
.B(n_181),
.C(n_161),
.D(n_171),
.E(n_166),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_184),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_186),
.B(n_185),
.Y(n_188)
);

AOI322xp5_ASAP7_75t_L g190 ( 
.A1(n_188),
.A2(n_189),
.A3(n_110),
.B1(n_87),
.B2(n_88),
.C1(n_85),
.C2(n_84),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_187),
.B(n_171),
.C(n_180),
.Y(n_189)
);

AOI221xp5_ASAP7_75t_L g191 ( 
.A1(n_190),
.A2(n_84),
.B1(n_74),
.B2(n_85),
.C(n_87),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_191),
.B(n_85),
.Y(n_192)
);


endmodule