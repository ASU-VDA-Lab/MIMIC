module fake_jpeg_25393_n_121 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_121);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_121;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_14),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_17),
.B(n_36),
.Y(n_42)
);

BUFx4f_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_8),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_18),
.Y(n_47)
);

BUFx4f_ASAP7_75t_SL g48 ( 
.A(n_7),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_29),
.B(n_0),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_10),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_9),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g53 ( 
.A(n_48),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_53),
.B(n_44),
.Y(n_64)
);

HAxp5_ASAP7_75t_SL g54 ( 
.A(n_45),
.B(n_0),
.CON(n_54),
.SN(n_54)
);

A2O1A1Ixp33_ASAP7_75t_L g71 ( 
.A1(n_54),
.A2(n_38),
.B(n_52),
.C(n_3),
.Y(n_71)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_49),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_55),
.B(n_60),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_56),
.Y(n_61)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_57),
.Y(n_68)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_50),
.Y(n_58)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_58),
.Y(n_65)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_59),
.Y(n_66)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_56),
.B(n_51),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_62),
.B(n_72),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_58),
.A2(n_47),
.B1(n_46),
.B2(n_40),
.Y(n_63)
);

OA22x2_ASAP7_75t_L g81 ( 
.A1(n_63),
.A2(n_69),
.B1(n_71),
.B2(n_4),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_64),
.B(n_2),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_54),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_67),
.B(n_3),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_59),
.A2(n_51),
.B1(n_38),
.B2(n_39),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_55),
.B(n_1),
.Y(n_72)
);

BUFx10_ASAP7_75t_L g73 ( 
.A(n_56),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_74),
.A2(n_75),
.B1(n_81),
.B2(n_82),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_72),
.B(n_2),
.Y(n_75)
);

CKINVDCx14_ASAP7_75t_R g94 ( 
.A(n_76),
.Y(n_94)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_66),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_77),
.B(n_22),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_65),
.B(n_25),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_78),
.B(n_84),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g79 ( 
.A(n_64),
.B(n_26),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_79),
.B(n_15),
.C(n_16),
.Y(n_88)
);

AND2x4_ASAP7_75t_L g82 ( 
.A(n_68),
.B(n_4),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_70),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_83),
.B(n_85),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_73),
.B(n_5),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_61),
.Y(n_85)
);

OA22x2_ASAP7_75t_L g86 ( 
.A1(n_67),
.A2(n_6),
.B1(n_11),
.B2(n_13),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_86),
.B(n_24),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_62),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_87),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_88),
.B(n_97),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_80),
.B(n_20),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_89),
.B(n_28),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_90),
.B(n_33),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_78),
.B(n_23),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_92),
.B(n_30),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_93),
.B(n_86),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_98),
.B(n_99),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_93),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_95),
.B(n_82),
.Y(n_101)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_101),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_102),
.B(n_103),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_104),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_100),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_105),
.B(n_96),
.Y(n_113)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_104),
.Y(n_109)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_109),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_106),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_112),
.B(n_113),
.C(n_108),
.Y(n_114)
);

OA21x2_ASAP7_75t_SL g115 ( 
.A1(n_114),
.A2(n_110),
.B(n_111),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_SL g116 ( 
.A(n_115),
.B(n_91),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_116),
.A2(n_94),
.B(n_107),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_117),
.B(n_110),
.Y(n_118)
);

INVxp67_ASAP7_75t_SL g119 ( 
.A(n_118),
.Y(n_119)
);

AO21x1_ASAP7_75t_L g120 ( 
.A1(n_119),
.A2(n_34),
.B(n_35),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_120),
.B(n_37),
.Y(n_121)
);


endmodule