module real_jpeg_29653_n_6 (n_5, n_4, n_0, n_1, n_2, n_3, n_6);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_3;

output n_6;

wire n_17;
wire n_8;
wire n_21;
wire n_33;
wire n_35;
wire n_29;
wire n_10;
wire n_31;
wire n_9;
wire n_12;
wire n_24;
wire n_34;
wire n_28;
wire n_23;
wire n_11;
wire n_14;
wire n_25;
wire n_7;
wire n_22;
wire n_18;
wire n_26;
wire n_27;
wire n_20;
wire n_19;
wire n_32;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_0),
.B(n_13),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_1),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_1),
.B(n_21),
.Y(n_20)
);

INVx1_ASAP7_75t_SL g18 ( 
.A(n_2),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g23 ( 
.A(n_2),
.B(n_10),
.Y(n_23)
);

HAxp5_ASAP7_75t_SL g12 ( 
.A(n_3),
.B(n_13),
.CON(n_12),
.SN(n_12)
);

INVx1_ASAP7_75t_L g9 ( 
.A(n_4),
.Y(n_9)
);

OAI21xp33_ASAP7_75t_L g29 ( 
.A1(n_4),
.A2(n_11),
.B(n_30),
.Y(n_29)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_5),
.B(n_11),
.Y(n_30)
);

AOI221xp5_ASAP7_75t_L g6 ( 
.A1(n_7),
.A2(n_16),
.B1(n_24),
.B2(n_28),
.C(n_31),
.Y(n_6)
);

CKINVDCx20_ASAP7_75t_R g7 ( 
.A(n_8),
.Y(n_7)
);

OAI21xp5_ASAP7_75t_L g8 ( 
.A1(n_9),
.A2(n_10),
.B(n_14),
.Y(n_8)
);

AND2x2_ASAP7_75t_SL g33 ( 
.A(n_9),
.B(n_15),
.Y(n_33)
);

OR2x2_ASAP7_75t_SL g35 ( 
.A(n_9),
.B(n_15),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g14 ( 
.A(n_10),
.B(n_15),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_SL g27 ( 
.A(n_10),
.B(n_18),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_10),
.A2(n_11),
.B1(n_33),
.B2(n_34),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_11),
.Y(n_10)
);

CKINVDCx5p33_ASAP7_75t_R g11 ( 
.A(n_12),
.Y(n_11)
);

BUFx24_ASAP7_75t_SL g36 ( 
.A(n_12),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_23),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_19),
.Y(n_17)
);

AOI21xp5_ASAP7_75t_L g25 ( 
.A1(n_18),
.A2(n_26),
.B(n_27),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_19),
.Y(n_26)
);

OR2x2_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_22),
.Y(n_19)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_29),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_32),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_35),
.Y(n_34)
);


endmodule