module real_jpeg_11538_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_322, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_322;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx2_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx4f_ASAP7_75t_L g50 ( 
.A(n_1),
.Y(n_50)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_2),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_3),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_4),
.A2(n_44),
.B1(n_45),
.B2(n_47),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_4),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_4),
.A2(n_47),
.B1(n_61),
.B2(n_62),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_4),
.A2(n_31),
.B1(n_34),
.B2(n_47),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_4),
.A2(n_47),
.B1(n_73),
.B2(n_74),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_5),
.A2(n_73),
.B1(n_74),
.B2(n_134),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_5),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_5),
.A2(n_61),
.B1(n_62),
.B2(n_134),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_5),
.A2(n_44),
.B1(n_45),
.B2(n_134),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_L g228 ( 
.A1(n_5),
.A2(n_31),
.B1(n_34),
.B2(n_134),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_6),
.A2(n_44),
.B1(n_45),
.B2(n_55),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_6),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_6),
.A2(n_55),
.B1(n_61),
.B2(n_62),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_6),
.A2(n_31),
.B1(n_34),
.B2(n_55),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_6),
.A2(n_55),
.B1(n_73),
.B2(n_74),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_7),
.A2(n_31),
.B1(n_33),
.B2(n_34),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_7),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_7),
.A2(n_33),
.B1(n_73),
.B2(n_74),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_7),
.A2(n_33),
.B1(n_44),
.B2(n_45),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_7),
.A2(n_33),
.B1(n_61),
.B2(n_62),
.Y(n_130)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_8),
.Y(n_62)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_9),
.Y(n_58)
);

O2A1O1Ixp33_ASAP7_75t_L g146 ( 
.A1(n_10),
.A2(n_72),
.B(n_73),
.C(n_147),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_10),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_10),
.A2(n_73),
.B1(n_74),
.B2(n_148),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_10),
.B(n_83),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_10),
.A2(n_44),
.B1(n_45),
.B2(n_148),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_10),
.A2(n_101),
.B1(n_102),
.B2(n_236),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_10),
.B(n_89),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_11),
.A2(n_73),
.B1(n_74),
.B2(n_157),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_11),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_11),
.A2(n_61),
.B1(n_62),
.B2(n_157),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_11),
.A2(n_44),
.B1(n_45),
.B2(n_157),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_11),
.A2(n_31),
.B1(n_34),
.B2(n_157),
.Y(n_236)
);

BUFx8_ASAP7_75t_L g72 ( 
.A(n_12),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_13),
.A2(n_31),
.B1(n_34),
.B2(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_13),
.A2(n_38),
.B1(n_61),
.B2(n_62),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_13),
.A2(n_38),
.B1(n_44),
.B2(n_45),
.Y(n_96)
);

OAI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_13),
.A2(n_38),
.B1(n_73),
.B2(n_74),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_14),
.A2(n_73),
.B1(n_74),
.B2(n_81),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_14),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_14),
.A2(n_61),
.B1(n_62),
.B2(n_81),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_14),
.A2(n_44),
.B1(n_45),
.B2(n_81),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_14),
.A2(n_31),
.B1(n_34),
.B2(n_81),
.Y(n_230)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_314),
.Y(n_16)
);

AOI21xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_306),
.B(n_313),
.Y(n_17)
);

OAI21xp5_ASAP7_75t_SL g18 ( 
.A1(n_19),
.A2(n_272),
.B(n_303),
.Y(n_18)
);

AOI21xp5_ASAP7_75t_SL g19 ( 
.A1(n_20),
.A2(n_135),
.B(n_271),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_115),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_21),
.B(n_115),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_85),
.B2(n_114),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_22),
.B(n_86),
.C(n_98),
.Y(n_301)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_56),
.C(n_68),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_24),
.A2(n_25),
.B1(n_118),
.B2(n_119),
.Y(n_117)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_40),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_26),
.A2(n_27),
.B1(n_40),
.B2(n_41),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

AND2x2_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_35),
.Y(n_27)
);

OAI21xp5_ASAP7_75t_L g245 ( 
.A1(n_28),
.A2(n_101),
.B(n_230),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_30),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_29),
.B(n_34),
.Y(n_39)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_29),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_29),
.A2(n_39),
.B1(n_125),
.B2(n_144),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_29),
.A2(n_39),
.B1(n_227),
.B2(n_229),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_30),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_30),
.A2(n_39),
.B(n_127),
.Y(n_201)
);

CKINVDCx6p67_ASAP7_75t_R g34 ( 
.A(n_31),
.Y(n_34)
);

OA22x2_ASAP7_75t_L g52 ( 
.A1(n_31),
.A2(n_34),
.B1(n_50),
.B2(n_51),
.Y(n_52)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_34),
.B(n_51),
.C(n_148),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_34),
.B(n_234),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_35),
.A2(n_102),
.B(n_145),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_36),
.B(n_39),
.Y(n_35)
);

INVxp67_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_37),
.B(n_102),
.Y(n_127)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_39),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g40 ( 
.A(n_41),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_48),
.B1(n_53),
.B2(n_54),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_43),
.A2(n_52),
.B(n_94),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_44),
.A2(n_45),
.B1(n_50),
.B2(n_51),
.Y(n_49)
);

OA22x2_ASAP7_75t_SL g57 ( 
.A1(n_44),
.A2(n_45),
.B1(n_58),
.B2(n_59),
.Y(n_57)
);

O2A1O1Ixp33_ASAP7_75t_SL g197 ( 
.A1(n_44),
.A2(n_58),
.B(n_198),
.C(n_200),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_44),
.B(n_220),
.Y(n_219)
);

INVx6_ASAP7_75t_SL g44 ( 
.A(n_45),
.Y(n_44)
);

NOR3xp33_ASAP7_75t_L g200 ( 
.A(n_45),
.B(n_59),
.C(n_61),
.Y(n_200)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_48),
.B(n_95),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_48),
.A2(n_54),
.B(n_106),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_48),
.A2(n_93),
.B(n_106),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_48),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_48),
.A2(n_53),
.B1(n_205),
.B2(n_213),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_48),
.A2(n_53),
.B1(n_222),
.B2(n_223),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_48),
.A2(n_53),
.B1(n_213),
.B2(n_223),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_48),
.A2(n_53),
.B(n_93),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_52),
.Y(n_48)
);

INVx13_ASAP7_75t_L g51 ( 
.A(n_50),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_52),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_52),
.B(n_96),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_52),
.B(n_148),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_53),
.B(n_93),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_56),
.B(n_68),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_60),
.B(n_63),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_57),
.B(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_57),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_57),
.B(n_67),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_57),
.A2(n_152),
.B1(n_185),
.B2(n_187),
.Y(n_184)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_58),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_58),
.A2(n_59),
.B1(n_61),
.B2(n_62),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_60),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_61),
.A2(n_62),
.B1(n_72),
.B2(n_77),
.Y(n_78)
);

OAI21xp33_ASAP7_75t_L g147 ( 
.A1(n_61),
.A2(n_77),
.B(n_148),
.Y(n_147)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

HAxp5_ASAP7_75t_SL g199 ( 
.A(n_62),
.B(n_148),
.CON(n_199),
.SN(n_199)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_63),
.B(n_153),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_64),
.B(n_66),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_64),
.A2(n_88),
.B1(n_89),
.B2(n_90),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_64),
.A2(n_130),
.B(n_131),
.Y(n_129)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_64),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_64),
.A2(n_89),
.B1(n_151),
.B2(n_170),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_64),
.A2(n_89),
.B1(n_186),
.B2(n_199),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_SL g308 ( 
.A1(n_64),
.A2(n_89),
.B(n_130),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_SL g68 ( 
.A1(n_69),
.A2(n_79),
.B(n_82),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_69),
.A2(n_111),
.B(n_112),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_69),
.A2(n_78),
.B1(n_155),
.B2(n_158),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g309 ( 
.A1(n_69),
.A2(n_112),
.B(n_310),
.Y(n_309)
);

CKINVDCx14_ASAP7_75t_R g69 ( 
.A(n_70),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_70),
.A2(n_80),
.B1(n_83),
.B2(n_133),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_70),
.A2(n_83),
.B1(n_156),
.B2(n_172),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_70),
.B(n_113),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_70),
.A2(n_83),
.B1(n_294),
.B2(n_295),
.Y(n_293)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_78),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_72),
.A2(n_73),
.B1(n_74),
.B2(n_77),
.Y(n_71)
);

INVx11_ASAP7_75t_L g77 ( 
.A(n_72),
.Y(n_77)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx13_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_78),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_78),
.A2(n_285),
.B(n_286),
.Y(n_284)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_80),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_82),
.B(n_286),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_84),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_83),
.B(n_113),
.Y(n_112)
);

CKINVDCx14_ASAP7_75t_R g111 ( 
.A(n_84),
.Y(n_111)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_85),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_SL g85 ( 
.A(n_86),
.B(n_98),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_91),
.B(n_97),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_87),
.B(n_91),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_89),
.B(n_130),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_90),
.Y(n_280)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_94),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_92),
.A2(n_203),
.B(n_204),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_97),
.B(n_275),
.C(n_288),
.Y(n_274)
);

FAx1_ASAP7_75t_SL g302 ( 
.A(n_97),
.B(n_275),
.CI(n_288),
.CON(n_302),
.SN(n_302)
);

XOR2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_107),
.Y(n_98)
);

AOI21xp33_ASAP7_75t_L g288 ( 
.A1(n_99),
.A2(n_100),
.B(n_109),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_104),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_100),
.A2(n_108),
.B1(n_109),
.B2(n_110),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_100),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_100),
.A2(n_104),
.B1(n_105),
.B2(n_108),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_101),
.A2(n_102),
.B(n_103),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_101),
.A2(n_124),
.B(n_126),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_101),
.A2(n_102),
.B1(n_228),
.B2(n_236),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_102),
.B(n_148),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_120),
.C(n_121),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_116),
.A2(n_117),
.B1(n_120),
.B2(n_269),
.Y(n_268)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_120),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_121),
.B(n_268),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_129),
.C(n_132),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_122),
.B(n_162),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_128),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_123),
.B(n_128),
.Y(n_173)
);

CKINVDCx14_ASAP7_75t_R g124 ( 
.A(n_125),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_129),
.B(n_132),
.Y(n_162)
);

INVxp33_ASAP7_75t_L g281 ( 
.A(n_131),
.Y(n_281)
);

CKINVDCx14_ASAP7_75t_R g158 ( 
.A(n_133),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_265),
.B(n_270),
.Y(n_135)
);

AOI221xp5_ASAP7_75t_SL g136 ( 
.A1(n_137),
.A2(n_174),
.B1(n_190),
.B2(n_264),
.C(n_322),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_138),
.B(n_163),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_138),
.B(n_163),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_159),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_139),
.B(n_160),
.C(n_161),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_149),
.C(n_154),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_140),
.A2(n_141),
.B1(n_165),
.B2(n_166),
.Y(n_164)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_146),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_142),
.A2(n_143),
.B1(n_146),
.B2(n_179),
.Y(n_178)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

CKINVDCx14_ASAP7_75t_R g144 ( 
.A(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_146),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_SL g166 ( 
.A(n_149),
.B(n_154),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_150),
.A2(n_152),
.B(n_153),
.Y(n_149)
);

CKINVDCx14_ASAP7_75t_R g150 ( 
.A(n_151),
.Y(n_150)
);

OAI21xp33_ASAP7_75t_L g279 ( 
.A1(n_152),
.A2(n_280),
.B(n_281),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_161),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_167),
.C(n_173),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_164),
.B(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_167),
.B(n_173),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_169),
.C(n_171),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_168),
.B(n_169),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_170),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_171),
.B(n_177),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_188),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_175),
.B(n_188),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_178),
.C(n_180),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_176),
.B(n_260),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_178),
.B(n_180),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_182),
.C(n_184),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_181),
.A2(n_182),
.B1(n_183),
.B2(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_181),
.Y(n_208)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_SL g206 ( 
.A(n_184),
.B(n_207),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_263),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_192),
.A2(n_258),
.B(n_262),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_193),
.A2(n_214),
.B(n_257),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_194),
.B(n_209),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_194),
.B(n_209),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_206),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_202),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_196),
.B(n_202),
.C(n_206),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_201),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_SL g210 ( 
.A(n_197),
.B(n_201),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_199),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_211),
.C(n_212),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_210),
.B(n_254),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_211),
.B(n_212),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_215),
.A2(n_252),
.B(n_256),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_216),
.A2(n_242),
.B(n_251),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_217),
.A2(n_231),
.B(n_241),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_218),
.B(n_226),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_218),
.B(n_226),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_219),
.A2(n_221),
.B1(n_224),
.B2(n_225),
.Y(n_218)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_219),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_221),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_221),
.B(n_224),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g229 ( 
.A(n_230),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_232),
.A2(n_237),
.B(n_240),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_235),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_238),
.B(n_239),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_238),
.B(n_239),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_244),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_243),
.B(n_244),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_246),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_245),
.B(n_247),
.C(n_250),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_247),
.A2(n_248),
.B1(n_249),
.B2(n_250),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_249),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_253),
.B(n_255),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_253),
.B(n_255),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_259),
.B(n_261),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_259),
.B(n_261),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_267),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_266),
.B(n_267),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_273),
.B(n_300),
.Y(n_272)
);

AOI21xp33_ASAP7_75t_L g303 ( 
.A1(n_273),
.A2(n_304),
.B(n_305),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_289),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_274),
.B(n_289),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_276),
.A2(n_277),
.B1(n_284),
.B2(n_287),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_278),
.A2(n_279),
.B1(n_282),
.B2(n_283),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_278),
.B(n_283),
.C(n_284),
.Y(n_290)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_282),
.A2(n_283),
.B1(n_297),
.B2(n_298),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_282),
.B(n_293),
.C(n_298),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_283),
.Y(n_282)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_284),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_284),
.A2(n_287),
.B1(n_292),
.B2(n_299),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_284),
.B(n_290),
.C(n_299),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_285),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_291),
.Y(n_289)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_292),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_296),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_295),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_297),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_302),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_301),
.B(n_302),
.Y(n_304)
);

BUFx24_ASAP7_75t_SL g320 ( 
.A(n_302),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_312),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_307),
.B(n_312),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_307),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_307),
.B(n_317),
.Y(n_319)
);

FAx1_ASAP7_75t_SL g307 ( 
.A(n_308),
.B(n_309),
.CI(n_311),
.CON(n_307),
.SN(n_307)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_319),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_318),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_317),
.Y(n_316)
);


endmodule