module fake_ibex_1541_n_1018 (n_151, n_147, n_85, n_167, n_128, n_84, n_64, n_3, n_73, n_152, n_171, n_145, n_65, n_103, n_95, n_139, n_55, n_130, n_63, n_98, n_129, n_161, n_29, n_143, n_106, n_177, n_148, n_2, n_76, n_8, n_118, n_183, n_67, n_9, n_164, n_38, n_124, n_37, n_110, n_47, n_169, n_108, n_10, n_82, n_21, n_27, n_165, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_175, n_137, n_48, n_57, n_59, n_28, n_125, n_39, n_178, n_5, n_62, n_71, n_153, n_173, n_120, n_93, n_168, n_155, n_162, n_13, n_180, n_122, n_116, n_61, n_14, n_0, n_94, n_134, n_12, n_42, n_77, n_112, n_150, n_88, n_133, n_44, n_142, n_51, n_46, n_80, n_172, n_49, n_40, n_66, n_17, n_74, n_90, n_176, n_58, n_43, n_140, n_22, n_136, n_4, n_119, n_33, n_30, n_6, n_100, n_179, n_72, n_166, n_163, n_26, n_188, n_114, n_34, n_97, n_102, n_181, n_15, n_131, n_123, n_24, n_52, n_189, n_99, n_135, n_105, n_156, n_126, n_187, n_1, n_154, n_182, n_111, n_25, n_36, n_104, n_41, n_45, n_141, n_18, n_89, n_83, n_32, n_53, n_107, n_115, n_149, n_186, n_50, n_11, n_92, n_144, n_170, n_101, n_190, n_113, n_138, n_96, n_185, n_68, n_117, n_79, n_81, n_35, n_159, n_158, n_132, n_174, n_157, n_160, n_184, n_31, n_56, n_23, n_146, n_91, n_54, n_19, n_1018);

input n_151;
input n_147;
input n_85;
input n_167;
input n_128;
input n_84;
input n_64;
input n_3;
input n_73;
input n_152;
input n_171;
input n_145;
input n_65;
input n_103;
input n_95;
input n_139;
input n_55;
input n_130;
input n_63;
input n_98;
input n_129;
input n_161;
input n_29;
input n_143;
input n_106;
input n_177;
input n_148;
input n_2;
input n_76;
input n_8;
input n_118;
input n_183;
input n_67;
input n_9;
input n_164;
input n_38;
input n_124;
input n_37;
input n_110;
input n_47;
input n_169;
input n_108;
input n_10;
input n_82;
input n_21;
input n_27;
input n_165;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_175;
input n_137;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_178;
input n_5;
input n_62;
input n_71;
input n_153;
input n_173;
input n_120;
input n_93;
input n_168;
input n_155;
input n_162;
input n_13;
input n_180;
input n_122;
input n_116;
input n_61;
input n_14;
input n_0;
input n_94;
input n_134;
input n_12;
input n_42;
input n_77;
input n_112;
input n_150;
input n_88;
input n_133;
input n_44;
input n_142;
input n_51;
input n_46;
input n_80;
input n_172;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_176;
input n_58;
input n_43;
input n_140;
input n_22;
input n_136;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_179;
input n_72;
input n_166;
input n_163;
input n_26;
input n_188;
input n_114;
input n_34;
input n_97;
input n_102;
input n_181;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_189;
input n_99;
input n_135;
input n_105;
input n_156;
input n_126;
input n_187;
input n_1;
input n_154;
input n_182;
input n_111;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_141;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_107;
input n_115;
input n_149;
input n_186;
input n_50;
input n_11;
input n_92;
input n_144;
input n_170;
input n_101;
input n_190;
input n_113;
input n_138;
input n_96;
input n_185;
input n_68;
input n_117;
input n_79;
input n_81;
input n_35;
input n_159;
input n_158;
input n_132;
input n_174;
input n_157;
input n_160;
input n_184;
input n_31;
input n_56;
input n_23;
input n_146;
input n_91;
input n_54;
input n_19;

output n_1018;

wire n_599;
wire n_822;
wire n_778;
wire n_507;
wire n_743;
wire n_540;
wire n_754;
wire n_395;
wire n_1011;
wire n_992;
wire n_756;
wire n_529;
wire n_389;
wire n_204;
wire n_626;
wire n_274;
wire n_387;
wire n_766;
wire n_688;
wire n_946;
wire n_707;
wire n_273;
wire n_330;
wire n_309;
wire n_926;
wire n_328;
wire n_372;
wire n_341;
wire n_293;
wire n_256;
wire n_418;
wire n_193;
wire n_510;
wire n_845;
wire n_972;
wire n_981;
wire n_446;
wire n_350;
wire n_601;
wire n_621;
wire n_610;
wire n_956;
wire n_790;
wire n_920;
wire n_452;
wire n_664;
wire n_255;
wire n_586;
wire n_773;
wire n_994;
wire n_638;
wire n_398;
wire n_304;
wire n_821;
wire n_191;
wire n_873;
wire n_962;
wire n_593;
wire n_909;
wire n_545;
wire n_862;
wire n_583;
wire n_887;
wire n_957;
wire n_1015;
wire n_678;
wire n_663;
wire n_969;
wire n_194;
wire n_249;
wire n_334;
wire n_634;
wire n_733;
wire n_961;
wire n_991;
wire n_312;
wire n_622;
wire n_578;
wire n_478;
wire n_239;
wire n_432;
wire n_371;
wire n_974;
wire n_403;
wire n_872;
wire n_423;
wire n_608;
wire n_864;
wire n_357;
wire n_412;
wire n_457;
wire n_494;
wire n_226;
wire n_930;
wire n_336;
wire n_959;
wire n_258;
wire n_861;
wire n_449;
wire n_547;
wire n_727;
wire n_216;
wire n_996;
wire n_915;
wire n_911;
wire n_652;
wire n_781;
wire n_421;
wire n_828;
wire n_738;
wire n_475;
wire n_802;
wire n_753;
wire n_645;
wire n_500;
wire n_747;
wire n_963;
wire n_542;
wire n_236;
wire n_900;
wire n_376;
wire n_377;
wire n_584;
wire n_531;
wire n_647;
wire n_761;
wire n_556;
wire n_748;
wire n_498;
wire n_698;
wire n_280;
wire n_375;
wire n_340;
wire n_317;
wire n_708;
wire n_901;
wire n_667;
wire n_884;
wire n_682;
wire n_850;
wire n_196;
wire n_327;
wire n_326;
wire n_879;
wire n_723;
wire n_270;
wire n_346;
wire n_383;
wire n_886;
wire n_840;
wire n_1010;
wire n_561;
wire n_883;
wire n_417;
wire n_471;
wire n_846;
wire n_739;
wire n_755;
wire n_265;
wire n_853;
wire n_504;
wire n_948;
wire n_859;
wire n_259;
wire n_276;
wire n_339;
wire n_470;
wire n_770;
wire n_965;
wire n_210;
wire n_348;
wire n_220;
wire n_875;
wire n_941;
wire n_674;
wire n_481;
wire n_243;
wire n_287;
wire n_497;
wire n_671;
wire n_228;
wire n_711;
wire n_876;
wire n_552;
wire n_384;
wire n_251;
wire n_632;
wire n_989;
wire n_373;
wire n_854;
wire n_1008;
wire n_458;
wire n_244;
wire n_343;
wire n_310;
wire n_714;
wire n_936;
wire n_703;
wire n_426;
wire n_323;
wire n_469;
wire n_829;
wire n_598;
wire n_825;
wire n_740;
wire n_386;
wire n_549;
wire n_224;
wire n_533;
wire n_508;
wire n_939;
wire n_453;
wire n_591;
wire n_928;
wire n_655;
wire n_333;
wire n_898;
wire n_967;
wire n_306;
wire n_400;
wire n_550;
wire n_736;
wire n_732;
wire n_673;
wire n_798;
wire n_832;
wire n_278;
wire n_242;
wire n_316;
wire n_404;
wire n_557;
wire n_641;
wire n_527;
wire n_893;
wire n_590;
wire n_465;
wire n_325;
wire n_301;
wire n_496;
wire n_617;
wire n_434;
wire n_296;
wire n_690;
wire n_914;
wire n_1013;
wire n_982;
wire n_835;
wire n_526;
wire n_785;
wire n_824;
wire n_929;
wire n_315;
wire n_441;
wire n_604;
wire n_637;
wire n_523;
wire n_694;
wire n_787;
wire n_977;
wire n_614;
wire n_370;
wire n_431;
wire n_719;
wire n_574;
wire n_289;
wire n_716;
wire n_865;
wire n_923;
wire n_515;
wire n_642;
wire n_286;
wire n_321;
wire n_569;
wire n_600;
wire n_907;
wire n_933;
wire n_215;
wire n_279;
wire n_374;
wire n_235;
wire n_464;
wire n_538;
wire n_669;
wire n_838;
wire n_987;
wire n_750;
wire n_746;
wire n_261;
wire n_742;
wire n_521;
wire n_665;
wire n_459;
wire n_518;
wire n_367;
wire n_221;
wire n_852;
wire n_789;
wire n_880;
wire n_654;
wire n_656;
wire n_1014;
wire n_724;
wire n_437;
wire n_731;
wire n_602;
wire n_904;
wire n_842;
wire n_938;
wire n_355;
wire n_767;
wire n_474;
wire n_878;
wire n_758;
wire n_594;
wire n_636;
wire n_720;
wire n_710;
wire n_407;
wire n_490;
wire n_568;
wire n_813;
wire n_448;
wire n_646;
wire n_595;
wire n_466;
wire n_269;
wire n_944;
wire n_1001;
wire n_570;
wire n_623;
wire n_585;
wire n_715;
wire n_791;
wire n_530;
wire n_356;
wire n_543;
wire n_420;
wire n_483;
wire n_580;
wire n_487;
wire n_769;
wire n_222;
wire n_660;
wire n_524;
wire n_349;
wire n_765;
wire n_849;
wire n_857;
wire n_980;
wire n_454;
wire n_777;
wire n_1017;
wire n_295;
wire n_730;
wire n_331;
wire n_576;
wire n_230;
wire n_759;
wire n_917;
wire n_388;
wire n_953;
wire n_625;
wire n_968;
wire n_619;
wire n_536;
wire n_611;
wire n_352;
wire n_290;
wire n_558;
wire n_931;
wire n_666;
wire n_467;
wire n_427;
wire n_607;
wire n_827;
wire n_219;
wire n_246;
wire n_442;
wire n_207;
wire n_922;
wire n_438;
wire n_851;
wire n_993;
wire n_1012;
wire n_689;
wire n_960;
wire n_793;
wire n_676;
wire n_937;
wire n_253;
wire n_208;
wire n_234;
wire n_300;
wire n_973;
wire n_358;
wire n_771;
wire n_205;
wire n_618;
wire n_488;
wire n_514;
wire n_705;
wire n_999;
wire n_560;
wire n_429;
wire n_275;
wire n_541;
wire n_613;
wire n_659;
wire n_267;
wire n_662;
wire n_910;
wire n_1009;
wire n_635;
wire n_979;
wire n_844;
wire n_245;
wire n_589;
wire n_571;
wire n_229;
wire n_209;
wire n_472;
wire n_648;
wire n_783;
wire n_347;
wire n_847;
wire n_830;
wire n_1004;
wire n_473;
wire n_445;
wire n_629;
wire n_335;
wire n_413;
wire n_263;
wire n_573;
wire n_353;
wire n_966;
wire n_359;
wire n_826;
wire n_262;
wire n_299;
wire n_433;
wire n_439;
wire n_704;
wire n_949;
wire n_1007;
wire n_924;
wire n_643;
wire n_679;
wire n_841;
wire n_772;
wire n_810;
wire n_768;
wire n_839;
wire n_338;
wire n_696;
wire n_796;
wire n_797;
wire n_837;
wire n_477;
wire n_640;
wire n_954;
wire n_363;
wire n_1006;
wire n_402;
wire n_725;
wire n_369;
wire n_976;
wire n_596;
wire n_201;
wire n_699;
wire n_351;
wire n_368;
wire n_456;
wire n_834;
wire n_257;
wire n_998;
wire n_935;
wire n_869;
wire n_925;
wire n_718;
wire n_801;
wire n_918;
wire n_672;
wire n_722;
wire n_401;
wire n_554;
wire n_553;
wire n_735;
wire n_305;
wire n_882;
wire n_942;
wire n_713;
wire n_307;
wire n_192;
wire n_804;
wire n_484;
wire n_566;
wire n_480;
wire n_416;
wire n_581;
wire n_721;
wire n_365;
wire n_651;
wire n_814;
wire n_955;
wire n_605;
wire n_539;
wire n_354;
wire n_206;
wire n_392;
wire n_630;
wire n_567;
wire n_548;
wire n_516;
wire n_943;
wire n_763;
wire n_745;
wire n_329;
wire n_447;
wire n_940;
wire n_444;
wire n_200;
wire n_564;
wire n_506;
wire n_562;
wire n_868;
wire n_546;
wire n_199;
wire n_788;
wire n_795;
wire n_592;
wire n_986;
wire n_495;
wire n_762;
wire n_410;
wire n_905;
wire n_308;
wire n_975;
wire n_675;
wire n_800;
wire n_463;
wire n_624;
wire n_706;
wire n_411;
wire n_520;
wire n_784;
wire n_684;
wire n_775;
wire n_934;
wire n_927;
wire n_658;
wire n_512;
wire n_615;
wire n_950;
wire n_685;
wire n_397;
wire n_366;
wire n_283;
wire n_803;
wire n_894;
wire n_692;
wire n_627;
wire n_990;
wire n_709;
wire n_322;
wire n_227;
wire n_499;
wire n_888;
wire n_757;
wire n_248;
wire n_702;
wire n_451;
wire n_712;
wire n_971;
wire n_906;
wire n_650;
wire n_776;
wire n_409;
wire n_582;
wire n_978;
wire n_818;
wire n_653;
wire n_214;
wire n_238;
wire n_579;
wire n_843;
wire n_899;
wire n_902;
wire n_332;
wire n_799;
wire n_517;
wire n_211;
wire n_744;
wire n_817;
wire n_218;
wire n_314;
wire n_691;
wire n_563;
wire n_277;
wire n_555;
wire n_337;
wire n_522;
wire n_700;
wire n_479;
wire n_534;
wire n_225;
wire n_360;
wire n_881;
wire n_272;
wire n_951;
wire n_511;
wire n_734;
wire n_468;
wire n_223;
wire n_381;
wire n_525;
wire n_815;
wire n_919;
wire n_780;
wire n_535;
wire n_1002;
wire n_382;
wire n_502;
wire n_681;
wire n_633;
wire n_532;
wire n_726;
wire n_405;
wire n_863;
wire n_415;
wire n_597;
wire n_288;
wire n_285;
wire n_247;
wire n_379;
wire n_320;
wire n_551;
wire n_612;
wire n_318;
wire n_291;
wire n_819;
wire n_237;
wire n_203;
wire n_268;
wire n_440;
wire n_858;
wire n_342;
wire n_385;
wire n_414;
wire n_233;
wire n_430;
wire n_729;
wire n_741;
wire n_603;
wire n_378;
wire n_486;
wire n_952;
wire n_422;
wire n_264;
wire n_198;
wire n_616;
wire n_782;
wire n_997;
wire n_833;
wire n_217;
wire n_324;
wire n_391;
wire n_831;
wire n_537;
wire n_728;
wire n_805;
wire n_670;
wire n_820;
wire n_892;
wire n_390;
wire n_544;
wire n_891;
wire n_913;
wire n_509;
wire n_695;
wire n_786;
wire n_639;
wire n_303;
wire n_362;
wire n_717;
wire n_505;
wire n_482;
wire n_240;
wire n_1016;
wire n_282;
wire n_680;
wire n_501;
wire n_809;
wire n_752;
wire n_856;
wire n_668;
wire n_779;
wire n_871;
wire n_266;
wire n_294;
wire n_866;
wire n_958;
wire n_485;
wire n_870;
wire n_284;
wire n_811;
wire n_808;
wire n_250;
wire n_945;
wire n_493;
wire n_460;
wire n_609;
wire n_476;
wire n_792;
wire n_461;
wire n_575;
wire n_313;
wire n_903;
wire n_519;
wire n_345;
wire n_408;
wire n_361;
wire n_455;
wire n_419;
wire n_774;
wire n_319;
wire n_195;
wire n_885;
wire n_513;
wire n_212;
wire n_588;
wire n_877;
wire n_693;
wire n_311;
wire n_860;
wire n_661;
wire n_848;
wire n_406;
wire n_606;
wire n_737;
wire n_896;
wire n_197;
wire n_528;
wire n_1005;
wire n_631;
wire n_683;
wire n_260;
wire n_620;
wire n_794;
wire n_836;
wire n_462;
wire n_302;
wire n_450;
wire n_443;
wire n_686;
wire n_985;
wire n_572;
wire n_867;
wire n_983;
wire n_1003;
wire n_644;
wire n_577;
wire n_344;
wire n_393;
wire n_889;
wire n_897;
wire n_436;
wire n_428;
wire n_970;
wire n_491;
wire n_297;
wire n_435;
wire n_628;
wire n_252;
wire n_396;
wire n_697;
wire n_816;
wire n_874;
wire n_912;
wire n_890;
wire n_921;
wire n_489;
wire n_677;
wire n_399;
wire n_254;
wire n_908;
wire n_213;
wire n_964;
wire n_565;
wire n_424;
wire n_916;
wire n_823;
wire n_701;
wire n_271;
wire n_995;
wire n_241;
wire n_503;
wire n_292;
wire n_807;
wire n_1000;
wire n_394;
wire n_984;
wire n_364;
wire n_687;
wire n_895;
wire n_988;
wire n_202;
wire n_231;
wire n_298;
wire n_587;
wire n_760;
wire n_751;
wire n_806;
wire n_932;
wire n_657;
wire n_764;
wire n_492;
wire n_649;
wire n_812;
wire n_855;
wire n_232;
wire n_380;
wire n_749;
wire n_281;
wire n_947;
wire n_559;
wire n_425;

INVx1_ASAP7_75t_L g191 ( 
.A(n_67),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_137),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_48),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_84),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_14),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_44),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_50),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g198 ( 
.A(n_153),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_180),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_56),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_100),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_105),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_4),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_80),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_73),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_59),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_176),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_79),
.Y(n_208)
);

BUFx3_ASAP7_75t_L g209 ( 
.A(n_186),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_179),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_38),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_89),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_125),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_54),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_113),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_143),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_21),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_40),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_51),
.Y(n_219)
);

BUFx3_ASAP7_75t_L g220 ( 
.A(n_102),
.Y(n_220)
);

NOR2xp67_ASAP7_75t_L g221 ( 
.A(n_126),
.B(n_2),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_101),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_158),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_38),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_31),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_4),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_182),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_74),
.Y(n_228)
);

INVxp67_ASAP7_75t_SL g229 ( 
.A(n_86),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_41),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_160),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_97),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_106),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_18),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_166),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_69),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g237 ( 
.A(n_161),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_124),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_81),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_8),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_15),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_95),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_30),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_149),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_173),
.Y(n_245)
);

CKINVDCx16_ASAP7_75t_R g246 ( 
.A(n_60),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_52),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_1),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_13),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_178),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_94),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_128),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_111),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_58),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_15),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_16),
.Y(n_256)
);

INVxp67_ASAP7_75t_SL g257 ( 
.A(n_107),
.Y(n_257)
);

BUFx3_ASAP7_75t_L g258 ( 
.A(n_99),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_22),
.Y(n_259)
);

OR2x2_ASAP7_75t_L g260 ( 
.A(n_162),
.B(n_40),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_12),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_145),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_68),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_148),
.Y(n_264)
);

NOR2xp67_ASAP7_75t_L g265 ( 
.A(n_35),
.B(n_189),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_114),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_157),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_108),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_72),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_39),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_117),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_168),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_66),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_53),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_92),
.Y(n_275)
);

BUFx3_ASAP7_75t_L g276 ( 
.A(n_0),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_78),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_13),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_12),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_64),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_6),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_151),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_144),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_75),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_109),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_23),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_120),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_20),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_110),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_133),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_122),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_65),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_45),
.Y(n_293)
);

INVx1_ASAP7_75t_SL g294 ( 
.A(n_121),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_35),
.Y(n_295)
);

NOR2xp67_ASAP7_75t_L g296 ( 
.A(n_187),
.B(n_116),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_19),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_115),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_88),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_163),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_188),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_131),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_47),
.Y(n_303)
);

BUFx5_ASAP7_75t_L g304 ( 
.A(n_190),
.Y(n_304)
);

BUFx3_ASAP7_75t_L g305 ( 
.A(n_150),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_156),
.Y(n_306)
);

BUFx6f_ASAP7_75t_L g307 ( 
.A(n_170),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_5),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_98),
.Y(n_309)
);

INVx3_ASAP7_75t_L g310 ( 
.A(n_16),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_129),
.Y(n_311)
);

INVxp33_ASAP7_75t_SL g312 ( 
.A(n_175),
.Y(n_312)
);

HB1xp67_ASAP7_75t_L g313 ( 
.A(n_310),
.Y(n_313)
);

INVx5_ASAP7_75t_L g314 ( 
.A(n_307),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_198),
.Y(n_315)
);

BUFx6f_ASAP7_75t_L g316 ( 
.A(n_307),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_237),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_246),
.Y(n_318)
);

BUFx3_ASAP7_75t_L g319 ( 
.A(n_209),
.Y(n_319)
);

BUFx6f_ASAP7_75t_L g320 ( 
.A(n_307),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_244),
.Y(n_321)
);

BUFx6f_ASAP7_75t_L g322 ( 
.A(n_307),
.Y(n_322)
);

INVx4_ASAP7_75t_L g323 ( 
.A(n_209),
.Y(n_323)
);

BUFx6f_ASAP7_75t_L g324 ( 
.A(n_220),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_304),
.Y(n_325)
);

BUFx3_ASAP7_75t_L g326 ( 
.A(n_220),
.Y(n_326)
);

AND2x4_ASAP7_75t_L g327 ( 
.A(n_310),
.B(n_3),
.Y(n_327)
);

BUFx3_ASAP7_75t_L g328 ( 
.A(n_258),
.Y(n_328)
);

INVx6_ASAP7_75t_L g329 ( 
.A(n_304),
.Y(n_329)
);

AND2x4_ASAP7_75t_L g330 ( 
.A(n_310),
.B(n_3),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_304),
.B(n_5),
.Y(n_331)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_276),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_304),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_276),
.Y(n_334)
);

OA21x2_ASAP7_75t_L g335 ( 
.A1(n_199),
.A2(n_215),
.B(n_207),
.Y(n_335)
);

BUFx6f_ASAP7_75t_L g336 ( 
.A(n_258),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_304),
.B(n_6),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_195),
.B(n_203),
.Y(n_338)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_304),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_224),
.Y(n_340)
);

HB1xp67_ASAP7_75t_L g341 ( 
.A(n_225),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_191),
.B(n_7),
.Y(n_342)
);

BUFx6f_ASAP7_75t_L g343 ( 
.A(n_305),
.Y(n_343)
);

BUFx6f_ASAP7_75t_L g344 ( 
.A(n_305),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_304),
.Y(n_345)
);

BUFx6f_ASAP7_75t_L g346 ( 
.A(n_199),
.Y(n_346)
);

NOR2x1_ASAP7_75t_L g347 ( 
.A(n_224),
.B(n_42),
.Y(n_347)
);

INVx2_ASAP7_75t_SL g348 ( 
.A(n_207),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_256),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_256),
.Y(n_350)
);

BUFx3_ASAP7_75t_L g351 ( 
.A(n_215),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_211),
.B(n_7),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_244),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_217),
.B(n_8),
.Y(n_354)
);

BUFx6f_ASAP7_75t_L g355 ( 
.A(n_226),
.Y(n_355)
);

NAND2xp33_ASAP7_75t_L g356 ( 
.A(n_226),
.B(n_43),
.Y(n_356)
);

INVx2_ASAP7_75t_SL g357 ( 
.A(n_222),
.Y(n_357)
);

AND2x2_ASAP7_75t_L g358 ( 
.A(n_218),
.B(n_9),
.Y(n_358)
);

AND2x2_ASAP7_75t_L g359 ( 
.A(n_234),
.B(n_9),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_222),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_228),
.Y(n_361)
);

BUFx6f_ASAP7_75t_L g362 ( 
.A(n_228),
.Y(n_362)
);

BUFx8_ASAP7_75t_L g363 ( 
.A(n_260),
.Y(n_363)
);

AND2x4_ASAP7_75t_L g364 ( 
.A(n_231),
.B(n_10),
.Y(n_364)
);

INVx4_ASAP7_75t_L g365 ( 
.A(n_193),
.Y(n_365)
);

AND2x4_ASAP7_75t_L g366 ( 
.A(n_250),
.B(n_10),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_249),
.B(n_11),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_250),
.Y(n_368)
);

HB1xp67_ASAP7_75t_L g369 ( 
.A(n_240),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_267),
.Y(n_370)
);

HB1xp67_ASAP7_75t_L g371 ( 
.A(n_241),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_245),
.Y(n_372)
);

BUFx2_ASAP7_75t_L g373 ( 
.A(n_243),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_255),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_259),
.Y(n_375)
);

AND2x4_ASAP7_75t_L g376 ( 
.A(n_268),
.B(n_11),
.Y(n_376)
);

BUFx6f_ASAP7_75t_L g377 ( 
.A(n_268),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_261),
.Y(n_378)
);

INVx3_ASAP7_75t_L g379 ( 
.A(n_226),
.Y(n_379)
);

INVx6_ASAP7_75t_L g380 ( 
.A(n_226),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_270),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_290),
.Y(n_382)
);

HB1xp67_ASAP7_75t_L g383 ( 
.A(n_248),
.Y(n_383)
);

INVx3_ASAP7_75t_L g384 ( 
.A(n_281),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_290),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_SL g386 ( 
.A1(n_279),
.A2(n_14),
.B1(n_17),
.B2(n_18),
.Y(n_386)
);

INVx6_ASAP7_75t_L g387 ( 
.A(n_223),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_300),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_327),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_315),
.Y(n_390)
);

AND2x2_ASAP7_75t_L g391 ( 
.A(n_313),
.B(n_200),
.Y(n_391)
);

BUFx6f_ASAP7_75t_L g392 ( 
.A(n_316),
.Y(n_392)
);

BUFx10_ASAP7_75t_L g393 ( 
.A(n_315),
.Y(n_393)
);

AO22x2_ASAP7_75t_L g394 ( 
.A1(n_327),
.A2(n_286),
.B1(n_295),
.B2(n_311),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_387),
.B(n_247),
.Y(n_395)
);

AND2x2_ASAP7_75t_L g396 ( 
.A(n_373),
.B(n_201),
.Y(n_396)
);

BUFx3_ASAP7_75t_L g397 ( 
.A(n_319),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_365),
.B(n_201),
.Y(n_398)
);

INVx2_ASAP7_75t_SL g399 ( 
.A(n_387),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_387),
.B(n_300),
.Y(n_400)
);

AND2x6_ASAP7_75t_L g401 ( 
.A(n_330),
.B(n_192),
.Y(n_401)
);

INVx3_ASAP7_75t_L g402 ( 
.A(n_330),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_365),
.B(n_332),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_346),
.Y(n_404)
);

INVx4_ASAP7_75t_L g405 ( 
.A(n_330),
.Y(n_405)
);

BUFx3_ASAP7_75t_L g406 ( 
.A(n_319),
.Y(n_406)
);

INVx3_ASAP7_75t_L g407 ( 
.A(n_364),
.Y(n_407)
);

BUFx10_ASAP7_75t_L g408 ( 
.A(n_318),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_346),
.Y(n_409)
);

AND2x2_ASAP7_75t_L g410 ( 
.A(n_341),
.B(n_202),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_364),
.Y(n_411)
);

BUFx4f_ASAP7_75t_L g412 ( 
.A(n_364),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_SL g413 ( 
.A(n_366),
.B(n_196),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_SL g414 ( 
.A(n_366),
.B(n_376),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_366),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_321),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_323),
.B(n_202),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_376),
.Y(n_418)
);

INVxp67_ASAP7_75t_L g419 ( 
.A(n_369),
.Y(n_419)
);

BUFx3_ASAP7_75t_L g420 ( 
.A(n_326),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_323),
.B(n_204),
.Y(n_421)
);

INVx4_ASAP7_75t_L g422 ( 
.A(n_329),
.Y(n_422)
);

INVx2_ASAP7_75t_SL g423 ( 
.A(n_371),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_362),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_376),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_323),
.B(n_204),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_326),
.B(n_205),
.Y(n_427)
);

AND2x6_ASAP7_75t_L g428 ( 
.A(n_347),
.B(n_197),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_362),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_334),
.Y(n_430)
);

BUFx3_ASAP7_75t_L g431 ( 
.A(n_328),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_377),
.Y(n_432)
);

OAI21xp33_ASAP7_75t_SL g433 ( 
.A1(n_348),
.A2(n_265),
.B(n_221),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_377),
.Y(n_434)
);

BUFx3_ASAP7_75t_L g435 ( 
.A(n_335),
.Y(n_435)
);

AND2x2_ASAP7_75t_L g436 ( 
.A(n_383),
.B(n_280),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_384),
.B(n_206),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_318),
.A2(n_312),
.B1(n_245),
.B2(n_289),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_358),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_374),
.B(n_208),
.Y(n_440)
);

INVx3_ASAP7_75t_L g441 ( 
.A(n_351),
.Y(n_441)
);

INVx3_ASAP7_75t_L g442 ( 
.A(n_351),
.Y(n_442)
);

BUFx6f_ASAP7_75t_L g443 ( 
.A(n_316),
.Y(n_443)
);

INVx3_ASAP7_75t_L g444 ( 
.A(n_360),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_358),
.Y(n_445)
);

AND2x2_ASAP7_75t_L g446 ( 
.A(n_375),
.B(n_301),
.Y(n_446)
);

BUFx10_ASAP7_75t_L g447 ( 
.A(n_329),
.Y(n_447)
);

INVx1_ASAP7_75t_SL g448 ( 
.A(n_321),
.Y(n_448)
);

HB1xp67_ASAP7_75t_L g449 ( 
.A(n_359),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_377),
.Y(n_450)
);

OR2x2_ASAP7_75t_L g451 ( 
.A(n_338),
.B(n_278),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_357),
.B(n_301),
.Y(n_452)
);

AOI22xp33_ASAP7_75t_L g453 ( 
.A1(n_359),
.A2(n_335),
.B1(n_361),
.B2(n_360),
.Y(n_453)
);

INVx3_ASAP7_75t_L g454 ( 
.A(n_361),
.Y(n_454)
);

BUFx6f_ASAP7_75t_L g455 ( 
.A(n_316),
.Y(n_455)
);

INVxp67_ASAP7_75t_R g456 ( 
.A(n_386),
.Y(n_456)
);

NAND2xp33_ASAP7_75t_L g457 ( 
.A(n_325),
.B(n_303),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_378),
.B(n_210),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_368),
.Y(n_459)
);

BUFx10_ASAP7_75t_L g460 ( 
.A(n_329),
.Y(n_460)
);

BUFx6f_ASAP7_75t_SL g461 ( 
.A(n_381),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_333),
.B(n_339),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_368),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_335),
.Y(n_464)
);

INVx2_ASAP7_75t_SL g465 ( 
.A(n_329),
.Y(n_465)
);

OR2x6_ASAP7_75t_L g466 ( 
.A(n_352),
.B(n_279),
.Y(n_466)
);

BUFx2_ASAP7_75t_L g467 ( 
.A(n_363),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_324),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_370),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_340),
.B(n_212),
.Y(n_470)
);

INVx4_ASAP7_75t_L g471 ( 
.A(n_324),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_370),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_349),
.B(n_213),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_350),
.B(n_306),
.Y(n_474)
);

CKINVDCx20_ASAP7_75t_R g475 ( 
.A(n_353),
.Y(n_475)
);

BUFx10_ASAP7_75t_L g476 ( 
.A(n_342),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_388),
.B(n_214),
.Y(n_477)
);

OAI22xp5_ASAP7_75t_L g478 ( 
.A1(n_317),
.A2(n_289),
.B1(n_252),
.B2(n_297),
.Y(n_478)
);

BUFx3_ASAP7_75t_L g479 ( 
.A(n_324),
.Y(n_479)
);

INVx2_ASAP7_75t_SL g480 ( 
.A(n_363),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_324),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_382),
.B(n_385),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_446),
.B(n_363),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_403),
.B(n_354),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_SL g485 ( 
.A(n_467),
.B(n_252),
.Y(n_485)
);

AOI21xp5_ASAP7_75t_L g486 ( 
.A1(n_464),
.A2(n_356),
.B(n_339),
.Y(n_486)
);

HB1xp67_ASAP7_75t_L g487 ( 
.A(n_449),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_397),
.Y(n_488)
);

AND2x2_ASAP7_75t_L g489 ( 
.A(n_391),
.B(n_449),
.Y(n_489)
);

AOI22xp5_ASAP7_75t_L g490 ( 
.A1(n_394),
.A2(n_288),
.B1(n_312),
.B2(n_367),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_397),
.Y(n_491)
);

O2A1O1Ixp5_ASAP7_75t_L g492 ( 
.A1(n_464),
.A2(n_337),
.B(n_331),
.C(n_333),
.Y(n_492)
);

OR2x2_ASAP7_75t_L g493 ( 
.A(n_419),
.B(n_353),
.Y(n_493)
);

AND2x2_ASAP7_75t_L g494 ( 
.A(n_396),
.B(n_451),
.Y(n_494)
);

AND2x4_ASAP7_75t_L g495 ( 
.A(n_480),
.B(n_382),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_441),
.Y(n_496)
);

OAI22xp33_ASAP7_75t_L g497 ( 
.A1(n_456),
.A2(n_308),
.B1(n_372),
.B2(n_388),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_442),
.B(n_194),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_398),
.B(n_219),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_SL g500 ( 
.A(n_412),
.B(n_238),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_395),
.B(n_385),
.Y(n_501)
);

OR2x2_ASAP7_75t_L g502 ( 
.A(n_466),
.B(n_372),
.Y(n_502)
);

NAND2xp33_ASAP7_75t_L g503 ( 
.A(n_401),
.B(n_239),
.Y(n_503)
);

O2A1O1Ixp33_ASAP7_75t_L g504 ( 
.A1(n_414),
.A2(n_345),
.B(n_356),
.C(n_275),
.Y(n_504)
);

AOI22xp33_ASAP7_75t_L g505 ( 
.A1(n_407),
.A2(n_345),
.B1(n_343),
.B2(n_344),
.Y(n_505)
);

OAI22xp5_ASAP7_75t_SL g506 ( 
.A1(n_475),
.A2(n_308),
.B1(n_257),
.B2(n_229),
.Y(n_506)
);

AOI22xp33_ASAP7_75t_L g507 ( 
.A1(n_407),
.A2(n_336),
.B1(n_343),
.B2(n_344),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_474),
.B(n_251),
.Y(n_508)
);

INVx8_ASAP7_75t_L g509 ( 
.A(n_401),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_SL g510 ( 
.A(n_412),
.B(n_264),
.Y(n_510)
);

NOR2x1p5_ASAP7_75t_L g511 ( 
.A(n_390),
.B(n_266),
.Y(n_511)
);

AOI21xp5_ASAP7_75t_L g512 ( 
.A1(n_414),
.A2(n_227),
.B(n_216),
.Y(n_512)
);

O2A1O1Ixp33_ASAP7_75t_L g513 ( 
.A1(n_439),
.A2(n_230),
.B(n_232),
.C(n_233),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_406),
.Y(n_514)
);

NAND2xp33_ASAP7_75t_L g515 ( 
.A(n_401),
.B(n_269),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_420),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_SL g517 ( 
.A(n_405),
.B(n_272),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_399),
.B(n_235),
.Y(n_518)
);

AOI22xp5_ASAP7_75t_L g519 ( 
.A1(n_394),
.A2(n_287),
.B1(n_242),
.B2(n_253),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_427),
.B(n_274),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_445),
.B(n_236),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_452),
.B(n_254),
.Y(n_522)
);

INVx4_ASAP7_75t_L g523 ( 
.A(n_461),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_420),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_431),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_402),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_431),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_402),
.Y(n_528)
);

AND2x2_ASAP7_75t_L g529 ( 
.A(n_410),
.B(n_294),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_436),
.B(n_284),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_475),
.Y(n_531)
);

NAND2x1p5_ASAP7_75t_L g532 ( 
.A(n_423),
.B(n_389),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_417),
.B(n_285),
.Y(n_533)
);

AOI21xp5_ASAP7_75t_L g534 ( 
.A1(n_413),
.A2(n_263),
.B(n_262),
.Y(n_534)
);

AOI22xp33_ASAP7_75t_L g535 ( 
.A1(n_411),
.A2(n_336),
.B1(n_343),
.B2(n_344),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_430),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_421),
.B(n_291),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_476),
.B(n_271),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_L g539 ( 
.A(n_476),
.B(n_273),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_479),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_426),
.B(n_292),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_413),
.B(n_298),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_479),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_SL g544 ( 
.A(n_447),
.B(n_309),
.Y(n_544)
);

OR2x6_ASAP7_75t_L g545 ( 
.A(n_466),
.B(n_296),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_415),
.B(n_277),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_418),
.B(n_282),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_425),
.B(n_283),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_L g549 ( 
.A(n_440),
.B(n_293),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_437),
.B(n_400),
.Y(n_550)
);

NOR3xp33_ASAP7_75t_L g551 ( 
.A(n_478),
.B(n_299),
.C(n_302),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_444),
.Y(n_552)
);

INVx2_ASAP7_75t_SL g553 ( 
.A(n_394),
.Y(n_553)
);

INVx2_ASAP7_75t_SL g554 ( 
.A(n_393),
.Y(n_554)
);

AOI22xp5_ASAP7_75t_L g555 ( 
.A1(n_457),
.A2(n_336),
.B1(n_343),
.B2(n_344),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_440),
.B(n_379),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_458),
.B(n_379),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_458),
.B(n_379),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_SL g559 ( 
.A(n_447),
.B(n_314),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_433),
.B(n_470),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_453),
.B(n_428),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_428),
.B(n_314),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_454),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_459),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_463),
.Y(n_565)
);

HB1xp67_ASAP7_75t_L g566 ( 
.A(n_435),
.Y(n_566)
);

OR2x2_ASAP7_75t_L g567 ( 
.A(n_466),
.B(n_17),
.Y(n_567)
);

A2O1A1Ixp33_ASAP7_75t_SL g568 ( 
.A1(n_477),
.A2(n_473),
.B(n_470),
.C(n_482),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_454),
.B(n_380),
.Y(n_569)
);

AND2x4_ASAP7_75t_L g570 ( 
.A(n_523),
.B(n_448),
.Y(n_570)
);

BUFx2_ASAP7_75t_L g571 ( 
.A(n_531),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_526),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_484),
.B(n_473),
.Y(n_573)
);

NOR2xp67_ASAP7_75t_SL g574 ( 
.A(n_566),
.B(n_390),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_494),
.B(n_469),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_528),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_560),
.B(n_472),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_552),
.Y(n_578)
);

OAI22xp5_ASAP7_75t_L g579 ( 
.A1(n_509),
.A2(n_438),
.B1(n_416),
.B2(n_477),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_560),
.B(n_482),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_487),
.B(n_393),
.Y(n_581)
);

AO22x1_ASAP7_75t_L g582 ( 
.A1(n_523),
.A2(n_408),
.B1(n_422),
.B2(n_471),
.Y(n_582)
);

INVx3_ASAP7_75t_L g583 ( 
.A(n_509),
.Y(n_583)
);

O2A1O1Ixp33_ASAP7_75t_L g584 ( 
.A1(n_568),
.A2(n_462),
.B(n_465),
.C(n_468),
.Y(n_584)
);

AND2x2_ASAP7_75t_L g585 ( 
.A(n_487),
.B(n_408),
.Y(n_585)
);

AND2x2_ASAP7_75t_L g586 ( 
.A(n_489),
.B(n_460),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_529),
.B(n_471),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_SL g588 ( 
.A(n_566),
.B(n_468),
.Y(n_588)
);

AOI21xp5_ASAP7_75t_L g589 ( 
.A1(n_486),
.A2(n_568),
.B(n_550),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_536),
.B(n_19),
.Y(n_590)
);

BUFx3_ASAP7_75t_L g591 ( 
.A(n_554),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_L g592 ( 
.A(n_483),
.B(n_20),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_L g593 ( 
.A(n_532),
.B(n_21),
.Y(n_593)
);

OAI21xp5_ASAP7_75t_L g594 ( 
.A1(n_492),
.A2(n_429),
.B(n_404),
.Y(n_594)
);

AOI21xp5_ASAP7_75t_L g595 ( 
.A1(n_561),
.A2(n_429),
.B(n_409),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_495),
.B(n_22),
.Y(n_596)
);

AND2x2_ASAP7_75t_L g597 ( 
.A(n_485),
.B(n_23),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_495),
.B(n_24),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_549),
.B(n_24),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_549),
.B(n_25),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_532),
.B(n_25),
.Y(n_601)
);

CKINVDCx16_ASAP7_75t_R g602 ( 
.A(n_493),
.Y(n_602)
);

CKINVDCx8_ASAP7_75t_R g603 ( 
.A(n_545),
.Y(n_603)
);

NAND2x1p5_ASAP7_75t_L g604 ( 
.A(n_519),
.B(n_567),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_564),
.Y(n_605)
);

OAI22xp5_ASAP7_75t_L g606 ( 
.A1(n_490),
.A2(n_380),
.B1(n_481),
.B2(n_450),
.Y(n_606)
);

OR2x2_ASAP7_75t_L g607 ( 
.A(n_502),
.B(n_26),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_522),
.B(n_538),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_563),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_522),
.B(n_27),
.Y(n_610)
);

AOI21xp5_ASAP7_75t_L g611 ( 
.A1(n_512),
.A2(n_548),
.B(n_547),
.Y(n_611)
);

CKINVDCx20_ASAP7_75t_R g612 ( 
.A(n_506),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_565),
.Y(n_613)
);

AOI21xp5_ASAP7_75t_L g614 ( 
.A1(n_533),
.A2(n_424),
.B(n_432),
.Y(n_614)
);

O2A1O1Ixp33_ASAP7_75t_L g615 ( 
.A1(n_551),
.A2(n_434),
.B(n_29),
.C(n_30),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_539),
.B(n_28),
.Y(n_616)
);

AOI21xp5_ASAP7_75t_L g617 ( 
.A1(n_537),
.A2(n_455),
.B(n_443),
.Y(n_617)
);

AOI21xp5_ASAP7_75t_L g618 ( 
.A1(n_541),
.A2(n_499),
.B(n_508),
.Y(n_618)
);

BUFx6f_ASAP7_75t_L g619 ( 
.A(n_488),
.Y(n_619)
);

OAI22xp5_ASAP7_75t_L g620 ( 
.A1(n_521),
.A2(n_355),
.B1(n_320),
.B2(n_322),
.Y(n_620)
);

BUFx2_ASAP7_75t_L g621 ( 
.A(n_545),
.Y(n_621)
);

AOI21xp5_ASAP7_75t_L g622 ( 
.A1(n_520),
.A2(n_455),
.B(n_443),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_521),
.B(n_29),
.Y(n_623)
);

NAND2x1p5_ASAP7_75t_L g624 ( 
.A(n_496),
.B(n_517),
.Y(n_624)
);

O2A1O1Ixp33_ASAP7_75t_L g625 ( 
.A1(n_551),
.A2(n_31),
.B(n_32),
.C(n_33),
.Y(n_625)
);

AOI22xp5_ASAP7_75t_L g626 ( 
.A1(n_546),
.A2(n_355),
.B1(n_322),
.B2(n_320),
.Y(n_626)
);

AND2x4_ASAP7_75t_L g627 ( 
.A(n_511),
.B(n_32),
.Y(n_627)
);

BUFx6f_ASAP7_75t_L g628 ( 
.A(n_491),
.Y(n_628)
);

NAND3xp33_ASAP7_75t_L g629 ( 
.A(n_513),
.B(n_355),
.C(n_322),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_546),
.B(n_33),
.Y(n_630)
);

INVx4_ASAP7_75t_L g631 ( 
.A(n_545),
.Y(n_631)
);

BUFx6f_ASAP7_75t_L g632 ( 
.A(n_514),
.Y(n_632)
);

AO22x1_ASAP7_75t_L g633 ( 
.A1(n_497),
.A2(n_34),
.B1(n_36),
.B2(n_37),
.Y(n_633)
);

NOR2xp33_ASAP7_75t_L g634 ( 
.A(n_530),
.B(n_36),
.Y(n_634)
);

OAI21xp33_ASAP7_75t_SL g635 ( 
.A1(n_501),
.A2(n_37),
.B(n_39),
.Y(n_635)
);

INVx4_ASAP7_75t_L g636 ( 
.A(n_516),
.Y(n_636)
);

AOI22xp33_ASAP7_75t_L g637 ( 
.A1(n_518),
.A2(n_322),
.B1(n_320),
.B2(n_316),
.Y(n_637)
);

OAI21xp5_ASAP7_75t_L g638 ( 
.A1(n_504),
.A2(n_392),
.B(n_322),
.Y(n_638)
);

AOI21xp5_ASAP7_75t_L g639 ( 
.A1(n_542),
.A2(n_392),
.B(n_320),
.Y(n_639)
);

BUFx6f_ASAP7_75t_L g640 ( 
.A(n_524),
.Y(n_640)
);

OAI22xp5_ASAP7_75t_L g641 ( 
.A1(n_556),
.A2(n_392),
.B1(n_49),
.B2(n_55),
.Y(n_641)
);

BUFx2_ASAP7_75t_L g642 ( 
.A(n_498),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_534),
.B(n_46),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_L g644 ( 
.A(n_500),
.B(n_57),
.Y(n_644)
);

BUFx4f_ASAP7_75t_L g645 ( 
.A(n_525),
.Y(n_645)
);

NOR2xp33_ASAP7_75t_L g646 ( 
.A(n_510),
.B(n_61),
.Y(n_646)
);

NOR2xp33_ASAP7_75t_L g647 ( 
.A(n_544),
.B(n_62),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_557),
.B(n_63),
.Y(n_648)
);

BUFx12f_ASAP7_75t_L g649 ( 
.A(n_503),
.Y(n_649)
);

A2O1A1Ixp33_ASAP7_75t_L g650 ( 
.A1(n_618),
.A2(n_558),
.B(n_555),
.C(n_515),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_605),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_613),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_576),
.Y(n_653)
);

A2O1A1Ixp33_ASAP7_75t_L g654 ( 
.A1(n_608),
.A2(n_527),
.B(n_505),
.C(n_569),
.Y(n_654)
);

BUFx3_ASAP7_75t_L g655 ( 
.A(n_571),
.Y(n_655)
);

NOR2xp33_ASAP7_75t_SL g656 ( 
.A(n_603),
.B(n_562),
.Y(n_656)
);

BUFx3_ASAP7_75t_L g657 ( 
.A(n_591),
.Y(n_657)
);

CKINVDCx6p67_ASAP7_75t_R g658 ( 
.A(n_602),
.Y(n_658)
);

OAI21x1_ASAP7_75t_L g659 ( 
.A1(n_594),
.A2(n_505),
.B(n_507),
.Y(n_659)
);

AO21x2_ASAP7_75t_L g660 ( 
.A1(n_589),
.A2(n_543),
.B(n_540),
.Y(n_660)
);

AO21x2_ASAP7_75t_L g661 ( 
.A1(n_638),
.A2(n_559),
.B(n_507),
.Y(n_661)
);

INVx4_ASAP7_75t_L g662 ( 
.A(n_570),
.Y(n_662)
);

AO31x2_ASAP7_75t_L g663 ( 
.A1(n_641),
.A2(n_535),
.A3(n_70),
.B(n_71),
.Y(n_663)
);

INVx1_ASAP7_75t_SL g664 ( 
.A(n_585),
.Y(n_664)
);

AOI21xp5_ASAP7_75t_L g665 ( 
.A1(n_617),
.A2(n_611),
.B(n_622),
.Y(n_665)
);

OAI22x1_ASAP7_75t_L g666 ( 
.A1(n_627),
.A2(n_76),
.B1(n_77),
.B2(n_82),
.Y(n_666)
);

AO31x2_ASAP7_75t_L g667 ( 
.A1(n_577),
.A2(n_83),
.A3(n_85),
.B(n_87),
.Y(n_667)
);

AOI221x1_ASAP7_75t_L g668 ( 
.A1(n_638),
.A2(n_90),
.B1(n_91),
.B2(n_93),
.C(n_96),
.Y(n_668)
);

INVx3_ASAP7_75t_L g669 ( 
.A(n_583),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_612),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_572),
.Y(n_671)
);

A2O1A1Ixp33_ASAP7_75t_L g672 ( 
.A1(n_616),
.A2(n_103),
.B(n_104),
.C(n_112),
.Y(n_672)
);

OAI21xp5_ASAP7_75t_L g673 ( 
.A1(n_580),
.A2(n_584),
.B(n_588),
.Y(n_673)
);

O2A1O1Ixp33_ASAP7_75t_L g674 ( 
.A1(n_635),
.A2(n_118),
.B(n_119),
.C(n_123),
.Y(n_674)
);

AO21x2_ASAP7_75t_L g675 ( 
.A1(n_639),
.A2(n_127),
.B(n_130),
.Y(n_675)
);

NAND2x1p5_ASAP7_75t_L g676 ( 
.A(n_574),
.B(n_132),
.Y(n_676)
);

AO31x2_ASAP7_75t_L g677 ( 
.A1(n_623),
.A2(n_134),
.A3(n_135),
.B(n_136),
.Y(n_677)
);

A2O1A1Ixp33_ASAP7_75t_L g678 ( 
.A1(n_634),
.A2(n_138),
.B(n_139),
.C(n_140),
.Y(n_678)
);

AOI21xp5_ASAP7_75t_L g679 ( 
.A1(n_614),
.A2(n_141),
.B(n_142),
.Y(n_679)
);

A2O1A1Ixp33_ASAP7_75t_L g680 ( 
.A1(n_592),
.A2(n_146),
.B(n_147),
.C(n_152),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_586),
.B(n_154),
.Y(n_681)
);

AOI221x1_ASAP7_75t_L g682 ( 
.A1(n_629),
.A2(n_155),
.B1(n_159),
.B2(n_164),
.C(n_165),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_590),
.Y(n_683)
);

OAI22xp5_ASAP7_75t_L g684 ( 
.A1(n_604),
.A2(n_167),
.B1(n_169),
.B2(n_171),
.Y(n_684)
);

AO31x2_ASAP7_75t_L g685 ( 
.A1(n_599),
.A2(n_172),
.A3(n_174),
.B(n_177),
.Y(n_685)
);

AO31x2_ASAP7_75t_L g686 ( 
.A1(n_600),
.A2(n_181),
.A3(n_183),
.B(n_184),
.Y(n_686)
);

AOI221xp5_ASAP7_75t_SL g687 ( 
.A1(n_615),
.A2(n_185),
.B1(n_610),
.B2(n_630),
.C(n_625),
.Y(n_687)
);

INVx3_ASAP7_75t_L g688 ( 
.A(n_583),
.Y(n_688)
);

BUFx6f_ASAP7_75t_L g689 ( 
.A(n_619),
.Y(n_689)
);

NOR2xp33_ASAP7_75t_SL g690 ( 
.A(n_631),
.B(n_649),
.Y(n_690)
);

NOR2x1_ASAP7_75t_SL g691 ( 
.A(n_581),
.B(n_607),
.Y(n_691)
);

BUFx4_ASAP7_75t_SL g692 ( 
.A(n_621),
.Y(n_692)
);

AND2x4_ASAP7_75t_L g693 ( 
.A(n_642),
.B(n_631),
.Y(n_693)
);

AND2x2_ASAP7_75t_L g694 ( 
.A(n_604),
.B(n_627),
.Y(n_694)
);

BUFx4f_ASAP7_75t_SL g695 ( 
.A(n_597),
.Y(n_695)
);

INVx3_ASAP7_75t_L g696 ( 
.A(n_636),
.Y(n_696)
);

INVxp67_ASAP7_75t_SL g697 ( 
.A(n_593),
.Y(n_697)
);

OR2x6_ASAP7_75t_L g698 ( 
.A(n_633),
.B(n_582),
.Y(n_698)
);

OR2x2_ASAP7_75t_L g699 ( 
.A(n_579),
.B(n_587),
.Y(n_699)
);

BUFx2_ASAP7_75t_SL g700 ( 
.A(n_636),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_596),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_598),
.B(n_624),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_578),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_609),
.Y(n_704)
);

OAI21x1_ASAP7_75t_L g705 ( 
.A1(n_637),
.A2(n_606),
.B(n_620),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_645),
.Y(n_706)
);

CKINVDCx8_ASAP7_75t_R g707 ( 
.A(n_619),
.Y(n_707)
);

AO31x2_ASAP7_75t_L g708 ( 
.A1(n_644),
.A2(n_646),
.A3(n_647),
.B(n_629),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_628),
.Y(n_709)
);

A2O1A1Ixp33_ASAP7_75t_L g710 ( 
.A1(n_626),
.A2(n_628),
.B(n_632),
.C(n_640),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_632),
.B(n_640),
.Y(n_711)
);

OAI21x1_ASAP7_75t_L g712 ( 
.A1(n_594),
.A2(n_589),
.B(n_595),
.Y(n_712)
);

AOI21xp5_ASAP7_75t_L g713 ( 
.A1(n_618),
.A2(n_566),
.B(n_589),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_605),
.Y(n_714)
);

OR2x2_ASAP7_75t_L g715 ( 
.A(n_602),
.B(n_493),
.Y(n_715)
);

AOI22xp5_ASAP7_75t_L g716 ( 
.A1(n_602),
.A2(n_353),
.B1(n_372),
.B2(n_321),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_605),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_605),
.Y(n_718)
);

BUFx2_ASAP7_75t_L g719 ( 
.A(n_585),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_605),
.Y(n_720)
);

BUFx3_ASAP7_75t_L g721 ( 
.A(n_571),
.Y(n_721)
);

AO31x2_ASAP7_75t_L g722 ( 
.A1(n_589),
.A2(n_641),
.A3(n_577),
.B(n_560),
.Y(n_722)
);

INVx3_ASAP7_75t_L g723 ( 
.A(n_583),
.Y(n_723)
);

AOI21xp5_ASAP7_75t_L g724 ( 
.A1(n_618),
.A2(n_566),
.B(n_589),
.Y(n_724)
);

INVx2_ASAP7_75t_SL g725 ( 
.A(n_591),
.Y(n_725)
);

A2O1A1Ixp33_ASAP7_75t_L g726 ( 
.A1(n_618),
.A2(n_608),
.B(n_611),
.C(n_616),
.Y(n_726)
);

OAI21x1_ASAP7_75t_L g727 ( 
.A1(n_594),
.A2(n_589),
.B(n_595),
.Y(n_727)
);

OAI21xp5_ASAP7_75t_L g728 ( 
.A1(n_589),
.A2(n_611),
.B(n_618),
.Y(n_728)
);

A2O1A1Ixp33_ASAP7_75t_L g729 ( 
.A1(n_618),
.A2(n_608),
.B(n_611),
.C(n_616),
.Y(n_729)
);

NOR2xp33_ASAP7_75t_SL g730 ( 
.A(n_603),
.B(n_485),
.Y(n_730)
);

O2A1O1Ixp33_ASAP7_75t_SL g731 ( 
.A1(n_648),
.A2(n_568),
.B(n_643),
.C(n_577),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_573),
.B(n_608),
.Y(n_732)
);

A2O1A1Ixp33_ASAP7_75t_L g733 ( 
.A1(n_618),
.A2(n_608),
.B(n_611),
.C(n_616),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_602),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_573),
.B(n_608),
.Y(n_735)
);

AOI21xp5_ASAP7_75t_L g736 ( 
.A1(n_618),
.A2(n_566),
.B(n_589),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_605),
.Y(n_737)
);

INVx1_ASAP7_75t_SL g738 ( 
.A(n_585),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_573),
.B(n_608),
.Y(n_739)
);

OAI21xp5_ASAP7_75t_L g740 ( 
.A1(n_589),
.A2(n_611),
.B(n_618),
.Y(n_740)
);

OAI22xp5_ASAP7_75t_L g741 ( 
.A1(n_608),
.A2(n_412),
.B1(n_553),
.B2(n_575),
.Y(n_741)
);

NOR2xp33_ASAP7_75t_L g742 ( 
.A(n_602),
.B(n_502),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_605),
.Y(n_743)
);

AOI21xp5_ASAP7_75t_L g744 ( 
.A1(n_618),
.A2(n_566),
.B(n_589),
.Y(n_744)
);

A2O1A1Ixp33_ASAP7_75t_L g745 ( 
.A1(n_618),
.A2(n_608),
.B(n_611),
.C(n_616),
.Y(n_745)
);

AO31x2_ASAP7_75t_L g746 ( 
.A1(n_589),
.A2(n_641),
.A3(n_577),
.B(n_560),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_605),
.Y(n_747)
);

BUFx2_ASAP7_75t_L g748 ( 
.A(n_585),
.Y(n_748)
);

OAI21x1_ASAP7_75t_L g749 ( 
.A1(n_594),
.A2(n_589),
.B(n_595),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_605),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_573),
.B(n_608),
.Y(n_751)
);

BUFx2_ASAP7_75t_L g752 ( 
.A(n_585),
.Y(n_752)
);

A2O1A1Ixp33_ASAP7_75t_L g753 ( 
.A1(n_732),
.A2(n_735),
.B(n_751),
.C(n_739),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_L g754 ( 
.A(n_715),
.B(n_664),
.Y(n_754)
);

AOI21xp5_ASAP7_75t_L g755 ( 
.A1(n_731),
.A2(n_733),
.B(n_726),
.Y(n_755)
);

AND2x4_ASAP7_75t_L g756 ( 
.A(n_694),
.B(n_693),
.Y(n_756)
);

AOI22xp5_ASAP7_75t_L g757 ( 
.A1(n_716),
.A2(n_738),
.B1(n_730),
.B2(n_697),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_720),
.Y(n_758)
);

AOI21xp5_ASAP7_75t_L g759 ( 
.A1(n_729),
.A2(n_745),
.B(n_744),
.Y(n_759)
);

OR2x2_ASAP7_75t_L g760 ( 
.A(n_658),
.B(n_719),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_720),
.Y(n_761)
);

NAND2x1_ASAP7_75t_L g762 ( 
.A(n_696),
.B(n_671),
.Y(n_762)
);

BUFx2_ASAP7_75t_L g763 ( 
.A(n_655),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_737),
.B(n_743),
.Y(n_764)
);

AOI21xp5_ASAP7_75t_L g765 ( 
.A1(n_713),
.A2(n_736),
.B(n_724),
.Y(n_765)
);

HB1xp67_ASAP7_75t_L g766 ( 
.A(n_721),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_737),
.B(n_743),
.Y(n_767)
);

AO31x2_ASAP7_75t_L g768 ( 
.A1(n_668),
.A2(n_710),
.A3(n_682),
.B(n_650),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_747),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_651),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_747),
.Y(n_771)
);

OAI21xp5_ASAP7_75t_L g772 ( 
.A1(n_654),
.A2(n_687),
.B(n_741),
.Y(n_772)
);

INVx2_ASAP7_75t_SL g773 ( 
.A(n_657),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_652),
.B(n_717),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_714),
.Y(n_775)
);

AOI22xp33_ASAP7_75t_L g776 ( 
.A1(n_699),
.A2(n_752),
.B1(n_748),
.B2(n_695),
.Y(n_776)
);

OR2x2_ASAP7_75t_L g777 ( 
.A(n_734),
.B(n_742),
.Y(n_777)
);

AND2x2_ASAP7_75t_L g778 ( 
.A(n_691),
.B(n_693),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_750),
.B(n_718),
.Y(n_779)
);

INVx1_ASAP7_75t_SL g780 ( 
.A(n_700),
.Y(n_780)
);

AOI21xp5_ASAP7_75t_SL g781 ( 
.A1(n_666),
.A2(n_676),
.B(n_698),
.Y(n_781)
);

INVx4_ASAP7_75t_L g782 ( 
.A(n_662),
.Y(n_782)
);

BUFx12f_ASAP7_75t_L g783 ( 
.A(n_725),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_671),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_653),
.B(n_683),
.Y(n_785)
);

INVx1_ASAP7_75t_SL g786 ( 
.A(n_692),
.Y(n_786)
);

O2A1O1Ixp33_ASAP7_75t_L g787 ( 
.A1(n_701),
.A2(n_674),
.B(n_702),
.C(n_681),
.Y(n_787)
);

CKINVDCx11_ASAP7_75t_R g788 ( 
.A(n_707),
.Y(n_788)
);

OAI21xp5_ASAP7_75t_L g789 ( 
.A1(n_673),
.A2(n_705),
.B(n_659),
.Y(n_789)
);

AO31x2_ASAP7_75t_L g790 ( 
.A1(n_672),
.A2(n_678),
.A3(n_680),
.B(n_679),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_704),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_704),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_703),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_706),
.Y(n_794)
);

OAI21x1_ASAP7_75t_L g795 ( 
.A1(n_709),
.A2(n_684),
.B(n_696),
.Y(n_795)
);

AOI21xp5_ASAP7_75t_L g796 ( 
.A1(n_660),
.A2(n_661),
.B(n_675),
.Y(n_796)
);

A2O1A1Ixp33_ASAP7_75t_L g797 ( 
.A1(n_669),
.A2(n_723),
.B(n_688),
.C(n_656),
.Y(n_797)
);

BUFx6f_ASAP7_75t_L g798 ( 
.A(n_689),
.Y(n_798)
);

AO31x2_ASAP7_75t_L g799 ( 
.A1(n_722),
.A2(n_746),
.A3(n_667),
.B(n_663),
.Y(n_799)
);

AO31x2_ASAP7_75t_L g800 ( 
.A1(n_722),
.A2(n_746),
.A3(n_667),
.B(n_663),
.Y(n_800)
);

OA21x2_ASAP7_75t_L g801 ( 
.A1(n_667),
.A2(n_677),
.B(n_685),
.Y(n_801)
);

NOR2xp33_ASAP7_75t_L g802 ( 
.A(n_690),
.B(n_670),
.Y(n_802)
);

BUFx3_ASAP7_75t_L g803 ( 
.A(n_689),
.Y(n_803)
);

OAI21x1_ASAP7_75t_SL g804 ( 
.A1(n_685),
.A2(n_686),
.B(n_677),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_685),
.Y(n_805)
);

OA21x2_ASAP7_75t_L g806 ( 
.A1(n_708),
.A2(n_727),
.B(n_712),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_708),
.B(n_732),
.Y(n_807)
);

OA21x2_ASAP7_75t_L g808 ( 
.A1(n_708),
.A2(n_727),
.B(n_712),
.Y(n_808)
);

AO31x2_ASAP7_75t_L g809 ( 
.A1(n_665),
.A2(n_729),
.A3(n_733),
.B(n_726),
.Y(n_809)
);

AO21x2_ASAP7_75t_L g810 ( 
.A1(n_728),
.A2(n_740),
.B(n_665),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_732),
.B(n_735),
.Y(n_811)
);

OAI21xp33_ASAP7_75t_SL g812 ( 
.A1(n_698),
.A2(n_553),
.B(n_732),
.Y(n_812)
);

BUFx8_ASAP7_75t_L g813 ( 
.A(n_655),
.Y(n_813)
);

INVx5_ASAP7_75t_L g814 ( 
.A(n_698),
.Y(n_814)
);

INVx1_ASAP7_75t_SL g815 ( 
.A(n_658),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_732),
.B(n_735),
.Y(n_816)
);

BUFx12f_ASAP7_75t_L g817 ( 
.A(n_734),
.Y(n_817)
);

AOI21xp33_ASAP7_75t_SL g818 ( 
.A1(n_670),
.A2(n_531),
.B(n_353),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_732),
.B(n_735),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_720),
.Y(n_820)
);

AO21x1_ASAP7_75t_SL g821 ( 
.A1(n_671),
.A2(n_711),
.B(n_601),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_732),
.B(n_735),
.Y(n_822)
);

CKINVDCx8_ASAP7_75t_R g823 ( 
.A(n_700),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_732),
.B(n_735),
.Y(n_824)
);

OA21x2_ASAP7_75t_L g825 ( 
.A1(n_712),
.A2(n_727),
.B(n_749),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_732),
.B(n_735),
.Y(n_826)
);

BUFx2_ASAP7_75t_L g827 ( 
.A(n_655),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_720),
.Y(n_828)
);

AOI21xp5_ASAP7_75t_L g829 ( 
.A1(n_731),
.A2(n_729),
.B(n_726),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_720),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_758),
.Y(n_831)
);

AO21x2_ASAP7_75t_L g832 ( 
.A1(n_804),
.A2(n_755),
.B(n_829),
.Y(n_832)
);

AO21x2_ASAP7_75t_L g833 ( 
.A1(n_796),
.A2(n_759),
.B(n_789),
.Y(n_833)
);

AO21x2_ASAP7_75t_L g834 ( 
.A1(n_765),
.A2(n_772),
.B(n_805),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_758),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_811),
.B(n_816),
.Y(n_836)
);

OR2x2_ASAP7_75t_L g837 ( 
.A(n_807),
.B(n_819),
.Y(n_837)
);

INVxp67_ASAP7_75t_L g838 ( 
.A(n_822),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_774),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_775),
.Y(n_840)
);

INVxp67_ASAP7_75t_SL g841 ( 
.A(n_784),
.Y(n_841)
);

INVx3_ASAP7_75t_L g842 ( 
.A(n_823),
.Y(n_842)
);

AND2x4_ASAP7_75t_L g843 ( 
.A(n_814),
.B(n_761),
.Y(n_843)
);

BUFx3_ASAP7_75t_L g844 ( 
.A(n_813),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_828),
.Y(n_845)
);

HB1xp67_ASAP7_75t_L g846 ( 
.A(n_780),
.Y(n_846)
);

OR2x2_ASAP7_75t_L g847 ( 
.A(n_824),
.B(n_826),
.Y(n_847)
);

HB1xp67_ASAP7_75t_L g848 ( 
.A(n_766),
.Y(n_848)
);

BUFx2_ASAP7_75t_L g849 ( 
.A(n_812),
.Y(n_849)
);

OR2x2_ASAP7_75t_L g850 ( 
.A(n_764),
.B(n_767),
.Y(n_850)
);

HB1xp67_ASAP7_75t_L g851 ( 
.A(n_763),
.Y(n_851)
);

OR2x2_ASAP7_75t_L g852 ( 
.A(n_792),
.B(n_753),
.Y(n_852)
);

HB1xp67_ASAP7_75t_L g853 ( 
.A(n_827),
.Y(n_853)
);

CKINVDCx20_ASAP7_75t_R g854 ( 
.A(n_788),
.Y(n_854)
);

INVx2_ASAP7_75t_SL g855 ( 
.A(n_813),
.Y(n_855)
);

BUFx2_ASAP7_75t_L g856 ( 
.A(n_798),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_810),
.Y(n_857)
);

AND2x2_ASAP7_75t_L g858 ( 
.A(n_792),
.B(n_791),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_785),
.B(n_754),
.Y(n_859)
);

INVx3_ASAP7_75t_L g860 ( 
.A(n_803),
.Y(n_860)
);

BUFx2_ASAP7_75t_L g861 ( 
.A(n_778),
.Y(n_861)
);

INVx2_ASAP7_75t_SL g862 ( 
.A(n_783),
.Y(n_862)
);

AND2x2_ASAP7_75t_L g863 ( 
.A(n_830),
.B(n_770),
.Y(n_863)
);

AO21x1_ASAP7_75t_SL g864 ( 
.A1(n_830),
.A2(n_781),
.B(n_814),
.Y(n_864)
);

INVxp67_ASAP7_75t_L g865 ( 
.A(n_760),
.Y(n_865)
);

CKINVDCx5p33_ASAP7_75t_R g866 ( 
.A(n_786),
.Y(n_866)
);

AND2x4_ASAP7_75t_L g867 ( 
.A(n_814),
.B(n_820),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_769),
.Y(n_868)
);

INVx2_ASAP7_75t_SL g869 ( 
.A(n_782),
.Y(n_869)
);

INVx1_ASAP7_75t_SL g870 ( 
.A(n_815),
.Y(n_870)
);

BUFx2_ASAP7_75t_L g871 ( 
.A(n_809),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_771),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_779),
.B(n_757),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_809),
.Y(n_874)
);

NOR2xp33_ASAP7_75t_L g875 ( 
.A(n_818),
.B(n_777),
.Y(n_875)
);

AOI21xp5_ASAP7_75t_SL g876 ( 
.A1(n_801),
.A2(n_787),
.B(n_797),
.Y(n_876)
);

BUFx3_ASAP7_75t_L g877 ( 
.A(n_773),
.Y(n_877)
);

HB1xp67_ASAP7_75t_L g878 ( 
.A(n_793),
.Y(n_878)
);

AND2x2_ASAP7_75t_L g879 ( 
.A(n_756),
.B(n_821),
.Y(n_879)
);

OAI21xp33_ASAP7_75t_SL g880 ( 
.A1(n_795),
.A2(n_776),
.B(n_782),
.Y(n_880)
);

AND2x2_ASAP7_75t_L g881 ( 
.A(n_756),
.B(n_794),
.Y(n_881)
);

INVx3_ASAP7_75t_L g882 ( 
.A(n_762),
.Y(n_882)
);

AND2x2_ASAP7_75t_L g883 ( 
.A(n_799),
.B(n_800),
.Y(n_883)
);

BUFx2_ASAP7_75t_L g884 ( 
.A(n_825),
.Y(n_884)
);

AND2x2_ASAP7_75t_L g885 ( 
.A(n_799),
.B(n_800),
.Y(n_885)
);

BUFx10_ASAP7_75t_L g886 ( 
.A(n_802),
.Y(n_886)
);

INVx2_ASAP7_75t_SL g887 ( 
.A(n_817),
.Y(n_887)
);

AND2x2_ASAP7_75t_L g888 ( 
.A(n_806),
.B(n_808),
.Y(n_888)
);

HB1xp67_ASAP7_75t_L g889 ( 
.A(n_768),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_831),
.Y(n_890)
);

AND2x2_ASAP7_75t_L g891 ( 
.A(n_835),
.B(n_790),
.Y(n_891)
);

HB1xp67_ASAP7_75t_L g892 ( 
.A(n_878),
.Y(n_892)
);

AND2x2_ASAP7_75t_L g893 ( 
.A(n_883),
.B(n_790),
.Y(n_893)
);

BUFx2_ASAP7_75t_L g894 ( 
.A(n_880),
.Y(n_894)
);

AND2x2_ASAP7_75t_L g895 ( 
.A(n_845),
.B(n_837),
.Y(n_895)
);

AND2x2_ASAP7_75t_L g896 ( 
.A(n_883),
.B(n_885),
.Y(n_896)
);

AND2x2_ASAP7_75t_L g897 ( 
.A(n_858),
.B(n_863),
.Y(n_897)
);

OAI21xp5_ASAP7_75t_L g898 ( 
.A1(n_838),
.A2(n_873),
.B(n_836),
.Y(n_898)
);

AND2x4_ASAP7_75t_L g899 ( 
.A(n_888),
.B(n_874),
.Y(n_899)
);

BUFx3_ASAP7_75t_L g900 ( 
.A(n_879),
.Y(n_900)
);

AND2x2_ASAP7_75t_L g901 ( 
.A(n_858),
.B(n_863),
.Y(n_901)
);

AND2x4_ASAP7_75t_L g902 ( 
.A(n_888),
.B(n_874),
.Y(n_902)
);

NOR2xp67_ASAP7_75t_L g903 ( 
.A(n_889),
.B(n_882),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_852),
.B(n_850),
.Y(n_904)
);

BUFx2_ASAP7_75t_SL g905 ( 
.A(n_869),
.Y(n_905)
);

AND2x2_ASAP7_75t_L g906 ( 
.A(n_885),
.B(n_871),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_852),
.B(n_850),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_868),
.B(n_872),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_839),
.B(n_847),
.Y(n_909)
);

HB1xp67_ASAP7_75t_L g910 ( 
.A(n_841),
.Y(n_910)
);

OR2x2_ASAP7_75t_SL g911 ( 
.A(n_851),
.B(n_853),
.Y(n_911)
);

AND2x2_ASAP7_75t_L g912 ( 
.A(n_861),
.B(n_847),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_840),
.B(n_849),
.Y(n_913)
);

AND2x2_ASAP7_75t_L g914 ( 
.A(n_832),
.B(n_834),
.Y(n_914)
);

OR2x2_ASAP7_75t_L g915 ( 
.A(n_859),
.B(n_848),
.Y(n_915)
);

AND2x2_ASAP7_75t_L g916 ( 
.A(n_832),
.B(n_881),
.Y(n_916)
);

AND2x2_ASAP7_75t_L g917 ( 
.A(n_832),
.B(n_881),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_912),
.B(n_846),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_890),
.Y(n_919)
);

INVxp67_ASAP7_75t_SL g920 ( 
.A(n_910),
.Y(n_920)
);

AND2x2_ASAP7_75t_L g921 ( 
.A(n_896),
.B(n_906),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_912),
.B(n_843),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_897),
.B(n_865),
.Y(n_923)
);

AND2x2_ASAP7_75t_L g924 ( 
.A(n_896),
.B(n_884),
.Y(n_924)
);

AND2x2_ASAP7_75t_L g925 ( 
.A(n_896),
.B(n_884),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_897),
.B(n_867),
.Y(n_926)
);

HB1xp67_ASAP7_75t_L g927 ( 
.A(n_892),
.Y(n_927)
);

AND2x2_ASAP7_75t_L g928 ( 
.A(n_906),
.B(n_916),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_892),
.Y(n_929)
);

AND2x4_ASAP7_75t_L g930 ( 
.A(n_899),
.B(n_902),
.Y(n_930)
);

AND2x2_ASAP7_75t_L g931 ( 
.A(n_906),
.B(n_833),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_901),
.B(n_895),
.Y(n_932)
);

HB1xp67_ASAP7_75t_L g933 ( 
.A(n_910),
.Y(n_933)
);

AND2x2_ASAP7_75t_L g934 ( 
.A(n_916),
.B(n_917),
.Y(n_934)
);

AOI22xp33_ASAP7_75t_L g935 ( 
.A1(n_917),
.A2(n_864),
.B1(n_875),
.B2(n_867),
.Y(n_935)
);

AND2x2_ASAP7_75t_L g936 ( 
.A(n_893),
.B(n_833),
.Y(n_936)
);

AND2x2_ASAP7_75t_SL g937 ( 
.A(n_894),
.B(n_867),
.Y(n_937)
);

AND2x2_ASAP7_75t_L g938 ( 
.A(n_893),
.B(n_857),
.Y(n_938)
);

AND2x2_ASAP7_75t_L g939 ( 
.A(n_934),
.B(n_893),
.Y(n_939)
);

AND2x2_ASAP7_75t_L g940 ( 
.A(n_934),
.B(n_928),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_921),
.B(n_901),
.Y(n_941)
);

INVx2_ASAP7_75t_L g942 ( 
.A(n_919),
.Y(n_942)
);

HB1xp67_ASAP7_75t_L g943 ( 
.A(n_933),
.Y(n_943)
);

INVx3_ASAP7_75t_L g944 ( 
.A(n_930),
.Y(n_944)
);

AND2x2_ASAP7_75t_L g945 ( 
.A(n_921),
.B(n_902),
.Y(n_945)
);

NAND4xp25_ASAP7_75t_L g946 ( 
.A(n_935),
.B(n_898),
.C(n_909),
.D(n_844),
.Y(n_946)
);

BUFx2_ASAP7_75t_L g947 ( 
.A(n_920),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_932),
.B(n_929),
.Y(n_948)
);

AND2x2_ASAP7_75t_L g949 ( 
.A(n_931),
.B(n_902),
.Y(n_949)
);

AND2x2_ASAP7_75t_L g950 ( 
.A(n_931),
.B(n_914),
.Y(n_950)
);

OR2x2_ASAP7_75t_L g951 ( 
.A(n_927),
.B(n_913),
.Y(n_951)
);

AND2x2_ASAP7_75t_L g952 ( 
.A(n_936),
.B(n_914),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_918),
.B(n_895),
.Y(n_953)
);

AND2x2_ASAP7_75t_L g954 ( 
.A(n_936),
.B(n_891),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_942),
.Y(n_955)
);

AND2x2_ASAP7_75t_L g956 ( 
.A(n_940),
.B(n_924),
.Y(n_956)
);

HB1xp67_ASAP7_75t_L g957 ( 
.A(n_947),
.Y(n_957)
);

OAI22xp5_ASAP7_75t_L g958 ( 
.A1(n_941),
.A2(n_911),
.B1(n_937),
.B2(n_900),
.Y(n_958)
);

INVx1_ASAP7_75t_SL g959 ( 
.A(n_947),
.Y(n_959)
);

INVx2_ASAP7_75t_L g960 ( 
.A(n_942),
.Y(n_960)
);

AND2x2_ASAP7_75t_L g961 ( 
.A(n_940),
.B(n_924),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_952),
.B(n_925),
.Y(n_962)
);

AND2x2_ASAP7_75t_L g963 ( 
.A(n_950),
.B(n_925),
.Y(n_963)
);

AOI22xp33_ASAP7_75t_SL g964 ( 
.A1(n_944),
.A2(n_937),
.B1(n_900),
.B2(n_905),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_952),
.B(n_938),
.Y(n_965)
);

HB1xp67_ASAP7_75t_L g966 ( 
.A(n_943),
.Y(n_966)
);

NOR2xp33_ASAP7_75t_L g967 ( 
.A(n_948),
.B(n_855),
.Y(n_967)
);

OR2x2_ASAP7_75t_L g968 ( 
.A(n_965),
.B(n_950),
.Y(n_968)
);

AOI21xp5_ASAP7_75t_L g969 ( 
.A1(n_958),
.A2(n_946),
.B(n_937),
.Y(n_969)
);

NOR2xp33_ASAP7_75t_SL g970 ( 
.A(n_959),
.B(n_844),
.Y(n_970)
);

AOI321xp33_ASAP7_75t_L g971 ( 
.A1(n_967),
.A2(n_926),
.A3(n_904),
.B1(n_907),
.B2(n_922),
.C(n_953),
.Y(n_971)
);

AND2x2_ASAP7_75t_L g972 ( 
.A(n_963),
.B(n_956),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_966),
.B(n_954),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_957),
.Y(n_974)
);

INVxp67_ASAP7_75t_SL g975 ( 
.A(n_960),
.Y(n_975)
);

AOI221xp5_ASAP7_75t_L g976 ( 
.A1(n_962),
.A2(n_946),
.B1(n_939),
.B2(n_923),
.C(n_898),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_SL g977 ( 
.A(n_964),
.B(n_944),
.Y(n_977)
);

AOI22xp5_ASAP7_75t_L g978 ( 
.A1(n_963),
.A2(n_944),
.B1(n_930),
.B2(n_949),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_956),
.Y(n_979)
);

INVx2_ASAP7_75t_SL g980 ( 
.A(n_961),
.Y(n_980)
);

HB1xp67_ASAP7_75t_L g981 ( 
.A(n_974),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_975),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_SL g983 ( 
.A(n_969),
.B(n_944),
.Y(n_983)
);

AND2x2_ASAP7_75t_L g984 ( 
.A(n_972),
.B(n_961),
.Y(n_984)
);

A2O1A1Ixp33_ASAP7_75t_L g985 ( 
.A1(n_970),
.A2(n_855),
.B(n_900),
.C(n_945),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_979),
.Y(n_986)
);

INVxp67_ASAP7_75t_L g987 ( 
.A(n_973),
.Y(n_987)
);

OAI211xp5_ASAP7_75t_SL g988 ( 
.A1(n_983),
.A2(n_976),
.B(n_977),
.C(n_971),
.Y(n_988)
);

AOI221xp5_ASAP7_75t_L g989 ( 
.A1(n_987),
.A2(n_977),
.B1(n_975),
.B2(n_980),
.C(n_978),
.Y(n_989)
);

AOI21xp33_ASAP7_75t_L g990 ( 
.A1(n_981),
.A2(n_915),
.B(n_870),
.Y(n_990)
);

AOI21xp5_ASAP7_75t_L g991 ( 
.A1(n_988),
.A2(n_985),
.B(n_982),
.Y(n_991)
);

AOI211xp5_ASAP7_75t_L g992 ( 
.A1(n_989),
.A2(n_866),
.B(n_982),
.C(n_887),
.Y(n_992)
);

NOR3xp33_ASAP7_75t_L g993 ( 
.A(n_992),
.B(n_887),
.C(n_862),
.Y(n_993)
);

NAND3xp33_ASAP7_75t_L g994 ( 
.A(n_991),
.B(n_866),
.C(n_990),
.Y(n_994)
);

AND2x4_ASAP7_75t_L g995 ( 
.A(n_993),
.B(n_862),
.Y(n_995)
);

NOR2xp33_ASAP7_75t_L g996 ( 
.A(n_994),
.B(n_854),
.Y(n_996)
);

OR2x2_ASAP7_75t_L g997 ( 
.A(n_995),
.B(n_986),
.Y(n_997)
);

INVx2_ASAP7_75t_L g998 ( 
.A(n_996),
.Y(n_998)
);

OAI22xp5_ASAP7_75t_SL g999 ( 
.A1(n_998),
.A2(n_854),
.B1(n_842),
.B2(n_877),
.Y(n_999)
);

INVx2_ASAP7_75t_L g1000 ( 
.A(n_997),
.Y(n_1000)
);

NOR2xp67_ASAP7_75t_L g1001 ( 
.A(n_998),
.B(n_842),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_SL g1002 ( 
.A(n_999),
.B(n_842),
.Y(n_1002)
);

OAI22xp5_ASAP7_75t_SL g1003 ( 
.A1(n_1000),
.A2(n_877),
.B1(n_911),
.B2(n_869),
.Y(n_1003)
);

XOR2xp5_ASAP7_75t_L g1004 ( 
.A(n_1001),
.B(n_915),
.Y(n_1004)
);

OR2x2_ASAP7_75t_L g1005 ( 
.A(n_1000),
.B(n_968),
.Y(n_1005)
);

OAI22xp5_ASAP7_75t_L g1006 ( 
.A1(n_999),
.A2(n_984),
.B1(n_951),
.B2(n_909),
.Y(n_1006)
);

AOI22xp33_ASAP7_75t_L g1007 ( 
.A1(n_1003),
.A2(n_886),
.B1(n_905),
.B2(n_864),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_1005),
.B(n_886),
.Y(n_1008)
);

AOI21xp33_ASAP7_75t_L g1009 ( 
.A1(n_1004),
.A2(n_860),
.B(n_908),
.Y(n_1009)
);

AOI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_1006),
.A2(n_907),
.B(n_904),
.Y(n_1010)
);

INVxp67_ASAP7_75t_L g1011 ( 
.A(n_1002),
.Y(n_1011)
);

OAI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_1011),
.A2(n_860),
.B(n_951),
.Y(n_1012)
);

AOI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_1008),
.A2(n_913),
.B(n_876),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_1009),
.B(n_955),
.Y(n_1014)
);

OR2x6_ASAP7_75t_L g1015 ( 
.A(n_1012),
.B(n_1010),
.Y(n_1015)
);

AO21x2_ASAP7_75t_L g1016 ( 
.A1(n_1014),
.A2(n_1007),
.B(n_903),
.Y(n_1016)
);

OR2x6_ASAP7_75t_L g1017 ( 
.A(n_1013),
.B(n_856),
.Y(n_1017)
);

AO21x2_ASAP7_75t_L g1018 ( 
.A1(n_1016),
.A2(n_1015),
.B(n_1017),
.Y(n_1018)
);


endmodule