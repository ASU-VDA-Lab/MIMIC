module fake_ariane_2930_n_1755 (n_83, n_8, n_56, n_60, n_170, n_160, n_64, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_158, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_169, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1755);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_160;
input n_64;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_158;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1755;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_1682;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_495;
wire n_267;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_238;
wire n_365;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1597;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1594;
wire n_680;
wire n_287;
wire n_1716;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_437;
wire n_337;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_824;
wire n_428;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1163;
wire n_186;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_1726;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_534;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1753;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_358;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_532;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1735;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_898;
wire n_857;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1285;
wire n_193;
wire n_761;
wire n_733;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1727;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1732;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_174;
wire n_275;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_866;
wire n_925;
wire n_246;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1252;
wire n_1129;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_548;
wire n_289;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1233;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_796;
wire n_573;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_167),
.Y(n_171)
);

INVx2_ASAP7_75t_SL g172 ( 
.A(n_169),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_138),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_28),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_74),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_165),
.Y(n_176)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_68),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_84),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_98),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_111),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_70),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_76),
.Y(n_182)
);

INVx1_ASAP7_75t_SL g183 ( 
.A(n_16),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_140),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_93),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_109),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_114),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_6),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_52),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_83),
.Y(n_190)
);

INVx1_ASAP7_75t_SL g191 ( 
.A(n_7),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_16),
.Y(n_192)
);

HB1xp67_ASAP7_75t_L g193 ( 
.A(n_80),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_21),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_145),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_30),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_66),
.Y(n_197)
);

BUFx10_ASAP7_75t_L g198 ( 
.A(n_9),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_117),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_37),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_88),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_153),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_38),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_142),
.Y(n_204)
);

BUFx2_ASAP7_75t_SL g205 ( 
.A(n_99),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_75),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_27),
.Y(n_207)
);

BUFx10_ASAP7_75t_L g208 ( 
.A(n_139),
.Y(n_208)
);

INVx1_ASAP7_75t_SL g209 ( 
.A(n_157),
.Y(n_209)
);

INVx1_ASAP7_75t_SL g210 ( 
.A(n_42),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_32),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_30),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_71),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_112),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_3),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_33),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_116),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_85),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_24),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_3),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_128),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_106),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_48),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_143),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_90),
.Y(n_225)
);

BUFx10_ASAP7_75t_L g226 ( 
.A(n_136),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_127),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_126),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_168),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_72),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_5),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_8),
.Y(n_232)
);

BUFx5_ASAP7_75t_L g233 ( 
.A(n_100),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_163),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_92),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_40),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_120),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_41),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_118),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_59),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_9),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_91),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_164),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_78),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_54),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_121),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_0),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_43),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_58),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_11),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_155),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_89),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_104),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_36),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_12),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_166),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_82),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_42),
.Y(n_258)
);

BUFx3_ASAP7_75t_L g259 ( 
.A(n_61),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_154),
.Y(n_260)
);

INVx2_ASAP7_75t_SL g261 ( 
.A(n_37),
.Y(n_261)
);

BUFx10_ASAP7_75t_L g262 ( 
.A(n_79),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_131),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_147),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_14),
.Y(n_265)
);

BUFx3_ASAP7_75t_L g266 ( 
.A(n_141),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_87),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_73),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_31),
.Y(n_269)
);

CKINVDCx16_ASAP7_75t_R g270 ( 
.A(n_94),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_22),
.Y(n_271)
);

INVx1_ASAP7_75t_SL g272 ( 
.A(n_52),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_95),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_20),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_108),
.Y(n_275)
);

INVx1_ASAP7_75t_SL g276 ( 
.A(n_14),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_148),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_34),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_25),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_7),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_39),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_64),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_44),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_15),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_12),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_115),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_50),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_33),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_67),
.Y(n_289)
);

BUFx2_ASAP7_75t_L g290 ( 
.A(n_28),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_102),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_53),
.Y(n_292)
);

BUFx10_ASAP7_75t_L g293 ( 
.A(n_161),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_13),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_113),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_6),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_134),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_144),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_25),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_23),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_55),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_159),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_146),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_47),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_35),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_96),
.Y(n_306)
);

BUFx2_ASAP7_75t_L g307 ( 
.A(n_137),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_31),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_21),
.Y(n_309)
);

BUFx10_ASAP7_75t_L g310 ( 
.A(n_81),
.Y(n_310)
);

BUFx2_ASAP7_75t_L g311 ( 
.A(n_62),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_35),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_0),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_39),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_38),
.Y(n_315)
);

BUFx3_ASAP7_75t_L g316 ( 
.A(n_26),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_43),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_32),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_46),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_51),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_132),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_49),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_170),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_5),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_162),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_20),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_46),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_26),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_135),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_150),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_57),
.Y(n_331)
);

INVx1_ASAP7_75t_SL g332 ( 
.A(n_123),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_160),
.Y(n_333)
);

BUFx8_ASAP7_75t_SL g334 ( 
.A(n_65),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_158),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_10),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_129),
.Y(n_337)
);

INVxp67_ASAP7_75t_SL g338 ( 
.A(n_316),
.Y(n_338)
);

INVxp33_ASAP7_75t_SL g339 ( 
.A(n_193),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_179),
.Y(n_340)
);

INVx2_ASAP7_75t_SL g341 ( 
.A(n_316),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_207),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_216),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_178),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_270),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_189),
.Y(n_346)
);

INVx1_ASAP7_75t_SL g347 ( 
.A(n_188),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_236),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_238),
.Y(n_349)
);

INVxp67_ASAP7_75t_L g350 ( 
.A(n_290),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_307),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_185),
.Y(n_352)
);

CKINVDCx16_ASAP7_75t_R g353 ( 
.A(n_198),
.Y(n_353)
);

INVxp33_ASAP7_75t_SL g354 ( 
.A(n_174),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_189),
.Y(n_355)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_259),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_259),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_266),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_325),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_196),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_274),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_311),
.Y(n_362)
);

INVxp67_ASAP7_75t_SL g363 ( 
.A(n_194),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_194),
.Y(n_364)
);

INVxp33_ASAP7_75t_SL g365 ( 
.A(n_174),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_211),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_211),
.Y(n_367)
);

BUFx6f_ASAP7_75t_L g368 ( 
.A(n_266),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_250),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_255),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_269),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_300),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_279),
.Y(n_373)
);

CKINVDCx14_ASAP7_75t_R g374 ( 
.A(n_208),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_294),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_208),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_312),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_336),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_215),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_313),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_314),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_318),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_208),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_226),
.Y(n_384)
);

INVxp33_ASAP7_75t_SL g385 ( 
.A(n_192),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_334),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_319),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_317),
.Y(n_388)
);

INVxp67_ASAP7_75t_L g389 ( 
.A(n_261),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_320),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_322),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_326),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_226),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_317),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_261),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_226),
.Y(n_396)
);

INVxp33_ASAP7_75t_SL g397 ( 
.A(n_192),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_262),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_262),
.Y(n_399)
);

HB1xp67_ASAP7_75t_L g400 ( 
.A(n_200),
.Y(n_400)
);

INVxp33_ASAP7_75t_SL g401 ( 
.A(n_200),
.Y(n_401)
);

INVxp67_ASAP7_75t_SL g402 ( 
.A(n_177),
.Y(n_402)
);

HB1xp67_ASAP7_75t_L g403 ( 
.A(n_203),
.Y(n_403)
);

CKINVDCx16_ASAP7_75t_R g404 ( 
.A(n_198),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_262),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_293),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_293),
.Y(n_407)
);

CKINVDCx16_ASAP7_75t_R g408 ( 
.A(n_198),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_293),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_310),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_310),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_310),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_175),
.Y(n_413)
);

XOR2xp5_ASAP7_75t_L g414 ( 
.A(n_203),
.B(n_1),
.Y(n_414)
);

CKINVDCx16_ASAP7_75t_R g415 ( 
.A(n_205),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_177),
.Y(n_416)
);

HB1xp67_ASAP7_75t_L g417 ( 
.A(n_212),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_199),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_199),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_206),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_206),
.Y(n_421)
);

INVxp33_ASAP7_75t_SL g422 ( 
.A(n_212),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_416),
.Y(n_423)
);

INVx3_ASAP7_75t_L g424 ( 
.A(n_368),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_416),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_418),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_360),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_418),
.Y(n_428)
);

AND2x4_ASAP7_75t_L g429 ( 
.A(n_413),
.B(n_172),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_419),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_399),
.B(n_182),
.Y(n_431)
);

NOR2x1_ASAP7_75t_L g432 ( 
.A(n_405),
.B(n_209),
.Y(n_432)
);

AND2x6_ASAP7_75t_L g433 ( 
.A(n_368),
.B(n_235),
.Y(n_433)
);

AND2x2_ASAP7_75t_L g434 ( 
.A(n_363),
.B(n_254),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_339),
.B(n_172),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_386),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_419),
.Y(n_437)
);

NOR2x1_ASAP7_75t_L g438 ( 
.A(n_406),
.B(n_332),
.Y(n_438)
);

INVx3_ASAP7_75t_L g439 ( 
.A(n_368),
.Y(n_439)
);

INVx3_ASAP7_75t_L g440 ( 
.A(n_368),
.Y(n_440)
);

XOR2xp5_ASAP7_75t_L g441 ( 
.A(n_361),
.B(n_254),
.Y(n_441)
);

BUFx8_ASAP7_75t_L g442 ( 
.A(n_407),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_420),
.Y(n_443)
);

AND2x4_ASAP7_75t_L g444 ( 
.A(n_402),
.B(n_235),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_409),
.B(n_197),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_372),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_420),
.Y(n_447)
);

CKINVDCx16_ASAP7_75t_R g448 ( 
.A(n_353),
.Y(n_448)
);

HB1xp67_ASAP7_75t_L g449 ( 
.A(n_347),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_421),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_421),
.Y(n_451)
);

BUFx6f_ASAP7_75t_L g452 ( 
.A(n_368),
.Y(n_452)
);

AND2x4_ASAP7_75t_L g453 ( 
.A(n_356),
.B(n_242),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_346),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_344),
.Y(n_455)
);

AND2x4_ASAP7_75t_L g456 ( 
.A(n_356),
.B(n_242),
.Y(n_456)
);

AND2x4_ASAP7_75t_L g457 ( 
.A(n_357),
.B(n_252),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_346),
.Y(n_458)
);

INVx1_ASAP7_75t_SL g459 ( 
.A(n_352),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_357),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_355),
.Y(n_461)
);

BUFx3_ASAP7_75t_L g462 ( 
.A(n_358),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_359),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_410),
.B(n_204),
.Y(n_464)
);

NOR2x1_ASAP7_75t_L g465 ( 
.A(n_358),
.B(n_218),
.Y(n_465)
);

BUFx10_ASAP7_75t_L g466 ( 
.A(n_340),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_355),
.Y(n_467)
);

CKINVDCx16_ASAP7_75t_R g468 ( 
.A(n_404),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_415),
.B(n_221),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_364),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_364),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_340),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_366),
.Y(n_473)
);

BUFx2_ASAP7_75t_L g474 ( 
.A(n_345),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_338),
.B(n_224),
.Y(n_475)
);

BUFx6f_ASAP7_75t_L g476 ( 
.A(n_366),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_367),
.Y(n_477)
);

INVx3_ASAP7_75t_L g478 ( 
.A(n_367),
.Y(n_478)
);

NOR2x1_ASAP7_75t_L g479 ( 
.A(n_395),
.B(n_244),
.Y(n_479)
);

INVx2_ASAP7_75t_SL g480 ( 
.A(n_376),
.Y(n_480)
);

INVx3_ASAP7_75t_L g481 ( 
.A(n_379),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_379),
.Y(n_482)
);

BUFx6f_ASAP7_75t_L g483 ( 
.A(n_388),
.Y(n_483)
);

BUFx6f_ASAP7_75t_L g484 ( 
.A(n_388),
.Y(n_484)
);

INVx3_ASAP7_75t_L g485 ( 
.A(n_394),
.Y(n_485)
);

AND2x4_ASAP7_75t_L g486 ( 
.A(n_341),
.B(n_252),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_345),
.Y(n_487)
);

HB1xp67_ASAP7_75t_L g488 ( 
.A(n_351),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_339),
.B(n_249),
.Y(n_489)
);

BUFx2_ASAP7_75t_L g490 ( 
.A(n_351),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_376),
.B(n_251),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_378),
.Y(n_492)
);

BUFx6f_ASAP7_75t_L g493 ( 
.A(n_342),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_343),
.Y(n_494)
);

INVx3_ASAP7_75t_L g495 ( 
.A(n_348),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_349),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_374),
.B(n_253),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_369),
.Y(n_498)
);

INVx3_ASAP7_75t_L g499 ( 
.A(n_370),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_371),
.Y(n_500)
);

INVx2_ASAP7_75t_SL g501 ( 
.A(n_432),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_430),
.Y(n_502)
);

OAI22xp33_ASAP7_75t_L g503 ( 
.A1(n_489),
.A2(n_362),
.B1(n_365),
.B2(n_354),
.Y(n_503)
);

OAI22xp33_ASAP7_75t_L g504 ( 
.A1(n_435),
.A2(n_362),
.B1(n_365),
.B2(n_354),
.Y(n_504)
);

NAND2xp33_ASAP7_75t_L g505 ( 
.A(n_480),
.B(n_383),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_444),
.B(n_383),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_430),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_450),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_SL g509 ( 
.A(n_480),
.B(n_384),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_450),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_SL g511 ( 
.A(n_491),
.B(n_384),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_444),
.B(n_429),
.Y(n_512)
);

INVx2_ASAP7_75t_SL g513 ( 
.A(n_432),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_436),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_450),
.Y(n_515)
);

INVx4_ASAP7_75t_L g516 ( 
.A(n_493),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_476),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_425),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_469),
.B(n_396),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_SL g520 ( 
.A(n_438),
.B(n_396),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_476),
.Y(n_521)
);

AOI22xp5_ASAP7_75t_L g522 ( 
.A1(n_438),
.A2(n_422),
.B1(n_385),
.B2(n_401),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_SL g523 ( 
.A(n_466),
.B(n_398),
.Y(n_523)
);

OR2x2_ASAP7_75t_L g524 ( 
.A(n_490),
.B(n_408),
.Y(n_524)
);

AOI22xp33_ASAP7_75t_L g525 ( 
.A1(n_444),
.A2(n_422),
.B1(n_385),
.B2(n_397),
.Y(n_525)
);

BUFx6f_ASAP7_75t_L g526 ( 
.A(n_452),
.Y(n_526)
);

BUFx2_ASAP7_75t_L g527 ( 
.A(n_490),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_425),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_476),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_SL g530 ( 
.A(n_442),
.B(n_466),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_426),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_444),
.B(n_398),
.Y(n_532)
);

INVx1_ASAP7_75t_SL g533 ( 
.A(n_449),
.Y(n_533)
);

AOI22xp33_ASAP7_75t_SL g534 ( 
.A1(n_442),
.A2(n_393),
.B1(n_411),
.B2(n_397),
.Y(n_534)
);

INVxp67_ASAP7_75t_SL g535 ( 
.A(n_462),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_476),
.Y(n_536)
);

HB1xp67_ASAP7_75t_L g537 ( 
.A(n_488),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_476),
.Y(n_538)
);

BUFx3_ASAP7_75t_L g539 ( 
.A(n_462),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_L g540 ( 
.A(n_497),
.B(n_412),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_475),
.B(n_412),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_476),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_SL g543 ( 
.A(n_466),
.B(n_401),
.Y(n_543)
);

INVx2_ASAP7_75t_SL g544 ( 
.A(n_434),
.Y(n_544)
);

AOI22xp5_ASAP7_75t_L g545 ( 
.A1(n_486),
.A2(n_183),
.B1(n_272),
.B2(n_191),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_483),
.Y(n_546)
);

BUFx2_ASAP7_75t_L g547 ( 
.A(n_474),
.Y(n_547)
);

BUFx16f_ASAP7_75t_R g548 ( 
.A(n_442),
.Y(n_548)
);

CKINVDCx16_ASAP7_75t_R g549 ( 
.A(n_448),
.Y(n_549)
);

OR2x2_ASAP7_75t_L g550 ( 
.A(n_448),
.B(n_350),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_483),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_483),
.Y(n_552)
);

BUFx3_ASAP7_75t_L g553 ( 
.A(n_462),
.Y(n_553)
);

INVx3_ASAP7_75t_L g554 ( 
.A(n_452),
.Y(n_554)
);

INVx4_ASAP7_75t_L g555 ( 
.A(n_493),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_426),
.Y(n_556)
);

BUFx6f_ASAP7_75t_L g557 ( 
.A(n_452),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_443),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_443),
.Y(n_559)
);

INVx3_ASAP7_75t_L g560 ( 
.A(n_452),
.Y(n_560)
);

INVx6_ASAP7_75t_L g561 ( 
.A(n_493),
.Y(n_561)
);

NOR2xp33_ASAP7_75t_L g562 ( 
.A(n_431),
.B(n_400),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_483),
.Y(n_563)
);

OAI22xp33_ASAP7_75t_L g564 ( 
.A1(n_468),
.A2(n_210),
.B1(n_276),
.B2(n_389),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_423),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_455),
.Y(n_566)
);

INVx8_ASAP7_75t_L g567 ( 
.A(n_433),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_SL g568 ( 
.A(n_466),
.B(n_403),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_423),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_483),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_483),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_463),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_484),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_484),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_484),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_445),
.B(n_417),
.Y(n_576)
);

OR2x6_ASAP7_75t_L g577 ( 
.A(n_486),
.B(n_429),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_484),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_428),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_429),
.B(n_341),
.Y(n_580)
);

INVx3_ASAP7_75t_L g581 ( 
.A(n_452),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_429),
.B(n_495),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_428),
.Y(n_583)
);

INVx1_ASAP7_75t_SL g584 ( 
.A(n_459),
.Y(n_584)
);

BUFx6f_ASAP7_75t_SL g585 ( 
.A(n_486),
.Y(n_585)
);

NOR2xp33_ASAP7_75t_L g586 ( 
.A(n_464),
.B(n_373),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_SL g587 ( 
.A(n_472),
.B(n_171),
.Y(n_587)
);

INVxp67_ASAP7_75t_L g588 ( 
.A(n_474),
.Y(n_588)
);

INVx3_ASAP7_75t_L g589 ( 
.A(n_452),
.Y(n_589)
);

INVx4_ASAP7_75t_L g590 ( 
.A(n_493),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_484),
.Y(n_591)
);

INVx3_ASAP7_75t_L g592 ( 
.A(n_484),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_461),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_461),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_461),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_SL g596 ( 
.A(n_487),
.B(n_171),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_437),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_471),
.Y(n_598)
);

OR2x6_ASAP7_75t_L g599 ( 
.A(n_486),
.B(n_375),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_492),
.Y(n_600)
);

NOR2x1p5_ASAP7_75t_L g601 ( 
.A(n_434),
.B(n_258),
.Y(n_601)
);

CKINVDCx14_ASAP7_75t_R g602 ( 
.A(n_427),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_437),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_471),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_447),
.Y(n_605)
);

BUFx3_ASAP7_75t_L g606 ( 
.A(n_424),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_446),
.Y(n_607)
);

BUFx10_ASAP7_75t_L g608 ( 
.A(n_453),
.Y(n_608)
);

NOR2xp33_ASAP7_75t_L g609 ( 
.A(n_499),
.B(n_377),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_447),
.Y(n_610)
);

INVx1_ASAP7_75t_SL g611 ( 
.A(n_441),
.Y(n_611)
);

INVx2_ASAP7_75t_SL g612 ( 
.A(n_453),
.Y(n_612)
);

BUFx2_ASAP7_75t_L g613 ( 
.A(n_468),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_451),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_SL g615 ( 
.A(n_493),
.B(n_173),
.Y(n_615)
);

AOI22xp33_ASAP7_75t_L g616 ( 
.A1(n_453),
.A2(n_381),
.B1(n_392),
.B2(n_391),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_SL g617 ( 
.A(n_493),
.B(n_173),
.Y(n_617)
);

AND3x1_ASAP7_75t_L g618 ( 
.A(n_479),
.B(n_382),
.C(n_380),
.Y(n_618)
);

INVx4_ASAP7_75t_L g619 ( 
.A(n_499),
.Y(n_619)
);

INVx3_ASAP7_75t_L g620 ( 
.A(n_424),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_471),
.Y(n_621)
);

AOI22xp33_ASAP7_75t_L g622 ( 
.A1(n_453),
.A2(n_390),
.B1(n_387),
.B2(n_414),
.Y(n_622)
);

NAND2xp33_ASAP7_75t_L g623 ( 
.A(n_499),
.B(n_176),
.Y(n_623)
);

BUFx3_ASAP7_75t_L g624 ( 
.A(n_424),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_451),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_478),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_478),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_460),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_460),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_478),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_478),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_481),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_481),
.Y(n_633)
);

AOI21x1_ASAP7_75t_L g634 ( 
.A1(n_465),
.A2(n_302),
.B(n_264),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_SL g635 ( 
.A(n_442),
.B(n_176),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_481),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_481),
.Y(n_637)
);

OAI22xp5_ASAP7_75t_L g638 ( 
.A1(n_499),
.A2(n_258),
.B1(n_328),
.B2(n_327),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_482),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_454),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_456),
.B(n_180),
.Y(n_641)
);

AND2x2_ASAP7_75t_SL g642 ( 
.A(n_456),
.B(n_264),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_482),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_485),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_485),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_485),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_454),
.Y(n_647)
);

INVx3_ASAP7_75t_L g648 ( 
.A(n_424),
.Y(n_648)
);

AOI22xp5_ASAP7_75t_L g649 ( 
.A1(n_494),
.A2(n_414),
.B1(n_287),
.B2(n_288),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_539),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_SL g651 ( 
.A(n_619),
.B(n_439),
.Y(n_651)
);

NOR2xp33_ASAP7_75t_L g652 ( 
.A(n_541),
.B(n_494),
.Y(n_652)
);

NOR2xp33_ASAP7_75t_L g653 ( 
.A(n_501),
.B(n_496),
.Y(n_653)
);

AND2x2_ASAP7_75t_L g654 ( 
.A(n_533),
.B(n_496),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_565),
.Y(n_655)
);

BUFx6f_ASAP7_75t_L g656 ( 
.A(n_567),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_539),
.Y(n_657)
);

HB1xp67_ASAP7_75t_L g658 ( 
.A(n_527),
.Y(n_658)
);

NOR2xp33_ASAP7_75t_L g659 ( 
.A(n_501),
.B(n_500),
.Y(n_659)
);

NAND3xp33_ASAP7_75t_L g660 ( 
.A(n_519),
.B(n_479),
.C(n_500),
.Y(n_660)
);

INVx2_ASAP7_75t_SL g661 ( 
.A(n_584),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_SL g662 ( 
.A(n_619),
.B(n_439),
.Y(n_662)
);

NOR3xp33_ASAP7_75t_L g663 ( 
.A(n_503),
.B(n_285),
.C(n_284),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_553),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_SL g665 ( 
.A(n_619),
.B(n_642),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_565),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_569),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_SL g668 ( 
.A(n_642),
.B(n_544),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_569),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_553),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_586),
.B(n_457),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_562),
.B(n_576),
.Y(n_672)
);

NOR2xp33_ASAP7_75t_SL g673 ( 
.A(n_530),
.B(n_284),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_642),
.B(n_457),
.Y(n_674)
);

O2A1O1Ixp33_ASAP7_75t_L g675 ( 
.A1(n_582),
.A2(n_498),
.B(n_485),
.C(n_477),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_540),
.B(n_457),
.Y(n_676)
);

NOR2xp33_ASAP7_75t_SL g677 ( 
.A(n_530),
.B(n_285),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_579),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_609),
.B(n_498),
.Y(n_679)
);

AND2x4_ASAP7_75t_L g680 ( 
.A(n_599),
.B(n_458),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_SL g681 ( 
.A(n_522),
.B(n_439),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_513),
.B(n_458),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_508),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_513),
.B(n_467),
.Y(n_684)
);

AOI21xp5_ASAP7_75t_L g685 ( 
.A1(n_632),
.A2(n_440),
.B(n_439),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_508),
.Y(n_686)
);

AOI221xp5_ASAP7_75t_L g687 ( 
.A1(n_504),
.A2(n_287),
.B1(n_328),
.B2(n_327),
.C(n_324),
.Y(n_687)
);

AOI22xp33_ASAP7_75t_L g688 ( 
.A1(n_579),
.A2(n_477),
.B1(n_473),
.B2(n_470),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_SL g689 ( 
.A(n_522),
.B(n_440),
.Y(n_689)
);

BUFx5_ASAP7_75t_L g690 ( 
.A(n_632),
.Y(n_690)
);

AND2x6_ASAP7_75t_L g691 ( 
.A(n_633),
.B(n_302),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_512),
.B(n_467),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_612),
.B(n_470),
.Y(n_693)
);

AND2x4_ASAP7_75t_L g694 ( 
.A(n_599),
.B(n_473),
.Y(n_694)
);

NAND2xp33_ASAP7_75t_L g695 ( 
.A(n_626),
.B(n_433),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_583),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_510),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_SL g698 ( 
.A(n_633),
.B(n_440),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_506),
.B(n_180),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_514),
.Y(n_700)
);

BUFx3_ASAP7_75t_L g701 ( 
.A(n_567),
.Y(n_701)
);

AOI22xp5_ASAP7_75t_L g702 ( 
.A1(n_601),
.A2(n_291),
.B1(n_202),
.B2(n_201),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_532),
.B(n_181),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_SL g704 ( 
.A(n_637),
.B(n_181),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_583),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_510),
.Y(n_706)
);

OAI22xp5_ASAP7_75t_L g707 ( 
.A1(n_525),
.A2(n_577),
.B1(n_603),
.B2(n_597),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_603),
.B(n_184),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_605),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_605),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_515),
.Y(n_711)
);

AND2x2_ASAP7_75t_L g712 ( 
.A(n_527),
.B(n_441),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_610),
.B(n_184),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_610),
.B(n_186),
.Y(n_714)
);

NOR2xp33_ASAP7_75t_L g715 ( 
.A(n_511),
.B(n_219),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_614),
.B(n_186),
.Y(n_716)
);

INVx3_ASAP7_75t_L g717 ( 
.A(n_608),
.Y(n_717)
);

NOR2xp33_ASAP7_75t_SL g718 ( 
.A(n_549),
.B(n_288),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_614),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_625),
.B(n_187),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_625),
.B(n_187),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_515),
.Y(n_722)
);

OAI22xp33_ASAP7_75t_L g723 ( 
.A1(n_649),
.A2(n_315),
.B1(n_299),
.B2(n_304),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_SL g724 ( 
.A(n_637),
.B(n_190),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_640),
.B(n_190),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_SL g726 ( 
.A(n_626),
.B(n_195),
.Y(n_726)
);

AND2x2_ASAP7_75t_L g727 ( 
.A(n_547),
.B(n_296),
.Y(n_727)
);

NOR2xp67_ASAP7_75t_L g728 ( 
.A(n_588),
.B(n_195),
.Y(n_728)
);

BUFx5_ASAP7_75t_L g729 ( 
.A(n_608),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_593),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_647),
.B(n_201),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_627),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_627),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_630),
.B(n_202),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_630),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_593),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_631),
.B(n_636),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_631),
.B(n_257),
.Y(n_738)
);

OR2x6_ASAP7_75t_L g739 ( 
.A(n_613),
.B(n_329),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_636),
.B(n_257),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_SL g741 ( 
.A(n_644),
.B(n_263),
.Y(n_741)
);

AND2x4_ASAP7_75t_L g742 ( 
.A(n_599),
.B(n_296),
.Y(n_742)
);

AOI22xp5_ASAP7_75t_L g743 ( 
.A1(n_601),
.A2(n_263),
.B1(n_335),
.B2(n_333),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_594),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_SL g745 ( 
.A(n_644),
.B(n_295),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_594),
.Y(n_746)
);

INVx2_ASAP7_75t_SL g747 ( 
.A(n_547),
.Y(n_747)
);

AND2x2_ASAP7_75t_L g748 ( 
.A(n_524),
.B(n_299),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_SL g749 ( 
.A(n_645),
.B(n_295),
.Y(n_749)
);

AND2x2_ASAP7_75t_L g750 ( 
.A(n_524),
.B(n_304),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_SL g751 ( 
.A(n_645),
.B(n_297),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_518),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_518),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_646),
.B(n_298),
.Y(n_754)
);

INVx2_ASAP7_75t_SL g755 ( 
.A(n_550),
.Y(n_755)
);

NOR2xp33_ASAP7_75t_L g756 ( 
.A(n_520),
.B(n_220),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_528),
.Y(n_757)
);

OR2x2_ASAP7_75t_L g758 ( 
.A(n_550),
.B(n_549),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_595),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_595),
.Y(n_760)
);

INVxp67_ASAP7_75t_L g761 ( 
.A(n_537),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_528),
.Y(n_762)
);

NOR2xp33_ASAP7_75t_L g763 ( 
.A(n_509),
.B(n_223),
.Y(n_763)
);

AOI22xp5_ASAP7_75t_L g764 ( 
.A1(n_599),
.A2(n_298),
.B1(n_335),
.B2(n_333),
.Y(n_764)
);

NOR3xp33_ASAP7_75t_L g765 ( 
.A(n_543),
.B(n_305),
.C(n_308),
.Y(n_765)
);

NOR2xp67_ASAP7_75t_L g766 ( 
.A(n_566),
.B(n_321),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_SL g767 ( 
.A(n_646),
.B(n_321),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_598),
.Y(n_768)
);

AND2x2_ASAP7_75t_L g769 ( 
.A(n_613),
.B(n_305),
.Y(n_769)
);

INVx5_ASAP7_75t_L g770 ( 
.A(n_567),
.Y(n_770)
);

NOR2xp33_ASAP7_75t_L g771 ( 
.A(n_587),
.B(n_231),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_535),
.B(n_331),
.Y(n_772)
);

NOR2xp33_ASAP7_75t_SL g773 ( 
.A(n_566),
.B(n_308),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_531),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_577),
.B(n_232),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_531),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_SL g777 ( 
.A(n_516),
.B(n_256),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_556),
.Y(n_778)
);

NOR2xp33_ASAP7_75t_L g779 ( 
.A(n_596),
.B(n_241),
.Y(n_779)
);

AOI22xp33_ASAP7_75t_L g780 ( 
.A1(n_556),
.A2(n_433),
.B1(n_337),
.B2(n_329),
.Y(n_780)
);

OR2x6_ASAP7_75t_L g781 ( 
.A(n_599),
.B(n_337),
.Y(n_781)
);

OAI221xp5_ASAP7_75t_L g782 ( 
.A1(n_545),
.A2(n_309),
.B1(n_315),
.B2(n_324),
.C(n_248),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_558),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_558),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_559),
.Y(n_785)
);

BUFx3_ASAP7_75t_L g786 ( 
.A(n_567),
.Y(n_786)
);

INVx2_ASAP7_75t_L g787 ( 
.A(n_604),
.Y(n_787)
);

NOR2xp33_ASAP7_75t_L g788 ( 
.A(n_635),
.B(n_585),
.Y(n_788)
);

OR2x2_ASAP7_75t_L g789 ( 
.A(n_607),
.B(n_309),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_559),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_604),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_628),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_SL g793 ( 
.A(n_516),
.B(n_260),
.Y(n_793)
);

BUFx3_ASAP7_75t_L g794 ( 
.A(n_567),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_628),
.Y(n_795)
);

INVx2_ASAP7_75t_SL g796 ( 
.A(n_607),
.Y(n_796)
);

NOR2xp33_ASAP7_75t_L g797 ( 
.A(n_585),
.B(n_247),
.Y(n_797)
);

OR2x2_ASAP7_75t_L g798 ( 
.A(n_572),
.B(n_600),
.Y(n_798)
);

AOI22xp33_ASAP7_75t_L g799 ( 
.A1(n_502),
.A2(n_507),
.B1(n_643),
.B2(n_639),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_577),
.B(n_265),
.Y(n_800)
);

AO22x1_ASAP7_75t_L g801 ( 
.A1(n_572),
.A2(n_271),
.B1(n_278),
.B2(n_280),
.Y(n_801)
);

NOR2xp33_ASAP7_75t_L g802 ( 
.A(n_585),
.B(n_281),
.Y(n_802)
);

NOR3xp33_ASAP7_75t_L g803 ( 
.A(n_505),
.B(n_283),
.C(n_292),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_629),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_629),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_621),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_672),
.B(n_580),
.Y(n_807)
);

BUFx6f_ASAP7_75t_L g808 ( 
.A(n_656),
.Y(n_808)
);

AOI22xp5_ASAP7_75t_SL g809 ( 
.A1(n_712),
.A2(n_514),
.B1(n_611),
.B2(n_602),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_655),
.Y(n_810)
);

NAND2xp33_ASAP7_75t_R g811 ( 
.A(n_700),
.B(n_548),
.Y(n_811)
);

BUFx6f_ASAP7_75t_L g812 ( 
.A(n_656),
.Y(n_812)
);

BUFx10_ASAP7_75t_L g813 ( 
.A(n_797),
.Y(n_813)
);

AND2x2_ASAP7_75t_L g814 ( 
.A(n_654),
.B(n_649),
.Y(n_814)
);

AOI22xp33_ASAP7_75t_L g815 ( 
.A1(n_723),
.A2(n_622),
.B1(n_545),
.B2(n_639),
.Y(n_815)
);

A2O1A1Ixp33_ASAP7_75t_L g816 ( 
.A1(n_652),
.A2(n_666),
.B(n_669),
.C(n_667),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_678),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_696),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_806),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_705),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_652),
.B(n_616),
.Y(n_821)
);

AOI22xp33_ASAP7_75t_L g822 ( 
.A1(n_723),
.A2(n_643),
.B1(n_507),
.B2(n_502),
.Y(n_822)
);

AND2x4_ASAP7_75t_L g823 ( 
.A(n_680),
.B(n_618),
.Y(n_823)
);

AOI22xp5_ASAP7_75t_L g824 ( 
.A1(n_668),
.A2(n_623),
.B1(n_618),
.B2(n_523),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_653),
.B(n_608),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_653),
.B(n_608),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_659),
.B(n_641),
.Y(n_827)
);

INVx2_ASAP7_75t_SL g828 ( 
.A(n_661),
.Y(n_828)
);

AOI22xp5_ASAP7_75t_L g829 ( 
.A1(n_668),
.A2(n_663),
.B1(n_665),
.B2(n_707),
.Y(n_829)
);

NOR2xp67_ASAP7_75t_L g830 ( 
.A(n_798),
.B(n_568),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_659),
.B(n_620),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_671),
.B(n_620),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_709),
.Y(n_833)
);

NAND3xp33_ASAP7_75t_L g834 ( 
.A(n_687),
.B(n_534),
.C(n_638),
.Y(n_834)
);

AND2x4_ASAP7_75t_L g835 ( 
.A(n_680),
.B(n_606),
.Y(n_835)
);

AOI22xp33_ASAP7_75t_L g836 ( 
.A1(n_674),
.A2(n_564),
.B1(n_555),
.B2(n_516),
.Y(n_836)
);

NOR2xp33_ASAP7_75t_L g837 ( 
.A(n_681),
.B(n_620),
.Y(n_837)
);

AOI22xp33_ASAP7_75t_L g838 ( 
.A1(n_782),
.A2(n_555),
.B1(n_590),
.B2(n_536),
.Y(n_838)
);

AOI22xp33_ASAP7_75t_L g839 ( 
.A1(n_663),
.A2(n_555),
.B1(n_590),
.B2(n_536),
.Y(n_839)
);

AND2x4_ASAP7_75t_L g840 ( 
.A(n_694),
.B(n_606),
.Y(n_840)
);

AOI22xp5_ASAP7_75t_L g841 ( 
.A1(n_665),
.A2(n_561),
.B1(n_617),
.B2(n_615),
.Y(n_841)
);

AOI22xp33_ASAP7_75t_SL g842 ( 
.A1(n_673),
.A2(n_677),
.B1(n_742),
.B2(n_718),
.Y(n_842)
);

INVx5_ASAP7_75t_L g843 ( 
.A(n_656),
.Y(n_843)
);

HB1xp67_ASAP7_75t_L g844 ( 
.A(n_658),
.Y(n_844)
);

BUFx4f_ASAP7_75t_L g845 ( 
.A(n_747),
.Y(n_845)
);

AND2x2_ASAP7_75t_L g846 ( 
.A(n_748),
.B(n_648),
.Y(n_846)
);

AND2x4_ASAP7_75t_L g847 ( 
.A(n_694),
.B(n_624),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_676),
.B(n_624),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_710),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_719),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_682),
.B(n_592),
.Y(n_851)
);

BUFx3_ASAP7_75t_L g852 ( 
.A(n_796),
.Y(n_852)
);

INVx3_ASAP7_75t_L g853 ( 
.A(n_656),
.Y(n_853)
);

INVx5_ASAP7_75t_L g854 ( 
.A(n_770),
.Y(n_854)
);

OAI21xp33_ASAP7_75t_L g855 ( 
.A1(n_773),
.A2(n_715),
.B(n_771),
.Y(n_855)
);

INVx2_ASAP7_75t_SL g856 ( 
.A(n_658),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_683),
.Y(n_857)
);

HB1xp67_ASAP7_75t_L g858 ( 
.A(n_781),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_SL g859 ( 
.A(n_729),
.B(n_590),
.Y(n_859)
);

INVx2_ASAP7_75t_SL g860 ( 
.A(n_758),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_792),
.Y(n_861)
);

BUFx2_ASAP7_75t_L g862 ( 
.A(n_755),
.Y(n_862)
);

INVxp67_ASAP7_75t_L g863 ( 
.A(n_681),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_795),
.Y(n_864)
);

INVx2_ASAP7_75t_L g865 ( 
.A(n_686),
.Y(n_865)
);

INVx2_ASAP7_75t_SL g866 ( 
.A(n_739),
.Y(n_866)
);

INVx2_ASAP7_75t_SL g867 ( 
.A(n_739),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_684),
.B(n_592),
.Y(n_868)
);

OAI21xp33_ASAP7_75t_L g869 ( 
.A1(n_715),
.A2(n_779),
.B(n_771),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_692),
.B(n_592),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_697),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_699),
.B(n_703),
.Y(n_872)
);

INVx2_ASAP7_75t_SL g873 ( 
.A(n_739),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_804),
.Y(n_874)
);

OR2x2_ASAP7_75t_L g875 ( 
.A(n_761),
.B(n_517),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_693),
.B(n_517),
.Y(n_876)
);

OR2x2_ASAP7_75t_L g877 ( 
.A(n_761),
.B(n_521),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_SL g878 ( 
.A(n_729),
.B(n_521),
.Y(n_878)
);

NAND2xp33_ASAP7_75t_SL g879 ( 
.A(n_717),
.B(n_529),
.Y(n_879)
);

CKINVDCx5p33_ASAP7_75t_R g880 ( 
.A(n_801),
.Y(n_880)
);

INVx2_ASAP7_75t_SL g881 ( 
.A(n_789),
.Y(n_881)
);

OAI21xp5_ASAP7_75t_L g882 ( 
.A1(n_737),
.A2(n_551),
.B(n_591),
.Y(n_882)
);

BUFx2_ASAP7_75t_L g883 ( 
.A(n_742),
.Y(n_883)
);

BUFx6f_ASAP7_75t_L g884 ( 
.A(n_701),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_805),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_679),
.B(n_529),
.Y(n_886)
);

NAND3xp33_ASAP7_75t_SL g887 ( 
.A(n_803),
.B(n_286),
.C(n_289),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_708),
.B(n_538),
.Y(n_888)
);

CKINVDCx5p33_ASAP7_75t_R g889 ( 
.A(n_769),
.Y(n_889)
);

NOR2xp33_ASAP7_75t_L g890 ( 
.A(n_689),
.B(n_538),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_752),
.Y(n_891)
);

AOI21xp5_ASAP7_75t_L g892 ( 
.A1(n_651),
.A2(n_554),
.B(n_560),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_SL g893 ( 
.A(n_729),
.B(n_542),
.Y(n_893)
);

BUFx3_ASAP7_75t_L g894 ( 
.A(n_786),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_713),
.B(n_542),
.Y(n_895)
);

BUFx2_ASAP7_75t_L g896 ( 
.A(n_727),
.Y(n_896)
);

OAI21xp5_ASAP7_75t_L g897 ( 
.A1(n_675),
.A2(n_573),
.B(n_591),
.Y(n_897)
);

AND2x4_ASAP7_75t_L g898 ( 
.A(n_781),
.B(n_546),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_753),
.Y(n_899)
);

CKINVDCx5p33_ASAP7_75t_R g900 ( 
.A(n_702),
.Y(n_900)
);

INVx3_ASAP7_75t_SL g901 ( 
.A(n_781),
.Y(n_901)
);

BUFx6f_ASAP7_75t_L g902 ( 
.A(n_786),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_706),
.Y(n_903)
);

INVx3_ASAP7_75t_L g904 ( 
.A(n_794),
.Y(n_904)
);

AND2x2_ASAP7_75t_L g905 ( 
.A(n_750),
.B(n_546),
.Y(n_905)
);

BUFx2_ASAP7_75t_L g906 ( 
.A(n_775),
.Y(n_906)
);

AOI22xp33_ASAP7_75t_L g907 ( 
.A1(n_757),
.A2(n_574),
.B1(n_551),
.B2(n_552),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_762),
.Y(n_908)
);

BUFx3_ASAP7_75t_L g909 ( 
.A(n_794),
.Y(n_909)
);

INVx3_ASAP7_75t_L g910 ( 
.A(n_717),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_711),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_774),
.Y(n_912)
);

NAND2x1p5_ASAP7_75t_L g913 ( 
.A(n_770),
.B(n_552),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_714),
.B(n_563),
.Y(n_914)
);

NOR2xp33_ASAP7_75t_L g915 ( 
.A(n_689),
.B(n_563),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_716),
.B(n_570),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_SL g917 ( 
.A(n_729),
.B(n_570),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_776),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_720),
.B(n_571),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_721),
.B(n_571),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_SL g921 ( 
.A(n_729),
.B(n_573),
.Y(n_921)
);

AOI22xp5_ASAP7_75t_L g922 ( 
.A1(n_803),
.A2(n_561),
.B1(n_574),
.B2(n_575),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_778),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_783),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_725),
.B(n_731),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_779),
.B(n_575),
.Y(n_926)
);

BUFx2_ASAP7_75t_L g927 ( 
.A(n_800),
.Y(n_927)
);

CKINVDCx5p33_ASAP7_75t_R g928 ( 
.A(n_743),
.Y(n_928)
);

INVx1_ASAP7_75t_SL g929 ( 
.A(n_797),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_763),
.B(n_728),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_784),
.Y(n_931)
);

HB1xp67_ASAP7_75t_L g932 ( 
.A(n_650),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_SL g933 ( 
.A(n_729),
.B(n_578),
.Y(n_933)
);

INVx4_ASAP7_75t_L g934 ( 
.A(n_770),
.Y(n_934)
);

NOR2xp33_ASAP7_75t_L g935 ( 
.A(n_660),
.B(n_561),
.Y(n_935)
);

BUFx3_ASAP7_75t_L g936 ( 
.A(n_657),
.Y(n_936)
);

AND2x2_ASAP7_75t_L g937 ( 
.A(n_802),
.B(n_634),
.Y(n_937)
);

INVx2_ASAP7_75t_L g938 ( 
.A(n_722),
.Y(n_938)
);

INVx2_ASAP7_75t_SL g939 ( 
.A(n_802),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_763),
.B(n_554),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_785),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_790),
.Y(n_942)
);

AND2x4_ASAP7_75t_L g943 ( 
.A(n_770),
.B(n_554),
.Y(n_943)
);

INVx5_ASAP7_75t_L g944 ( 
.A(n_691),
.Y(n_944)
);

OR2x2_ASAP7_75t_L g945 ( 
.A(n_765),
.B(n_560),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_730),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_736),
.Y(n_947)
);

AND2x2_ASAP7_75t_L g948 ( 
.A(n_766),
.B(n_634),
.Y(n_948)
);

INVx2_ASAP7_75t_L g949 ( 
.A(n_744),
.Y(n_949)
);

AND2x2_ASAP7_75t_L g950 ( 
.A(n_765),
.B(n_561),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_SL g951 ( 
.A(n_690),
.B(n_732),
.Y(n_951)
);

INVx2_ASAP7_75t_L g952 ( 
.A(n_746),
.Y(n_952)
);

HB1xp67_ASAP7_75t_L g953 ( 
.A(n_664),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_733),
.Y(n_954)
);

AOI21xp5_ASAP7_75t_L g955 ( 
.A1(n_651),
.A2(n_589),
.B(n_581),
.Y(n_955)
);

AND2x2_ASAP7_75t_L g956 ( 
.A(n_756),
.B(n_581),
.Y(n_956)
);

INVx5_ASAP7_75t_L g957 ( 
.A(n_691),
.Y(n_957)
);

AOI22xp33_ASAP7_75t_L g958 ( 
.A1(n_759),
.A2(n_433),
.B1(n_301),
.B2(n_303),
.Y(n_958)
);

INVx2_ASAP7_75t_SL g959 ( 
.A(n_670),
.Y(n_959)
);

INVx2_ASAP7_75t_L g960 ( 
.A(n_760),
.Y(n_960)
);

INVxp67_ASAP7_75t_L g961 ( 
.A(n_726),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_735),
.Y(n_962)
);

INVx2_ASAP7_75t_L g963 ( 
.A(n_768),
.Y(n_963)
);

INVx4_ASAP7_75t_L g964 ( 
.A(n_691),
.Y(n_964)
);

OR2x6_ASAP7_75t_L g965 ( 
.A(n_788),
.B(n_589),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_756),
.B(n_526),
.Y(n_966)
);

AOI221xp5_ASAP7_75t_SL g967 ( 
.A1(n_688),
.A2(n_724),
.B1(n_704),
.B2(n_726),
.C(n_745),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_787),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_688),
.B(n_526),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_791),
.Y(n_970)
);

INVx3_ASAP7_75t_L g971 ( 
.A(n_690),
.Y(n_971)
);

NOR2xp33_ASAP7_75t_L g972 ( 
.A(n_764),
.B(n_526),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_772),
.B(n_526),
.Y(n_973)
);

INVx2_ASAP7_75t_SL g974 ( 
.A(n_741),
.Y(n_974)
);

AOI21xp5_ASAP7_75t_L g975 ( 
.A1(n_662),
.A2(n_557),
.B(n_526),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_698),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_SL g977 ( 
.A(n_690),
.B(n_557),
.Y(n_977)
);

INVx2_ASAP7_75t_SL g978 ( 
.A(n_741),
.Y(n_978)
);

BUFx6f_ASAP7_75t_L g979 ( 
.A(n_691),
.Y(n_979)
);

INVx3_ASAP7_75t_L g980 ( 
.A(n_690),
.Y(n_980)
);

INVx2_ASAP7_75t_L g981 ( 
.A(n_690),
.Y(n_981)
);

OAI21xp5_ASAP7_75t_L g982 ( 
.A1(n_837),
.A2(n_698),
.B(n_685),
.Y(n_982)
);

BUFx6f_ASAP7_75t_L g983 ( 
.A(n_835),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_810),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_817),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_SL g986 ( 
.A(n_845),
.B(n_788),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_818),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_SL g988 ( 
.A(n_845),
.B(n_690),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_807),
.B(n_704),
.Y(n_989)
);

HB1xp67_ASAP7_75t_L g990 ( 
.A(n_844),
.Y(n_990)
);

BUFx3_ASAP7_75t_L g991 ( 
.A(n_862),
.Y(n_991)
);

OAI22xp5_ASAP7_75t_L g992 ( 
.A1(n_825),
.A2(n_740),
.B1(n_734),
.B2(n_738),
.Y(n_992)
);

NOR3xp33_ASAP7_75t_SL g993 ( 
.A(n_811),
.B(n_724),
.C(n_751),
.Y(n_993)
);

AOI22x1_ASAP7_75t_L g994 ( 
.A1(n_981),
.A2(n_557),
.B1(n_662),
.B2(n_691),
.Y(n_994)
);

HB1xp67_ASAP7_75t_L g995 ( 
.A(n_844),
.Y(n_995)
);

INVx5_ASAP7_75t_L g996 ( 
.A(n_979),
.Y(n_996)
);

INVx3_ASAP7_75t_SL g997 ( 
.A(n_880),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_820),
.Y(n_998)
);

INVx5_ASAP7_75t_L g999 ( 
.A(n_979),
.Y(n_999)
);

BUFx6f_ASAP7_75t_L g1000 ( 
.A(n_835),
.Y(n_1000)
);

AOI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_826),
.A2(n_831),
.B(n_827),
.Y(n_1001)
);

AOI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_872),
.A2(n_695),
.B(n_754),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_833),
.Y(n_1003)
);

AOI21xp5_ASAP7_75t_L g1004 ( 
.A1(n_977),
.A2(n_749),
.B(n_745),
.Y(n_1004)
);

AOI21xp5_ASAP7_75t_L g1005 ( 
.A1(n_816),
.A2(n_767),
.B(n_793),
.Y(n_1005)
);

AOI22xp5_ASAP7_75t_L g1006 ( 
.A1(n_869),
.A2(n_767),
.B1(n_793),
.B2(n_777),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_SL g1007 ( 
.A(n_855),
.B(n_799),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_849),
.Y(n_1008)
);

AND2x4_ASAP7_75t_L g1009 ( 
.A(n_840),
.B(n_799),
.Y(n_1009)
);

NOR2xp33_ASAP7_75t_R g1010 ( 
.A(n_811),
.B(n_780),
.Y(n_1010)
);

CKINVDCx11_ASAP7_75t_R g1011 ( 
.A(n_813),
.Y(n_1011)
);

NAND2xp33_ASAP7_75t_SL g1012 ( 
.A(n_930),
.B(n_557),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_821),
.B(n_780),
.Y(n_1013)
);

NOR3xp33_ASAP7_75t_SL g1014 ( 
.A(n_889),
.B(n_928),
.C(n_900),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_814),
.B(n_557),
.Y(n_1015)
);

BUFx2_ASAP7_75t_L g1016 ( 
.A(n_856),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_SL g1017 ( 
.A(n_929),
.B(n_213),
.Y(n_1017)
);

AO21x1_ASAP7_75t_L g1018 ( 
.A1(n_890),
.A2(n_330),
.B(n_323),
.Y(n_1018)
);

O2A1O1Ixp33_ASAP7_75t_L g1019 ( 
.A1(n_925),
.A2(n_306),
.B(n_2),
.C(n_4),
.Y(n_1019)
);

OA22x2_ASAP7_75t_L g1020 ( 
.A1(n_881),
.A2(n_239),
.B1(n_282),
.B2(n_277),
.Y(n_1020)
);

AO221x2_ASAP7_75t_L g1021 ( 
.A1(n_834),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.C(n_10),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_850),
.Y(n_1022)
);

AOI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_816),
.A2(n_214),
.B(n_275),
.Y(n_1023)
);

INVx2_ASAP7_75t_L g1024 ( 
.A(n_819),
.Y(n_1024)
);

BUFx6f_ASAP7_75t_L g1025 ( 
.A(n_840),
.Y(n_1025)
);

OAI22x1_ASAP7_75t_L g1026 ( 
.A1(n_883),
.A2(n_217),
.B1(n_222),
.B2(n_225),
.Y(n_1026)
);

NOR2x1_ASAP7_75t_L g1027 ( 
.A(n_852),
.B(n_433),
.Y(n_1027)
);

NOR2xp33_ASAP7_75t_L g1028 ( 
.A(n_939),
.B(n_227),
.Y(n_1028)
);

NAND3xp33_ASAP7_75t_SL g1029 ( 
.A(n_842),
.B(n_228),
.C(n_229),
.Y(n_1029)
);

AOI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_832),
.A2(n_230),
.B(n_273),
.Y(n_1030)
);

HB1xp67_ASAP7_75t_L g1031 ( 
.A(n_896),
.Y(n_1031)
);

INVx3_ASAP7_75t_SL g1032 ( 
.A(n_809),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_SL g1033 ( 
.A(n_842),
.B(n_243),
.Y(n_1033)
);

O2A1O1Ixp33_ASAP7_75t_L g1034 ( 
.A1(n_887),
.A2(n_13),
.B(n_15),
.C(n_17),
.Y(n_1034)
);

HB1xp67_ASAP7_75t_L g1035 ( 
.A(n_860),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_SL g1036 ( 
.A(n_830),
.B(n_245),
.Y(n_1036)
);

BUFx2_ASAP7_75t_L g1037 ( 
.A(n_823),
.Y(n_1037)
);

AOI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_886),
.A2(n_234),
.B(n_268),
.Y(n_1038)
);

OAI22xp5_ASAP7_75t_L g1039 ( 
.A1(n_829),
.A2(n_237),
.B1(n_240),
.B2(n_246),
.Y(n_1039)
);

OAI22xp5_ASAP7_75t_L g1040 ( 
.A1(n_824),
.A2(n_267),
.B1(n_19),
.B2(n_22),
.Y(n_1040)
);

INVx4_ASAP7_75t_L g1041 ( 
.A(n_847),
.Y(n_1041)
);

A2O1A1Ixp33_ASAP7_75t_L g1042 ( 
.A1(n_837),
.A2(n_433),
.B(n_233),
.C(n_23),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_861),
.Y(n_1043)
);

AOI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_848),
.A2(n_86),
.B(n_103),
.Y(n_1044)
);

OAI21x1_ASAP7_75t_SL g1045 ( 
.A1(n_981),
.A2(n_18),
.B(n_19),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_815),
.B(n_18),
.Y(n_1046)
);

AND2x4_ASAP7_75t_L g1047 ( 
.A(n_847),
.B(n_433),
.Y(n_1047)
);

OAI21xp33_ASAP7_75t_SL g1048 ( 
.A1(n_864),
.A2(n_24),
.B(n_27),
.Y(n_1048)
);

NOR2xp33_ASAP7_75t_SL g1049 ( 
.A(n_901),
.B(n_828),
.Y(n_1049)
);

AOI22xp5_ASAP7_75t_L g1050 ( 
.A1(n_887),
.A2(n_233),
.B1(n_34),
.B2(n_36),
.Y(n_1050)
);

INVx1_ASAP7_75t_SL g1051 ( 
.A(n_852),
.Y(n_1051)
);

NAND3xp33_ASAP7_75t_SL g1052 ( 
.A(n_815),
.B(n_29),
.C(n_40),
.Y(n_1052)
);

BUFx2_ASAP7_75t_L g1053 ( 
.A(n_823),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_SL g1054 ( 
.A(n_813),
.B(n_233),
.Y(n_1054)
);

AND2x2_ASAP7_75t_L g1055 ( 
.A(n_901),
.B(n_29),
.Y(n_1055)
);

AOI22xp5_ASAP7_75t_L g1056 ( 
.A1(n_863),
.A2(n_233),
.B1(n_45),
.B2(n_47),
.Y(n_1056)
);

AOI22xp5_ASAP7_75t_L g1057 ( 
.A1(n_863),
.A2(n_233),
.B1(n_45),
.B2(n_48),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_874),
.Y(n_1058)
);

INVx2_ASAP7_75t_L g1059 ( 
.A(n_819),
.Y(n_1059)
);

O2A1O1Ixp33_ASAP7_75t_L g1060 ( 
.A1(n_961),
.A2(n_41),
.B(n_49),
.C(n_50),
.Y(n_1060)
);

A2O1A1Ixp33_ASAP7_75t_L g1061 ( 
.A1(n_961),
.A2(n_233),
.B(n_51),
.C(n_60),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_885),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_846),
.B(n_233),
.Y(n_1063)
);

O2A1O1Ixp33_ASAP7_75t_L g1064 ( 
.A1(n_945),
.A2(n_56),
.B(n_63),
.C(n_69),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_905),
.B(n_77),
.Y(n_1065)
);

NAND2xp33_ASAP7_75t_SL g1066 ( 
.A(n_964),
.B(n_97),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_906),
.B(n_101),
.Y(n_1067)
);

NOR2xp33_ASAP7_75t_SL g1068 ( 
.A(n_964),
.B(n_105),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_927),
.B(n_107),
.Y(n_1069)
);

OAI22xp5_ASAP7_75t_L g1070 ( 
.A1(n_891),
.A2(n_110),
.B1(n_119),
.B2(n_122),
.Y(n_1070)
);

OAI22xp5_ASAP7_75t_L g1071 ( 
.A1(n_899),
.A2(n_124),
.B1(n_125),
.B2(n_130),
.Y(n_1071)
);

AOI21xp5_ASAP7_75t_L g1072 ( 
.A1(n_973),
.A2(n_951),
.B(n_870),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_SL g1073 ( 
.A(n_843),
.B(n_133),
.Y(n_1073)
);

BUFx2_ASAP7_75t_L g1074 ( 
.A(n_858),
.Y(n_1074)
);

AOI22xp33_ASAP7_75t_L g1075 ( 
.A1(n_866),
.A2(n_149),
.B1(n_151),
.B2(n_152),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_908),
.B(n_156),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_912),
.Y(n_1077)
);

BUFx6f_ASAP7_75t_L g1078 ( 
.A(n_884),
.Y(n_1078)
);

NOR2xp33_ASAP7_75t_L g1079 ( 
.A(n_858),
.B(n_932),
.Y(n_1079)
);

O2A1O1Ixp33_ASAP7_75t_L g1080 ( 
.A1(n_918),
.A2(n_923),
.B(n_931),
.C(n_941),
.Y(n_1080)
);

INVx3_ASAP7_75t_L g1081 ( 
.A(n_894),
.Y(n_1081)
);

NAND3xp33_ASAP7_75t_L g1082 ( 
.A(n_967),
.B(n_935),
.C(n_839),
.Y(n_1082)
);

O2A1O1Ixp5_ASAP7_75t_L g1083 ( 
.A1(n_940),
.A2(n_921),
.B(n_878),
.C(n_893),
.Y(n_1083)
);

NAND2x1_ASAP7_75t_L g1084 ( 
.A(n_934),
.B(n_904),
.Y(n_1084)
);

OAI21x1_ASAP7_75t_L g1085 ( 
.A1(n_882),
.A2(n_975),
.B(n_897),
.Y(n_1085)
);

AOI21xp5_ASAP7_75t_L g1086 ( 
.A1(n_951),
.A2(n_921),
.B(n_878),
.Y(n_1086)
);

AND2x2_ASAP7_75t_L g1087 ( 
.A(n_867),
.B(n_873),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_924),
.B(n_942),
.Y(n_1088)
);

NOR3xp33_ASAP7_75t_SL g1089 ( 
.A(n_935),
.B(n_892),
.C(n_955),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_SL g1090 ( 
.A(n_843),
.B(n_909),
.Y(n_1090)
);

NOR2xp33_ASAP7_75t_R g1091 ( 
.A(n_909),
.B(n_843),
.Y(n_1091)
);

AND2x2_ASAP7_75t_L g1092 ( 
.A(n_875),
.B(n_877),
.Y(n_1092)
);

BUFx3_ASAP7_75t_L g1093 ( 
.A(n_936),
.Y(n_1093)
);

NOR2xp33_ASAP7_75t_L g1094 ( 
.A(n_932),
.B(n_953),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_954),
.Y(n_1095)
);

AO32x1_ASAP7_75t_L g1096 ( 
.A1(n_937),
.A2(n_948),
.A3(n_978),
.B1(n_974),
.B2(n_956),
.Y(n_1096)
);

OAI22xp33_ASAP7_75t_L g1097 ( 
.A1(n_969),
.A2(n_957),
.B1(n_944),
.B2(n_953),
.Y(n_1097)
);

AOI22xp5_ASAP7_75t_L g1098 ( 
.A1(n_836),
.A2(n_950),
.B1(n_972),
.B2(n_822),
.Y(n_1098)
);

AOI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_893),
.A2(n_917),
.B(n_933),
.Y(n_1099)
);

BUFx8_ASAP7_75t_L g1100 ( 
.A(n_979),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_962),
.Y(n_1101)
);

AND2x4_ASAP7_75t_L g1102 ( 
.A(n_898),
.B(n_843),
.Y(n_1102)
);

BUFx6f_ASAP7_75t_L g1103 ( 
.A(n_884),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_936),
.B(n_822),
.Y(n_1104)
);

AOI21xp5_ASAP7_75t_L g1105 ( 
.A1(n_917),
.A2(n_933),
.B(n_879),
.Y(n_1105)
);

INVx4_ASAP7_75t_L g1106 ( 
.A(n_884),
.Y(n_1106)
);

OAI21xp33_ASAP7_75t_L g1107 ( 
.A1(n_972),
.A2(n_839),
.B(n_851),
.Y(n_1107)
);

NOR2xp33_ASAP7_75t_L g1108 ( 
.A(n_959),
.B(n_910),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_910),
.B(n_898),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_968),
.B(n_970),
.Y(n_1110)
);

AOI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_879),
.A2(n_916),
.B(n_888),
.Y(n_1111)
);

AOI21xp5_ASAP7_75t_L g1112 ( 
.A1(n_895),
.A2(n_919),
.B(n_920),
.Y(n_1112)
);

NOR2xp33_ASAP7_75t_L g1113 ( 
.A(n_926),
.B(n_976),
.Y(n_1113)
);

O2A1O1Ixp33_ASAP7_75t_L g1114 ( 
.A1(n_914),
.A2(n_868),
.B(n_966),
.C(n_876),
.Y(n_1114)
);

OAI21xp33_ASAP7_75t_SL g1115 ( 
.A1(n_971),
.A2(n_980),
.B(n_841),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_857),
.Y(n_1116)
);

OR2x2_ASAP7_75t_L g1117 ( 
.A(n_965),
.B(n_903),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_890),
.B(n_915),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_915),
.B(n_946),
.Y(n_1119)
);

BUFx2_ASAP7_75t_L g1120 ( 
.A(n_965),
.Y(n_1120)
);

NOR2xp33_ASAP7_75t_L g1121 ( 
.A(n_871),
.B(n_938),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_911),
.Y(n_1122)
);

AOI21xp5_ASAP7_75t_L g1123 ( 
.A1(n_859),
.A2(n_980),
.B(n_971),
.Y(n_1123)
);

OAI21xp33_ASAP7_75t_SL g1124 ( 
.A1(n_907),
.A2(n_922),
.B(n_838),
.Y(n_1124)
);

NOR2xp33_ASAP7_75t_L g1125 ( 
.A(n_865),
.B(n_946),
.Y(n_1125)
);

AO21x1_ASAP7_75t_L g1126 ( 
.A1(n_1007),
.A2(n_913),
.B(n_943),
.Y(n_1126)
);

HB1xp67_ASAP7_75t_L g1127 ( 
.A(n_1031),
.Y(n_1127)
);

OAI21x1_ASAP7_75t_L g1128 ( 
.A1(n_1085),
.A2(n_913),
.B(n_907),
.Y(n_1128)
);

AND2x4_ASAP7_75t_L g1129 ( 
.A(n_1041),
.B(n_902),
.Y(n_1129)
);

AOI21xp5_ASAP7_75t_L g1130 ( 
.A1(n_1001),
.A2(n_854),
.B(n_957),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_SL g1131 ( 
.A(n_1009),
.B(n_979),
.Y(n_1131)
);

AND2x6_ASAP7_75t_L g1132 ( 
.A(n_1009),
.B(n_902),
.Y(n_1132)
);

BUFx8_ASAP7_75t_L g1133 ( 
.A(n_1016),
.Y(n_1133)
);

BUFx3_ASAP7_75t_L g1134 ( 
.A(n_991),
.Y(n_1134)
);

AOI21xp5_ASAP7_75t_L g1135 ( 
.A1(n_1111),
.A2(n_854),
.B(n_957),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_1118),
.B(n_865),
.Y(n_1136)
);

A2O1A1Ixp33_ASAP7_75t_L g1137 ( 
.A1(n_1098),
.A2(n_838),
.B(n_957),
.C(n_944),
.Y(n_1137)
);

OAI21x1_ASAP7_75t_L g1138 ( 
.A1(n_1099),
.A2(n_853),
.B(n_963),
.Y(n_1138)
);

OAI21xp5_ASAP7_75t_L g1139 ( 
.A1(n_1082),
.A2(n_947),
.B(n_952),
.Y(n_1139)
);

INVxp67_ASAP7_75t_L g1140 ( 
.A(n_1035),
.Y(n_1140)
);

AND2x2_ASAP7_75t_L g1141 ( 
.A(n_990),
.B(n_995),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_1113),
.B(n_952),
.Y(n_1142)
);

OAI21x1_ASAP7_75t_L g1143 ( 
.A1(n_1086),
.A2(n_960),
.B(n_949),
.Y(n_1143)
);

INVx3_ASAP7_75t_L g1144 ( 
.A(n_1100),
.Y(n_1144)
);

OAI21x1_ASAP7_75t_L g1145 ( 
.A1(n_1072),
.A2(n_960),
.B(n_949),
.Y(n_1145)
);

AOI21xp5_ASAP7_75t_L g1146 ( 
.A1(n_1002),
.A2(n_854),
.B(n_934),
.Y(n_1146)
);

BUFx12f_ASAP7_75t_L g1147 ( 
.A(n_1011),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_1092),
.B(n_808),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_984),
.Y(n_1149)
);

NOR2xp33_ASAP7_75t_SL g1150 ( 
.A(n_1068),
.B(n_808),
.Y(n_1150)
);

OAI21x1_ASAP7_75t_SL g1151 ( 
.A1(n_982),
.A2(n_958),
.B(n_808),
.Y(n_1151)
);

AO31x2_ASAP7_75t_L g1152 ( 
.A1(n_1018),
.A2(n_1112),
.A3(n_1119),
.B(n_1125),
.Y(n_1152)
);

OAI21xp33_ASAP7_75t_L g1153 ( 
.A1(n_1050),
.A2(n_812),
.B(n_1056),
.Y(n_1153)
);

BUFx2_ASAP7_75t_L g1154 ( 
.A(n_983),
.Y(n_1154)
);

OAI22x1_ASAP7_75t_L g1155 ( 
.A1(n_1056),
.A2(n_812),
.B1(n_1057),
.B2(n_1050),
.Y(n_1155)
);

AOI21xp5_ASAP7_75t_L g1156 ( 
.A1(n_1114),
.A2(n_1107),
.B(n_1012),
.Y(n_1156)
);

AOI21xp5_ASAP7_75t_L g1157 ( 
.A1(n_1107),
.A2(n_1105),
.B(n_992),
.Y(n_1157)
);

OAI21x1_ASAP7_75t_L g1158 ( 
.A1(n_1123),
.A2(n_1083),
.B(n_994),
.Y(n_1158)
);

OAI21x1_ASAP7_75t_L g1159 ( 
.A1(n_1044),
.A2(n_1063),
.B(n_1076),
.Y(n_1159)
);

OAI21x1_ASAP7_75t_L g1160 ( 
.A1(n_1064),
.A2(n_1084),
.B(n_1027),
.Y(n_1160)
);

OAI22xp5_ASAP7_75t_L g1161 ( 
.A1(n_1057),
.A2(n_1046),
.B1(n_989),
.B2(n_1088),
.Y(n_1161)
);

OAI21x1_ASAP7_75t_L g1162 ( 
.A1(n_1065),
.A2(n_1104),
.B(n_1080),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_985),
.Y(n_1163)
);

INVxp67_ASAP7_75t_SL g1164 ( 
.A(n_1094),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_1079),
.B(n_1041),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_L g1166 ( 
.A(n_1037),
.B(n_1053),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_1051),
.B(n_1028),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_987),
.B(n_998),
.Y(n_1168)
);

INVx1_ASAP7_75t_SL g1169 ( 
.A(n_1093),
.Y(n_1169)
);

HB1xp67_ASAP7_75t_L g1170 ( 
.A(n_1074),
.Y(n_1170)
);

AOI221x1_ASAP7_75t_L g1171 ( 
.A1(n_1052),
.A2(n_1061),
.B1(n_1042),
.B2(n_1045),
.C(n_1039),
.Y(n_1171)
);

OAI21x1_ASAP7_75t_SL g1172 ( 
.A1(n_1006),
.A2(n_1109),
.B(n_1015),
.Y(n_1172)
);

OAI21xp5_ASAP7_75t_SL g1173 ( 
.A1(n_1034),
.A2(n_1060),
.B(n_1019),
.Y(n_1173)
);

OAI21x1_ASAP7_75t_L g1174 ( 
.A1(n_1073),
.A2(n_1059),
.B(n_1024),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_SL g1175 ( 
.A(n_996),
.B(n_999),
.Y(n_1175)
);

NOR2xp33_ASAP7_75t_L g1176 ( 
.A(n_983),
.B(n_1000),
.Y(n_1176)
);

CKINVDCx11_ASAP7_75t_R g1177 ( 
.A(n_997),
.Y(n_1177)
);

O2A1O1Ixp5_ASAP7_75t_L g1178 ( 
.A1(n_1066),
.A2(n_988),
.B(n_1023),
.C(n_986),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_SL g1179 ( 
.A(n_996),
.B(n_999),
.Y(n_1179)
);

BUFx3_ASAP7_75t_L g1180 ( 
.A(n_1100),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_1003),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_1008),
.B(n_1077),
.Y(n_1182)
);

O2A1O1Ixp33_ASAP7_75t_SL g1183 ( 
.A1(n_1017),
.A2(n_1090),
.B(n_1069),
.C(n_1067),
.Y(n_1183)
);

OAI21x1_ASAP7_75t_SL g1184 ( 
.A1(n_1006),
.A2(n_1058),
.B(n_1043),
.Y(n_1184)
);

OAI21x1_ASAP7_75t_L g1185 ( 
.A1(n_1110),
.A2(n_1070),
.B(n_1071),
.Y(n_1185)
);

OAI21x1_ASAP7_75t_L g1186 ( 
.A1(n_1095),
.A2(n_1101),
.B(n_1117),
.Y(n_1186)
);

BUFx6f_ASAP7_75t_L g1187 ( 
.A(n_1000),
.Y(n_1187)
);

AOI21x1_ASAP7_75t_L g1188 ( 
.A1(n_1120),
.A2(n_1013),
.B(n_1030),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_1022),
.B(n_1062),
.Y(n_1189)
);

INVx5_ASAP7_75t_L g1190 ( 
.A(n_1000),
.Y(n_1190)
);

INVx2_ASAP7_75t_SL g1191 ( 
.A(n_1025),
.Y(n_1191)
);

INVx5_ASAP7_75t_L g1192 ( 
.A(n_1025),
.Y(n_1192)
);

AO31x2_ASAP7_75t_L g1193 ( 
.A1(n_1121),
.A2(n_1096),
.A3(n_1122),
.B(n_1116),
.Y(n_1193)
);

O2A1O1Ixp5_ASAP7_75t_L g1194 ( 
.A1(n_1036),
.A2(n_1108),
.B(n_1033),
.C(n_1038),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_SL g1195 ( 
.A(n_1091),
.B(n_993),
.Y(n_1195)
);

OAI21x1_ASAP7_75t_L g1196 ( 
.A1(n_1081),
.A2(n_1089),
.B(n_1075),
.Y(n_1196)
);

OAI21xp5_ASAP7_75t_SL g1197 ( 
.A1(n_1029),
.A2(n_1021),
.B(n_1055),
.Y(n_1197)
);

OAI21x1_ASAP7_75t_SL g1198 ( 
.A1(n_1106),
.A2(n_1021),
.B(n_1124),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_L g1199 ( 
.A(n_1025),
.B(n_1032),
.Y(n_1199)
);

O2A1O1Ixp5_ASAP7_75t_L g1200 ( 
.A1(n_1097),
.A2(n_1102),
.B(n_1047),
.C(n_1087),
.Y(n_1200)
);

AOI21xp5_ASAP7_75t_L g1201 ( 
.A1(n_1115),
.A2(n_1124),
.B(n_1096),
.Y(n_1201)
);

OR2x2_ASAP7_75t_L g1202 ( 
.A(n_1102),
.B(n_1026),
.Y(n_1202)
);

AOI21xp5_ASAP7_75t_L g1203 ( 
.A1(n_1115),
.A2(n_1096),
.B(n_1048),
.Y(n_1203)
);

HB1xp67_ASAP7_75t_L g1204 ( 
.A(n_1078),
.Y(n_1204)
);

AO31x2_ASAP7_75t_L g1205 ( 
.A1(n_1048),
.A2(n_1020),
.A3(n_1010),
.B(n_1078),
.Y(n_1205)
);

CKINVDCx5p33_ASAP7_75t_R g1206 ( 
.A(n_1014),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_1078),
.B(n_1103),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_1103),
.B(n_1047),
.Y(n_1208)
);

AOI221xp5_ASAP7_75t_L g1209 ( 
.A1(n_1049),
.A2(n_672),
.B1(n_723),
.B2(n_489),
.C(n_435),
.Y(n_1209)
);

OAI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_1103),
.A2(n_1082),
.B(n_816),
.Y(n_1210)
);

AO21x1_ASAP7_75t_L g1211 ( 
.A1(n_1007),
.A2(n_672),
.B(n_1005),
.Y(n_1211)
);

OAI21xp5_ASAP7_75t_L g1212 ( 
.A1(n_1082),
.A2(n_816),
.B(n_869),
.Y(n_1212)
);

O2A1O1Ixp5_ASAP7_75t_L g1213 ( 
.A1(n_1054),
.A2(n_672),
.B(n_930),
.C(n_1012),
.Y(n_1213)
);

INVx1_ASAP7_75t_SL g1214 ( 
.A(n_1016),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_1118),
.B(n_1009),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_1092),
.B(n_672),
.Y(n_1216)
);

AND2x2_ASAP7_75t_L g1217 ( 
.A(n_990),
.B(n_814),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_L g1218 ( 
.A(n_1092),
.B(n_672),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_SL g1219 ( 
.A(n_1009),
.B(n_869),
.Y(n_1219)
);

INVx3_ASAP7_75t_L g1220 ( 
.A(n_1100),
.Y(n_1220)
);

INVxp67_ASAP7_75t_L g1221 ( 
.A(n_1031),
.Y(n_1221)
);

INVx3_ASAP7_75t_L g1222 ( 
.A(n_1100),
.Y(n_1222)
);

NOR4xp25_ASAP7_75t_L g1223 ( 
.A(n_1048),
.B(n_1052),
.C(n_869),
.D(n_855),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_L g1224 ( 
.A(n_1092),
.B(n_672),
.Y(n_1224)
);

NOR2x1_ASAP7_75t_SL g1225 ( 
.A(n_996),
.B(n_965),
.Y(n_1225)
);

NOR2xp33_ASAP7_75t_L g1226 ( 
.A(n_991),
.B(n_672),
.Y(n_1226)
);

AO21x1_ASAP7_75t_L g1227 ( 
.A1(n_1007),
.A2(n_672),
.B(n_1005),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_984),
.Y(n_1228)
);

OAI22xp5_ASAP7_75t_L g1229 ( 
.A1(n_1098),
.A2(n_672),
.B1(n_821),
.B2(n_869),
.Y(n_1229)
);

AOI21xp5_ASAP7_75t_L g1230 ( 
.A1(n_1001),
.A2(n_826),
.B(n_825),
.Y(n_1230)
);

CKINVDCx5p33_ASAP7_75t_R g1231 ( 
.A(n_1011),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_1092),
.B(n_672),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_L g1233 ( 
.A(n_1092),
.B(n_672),
.Y(n_1233)
);

NAND2xp33_ASAP7_75t_R g1234 ( 
.A(n_1091),
.B(n_566),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_1092),
.B(n_672),
.Y(n_1235)
);

OAI21xp33_ASAP7_75t_SL g1236 ( 
.A1(n_1050),
.A2(n_1057),
.B(n_1056),
.Y(n_1236)
);

AND2x4_ASAP7_75t_L g1237 ( 
.A(n_1041),
.B(n_835),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_1118),
.B(n_1009),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_984),
.Y(n_1239)
);

OAI21x1_ASAP7_75t_SL g1240 ( 
.A1(n_1005),
.A2(n_982),
.B(n_1004),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_L g1241 ( 
.A(n_1118),
.B(n_1009),
.Y(n_1241)
);

OAI21x1_ASAP7_75t_L g1242 ( 
.A1(n_1085),
.A2(n_1099),
.B(n_1086),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_L g1243 ( 
.A(n_1118),
.B(n_1009),
.Y(n_1243)
);

BUFx6f_ASAP7_75t_L g1244 ( 
.A(n_983),
.Y(n_1244)
);

AOI21xp33_ASAP7_75t_L g1245 ( 
.A1(n_1098),
.A2(n_672),
.B(n_869),
.Y(n_1245)
);

OAI21x1_ASAP7_75t_L g1246 ( 
.A1(n_1085),
.A2(n_1099),
.B(n_1086),
.Y(n_1246)
);

AOI21xp5_ASAP7_75t_L g1247 ( 
.A1(n_1001),
.A2(n_826),
.B(n_825),
.Y(n_1247)
);

OAI21x1_ASAP7_75t_L g1248 ( 
.A1(n_1085),
.A2(n_1099),
.B(n_1086),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_L g1249 ( 
.A(n_1118),
.B(n_1009),
.Y(n_1249)
);

OR2x2_ASAP7_75t_L g1250 ( 
.A(n_990),
.B(n_844),
.Y(n_1250)
);

OAI21x1_ASAP7_75t_L g1251 ( 
.A1(n_1085),
.A2(n_1099),
.B(n_1086),
.Y(n_1251)
);

O2A1O1Ixp33_ASAP7_75t_L g1252 ( 
.A1(n_1040),
.A2(n_672),
.B(n_869),
.C(n_855),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_984),
.Y(n_1253)
);

NOR3xp33_ASAP7_75t_L g1254 ( 
.A(n_1052),
.B(n_672),
.C(n_869),
.Y(n_1254)
);

AOI21xp5_ASAP7_75t_L g1255 ( 
.A1(n_1001),
.A2(n_826),
.B(n_825),
.Y(n_1255)
);

A2O1A1Ixp33_ASAP7_75t_L g1256 ( 
.A1(n_1098),
.A2(n_869),
.B(n_855),
.C(n_672),
.Y(n_1256)
);

OAI22xp5_ASAP7_75t_L g1257 ( 
.A1(n_1098),
.A2(n_672),
.B1(n_821),
.B2(n_869),
.Y(n_1257)
);

OAI21x1_ASAP7_75t_L g1258 ( 
.A1(n_1085),
.A2(n_1099),
.B(n_1086),
.Y(n_1258)
);

INVx2_ASAP7_75t_SL g1259 ( 
.A(n_991),
.Y(n_1259)
);

INVx3_ASAP7_75t_L g1260 ( 
.A(n_1100),
.Y(n_1260)
);

A2O1A1Ixp33_ASAP7_75t_L g1261 ( 
.A1(n_1098),
.A2(n_869),
.B(n_855),
.C(n_672),
.Y(n_1261)
);

AO31x2_ASAP7_75t_L g1262 ( 
.A1(n_1018),
.A2(n_1112),
.A3(n_1111),
.B(n_1072),
.Y(n_1262)
);

NOR2xp33_ASAP7_75t_L g1263 ( 
.A(n_991),
.B(n_672),
.Y(n_1263)
);

OAI21xp5_ASAP7_75t_L g1264 ( 
.A1(n_1082),
.A2(n_816),
.B(n_869),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_L g1265 ( 
.A(n_1092),
.B(n_672),
.Y(n_1265)
);

CKINVDCx20_ASAP7_75t_R g1266 ( 
.A(n_1011),
.Y(n_1266)
);

AOI21xp5_ASAP7_75t_L g1267 ( 
.A1(n_1001),
.A2(n_826),
.B(n_825),
.Y(n_1267)
);

A2O1A1Ixp33_ASAP7_75t_L g1268 ( 
.A1(n_1098),
.A2(n_869),
.B(n_855),
.C(n_672),
.Y(n_1268)
);

INVx2_ASAP7_75t_SL g1269 ( 
.A(n_1180),
.Y(n_1269)
);

AND2x4_ASAP7_75t_L g1270 ( 
.A(n_1131),
.B(n_1132),
.Y(n_1270)
);

OAI221xp5_ASAP7_75t_L g1271 ( 
.A1(n_1209),
.A2(n_1236),
.B1(n_1173),
.B2(n_1197),
.C(n_1245),
.Y(n_1271)
);

A2O1A1Ixp33_ASAP7_75t_L g1272 ( 
.A1(n_1245),
.A2(n_1268),
.B(n_1256),
.C(n_1261),
.Y(n_1272)
);

AO31x2_ASAP7_75t_L g1273 ( 
.A1(n_1203),
.A2(n_1201),
.A3(n_1227),
.B(n_1211),
.Y(n_1273)
);

AO32x2_ASAP7_75t_L g1274 ( 
.A1(n_1229),
.A2(n_1257),
.A3(n_1161),
.B1(n_1223),
.B2(n_1191),
.Y(n_1274)
);

AOI22xp33_ASAP7_75t_L g1275 ( 
.A1(n_1229),
.A2(n_1257),
.B1(n_1155),
.B2(n_1254),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1168),
.Y(n_1276)
);

AOI21x1_ASAP7_75t_L g1277 ( 
.A1(n_1156),
.A2(n_1157),
.B(n_1188),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1182),
.Y(n_1278)
);

OAI21x1_ASAP7_75t_L g1279 ( 
.A1(n_1158),
.A2(n_1246),
.B(n_1242),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1189),
.Y(n_1280)
);

OAI21x1_ASAP7_75t_L g1281 ( 
.A1(n_1248),
.A2(n_1258),
.B(n_1251),
.Y(n_1281)
);

OAI221xp5_ASAP7_75t_L g1282 ( 
.A1(n_1173),
.A2(n_1197),
.B1(n_1252),
.B2(n_1223),
.C(n_1167),
.Y(n_1282)
);

OAI21x1_ASAP7_75t_SL g1283 ( 
.A1(n_1212),
.A2(n_1264),
.B(n_1198),
.Y(n_1283)
);

OAI21x1_ASAP7_75t_SL g1284 ( 
.A1(n_1212),
.A2(n_1264),
.B(n_1184),
.Y(n_1284)
);

O2A1O1Ixp33_ASAP7_75t_L g1285 ( 
.A1(n_1161),
.A2(n_1226),
.B(n_1263),
.C(n_1265),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1149),
.Y(n_1286)
);

OAI21x1_ASAP7_75t_L g1287 ( 
.A1(n_1240),
.A2(n_1128),
.B(n_1159),
.Y(n_1287)
);

OAI222xp33_ASAP7_75t_L g1288 ( 
.A1(n_1219),
.A2(n_1241),
.B1(n_1249),
.B2(n_1215),
.C1(n_1243),
.C2(n_1238),
.Y(n_1288)
);

BUFx2_ASAP7_75t_L g1289 ( 
.A(n_1133),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_L g1290 ( 
.A(n_1216),
.B(n_1218),
.Y(n_1290)
);

OAI21x1_ASAP7_75t_L g1291 ( 
.A1(n_1145),
.A2(n_1143),
.B(n_1138),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1163),
.Y(n_1292)
);

AOI22xp33_ASAP7_75t_L g1293 ( 
.A1(n_1153),
.A2(n_1215),
.B1(n_1249),
.B2(n_1243),
.Y(n_1293)
);

BUFx3_ASAP7_75t_L g1294 ( 
.A(n_1134),
.Y(n_1294)
);

OR2x2_ASAP7_75t_L g1295 ( 
.A(n_1164),
.B(n_1250),
.Y(n_1295)
);

OAI21x1_ASAP7_75t_L g1296 ( 
.A1(n_1135),
.A2(n_1146),
.B(n_1130),
.Y(n_1296)
);

NAND2x1p5_ASAP7_75t_L g1297 ( 
.A(n_1190),
.B(n_1192),
.Y(n_1297)
);

BUFx2_ASAP7_75t_L g1298 ( 
.A(n_1133),
.Y(n_1298)
);

AND2x2_ASAP7_75t_SL g1299 ( 
.A(n_1150),
.B(n_1238),
.Y(n_1299)
);

CKINVDCx20_ASAP7_75t_R g1300 ( 
.A(n_1266),
.Y(n_1300)
);

O2A1O1Ixp33_ASAP7_75t_L g1301 ( 
.A1(n_1224),
.A2(n_1232),
.B(n_1233),
.C(n_1235),
.Y(n_1301)
);

OAI21x1_ASAP7_75t_L g1302 ( 
.A1(n_1230),
.A2(n_1267),
.B(n_1255),
.Y(n_1302)
);

AO21x2_ASAP7_75t_L g1303 ( 
.A1(n_1172),
.A2(n_1151),
.B(n_1137),
.Y(n_1303)
);

OAI21x1_ASAP7_75t_L g1304 ( 
.A1(n_1247),
.A2(n_1196),
.B(n_1210),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1181),
.Y(n_1305)
);

OAI21xp5_ASAP7_75t_L g1306 ( 
.A1(n_1213),
.A2(n_1162),
.B(n_1171),
.Y(n_1306)
);

AND2x4_ASAP7_75t_L g1307 ( 
.A(n_1132),
.B(n_1225),
.Y(n_1307)
);

OAI21xp5_ASAP7_75t_L g1308 ( 
.A1(n_1178),
.A2(n_1210),
.B(n_1185),
.Y(n_1308)
);

OAI21x1_ASAP7_75t_L g1309 ( 
.A1(n_1160),
.A2(n_1174),
.B(n_1139),
.Y(n_1309)
);

AOI21x1_ASAP7_75t_L g1310 ( 
.A1(n_1126),
.A2(n_1142),
.B(n_1136),
.Y(n_1310)
);

INVxp67_ASAP7_75t_L g1311 ( 
.A(n_1127),
.Y(n_1311)
);

O2A1O1Ixp33_ASAP7_75t_L g1312 ( 
.A1(n_1183),
.A2(n_1214),
.B(n_1195),
.C(n_1165),
.Y(n_1312)
);

OAI21x1_ASAP7_75t_L g1313 ( 
.A1(n_1136),
.A2(n_1186),
.B(n_1142),
.Y(n_1313)
);

CKINVDCx5p33_ASAP7_75t_R g1314 ( 
.A(n_1234),
.Y(n_1314)
);

OAI21x1_ASAP7_75t_L g1315 ( 
.A1(n_1200),
.A2(n_1241),
.B(n_1207),
.Y(n_1315)
);

OR2x6_ASAP7_75t_L g1316 ( 
.A(n_1199),
.B(n_1202),
.Y(n_1316)
);

OAI21xp33_ASAP7_75t_SL g1317 ( 
.A1(n_1175),
.A2(n_1179),
.B(n_1150),
.Y(n_1317)
);

OAI21xp5_ASAP7_75t_L g1318 ( 
.A1(n_1194),
.A2(n_1140),
.B(n_1221),
.Y(n_1318)
);

INVxp67_ASAP7_75t_L g1319 ( 
.A(n_1170),
.Y(n_1319)
);

OAI21x1_ASAP7_75t_L g1320 ( 
.A1(n_1228),
.A2(n_1253),
.B(n_1239),
.Y(n_1320)
);

AOI21x1_ASAP7_75t_L g1321 ( 
.A1(n_1204),
.A2(n_1148),
.B(n_1217),
.Y(n_1321)
);

AO21x1_ASAP7_75t_L g1322 ( 
.A1(n_1166),
.A2(n_1141),
.B(n_1208),
.Y(n_1322)
);

OAI21x1_ASAP7_75t_L g1323 ( 
.A1(n_1262),
.A2(n_1208),
.B(n_1222),
.Y(n_1323)
);

A2O1A1Ixp33_ASAP7_75t_L g1324 ( 
.A1(n_1206),
.A2(n_1129),
.B(n_1237),
.C(n_1176),
.Y(n_1324)
);

AO31x2_ASAP7_75t_L g1325 ( 
.A1(n_1152),
.A2(n_1262),
.A3(n_1193),
.B(n_1154),
.Y(n_1325)
);

AO21x2_ASAP7_75t_L g1326 ( 
.A1(n_1152),
.A2(n_1262),
.B(n_1193),
.Y(n_1326)
);

HB1xp67_ASAP7_75t_L g1327 ( 
.A(n_1152),
.Y(n_1327)
);

HB1xp67_ASAP7_75t_L g1328 ( 
.A(n_1205),
.Y(n_1328)
);

OAI21xp5_ASAP7_75t_L g1329 ( 
.A1(n_1259),
.A2(n_1169),
.B(n_1237),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1205),
.Y(n_1330)
);

BUFx2_ASAP7_75t_L g1331 ( 
.A(n_1144),
.Y(n_1331)
);

NAND2x1p5_ASAP7_75t_L g1332 ( 
.A(n_1190),
.B(n_1192),
.Y(n_1332)
);

BUFx3_ASAP7_75t_L g1333 ( 
.A(n_1187),
.Y(n_1333)
);

CKINVDCx6p67_ASAP7_75t_R g1334 ( 
.A(n_1147),
.Y(n_1334)
);

BUFx12f_ASAP7_75t_L g1335 ( 
.A(n_1177),
.Y(n_1335)
);

AO21x2_ASAP7_75t_L g1336 ( 
.A1(n_1132),
.A2(n_1190),
.B(n_1192),
.Y(n_1336)
);

OAI21x1_ASAP7_75t_L g1337 ( 
.A1(n_1220),
.A2(n_1222),
.B(n_1260),
.Y(n_1337)
);

A2O1A1Ixp33_ASAP7_75t_L g1338 ( 
.A1(n_1220),
.A2(n_869),
.B(n_1236),
.C(n_855),
.Y(n_1338)
);

OAI21x1_ASAP7_75t_L g1339 ( 
.A1(n_1244),
.A2(n_1246),
.B(n_1242),
.Y(n_1339)
);

AO21x2_ASAP7_75t_L g1340 ( 
.A1(n_1244),
.A2(n_1156),
.B(n_1172),
.Y(n_1340)
);

NOR2xp33_ASAP7_75t_L g1341 ( 
.A(n_1244),
.B(n_1231),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1168),
.Y(n_1342)
);

BUFx3_ASAP7_75t_L g1343 ( 
.A(n_1134),
.Y(n_1343)
);

NAND3xp33_ASAP7_75t_L g1344 ( 
.A(n_1209),
.B(n_672),
.C(n_869),
.Y(n_1344)
);

OA21x2_ASAP7_75t_L g1345 ( 
.A1(n_1157),
.A2(n_1203),
.B(n_1156),
.Y(n_1345)
);

NAND2xp5_ASAP7_75t_L g1346 ( 
.A(n_1216),
.B(n_1218),
.Y(n_1346)
);

INVx2_ASAP7_75t_SL g1347 ( 
.A(n_1180),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1168),
.Y(n_1348)
);

OR2x6_ASAP7_75t_L g1349 ( 
.A(n_1131),
.B(n_1155),
.Y(n_1349)
);

CKINVDCx8_ASAP7_75t_R g1350 ( 
.A(n_1231),
.Y(n_1350)
);

OR2x6_ASAP7_75t_L g1351 ( 
.A(n_1131),
.B(n_1155),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1168),
.Y(n_1352)
);

OAI22xp5_ASAP7_75t_L g1353 ( 
.A1(n_1209),
.A2(n_672),
.B1(n_869),
.B2(n_1226),
.Y(n_1353)
);

BUFx3_ASAP7_75t_L g1354 ( 
.A(n_1134),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1168),
.Y(n_1355)
);

OR2x2_ASAP7_75t_L g1356 ( 
.A(n_1164),
.B(n_1250),
.Y(n_1356)
);

O2A1O1Ixp33_ASAP7_75t_L g1357 ( 
.A1(n_1256),
.A2(n_672),
.B(n_869),
.C(n_855),
.Y(n_1357)
);

OR2x2_ASAP7_75t_L g1358 ( 
.A(n_1164),
.B(n_1250),
.Y(n_1358)
);

OAI21x1_ASAP7_75t_L g1359 ( 
.A1(n_1242),
.A2(n_1248),
.B(n_1246),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_SL g1360 ( 
.A(n_1229),
.B(n_1257),
.Y(n_1360)
);

CKINVDCx5p33_ASAP7_75t_R g1361 ( 
.A(n_1234),
.Y(n_1361)
);

AOI221xp5_ASAP7_75t_L g1362 ( 
.A1(n_1236),
.A2(n_672),
.B1(n_723),
.B2(n_869),
.C(n_489),
.Y(n_1362)
);

AND2x4_ASAP7_75t_L g1363 ( 
.A(n_1131),
.B(n_1132),
.Y(n_1363)
);

AOI22xp33_ASAP7_75t_L g1364 ( 
.A1(n_1236),
.A2(n_1021),
.B1(n_1257),
.B2(n_1229),
.Y(n_1364)
);

OAI21x1_ASAP7_75t_L g1365 ( 
.A1(n_1242),
.A2(n_1248),
.B(n_1246),
.Y(n_1365)
);

OAI22xp5_ASAP7_75t_L g1366 ( 
.A1(n_1209),
.A2(n_672),
.B1(n_869),
.B2(n_1226),
.Y(n_1366)
);

AOI21xp5_ASAP7_75t_L g1367 ( 
.A1(n_1157),
.A2(n_1267),
.B(n_1247),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_L g1368 ( 
.A(n_1216),
.B(n_1218),
.Y(n_1368)
);

OR2x2_ASAP7_75t_L g1369 ( 
.A(n_1164),
.B(n_1250),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1216),
.B(n_1218),
.Y(n_1370)
);

OAI21x1_ASAP7_75t_L g1371 ( 
.A1(n_1242),
.A2(n_1248),
.B(n_1246),
.Y(n_1371)
);

OAI21xp5_ASAP7_75t_L g1372 ( 
.A1(n_1209),
.A2(n_672),
.B(n_869),
.Y(n_1372)
);

BUFx3_ASAP7_75t_L g1373 ( 
.A(n_1134),
.Y(n_1373)
);

A2O1A1Ixp33_ASAP7_75t_L g1374 ( 
.A1(n_1236),
.A2(n_869),
.B(n_855),
.C(n_1245),
.Y(n_1374)
);

OAI21x1_ASAP7_75t_L g1375 ( 
.A1(n_1158),
.A2(n_1246),
.B(n_1242),
.Y(n_1375)
);

OAI21x1_ASAP7_75t_L g1376 ( 
.A1(n_1158),
.A2(n_1246),
.B(n_1242),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1168),
.Y(n_1377)
);

NOR2xp33_ASAP7_75t_L g1378 ( 
.A(n_1226),
.B(n_869),
.Y(n_1378)
);

O2A1O1Ixp33_ASAP7_75t_L g1379 ( 
.A1(n_1256),
.A2(n_672),
.B(n_869),
.C(n_855),
.Y(n_1379)
);

BUFx2_ASAP7_75t_L g1380 ( 
.A(n_1133),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1168),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_L g1382 ( 
.A(n_1216),
.B(n_1218),
.Y(n_1382)
);

OAI21x1_ASAP7_75t_L g1383 ( 
.A1(n_1242),
.A2(n_1248),
.B(n_1246),
.Y(n_1383)
);

AO21x1_ASAP7_75t_L g1384 ( 
.A1(n_1229),
.A2(n_1257),
.B(n_1245),
.Y(n_1384)
);

AND2x2_ASAP7_75t_L g1385 ( 
.A(n_1217),
.B(n_1226),
.Y(n_1385)
);

OAI22xp5_ASAP7_75t_L g1386 ( 
.A1(n_1209),
.A2(n_672),
.B1(n_869),
.B2(n_1226),
.Y(n_1386)
);

AND2x2_ASAP7_75t_L g1387 ( 
.A(n_1217),
.B(n_1226),
.Y(n_1387)
);

OAI21x1_ASAP7_75t_L g1388 ( 
.A1(n_1242),
.A2(n_1248),
.B(n_1246),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_L g1389 ( 
.A(n_1295),
.B(n_1356),
.Y(n_1389)
);

OR2x2_ASAP7_75t_L g1390 ( 
.A(n_1358),
.B(n_1369),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_1276),
.B(n_1278),
.Y(n_1391)
);

AOI21xp5_ASAP7_75t_L g1392 ( 
.A1(n_1367),
.A2(n_1360),
.B(n_1272),
.Y(n_1392)
);

OAI22xp5_ASAP7_75t_L g1393 ( 
.A1(n_1364),
.A2(n_1362),
.B1(n_1271),
.B2(n_1344),
.Y(n_1393)
);

AOI21xp5_ASAP7_75t_SL g1394 ( 
.A1(n_1374),
.A2(n_1360),
.B(n_1357),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1320),
.Y(n_1395)
);

CKINVDCx14_ASAP7_75t_R g1396 ( 
.A(n_1300),
.Y(n_1396)
);

AND2x2_ASAP7_75t_L g1397 ( 
.A(n_1385),
.B(n_1387),
.Y(n_1397)
);

AOI21xp5_ASAP7_75t_SL g1398 ( 
.A1(n_1374),
.A2(n_1379),
.B(n_1338),
.Y(n_1398)
);

AND2x2_ASAP7_75t_L g1399 ( 
.A(n_1378),
.B(n_1319),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1320),
.Y(n_1400)
);

AOI21xp5_ASAP7_75t_SL g1401 ( 
.A1(n_1338),
.A2(n_1272),
.B(n_1324),
.Y(n_1401)
);

O2A1O1Ixp5_ASAP7_75t_L g1402 ( 
.A1(n_1372),
.A2(n_1384),
.B(n_1386),
.C(n_1366),
.Y(n_1402)
);

OR2x2_ASAP7_75t_L g1403 ( 
.A(n_1311),
.B(n_1286),
.Y(n_1403)
);

AND2x2_ASAP7_75t_L g1404 ( 
.A(n_1378),
.B(n_1329),
.Y(n_1404)
);

AND2x2_ASAP7_75t_L g1405 ( 
.A(n_1364),
.B(n_1280),
.Y(n_1405)
);

AND2x2_ASAP7_75t_L g1406 ( 
.A(n_1342),
.B(n_1348),
.Y(n_1406)
);

OA21x2_ASAP7_75t_L g1407 ( 
.A1(n_1302),
.A2(n_1306),
.B(n_1308),
.Y(n_1407)
);

AND2x2_ASAP7_75t_L g1408 ( 
.A(n_1274),
.B(n_1292),
.Y(n_1408)
);

NAND2xp5_ASAP7_75t_L g1409 ( 
.A(n_1352),
.B(n_1355),
.Y(n_1409)
);

CKINVDCx16_ASAP7_75t_R g1410 ( 
.A(n_1300),
.Y(n_1410)
);

AND2x4_ASAP7_75t_L g1411 ( 
.A(n_1323),
.B(n_1307),
.Y(n_1411)
);

OA21x2_ASAP7_75t_L g1412 ( 
.A1(n_1302),
.A2(n_1304),
.B(n_1375),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_L g1413 ( 
.A(n_1377),
.B(n_1381),
.Y(n_1413)
);

O2A1O1Ixp33_ASAP7_75t_L g1414 ( 
.A1(n_1353),
.A2(n_1282),
.B(n_1285),
.C(n_1275),
.Y(n_1414)
);

AND2x2_ASAP7_75t_L g1415 ( 
.A(n_1331),
.B(n_1305),
.Y(n_1415)
);

INVx3_ASAP7_75t_L g1416 ( 
.A(n_1340),
.Y(n_1416)
);

OA21x2_ASAP7_75t_L g1417 ( 
.A1(n_1304),
.A2(n_1279),
.B(n_1376),
.Y(n_1417)
);

AOI21xp5_ASAP7_75t_L g1418 ( 
.A1(n_1275),
.A2(n_1296),
.B(n_1345),
.Y(n_1418)
);

AND2x2_ASAP7_75t_L g1419 ( 
.A(n_1274),
.B(n_1325),
.Y(n_1419)
);

AOI21xp5_ASAP7_75t_SL g1420 ( 
.A1(n_1324),
.A2(n_1312),
.B(n_1336),
.Y(n_1420)
);

OA21x2_ASAP7_75t_L g1421 ( 
.A1(n_1281),
.A2(n_1388),
.B(n_1383),
.Y(n_1421)
);

OA21x2_ASAP7_75t_L g1422 ( 
.A1(n_1281),
.A2(n_1365),
.B(n_1371),
.Y(n_1422)
);

NAND2xp5_ASAP7_75t_L g1423 ( 
.A(n_1290),
.B(n_1346),
.Y(n_1423)
);

OAI22xp5_ASAP7_75t_L g1424 ( 
.A1(n_1368),
.A2(n_1382),
.B1(n_1370),
.B2(n_1293),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1313),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_L g1426 ( 
.A(n_1301),
.B(n_1293),
.Y(n_1426)
);

AND2x2_ASAP7_75t_L g1427 ( 
.A(n_1318),
.B(n_1316),
.Y(n_1427)
);

AOI21xp5_ASAP7_75t_L g1428 ( 
.A1(n_1345),
.A2(n_1299),
.B(n_1284),
.Y(n_1428)
);

INVx3_ASAP7_75t_L g1429 ( 
.A(n_1340),
.Y(n_1429)
);

AND2x2_ASAP7_75t_L g1430 ( 
.A(n_1274),
.B(n_1325),
.Y(n_1430)
);

OR2x2_ASAP7_75t_L g1431 ( 
.A(n_1316),
.B(n_1349),
.Y(n_1431)
);

AOI21x1_ASAP7_75t_SL g1432 ( 
.A1(n_1327),
.A2(n_1274),
.B(n_1334),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_L g1433 ( 
.A(n_1343),
.B(n_1354),
.Y(n_1433)
);

BUFx3_ASAP7_75t_L g1434 ( 
.A(n_1354),
.Y(n_1434)
);

O2A1O1Ixp33_ASAP7_75t_L g1435 ( 
.A1(n_1283),
.A2(n_1269),
.B(n_1347),
.C(n_1288),
.Y(n_1435)
);

AND2x2_ASAP7_75t_L g1436 ( 
.A(n_1373),
.B(n_1337),
.Y(n_1436)
);

O2A1O1Ixp33_ASAP7_75t_L g1437 ( 
.A1(n_1341),
.A2(n_1327),
.B(n_1317),
.C(n_1380),
.Y(n_1437)
);

AND2x2_ASAP7_75t_L g1438 ( 
.A(n_1326),
.B(n_1273),
.Y(n_1438)
);

OAI22xp5_ASAP7_75t_L g1439 ( 
.A1(n_1314),
.A2(n_1361),
.B1(n_1351),
.B2(n_1349),
.Y(n_1439)
);

AOI21xp5_ASAP7_75t_SL g1440 ( 
.A1(n_1336),
.A2(n_1307),
.B(n_1332),
.Y(n_1440)
);

AOI21xp5_ASAP7_75t_SL g1441 ( 
.A1(n_1297),
.A2(n_1332),
.B(n_1303),
.Y(n_1441)
);

OAI22xp5_ASAP7_75t_L g1442 ( 
.A1(n_1349),
.A2(n_1351),
.B1(n_1298),
.B2(n_1289),
.Y(n_1442)
);

AND2x2_ASAP7_75t_L g1443 ( 
.A(n_1337),
.B(n_1333),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_L g1444 ( 
.A(n_1322),
.B(n_1321),
.Y(n_1444)
);

BUFx12f_ASAP7_75t_L g1445 ( 
.A(n_1335),
.Y(n_1445)
);

A2O1A1Ixp33_ASAP7_75t_L g1446 ( 
.A1(n_1328),
.A2(n_1315),
.B(n_1363),
.C(n_1270),
.Y(n_1446)
);

A2O1A1Ixp33_ASAP7_75t_L g1447 ( 
.A1(n_1328),
.A2(n_1315),
.B(n_1363),
.C(n_1270),
.Y(n_1447)
);

OA21x2_ASAP7_75t_L g1448 ( 
.A1(n_1359),
.A2(n_1291),
.B(n_1287),
.Y(n_1448)
);

INVx3_ASAP7_75t_L g1449 ( 
.A(n_1273),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1310),
.Y(n_1450)
);

OAI22xp5_ASAP7_75t_L g1451 ( 
.A1(n_1350),
.A2(n_1297),
.B1(n_1277),
.B2(n_1330),
.Y(n_1451)
);

HB1xp67_ASAP7_75t_L g1452 ( 
.A(n_1339),
.Y(n_1452)
);

AND2x2_ASAP7_75t_L g1453 ( 
.A(n_1309),
.B(n_1274),
.Y(n_1453)
);

BUFx2_ASAP7_75t_L g1454 ( 
.A(n_1294),
.Y(n_1454)
);

O2A1O1Ixp33_ASAP7_75t_L g1455 ( 
.A1(n_1353),
.A2(n_672),
.B(n_1386),
.C(n_1366),
.Y(n_1455)
);

NAND2xp5_ASAP7_75t_L g1456 ( 
.A(n_1295),
.B(n_1164),
.Y(n_1456)
);

OAI22xp5_ASAP7_75t_L g1457 ( 
.A1(n_1364),
.A2(n_1362),
.B1(n_1271),
.B2(n_1344),
.Y(n_1457)
);

OAI22xp5_ASAP7_75t_L g1458 ( 
.A1(n_1364),
.A2(n_1362),
.B1(n_1271),
.B2(n_1344),
.Y(n_1458)
);

O2A1O1Ixp33_ASAP7_75t_L g1459 ( 
.A1(n_1353),
.A2(n_672),
.B(n_1386),
.C(n_1366),
.Y(n_1459)
);

INVx1_ASAP7_75t_SL g1460 ( 
.A(n_1294),
.Y(n_1460)
);

A2O1A1Ixp33_ASAP7_75t_L g1461 ( 
.A1(n_1362),
.A2(n_1236),
.B(n_869),
.C(n_855),
.Y(n_1461)
);

INVx2_ASAP7_75t_L g1462 ( 
.A(n_1313),
.Y(n_1462)
);

OR2x2_ASAP7_75t_L g1463 ( 
.A(n_1295),
.B(n_1356),
.Y(n_1463)
);

AND2x2_ASAP7_75t_L g1464 ( 
.A(n_1385),
.B(n_1387),
.Y(n_1464)
);

BUFx2_ASAP7_75t_L g1465 ( 
.A(n_1411),
.Y(n_1465)
);

OR2x2_ASAP7_75t_L g1466 ( 
.A(n_1390),
.B(n_1463),
.Y(n_1466)
);

NAND2xp5_ASAP7_75t_L g1467 ( 
.A(n_1408),
.B(n_1392),
.Y(n_1467)
);

OR2x2_ASAP7_75t_L g1468 ( 
.A(n_1389),
.B(n_1408),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_L g1469 ( 
.A(n_1419),
.B(n_1430),
.Y(n_1469)
);

HB1xp67_ASAP7_75t_L g1470 ( 
.A(n_1415),
.Y(n_1470)
);

AO21x2_ASAP7_75t_L g1471 ( 
.A1(n_1418),
.A2(n_1444),
.B(n_1450),
.Y(n_1471)
);

HB1xp67_ASAP7_75t_L g1472 ( 
.A(n_1395),
.Y(n_1472)
);

AND2x2_ASAP7_75t_L g1473 ( 
.A(n_1419),
.B(n_1430),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1405),
.B(n_1456),
.Y(n_1474)
);

AOI21x1_ASAP7_75t_L g1475 ( 
.A1(n_1452),
.A2(n_1428),
.B(n_1451),
.Y(n_1475)
);

OR2x6_ASAP7_75t_L g1476 ( 
.A(n_1440),
.B(n_1401),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_L g1477 ( 
.A(n_1455),
.B(n_1459),
.Y(n_1477)
);

AND2x2_ASAP7_75t_L g1478 ( 
.A(n_1453),
.B(n_1438),
.Y(n_1478)
);

OR2x6_ASAP7_75t_L g1479 ( 
.A(n_1440),
.B(n_1401),
.Y(n_1479)
);

AND2x2_ASAP7_75t_L g1480 ( 
.A(n_1453),
.B(n_1438),
.Y(n_1480)
);

AND2x4_ASAP7_75t_L g1481 ( 
.A(n_1411),
.B(n_1443),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1400),
.Y(n_1482)
);

AOI22xp33_ASAP7_75t_L g1483 ( 
.A1(n_1393),
.A2(n_1458),
.B1(n_1457),
.B2(n_1426),
.Y(n_1483)
);

AND2x2_ASAP7_75t_L g1484 ( 
.A(n_1436),
.B(n_1411),
.Y(n_1484)
);

AOI21xp5_ASAP7_75t_L g1485 ( 
.A1(n_1398),
.A2(n_1394),
.B(n_1402),
.Y(n_1485)
);

AND2x4_ASAP7_75t_L g1486 ( 
.A(n_1446),
.B(n_1447),
.Y(n_1486)
);

HB1xp67_ASAP7_75t_L g1487 ( 
.A(n_1403),
.Y(n_1487)
);

AND2x4_ASAP7_75t_L g1488 ( 
.A(n_1446),
.B(n_1447),
.Y(n_1488)
);

AOI22xp33_ASAP7_75t_L g1489 ( 
.A1(n_1439),
.A2(n_1427),
.B1(n_1424),
.B2(n_1431),
.Y(n_1489)
);

AND2x2_ASAP7_75t_L g1490 ( 
.A(n_1399),
.B(n_1407),
.Y(n_1490)
);

AND2x2_ASAP7_75t_L g1491 ( 
.A(n_1404),
.B(n_1449),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1425),
.Y(n_1492)
);

AO21x2_ASAP7_75t_L g1493 ( 
.A1(n_1462),
.A2(n_1461),
.B(n_1398),
.Y(n_1493)
);

INVx3_ASAP7_75t_L g1494 ( 
.A(n_1421),
.Y(n_1494)
);

AND2x2_ASAP7_75t_L g1495 ( 
.A(n_1464),
.B(n_1397),
.Y(n_1495)
);

HB1xp67_ASAP7_75t_L g1496 ( 
.A(n_1454),
.Y(n_1496)
);

OR2x2_ASAP7_75t_L g1497 ( 
.A(n_1391),
.B(n_1413),
.Y(n_1497)
);

OR2x6_ASAP7_75t_L g1498 ( 
.A(n_1420),
.B(n_1441),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1409),
.Y(n_1499)
);

NOR2xp33_ASAP7_75t_L g1500 ( 
.A(n_1410),
.B(n_1396),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1406),
.Y(n_1501)
);

OAI21x1_ASAP7_75t_L g1502 ( 
.A1(n_1416),
.A2(n_1429),
.B(n_1422),
.Y(n_1502)
);

INVxp67_ASAP7_75t_L g1503 ( 
.A(n_1490),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1482),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1492),
.Y(n_1505)
);

OR2x2_ASAP7_75t_L g1506 ( 
.A(n_1469),
.B(n_1429),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1490),
.B(n_1412),
.Y(n_1507)
);

OR2x2_ASAP7_75t_L g1508 ( 
.A(n_1469),
.B(n_1460),
.Y(n_1508)
);

AND2x2_ASAP7_75t_L g1509 ( 
.A(n_1478),
.B(n_1412),
.Y(n_1509)
);

AND2x2_ASAP7_75t_L g1510 ( 
.A(n_1480),
.B(n_1417),
.Y(n_1510)
);

OR2x2_ASAP7_75t_L g1511 ( 
.A(n_1467),
.B(n_1417),
.Y(n_1511)
);

BUFx2_ASAP7_75t_L g1512 ( 
.A(n_1465),
.Y(n_1512)
);

AND2x2_ASAP7_75t_L g1513 ( 
.A(n_1480),
.B(n_1417),
.Y(n_1513)
);

AND2x2_ASAP7_75t_L g1514 ( 
.A(n_1473),
.B(n_1448),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1491),
.B(n_1414),
.Y(n_1515)
);

HB1xp67_ASAP7_75t_L g1516 ( 
.A(n_1472),
.Y(n_1516)
);

HB1xp67_ASAP7_75t_L g1517 ( 
.A(n_1472),
.Y(n_1517)
);

NAND2xp5_ASAP7_75t_L g1518 ( 
.A(n_1491),
.B(n_1423),
.Y(n_1518)
);

AO21x2_ASAP7_75t_L g1519 ( 
.A1(n_1502),
.A2(n_1461),
.B(n_1420),
.Y(n_1519)
);

INVxp67_ASAP7_75t_L g1520 ( 
.A(n_1471),
.Y(n_1520)
);

INVxp67_ASAP7_75t_SL g1521 ( 
.A(n_1494),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1473),
.B(n_1448),
.Y(n_1522)
);

OAI22xp5_ASAP7_75t_L g1523 ( 
.A1(n_1483),
.A2(n_1396),
.B1(n_1442),
.B2(n_1435),
.Y(n_1523)
);

NOR2x1_ASAP7_75t_SL g1524 ( 
.A(n_1476),
.B(n_1434),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_L g1525 ( 
.A(n_1499),
.B(n_1497),
.Y(n_1525)
);

BUFx2_ASAP7_75t_L g1526 ( 
.A(n_1481),
.Y(n_1526)
);

OAI22xp5_ASAP7_75t_SL g1527 ( 
.A1(n_1476),
.A2(n_1445),
.B1(n_1432),
.B2(n_1433),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1504),
.Y(n_1528)
);

AOI22xp5_ASAP7_75t_L g1529 ( 
.A1(n_1523),
.A2(n_1485),
.B1(n_1477),
.B2(n_1488),
.Y(n_1529)
);

HB1xp67_ASAP7_75t_L g1530 ( 
.A(n_1516),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1504),
.Y(n_1531)
);

INVx4_ASAP7_75t_L g1532 ( 
.A(n_1519),
.Y(n_1532)
);

AO21x2_ASAP7_75t_L g1533 ( 
.A1(n_1520),
.A2(n_1519),
.B(n_1502),
.Y(n_1533)
);

AOI221xp5_ASAP7_75t_L g1534 ( 
.A1(n_1523),
.A2(n_1485),
.B1(n_1477),
.B2(n_1486),
.C(n_1488),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_L g1535 ( 
.A(n_1511),
.B(n_1471),
.Y(n_1535)
);

AOI22xp33_ASAP7_75t_L g1536 ( 
.A1(n_1519),
.A2(n_1486),
.B1(n_1476),
.B2(n_1479),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1505),
.Y(n_1537)
);

OAI33xp33_ASAP7_75t_L g1538 ( 
.A1(n_1515),
.A2(n_1474),
.A3(n_1499),
.B1(n_1497),
.B2(n_1466),
.B3(n_1501),
.Y(n_1538)
);

NOR2x1_ASAP7_75t_L g1539 ( 
.A(n_1511),
.B(n_1479),
.Y(n_1539)
);

AO21x2_ASAP7_75t_L g1540 ( 
.A1(n_1519),
.A2(n_1471),
.B(n_1475),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1505),
.Y(n_1541)
);

AND2x2_ASAP7_75t_L g1542 ( 
.A(n_1526),
.B(n_1470),
.Y(n_1542)
);

NAND4xp25_ASAP7_75t_SL g1543 ( 
.A(n_1515),
.B(n_1437),
.C(n_1489),
.D(n_1495),
.Y(n_1543)
);

AND2x4_ASAP7_75t_L g1544 ( 
.A(n_1524),
.B(n_1481),
.Y(n_1544)
);

AOI22xp33_ASAP7_75t_L g1545 ( 
.A1(n_1508),
.A2(n_1479),
.B1(n_1474),
.B2(n_1493),
.Y(n_1545)
);

AND2x6_ASAP7_75t_SL g1546 ( 
.A(n_1518),
.B(n_1500),
.Y(n_1546)
);

OAI31xp33_ASAP7_75t_L g1547 ( 
.A1(n_1527),
.A2(n_1487),
.A3(n_1466),
.B(n_1495),
.Y(n_1547)
);

OAI22xp5_ASAP7_75t_L g1548 ( 
.A1(n_1508),
.A2(n_1498),
.B1(n_1468),
.B2(n_1501),
.Y(n_1548)
);

OR2x2_ASAP7_75t_L g1549 ( 
.A(n_1506),
.B(n_1496),
.Y(n_1549)
);

BUFx3_ASAP7_75t_L g1550 ( 
.A(n_1512),
.Y(n_1550)
);

AND2x2_ASAP7_75t_L g1551 ( 
.A(n_1526),
.B(n_1484),
.Y(n_1551)
);

HB1xp67_ASAP7_75t_L g1552 ( 
.A(n_1516),
.Y(n_1552)
);

INVxp67_ASAP7_75t_SL g1553 ( 
.A(n_1517),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1528),
.Y(n_1554)
);

INVx2_ASAP7_75t_L g1555 ( 
.A(n_1540),
.Y(n_1555)
);

INVx2_ASAP7_75t_L g1556 ( 
.A(n_1540),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1528),
.Y(n_1557)
);

INVx2_ASAP7_75t_L g1558 ( 
.A(n_1540),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1551),
.B(n_1503),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1531),
.Y(n_1560)
);

AND2x2_ASAP7_75t_L g1561 ( 
.A(n_1551),
.B(n_1503),
.Y(n_1561)
);

AND2x2_ASAP7_75t_L g1562 ( 
.A(n_1550),
.B(n_1514),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1550),
.B(n_1514),
.Y(n_1563)
);

INVxp67_ASAP7_75t_L g1564 ( 
.A(n_1530),
.Y(n_1564)
);

INVx5_ASAP7_75t_L g1565 ( 
.A(n_1532),
.Y(n_1565)
);

HB1xp67_ASAP7_75t_L g1566 ( 
.A(n_1552),
.Y(n_1566)
);

OA21x2_ASAP7_75t_L g1567 ( 
.A1(n_1535),
.A2(n_1521),
.B(n_1507),
.Y(n_1567)
);

BUFx2_ASAP7_75t_L g1568 ( 
.A(n_1544),
.Y(n_1568)
);

INVx4_ASAP7_75t_L g1569 ( 
.A(n_1546),
.Y(n_1569)
);

INVxp67_ASAP7_75t_L g1570 ( 
.A(n_1543),
.Y(n_1570)
);

INVx4_ASAP7_75t_SL g1571 ( 
.A(n_1544),
.Y(n_1571)
);

BUFx12f_ASAP7_75t_L g1572 ( 
.A(n_1546),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1537),
.Y(n_1573)
);

AND2x2_ASAP7_75t_L g1574 ( 
.A(n_1542),
.B(n_1522),
.Y(n_1574)
);

INVx2_ASAP7_75t_SL g1575 ( 
.A(n_1544),
.Y(n_1575)
);

HB1xp67_ASAP7_75t_L g1576 ( 
.A(n_1553),
.Y(n_1576)
);

INVx2_ASAP7_75t_L g1577 ( 
.A(n_1533),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1537),
.Y(n_1578)
);

AND2x2_ASAP7_75t_L g1579 ( 
.A(n_1542),
.B(n_1522),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1541),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_L g1581 ( 
.A(n_1569),
.B(n_1534),
.Y(n_1581)
);

INVx1_ASAP7_75t_SL g1582 ( 
.A(n_1572),
.Y(n_1582)
);

OAI21xp33_ASAP7_75t_L g1583 ( 
.A1(n_1570),
.A2(n_1529),
.B(n_1543),
.Y(n_1583)
);

OR2x2_ASAP7_75t_L g1584 ( 
.A(n_1564),
.B(n_1535),
.Y(n_1584)
);

OAI221xp5_ASAP7_75t_L g1585 ( 
.A1(n_1570),
.A2(n_1529),
.B1(n_1547),
.B2(n_1545),
.C(n_1532),
.Y(n_1585)
);

INVx2_ASAP7_75t_SL g1586 ( 
.A(n_1568),
.Y(n_1586)
);

OR2x2_ASAP7_75t_L g1587 ( 
.A(n_1564),
.B(n_1549),
.Y(n_1587)
);

AND2x2_ASAP7_75t_L g1588 ( 
.A(n_1571),
.B(n_1568),
.Y(n_1588)
);

INVx1_ASAP7_75t_SL g1589 ( 
.A(n_1572),
.Y(n_1589)
);

OR2x2_ASAP7_75t_L g1590 ( 
.A(n_1566),
.B(n_1576),
.Y(n_1590)
);

CKINVDCx16_ASAP7_75t_R g1591 ( 
.A(n_1572),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1554),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1554),
.Y(n_1593)
);

INVx2_ASAP7_75t_L g1594 ( 
.A(n_1567),
.Y(n_1594)
);

INVx1_ASAP7_75t_SL g1595 ( 
.A(n_1572),
.Y(n_1595)
);

CKINVDCx16_ASAP7_75t_R g1596 ( 
.A(n_1569),
.Y(n_1596)
);

NOR2xp67_ASAP7_75t_L g1597 ( 
.A(n_1575),
.B(n_1532),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_L g1598 ( 
.A(n_1569),
.B(n_1518),
.Y(n_1598)
);

AND2x4_ASAP7_75t_L g1599 ( 
.A(n_1571),
.B(n_1532),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1554),
.Y(n_1600)
);

BUFx2_ASAP7_75t_L g1601 ( 
.A(n_1569),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_L g1602 ( 
.A(n_1569),
.B(n_1510),
.Y(n_1602)
);

OR2x2_ASAP7_75t_L g1603 ( 
.A(n_1566),
.B(n_1549),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1576),
.B(n_1510),
.Y(n_1604)
);

AND2x2_ASAP7_75t_L g1605 ( 
.A(n_1568),
.B(n_1513),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_L g1606 ( 
.A(n_1559),
.B(n_1509),
.Y(n_1606)
);

AND2x2_ASAP7_75t_L g1607 ( 
.A(n_1559),
.B(n_1509),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1580),
.Y(n_1608)
);

INVx6_ASAP7_75t_L g1609 ( 
.A(n_1565),
.Y(n_1609)
);

AND2x2_ASAP7_75t_L g1610 ( 
.A(n_1561),
.B(n_1509),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1580),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1575),
.B(n_1512),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1562),
.B(n_1525),
.Y(n_1613)
);

NOR2xp67_ASAP7_75t_L g1614 ( 
.A(n_1565),
.B(n_1548),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_1588),
.B(n_1562),
.Y(n_1615)
);

HB1xp67_ASAP7_75t_L g1616 ( 
.A(n_1590),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1592),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1592),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_L g1619 ( 
.A(n_1583),
.B(n_1574),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_L g1620 ( 
.A(n_1583),
.B(n_1574),
.Y(n_1620)
);

INVx2_ASAP7_75t_L g1621 ( 
.A(n_1594),
.Y(n_1621)
);

AOI22xp5_ASAP7_75t_L g1622 ( 
.A1(n_1585),
.A2(n_1538),
.B1(n_1539),
.B2(n_1536),
.Y(n_1622)
);

HB1xp67_ASAP7_75t_L g1623 ( 
.A(n_1590),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1588),
.B(n_1562),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_L g1625 ( 
.A(n_1581),
.B(n_1574),
.Y(n_1625)
);

NAND2xp33_ASAP7_75t_L g1626 ( 
.A(n_1582),
.B(n_1565),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1593),
.Y(n_1627)
);

AND2x2_ASAP7_75t_L g1628 ( 
.A(n_1586),
.B(n_1563),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1593),
.Y(n_1629)
);

OR2x2_ASAP7_75t_L g1630 ( 
.A(n_1603),
.B(n_1557),
.Y(n_1630)
);

AND2x4_ASAP7_75t_SL g1631 ( 
.A(n_1599),
.B(n_1563),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_L g1632 ( 
.A(n_1598),
.B(n_1579),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1600),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1600),
.Y(n_1634)
);

INVxp33_ASAP7_75t_L g1635 ( 
.A(n_1601),
.Y(n_1635)
);

BUFx3_ASAP7_75t_L g1636 ( 
.A(n_1601),
.Y(n_1636)
);

INVx2_ASAP7_75t_L g1637 ( 
.A(n_1594),
.Y(n_1637)
);

O2A1O1Ixp5_ASAP7_75t_SL g1638 ( 
.A1(n_1608),
.A2(n_1580),
.B(n_1578),
.C(n_1573),
.Y(n_1638)
);

OR2x2_ASAP7_75t_L g1639 ( 
.A(n_1603),
.B(n_1587),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_SL g1640 ( 
.A(n_1596),
.B(n_1565),
.Y(n_1640)
);

INVx1_ASAP7_75t_SL g1641 ( 
.A(n_1591),
.Y(n_1641)
);

OAI21xp5_ASAP7_75t_L g1642 ( 
.A1(n_1594),
.A2(n_1547),
.B(n_1567),
.Y(n_1642)
);

NAND2x1p5_ASAP7_75t_L g1643 ( 
.A(n_1586),
.B(n_1539),
.Y(n_1643)
);

OR2x2_ASAP7_75t_L g1644 ( 
.A(n_1587),
.B(n_1584),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1608),
.Y(n_1645)
);

O2A1O1Ixp33_ASAP7_75t_L g1646 ( 
.A1(n_1582),
.A2(n_1555),
.B(n_1558),
.C(n_1556),
.Y(n_1646)
);

OR2x2_ASAP7_75t_L g1647 ( 
.A(n_1584),
.B(n_1557),
.Y(n_1647)
);

OR2x2_ASAP7_75t_L g1648 ( 
.A(n_1613),
.B(n_1560),
.Y(n_1648)
);

HB1xp67_ASAP7_75t_L g1649 ( 
.A(n_1602),
.Y(n_1649)
);

INVx2_ASAP7_75t_L g1650 ( 
.A(n_1605),
.Y(n_1650)
);

INVx2_ASAP7_75t_SL g1651 ( 
.A(n_1631),
.Y(n_1651)
);

OR2x2_ASAP7_75t_L g1652 ( 
.A(n_1639),
.B(n_1596),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_L g1653 ( 
.A(n_1616),
.B(n_1589),
.Y(n_1653)
);

INVx2_ASAP7_75t_L g1654 ( 
.A(n_1621),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1615),
.B(n_1589),
.Y(n_1655)
);

NOR2xp33_ASAP7_75t_L g1656 ( 
.A(n_1641),
.B(n_1591),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1617),
.Y(n_1657)
);

INVx2_ASAP7_75t_L g1658 ( 
.A(n_1621),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1618),
.Y(n_1659)
);

AND2x2_ASAP7_75t_L g1660 ( 
.A(n_1615),
.B(n_1595),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_L g1661 ( 
.A(n_1623),
.B(n_1607),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1627),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1629),
.Y(n_1663)
);

INVx2_ASAP7_75t_L g1664 ( 
.A(n_1637),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1633),
.Y(n_1665)
);

HB1xp67_ASAP7_75t_L g1666 ( 
.A(n_1636),
.Y(n_1666)
);

AND2x2_ASAP7_75t_L g1667 ( 
.A(n_1624),
.B(n_1612),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_L g1668 ( 
.A(n_1619),
.B(n_1607),
.Y(n_1668)
);

INVx1_ASAP7_75t_SL g1669 ( 
.A(n_1639),
.Y(n_1669)
);

INVx1_ASAP7_75t_SL g1670 ( 
.A(n_1636),
.Y(n_1670)
);

NAND2xp5_ASAP7_75t_L g1671 ( 
.A(n_1620),
.B(n_1610),
.Y(n_1671)
);

INVxp67_ASAP7_75t_L g1672 ( 
.A(n_1644),
.Y(n_1672)
);

OR2x2_ASAP7_75t_L g1673 ( 
.A(n_1644),
.B(n_1611),
.Y(n_1673)
);

INVx1_ASAP7_75t_SL g1674 ( 
.A(n_1635),
.Y(n_1674)
);

INVx1_ASAP7_75t_SL g1675 ( 
.A(n_1628),
.Y(n_1675)
);

HB1xp67_ASAP7_75t_L g1676 ( 
.A(n_1649),
.Y(n_1676)
);

INVxp67_ASAP7_75t_SL g1677 ( 
.A(n_1656),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1673),
.Y(n_1678)
);

INVxp67_ASAP7_75t_L g1679 ( 
.A(n_1655),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1673),
.Y(n_1680)
);

OAI21xp5_ASAP7_75t_SL g1681 ( 
.A1(n_1669),
.A2(n_1642),
.B(n_1631),
.Y(n_1681)
);

NAND2xp5_ASAP7_75t_L g1682 ( 
.A(n_1672),
.B(n_1638),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1657),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1657),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_L g1685 ( 
.A(n_1676),
.B(n_1674),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1659),
.Y(n_1686)
);

AOI22xp5_ASAP7_75t_L g1687 ( 
.A1(n_1654),
.A2(n_1622),
.B1(n_1625),
.B2(n_1637),
.Y(n_1687)
);

OAI211xp5_ASAP7_75t_SL g1688 ( 
.A1(n_1652),
.A2(n_1626),
.B(n_1640),
.C(n_1650),
.Y(n_1688)
);

AND2x4_ASAP7_75t_L g1689 ( 
.A(n_1660),
.B(n_1628),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1670),
.B(n_1635),
.Y(n_1690)
);

NOR2xp33_ASAP7_75t_L g1691 ( 
.A(n_1652),
.B(n_1640),
.Y(n_1691)
);

INVx2_ASAP7_75t_SL g1692 ( 
.A(n_1655),
.Y(n_1692)
);

HB1xp67_ASAP7_75t_L g1693 ( 
.A(n_1660),
.Y(n_1693)
);

NAND3xp33_ASAP7_75t_L g1694 ( 
.A(n_1666),
.B(n_1638),
.C(n_1626),
.Y(n_1694)
);

AND2x2_ASAP7_75t_L g1695 ( 
.A(n_1667),
.B(n_1675),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1659),
.Y(n_1696)
);

INVx2_ASAP7_75t_L g1697 ( 
.A(n_1689),
.Y(n_1697)
);

OR2x2_ASAP7_75t_L g1698 ( 
.A(n_1693),
.B(n_1674),
.Y(n_1698)
);

INVx2_ASAP7_75t_L g1699 ( 
.A(n_1689),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_SL g1700 ( 
.A(n_1694),
.B(n_1692),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1685),
.Y(n_1701)
);

AND2x2_ASAP7_75t_L g1702 ( 
.A(n_1695),
.B(n_1651),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_L g1703 ( 
.A(n_1679),
.B(n_1670),
.Y(n_1703)
);

AND2x2_ASAP7_75t_L g1704 ( 
.A(n_1677),
.B(n_1651),
.Y(n_1704)
);

INVx1_ASAP7_75t_SL g1705 ( 
.A(n_1685),
.Y(n_1705)
);

NAND2xp5_ASAP7_75t_SL g1706 ( 
.A(n_1682),
.B(n_1690),
.Y(n_1706)
);

AOI222xp33_ASAP7_75t_L g1707 ( 
.A1(n_1682),
.A2(n_1664),
.B1(n_1654),
.B2(n_1658),
.C1(n_1577),
.C2(n_1653),
.Y(n_1707)
);

INVx2_ASAP7_75t_SL g1708 ( 
.A(n_1678),
.Y(n_1708)
);

INVx2_ASAP7_75t_L g1709 ( 
.A(n_1680),
.Y(n_1709)
);

NAND4xp25_ASAP7_75t_L g1710 ( 
.A(n_1702),
.B(n_1681),
.C(n_1691),
.D(n_1688),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1698),
.Y(n_1711)
);

AOI21xp5_ASAP7_75t_L g1712 ( 
.A1(n_1700),
.A2(n_1706),
.B(n_1705),
.Y(n_1712)
);

AOI211xp5_ASAP7_75t_L g1713 ( 
.A1(n_1700),
.A2(n_1687),
.B(n_1696),
.C(n_1686),
.Y(n_1713)
);

OAI211xp5_ASAP7_75t_SL g1714 ( 
.A1(n_1706),
.A2(n_1684),
.B(n_1683),
.C(n_1661),
.Y(n_1714)
);

NAND4xp75_ASAP7_75t_L g1715 ( 
.A(n_1704),
.B(n_1664),
.C(n_1654),
.D(n_1658),
.Y(n_1715)
);

OAI22xp5_ASAP7_75t_L g1716 ( 
.A1(n_1699),
.A2(n_1650),
.B1(n_1668),
.B2(n_1671),
.Y(n_1716)
);

NAND2xp5_ASAP7_75t_L g1717 ( 
.A(n_1699),
.B(n_1667),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_SL g1718 ( 
.A(n_1697),
.B(n_1643),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1703),
.Y(n_1719)
);

NAND3xp33_ASAP7_75t_L g1720 ( 
.A(n_1707),
.B(n_1664),
.C(n_1658),
.Y(n_1720)
);

AOI22xp5_ASAP7_75t_SL g1721 ( 
.A1(n_1712),
.A2(n_1701),
.B1(n_1703),
.B2(n_1708),
.Y(n_1721)
);

OAI21xp33_ASAP7_75t_L g1722 ( 
.A1(n_1710),
.A2(n_1709),
.B(n_1663),
.Y(n_1722)
);

OAI21xp5_ASAP7_75t_L g1723 ( 
.A1(n_1713),
.A2(n_1643),
.B(n_1597),
.Y(n_1723)
);

AOI22xp5_ASAP7_75t_L g1724 ( 
.A1(n_1720),
.A2(n_1614),
.B1(n_1663),
.B2(n_1662),
.Y(n_1724)
);

AOI21xp5_ASAP7_75t_L g1725 ( 
.A1(n_1714),
.A2(n_1665),
.B(n_1662),
.Y(n_1725)
);

A2O1A1Ixp33_ASAP7_75t_L g1726 ( 
.A1(n_1719),
.A2(n_1646),
.B(n_1665),
.C(n_1614),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1721),
.Y(n_1727)
);

NOR2xp33_ASAP7_75t_L g1728 ( 
.A(n_1722),
.B(n_1715),
.Y(n_1728)
);

NAND3xp33_ASAP7_75t_L g1729 ( 
.A(n_1725),
.B(n_1711),
.C(n_1717),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1724),
.Y(n_1730)
);

AND2x2_ASAP7_75t_L g1731 ( 
.A(n_1723),
.B(n_1716),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1726),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1721),
.Y(n_1733)
);

OR2x2_ASAP7_75t_L g1734 ( 
.A(n_1727),
.B(n_1630),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1733),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1729),
.Y(n_1736)
);

NOR2x1p5_ASAP7_75t_L g1737 ( 
.A(n_1732),
.B(n_1630),
.Y(n_1737)
);

NAND2xp33_ASAP7_75t_SL g1738 ( 
.A(n_1731),
.B(n_1718),
.Y(n_1738)
);

NOR2x1_ASAP7_75t_L g1739 ( 
.A(n_1736),
.B(n_1728),
.Y(n_1739)
);

AND2x2_ASAP7_75t_L g1740 ( 
.A(n_1737),
.B(n_1728),
.Y(n_1740)
);

NOR2x1_ASAP7_75t_L g1741 ( 
.A(n_1735),
.B(n_1730),
.Y(n_1741)
);

HB1xp67_ASAP7_75t_L g1742 ( 
.A(n_1741),
.Y(n_1742)
);

NOR3xp33_ASAP7_75t_L g1743 ( 
.A(n_1742),
.B(n_1739),
.C(n_1740),
.Y(n_1743)
);

BUFx2_ASAP7_75t_L g1744 ( 
.A(n_1743),
.Y(n_1744)
);

INVx2_ASAP7_75t_SL g1745 ( 
.A(n_1743),
.Y(n_1745)
);

OAI22x1_ASAP7_75t_L g1746 ( 
.A1(n_1744),
.A2(n_1734),
.B1(n_1738),
.B2(n_1645),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1745),
.Y(n_1747)
);

OAI21xp5_ASAP7_75t_L g1748 ( 
.A1(n_1747),
.A2(n_1647),
.B(n_1624),
.Y(n_1748)
);

OAI22xp5_ASAP7_75t_SL g1749 ( 
.A1(n_1746),
.A2(n_1609),
.B1(n_1599),
.B2(n_1632),
.Y(n_1749)
);

NAND2xp33_ASAP7_75t_SL g1750 ( 
.A(n_1749),
.B(n_1647),
.Y(n_1750)
);

HB1xp67_ASAP7_75t_L g1751 ( 
.A(n_1750),
.Y(n_1751)
);

OAI21xp5_ASAP7_75t_L g1752 ( 
.A1(n_1751),
.A2(n_1748),
.B(n_1634),
.Y(n_1752)
);

AO221x2_ASAP7_75t_L g1753 ( 
.A1(n_1752),
.A2(n_1609),
.B1(n_1611),
.B2(n_1604),
.C(n_1606),
.Y(n_1753)
);

AOI22xp33_ASAP7_75t_SL g1754 ( 
.A1(n_1753),
.A2(n_1609),
.B1(n_1599),
.B2(n_1565),
.Y(n_1754)
);

AOI211xp5_ASAP7_75t_L g1755 ( 
.A1(n_1754),
.A2(n_1597),
.B(n_1599),
.C(n_1648),
.Y(n_1755)
);


endmodule