module fake_jpeg_12443_n_90 (n_13, n_21, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_90);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_90;

wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_24;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

INVx2_ASAP7_75t_R g22 ( 
.A(n_0),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_18),
.Y(n_24)
);

CKINVDCx16_ASAP7_75t_R g25 ( 
.A(n_19),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx2_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

INVx6_ASAP7_75t_SL g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_20),
.Y(n_31)
);

OR2x2_ASAP7_75t_L g32 ( 
.A(n_14),
.B(n_8),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_30),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_37),
.Y(n_43)
);

INVx1_ASAP7_75t_SL g34 ( 
.A(n_31),
.Y(n_34)
);

INVx13_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_36),
.B(n_25),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_38),
.B(n_31),
.Y(n_45)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_38),
.B(n_26),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_41),
.B(n_42),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_35),
.A2(n_23),
.B1(n_28),
.B2(n_32),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_34),
.A2(n_23),
.B1(n_28),
.B2(n_32),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_44),
.B(n_45),
.Y(n_54)
);

INVx4_ASAP7_75t_SL g47 ( 
.A(n_39),
.Y(n_47)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_47),
.Y(n_55)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_46),
.Y(n_48)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_48),
.Y(n_57)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_46),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_49),
.B(n_50),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_22),
.Y(n_50)
);

INVx2_ASAP7_75t_SL g52 ( 
.A(n_39),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_52),
.B(n_47),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_56),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_48),
.A2(n_49),
.B1(n_52),
.B2(n_36),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_58),
.B(n_59),
.Y(n_66)
);

NOR3xp33_ASAP7_75t_SL g59 ( 
.A(n_51),
.B(n_27),
.C(n_22),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_53),
.B(n_43),
.C(n_24),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_60),
.B(n_2),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_54),
.B(n_33),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_61),
.B(n_62),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_53),
.B(n_1),
.Y(n_62)
);

BUFx24_ASAP7_75t_SL g64 ( 
.A(n_63),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_64),
.Y(n_73)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_55),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_67),
.B(n_68),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_57),
.A2(n_37),
.B1(n_36),
.B2(n_3),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_59),
.B(n_1),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_69),
.B(n_70),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_58),
.B(n_2),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_L g75 ( 
.A1(n_72),
.A2(n_66),
.B(n_65),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_75),
.Y(n_82)
);

AOI322xp5_ASAP7_75t_L g77 ( 
.A1(n_65),
.A2(n_4),
.A3(n_5),
.B1(n_6),
.B2(n_21),
.C1(n_10),
.C2(n_12),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_77),
.B(n_79),
.C(n_16),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_71),
.Y(n_78)
);

CKINVDCx14_ASAP7_75t_R g81 ( 
.A(n_78),
.Y(n_81)
);

BUFx10_ASAP7_75t_L g79 ( 
.A(n_65),
.Y(n_79)
);

XOR2xp5_ASAP7_75t_L g83 ( 
.A(n_80),
.B(n_74),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_83),
.B(n_82),
.C(n_79),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_84),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_85),
.B(n_73),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_86),
.A2(n_81),
.B1(n_76),
.B2(n_77),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g88 ( 
.A1(n_87),
.A2(n_6),
.B(n_9),
.Y(n_88)
);

OAI21x1_ASAP7_75t_L g89 ( 
.A1(n_88),
.A2(n_13),
.B(n_15),
.Y(n_89)
);

XOR2xp5_ASAP7_75t_L g90 ( 
.A(n_89),
.B(n_17),
.Y(n_90)
);


endmodule