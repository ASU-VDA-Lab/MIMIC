module fake_netlist_6_2802_n_2714 (n_52, n_591, n_435, n_1, n_91, n_326, n_256, n_440, n_587, n_507, n_580, n_209, n_367, n_465, n_590, n_625, n_63, n_223, n_278, n_341, n_362, n_148, n_226, n_161, n_22, n_208, n_462, n_68, n_607, n_316, n_419, n_28, n_304, n_212, n_50, n_7, n_578, n_144, n_365, n_125, n_168, n_384, n_297, n_595, n_627, n_524, n_342, n_77, n_106, n_358, n_160, n_449, n_131, n_188, n_310, n_509, n_186, n_245, n_0, n_368, n_575, n_396, n_495, n_350, n_78, n_84, n_585, n_568, n_392, n_442, n_480, n_142, n_143, n_382, n_180, n_62, n_628, n_557, n_349, n_233, n_617, n_255, n_284, n_400, n_140, n_337, n_214, n_485, n_67, n_15, n_443, n_246, n_38, n_471, n_289, n_421, n_424, n_615, n_59, n_181, n_182, n_238, n_573, n_202, n_320, n_108, n_327, n_369, n_597, n_280, n_287, n_353, n_610, n_555, n_389, n_415, n_65, n_230, n_605, n_461, n_141, n_383, n_200, n_447, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_517, n_71, n_74, n_229, n_542, n_621, n_305, n_72, n_532, n_173, n_535, n_250, n_372, n_468, n_544, n_111, n_504, n_314, n_378, n_413, n_377, n_35, n_183, n_510, n_79, n_375, n_601, n_338, n_522, n_466, n_506, n_56, n_360, n_603, n_119, n_235, n_536, n_622, n_147, n_191, n_340, n_387, n_452, n_616, n_39, n_344, n_73, n_581, n_428, n_609, n_432, n_101, n_167, n_631, n_174, n_127, n_516, n_153, n_525, n_611, n_156, n_491, n_145, n_42, n_133, n_96, n_8, n_371, n_567, n_189, n_405, n_213, n_538, n_294, n_302, n_499, n_380, n_129, n_197, n_11, n_137, n_17, n_343, n_448, n_20, n_494, n_539, n_493, n_397, n_155, n_109, n_614, n_529, n_445, n_425, n_122, n_45, n_454, n_34, n_218, n_70, n_234, n_37, n_486, n_381, n_82, n_27, n_236, n_112, n_172, n_576, n_472, n_270, n_239, n_126, n_414, n_97, n_563, n_58, n_490, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_402, n_352, n_478, n_626, n_574, n_9, n_460, n_107, n_6, n_417, n_14, n_446, n_498, n_89, n_374, n_366, n_407, n_450, n_103, n_272, n_526, n_185, n_348, n_579, n_69, n_376, n_390, n_473, n_293, n_31, n_334, n_559, n_53, n_370, n_44, n_458, n_232, n_16, n_163, n_46, n_330, n_470, n_475, n_298, n_18, n_492, n_281, n_258, n_551, n_154, n_456, n_564, n_98, n_260, n_265, n_313, n_451, n_624, n_279, n_252, n_228, n_565, n_594, n_356, n_577, n_166, n_184, n_552, n_619, n_216, n_455, n_83, n_521, n_363, n_572, n_395, n_592, n_323, n_606, n_393, n_411, n_503, n_152, n_623, n_92, n_599, n_513, n_321, n_331, n_105, n_227, n_132, n_570, n_406, n_483, n_102, n_204, n_482, n_474, n_527, n_261, n_608, n_620, n_420, n_630, n_312, n_394, n_32, n_66, n_130, n_519, n_541, n_512, n_164, n_292, n_100, n_121, n_307, n_469, n_433, n_500, n_23, n_476, n_2, n_291, n_219, n_543, n_357, n_150, n_264, n_263, n_589, n_481, n_325, n_329, n_464, n_600, n_561, n_33, n_477, n_549, n_533, n_408, n_61, n_237, n_584, n_244, n_399, n_76, n_243, n_124, n_548, n_94, n_282, n_436, n_116, n_211, n_523, n_117, n_175, n_322, n_345, n_409, n_231, n_354, n_40, n_505, n_240, n_139, n_319, n_41, n_134, n_547, n_537, n_273, n_558, n_95, n_311, n_10, n_403, n_253, n_583, n_596, n_123, n_136, n_546, n_562, n_249, n_201, n_386, n_556, n_159, n_157, n_162, n_115, n_487, n_550, n_128, n_241, n_30, n_275, n_553, n_43, n_560, n_276, n_569, n_441, n_221, n_444, n_586, n_423, n_146, n_318, n_303, n_511, n_467, n_306, n_21, n_193, n_269, n_359, n_346, n_88, n_3, n_416, n_530, n_277, n_520, n_418, n_113, n_618, n_582, n_4, n_199, n_138, n_266, n_296, n_571, n_268, n_271, n_404, n_439, n_158, n_217, n_49, n_210, n_299, n_518, n_206, n_5, n_453, n_612, n_633, n_333, n_588, n_215, n_178, n_247, n_225, n_308, n_309, n_355, n_426, n_317, n_149, n_632, n_431, n_90, n_347, n_24, n_459, n_54, n_502, n_328, n_534, n_488, n_429, n_373, n_87, n_195, n_285, n_497, n_85, n_99, n_257, n_13, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_29, n_75, n_401, n_324, n_335, n_430, n_463, n_545, n_489, n_205, n_604, n_120, n_251, n_301, n_274, n_110, n_151, n_412, n_81, n_36, n_26, n_55, n_267, n_438, n_339, n_315, n_434, n_515, n_64, n_288, n_427, n_479, n_496, n_598, n_422, n_135, n_165, n_351, n_437, n_259, n_177, n_540, n_593, n_514, n_528, n_391, n_457, n_364, n_295, n_385, n_629, n_388, n_190, n_262, n_484, n_613, n_187, n_501, n_531, n_60, n_361, n_508, n_379, n_170, n_332, n_336, n_12, n_398, n_410, n_566, n_554, n_602, n_194, n_171, n_192, n_57, n_169, n_51, n_283, n_2714);

input n_52;
input n_591;
input n_435;
input n_1;
input n_91;
input n_326;
input n_256;
input n_440;
input n_587;
input n_507;
input n_580;
input n_209;
input n_367;
input n_465;
input n_590;
input n_625;
input n_63;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_462;
input n_68;
input n_607;
input n_316;
input n_419;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_578;
input n_144;
input n_365;
input n_125;
input n_168;
input n_384;
input n_297;
input n_595;
input n_627;
input n_524;
input n_342;
input n_77;
input n_106;
input n_358;
input n_160;
input n_449;
input n_131;
input n_188;
input n_310;
input n_509;
input n_186;
input n_245;
input n_0;
input n_368;
input n_575;
input n_396;
input n_495;
input n_350;
input n_78;
input n_84;
input n_585;
input n_568;
input n_392;
input n_442;
input n_480;
input n_142;
input n_143;
input n_382;
input n_180;
input n_62;
input n_628;
input n_557;
input n_349;
input n_233;
input n_617;
input n_255;
input n_284;
input n_400;
input n_140;
input n_337;
input n_214;
input n_485;
input n_67;
input n_15;
input n_443;
input n_246;
input n_38;
input n_471;
input n_289;
input n_421;
input n_424;
input n_615;
input n_59;
input n_181;
input n_182;
input n_238;
input n_573;
input n_202;
input n_320;
input n_108;
input n_327;
input n_369;
input n_597;
input n_280;
input n_287;
input n_353;
input n_610;
input n_555;
input n_389;
input n_415;
input n_65;
input n_230;
input n_605;
input n_461;
input n_141;
input n_383;
input n_200;
input n_447;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_517;
input n_71;
input n_74;
input n_229;
input n_542;
input n_621;
input n_305;
input n_72;
input n_532;
input n_173;
input n_535;
input n_250;
input n_372;
input n_468;
input n_544;
input n_111;
input n_504;
input n_314;
input n_378;
input n_413;
input n_377;
input n_35;
input n_183;
input n_510;
input n_79;
input n_375;
input n_601;
input n_338;
input n_522;
input n_466;
input n_506;
input n_56;
input n_360;
input n_603;
input n_119;
input n_235;
input n_536;
input n_622;
input n_147;
input n_191;
input n_340;
input n_387;
input n_452;
input n_616;
input n_39;
input n_344;
input n_73;
input n_581;
input n_428;
input n_609;
input n_432;
input n_101;
input n_167;
input n_631;
input n_174;
input n_127;
input n_516;
input n_153;
input n_525;
input n_611;
input n_156;
input n_491;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_371;
input n_567;
input n_189;
input n_405;
input n_213;
input n_538;
input n_294;
input n_302;
input n_499;
input n_380;
input n_129;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_448;
input n_20;
input n_494;
input n_539;
input n_493;
input n_397;
input n_155;
input n_109;
input n_614;
input n_529;
input n_445;
input n_425;
input n_122;
input n_45;
input n_454;
input n_34;
input n_218;
input n_70;
input n_234;
input n_37;
input n_486;
input n_381;
input n_82;
input n_27;
input n_236;
input n_112;
input n_172;
input n_576;
input n_472;
input n_270;
input n_239;
input n_126;
input n_414;
input n_97;
input n_563;
input n_58;
input n_490;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_402;
input n_352;
input n_478;
input n_626;
input n_574;
input n_9;
input n_460;
input n_107;
input n_6;
input n_417;
input n_14;
input n_446;
input n_498;
input n_89;
input n_374;
input n_366;
input n_407;
input n_450;
input n_103;
input n_272;
input n_526;
input n_185;
input n_348;
input n_579;
input n_69;
input n_376;
input n_390;
input n_473;
input n_293;
input n_31;
input n_334;
input n_559;
input n_53;
input n_370;
input n_44;
input n_458;
input n_232;
input n_16;
input n_163;
input n_46;
input n_330;
input n_470;
input n_475;
input n_298;
input n_18;
input n_492;
input n_281;
input n_258;
input n_551;
input n_154;
input n_456;
input n_564;
input n_98;
input n_260;
input n_265;
input n_313;
input n_451;
input n_624;
input n_279;
input n_252;
input n_228;
input n_565;
input n_594;
input n_356;
input n_577;
input n_166;
input n_184;
input n_552;
input n_619;
input n_216;
input n_455;
input n_83;
input n_521;
input n_363;
input n_572;
input n_395;
input n_592;
input n_323;
input n_606;
input n_393;
input n_411;
input n_503;
input n_152;
input n_623;
input n_92;
input n_599;
input n_513;
input n_321;
input n_331;
input n_105;
input n_227;
input n_132;
input n_570;
input n_406;
input n_483;
input n_102;
input n_204;
input n_482;
input n_474;
input n_527;
input n_261;
input n_608;
input n_620;
input n_420;
input n_630;
input n_312;
input n_394;
input n_32;
input n_66;
input n_130;
input n_519;
input n_541;
input n_512;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_469;
input n_433;
input n_500;
input n_23;
input n_476;
input n_2;
input n_291;
input n_219;
input n_543;
input n_357;
input n_150;
input n_264;
input n_263;
input n_589;
input n_481;
input n_325;
input n_329;
input n_464;
input n_600;
input n_561;
input n_33;
input n_477;
input n_549;
input n_533;
input n_408;
input n_61;
input n_237;
input n_584;
input n_244;
input n_399;
input n_76;
input n_243;
input n_124;
input n_548;
input n_94;
input n_282;
input n_436;
input n_116;
input n_211;
input n_523;
input n_117;
input n_175;
input n_322;
input n_345;
input n_409;
input n_231;
input n_354;
input n_40;
input n_505;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_547;
input n_537;
input n_273;
input n_558;
input n_95;
input n_311;
input n_10;
input n_403;
input n_253;
input n_583;
input n_596;
input n_123;
input n_136;
input n_546;
input n_562;
input n_249;
input n_201;
input n_386;
input n_556;
input n_159;
input n_157;
input n_162;
input n_115;
input n_487;
input n_550;
input n_128;
input n_241;
input n_30;
input n_275;
input n_553;
input n_43;
input n_560;
input n_276;
input n_569;
input n_441;
input n_221;
input n_444;
input n_586;
input n_423;
input n_146;
input n_318;
input n_303;
input n_511;
input n_467;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_346;
input n_88;
input n_3;
input n_416;
input n_530;
input n_277;
input n_520;
input n_418;
input n_113;
input n_618;
input n_582;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_571;
input n_268;
input n_271;
input n_404;
input n_439;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_518;
input n_206;
input n_5;
input n_453;
input n_612;
input n_633;
input n_333;
input n_588;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_355;
input n_426;
input n_317;
input n_149;
input n_632;
input n_431;
input n_90;
input n_347;
input n_24;
input n_459;
input n_54;
input n_502;
input n_328;
input n_534;
input n_488;
input n_429;
input n_373;
input n_87;
input n_195;
input n_285;
input n_497;
input n_85;
input n_99;
input n_257;
input n_13;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_29;
input n_75;
input n_401;
input n_324;
input n_335;
input n_430;
input n_463;
input n_545;
input n_489;
input n_205;
input n_604;
input n_120;
input n_251;
input n_301;
input n_274;
input n_110;
input n_151;
input n_412;
input n_81;
input n_36;
input n_26;
input n_55;
input n_267;
input n_438;
input n_339;
input n_315;
input n_434;
input n_515;
input n_64;
input n_288;
input n_427;
input n_479;
input n_496;
input n_598;
input n_422;
input n_135;
input n_165;
input n_351;
input n_437;
input n_259;
input n_177;
input n_540;
input n_593;
input n_514;
input n_528;
input n_391;
input n_457;
input n_364;
input n_295;
input n_385;
input n_629;
input n_388;
input n_190;
input n_262;
input n_484;
input n_613;
input n_187;
input n_501;
input n_531;
input n_60;
input n_361;
input n_508;
input n_379;
input n_170;
input n_332;
input n_336;
input n_12;
input n_398;
input n_410;
input n_566;
input n_554;
input n_602;
input n_194;
input n_171;
input n_192;
input n_57;
input n_169;
input n_51;
input n_283;

output n_2714;

wire n_992;
wire n_2542;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_2576;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_1189;
wire n_1212;
wire n_726;
wire n_2157;
wire n_2332;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_1581;
wire n_1003;
wire n_1237;
wire n_1061;
wire n_2353;
wire n_2534;
wire n_1357;
wire n_1853;
wire n_783;
wire n_2451;
wire n_1738;
wire n_2243;
wire n_798;
wire n_1575;
wire n_1854;
wire n_2324;
wire n_1923;
wire n_1342;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_2260;
wire n_1708;
wire n_677;
wire n_805;
wire n_1151;
wire n_1739;
wire n_2051;
wire n_2317;
wire n_1380;
wire n_2359;
wire n_1402;
wire n_2557;
wire n_1688;
wire n_1691;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_2405;
wire n_1160;
wire n_883;
wire n_2647;
wire n_1238;
wire n_1991;
wire n_2570;
wire n_2179;
wire n_2386;
wire n_1724;
wire n_1032;
wire n_2336;
wire n_1247;
wire n_1547;
wire n_2521;
wire n_1553;
wire n_893;
wire n_1099;
wire n_2491;
wire n_1264;
wire n_1192;
wire n_1844;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_2211;
wire n_1370;
wire n_1786;
wire n_2382;
wire n_2672;
wire n_2291;
wire n_830;
wire n_2299;
wire n_873;
wire n_1285;
wire n_1371;
wire n_1985;
wire n_2184;
wire n_1803;
wire n_1172;
wire n_852;
wire n_2509;
wire n_2513;
wire n_1590;
wire n_2645;
wire n_1532;
wire n_2313;
wire n_2628;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_1711;
wire n_2247;
wire n_1140;
wire n_2630;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_2344;
wire n_1579;
wire n_2365;
wire n_2470;
wire n_2321;
wire n_1263;
wire n_2019;
wire n_836;
wire n_2074;
wire n_2447;
wire n_2129;
wire n_2340;
wire n_1261;
wire n_945;
wire n_2286;
wire n_1649;
wire n_2094;
wire n_2018;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_2356;
wire n_2399;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_658;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_2510;
wire n_1541;
wire n_1300;
wire n_641;
wire n_2480;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_2212;
wire n_758;
wire n_1455;
wire n_2418;
wire n_1163;
wire n_1180;
wire n_2256;
wire n_2582;
wire n_943;
wire n_1798;
wire n_1550;
wire n_2703;
wire n_1591;
wire n_772;
wire n_1344;
wire n_2495;
wire n_666;
wire n_940;
wire n_770;
wire n_1781;
wire n_1971;
wire n_2058;
wire n_2090;
wire n_2603;
wire n_2660;
wire n_2173;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_2394;
wire n_2108;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_2378;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_2655;
wire n_1400;
wire n_2625;
wire n_1467;
wire n_976;
wire n_2155;
wire n_2686;
wire n_1445;
wire n_2364;
wire n_2551;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_2599;
wire n_1978;
wire n_2085;
wire n_917;
wire n_2370;
wire n_2612;
wire n_907;
wire n_1446;
wire n_2591;
wire n_659;
wire n_1815;
wire n_2214;
wire n_913;
wire n_1658;
wire n_2593;
wire n_808;
wire n_867;
wire n_1230;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_2613;
wire n_1333;
wire n_2496;
wire n_2708;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_2277;
wire n_1558;
wire n_1732;
wire n_2300;
wire n_699;
wire n_1986;
wire n_2397;
wire n_824;
wire n_686;
wire n_757;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_2190;
wire n_1843;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_813;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_2104;
wire n_645;
wire n_1381;
wire n_1699;
wire n_916;
wire n_2093;
wire n_2633;
wire n_2207;
wire n_1970;
wire n_2101;
wire n_2696;
wire n_2059;
wire n_2198;
wire n_2669;
wire n_2073;
wire n_2273;
wire n_2546;
wire n_792;
wire n_2522;
wire n_1328;
wire n_1957;
wire n_2616;
wire n_1907;
wire n_2529;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_982;
wire n_2674;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_932;
wire n_1876;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_993;
wire n_2692;
wire n_689;
wire n_2031;
wire n_2130;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_2228;
wire n_1988;
wire n_1278;
wire n_2455;
wire n_2654;
wire n_2469;
wire n_1064;
wire n_1396;
wire n_634;
wire n_2355;
wire n_966;
wire n_764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_2245;
wire n_2068;
wire n_1107;
wire n_2457;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_2580;
wire n_882;
wire n_2176;
wire n_2072;
wire n_1354;
wire n_1875;
wire n_1865;
wire n_1701;
wire n_2459;
wire n_1111;
wire n_1713;
wire n_715;
wire n_2678;
wire n_1251;
wire n_1265;
wire n_2711;
wire n_1726;
wire n_1950;
wire n_1563;
wire n_1912;
wire n_2434;
wire n_1982;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_2428;
wire n_674;
wire n_871;
wire n_922;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_2664;
wire n_1664;
wire n_1722;
wire n_2641;
wire n_1165;
wire n_702;
wire n_2008;
wire n_2192;
wire n_2254;
wire n_2345;
wire n_1926;
wire n_1175;
wire n_1386;
wire n_2311;
wire n_1896;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_2624;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_2350;
wire n_2453;
wire n_2193;
wire n_2676;
wire n_1655;
wire n_835;
wire n_928;
wire n_1214;
wire n_1801;
wire n_690;
wire n_850;
wire n_1886;
wire n_2092;
wire n_2347;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_2514;
wire n_2206;
wire n_2319;
wire n_2519;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_2467;
wire n_2602;
wire n_2468;
wire n_1124;
wire n_1624;
wire n_2096;
wire n_1965;
wire n_2476;
wire n_696;
wire n_1515;
wire n_961;
wire n_1082;
wire n_1317;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_2377;
wire n_701;
wire n_2178;
wire n_950;
wire n_2644;
wire n_2036;
wire n_2152;
wire n_1709;
wire n_2652;
wire n_2411;
wire n_2525;
wire n_1825;
wire n_2393;
wire n_1757;
wire n_1796;
wire n_2657;
wire n_1792;
wire n_891;
wire n_2067;
wire n_2136;
wire n_2409;
wire n_2082;
wire n_2252;
wire n_1412;
wire n_2497;
wire n_2687;
wire n_949;
wire n_1630;
wire n_678;
wire n_2075;
wire n_2194;
wire n_2619;
wire n_1987;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_2271;
wire n_1008;
wire n_760;
wire n_1546;
wire n_2583;
wire n_2606;
wire n_2279;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_2663;
wire n_1990;
wire n_2391;
wire n_2431;
wire n_694;
wire n_2150;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_2078;
wire n_1767;
wire n_1779;
wire n_1465;
wire n_2622;
wire n_1858;
wire n_1044;
wire n_2658;
wire n_2665;
wire n_2165;
wire n_2133;
wire n_1712;
wire n_1391;
wire n_1523;
wire n_2558;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_2349;
wire n_2684;
wire n_2712;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_815;
wire n_1100;
wire n_1487;
wire n_2691;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_2493;
wire n_673;
wire n_2230;
wire n_2705;
wire n_1969;
wire n_2690;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_2145;
wire n_1968;
wire n_898;
wire n_1952;
wire n_865;
wire n_2573;
wire n_2646;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_2535;
wire n_2631;
wire n_1364;
wire n_2436;
wire n_1249;
wire n_2706;
wire n_1293;
wire n_2693;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_1451;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_2341;
wire n_685;
wire n_1765;
wire n_2707;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_2537;
wire n_2554;
wire n_996;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_1513;
wire n_791;
wire n_1913;
wire n_837;
wire n_2097;
wire n_2170;
wire n_1488;
wire n_1808;
wire n_948;
wire n_2517;
wire n_2713;
wire n_704;
wire n_2148;
wire n_977;
wire n_2339;
wire n_1005;
wire n_1947;
wire n_1788;
wire n_1999;
wire n_2590;
wire n_2643;
wire n_1469;
wire n_2060;
wire n_2608;
wire n_1838;
wire n_2638;
wire n_1835;
wire n_1776;
wire n_1766;
wire n_1959;
wire n_2002;
wire n_2650;
wire n_2138;
wire n_765;
wire n_1492;
wire n_987;
wire n_2414;
wire n_1340;
wire n_1771;
wire n_2316;
wire n_720;
wire n_842;
wire n_2262;
wire n_1707;
wire n_2239;
wire n_1432;
wire n_2208;
wire n_843;
wire n_656;
wire n_989;
wire n_2604;
wire n_2407;
wire n_1277;
wire n_797;
wire n_2689;
wire n_1473;
wire n_2191;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_2574;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_2675;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_2134;
wire n_1529;
wire n_2335;
wire n_2473;
wire n_1022;
wire n_2069;
wire n_2307;
wire n_2362;
wire n_684;
wire n_2539;
wire n_2667;
wire n_2698;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_2297;
wire n_1181;
wire n_2119;
wire n_1822;
wire n_947;
wire n_1117;
wire n_2489;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_2445;
wire n_2057;
wire n_2103;
wire n_2605;
wire n_1666;
wire n_1505;
wire n_803;
wire n_1717;
wire n_926;
wire n_1817;
wire n_2449;
wire n_927;
wire n_2610;
wire n_1849;
wire n_919;
wire n_1698;
wire n_2231;
wire n_929;
wire n_2520;
wire n_1228;
wire n_1568;
wire n_1490;
wire n_2372;
wire n_777;
wire n_1299;
wire n_2639;
wire n_1183;
wire n_1436;
wire n_2251;
wire n_1384;
wire n_2494;
wire n_2501;
wire n_2238;
wire n_2368;
wire n_1070;
wire n_2403;
wire n_998;
wire n_717;
wire n_1665;
wire n_2524;
wire n_1383;
wire n_2460;
wire n_1178;
wire n_2127;
wire n_1424;
wire n_2338;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_2137;
wire n_1626;
wire n_1507;
wire n_2482;
wire n_2532;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_2481;
wire n_912;
wire n_1857;
wire n_1519;
wire n_2144;
wire n_745;
wire n_1284;
wire n_1604;
wire n_2296;
wire n_2424;
wire n_1142;
wire n_716;
wire n_1475;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_2354;
wire n_2682;
wire n_2589;
wire n_1395;
wire n_2110;
wire n_2199;
wire n_2661;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_811;
wire n_683;
wire n_1207;
wire n_2442;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_1250;
wire n_958;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_2053;
wire n_2259;
wire n_2121;
wire n_2545;
wire n_889;
wire n_2432;
wire n_2710;
wire n_1478;
wire n_1310;
wire n_819;
wire n_2294;
wire n_1363;
wire n_2581;
wire n_1334;
wire n_1966;
wire n_1942;
wire n_767;
wire n_1314;
wire n_964;
wire n_831;
wire n_1837;
wire n_2218;
wire n_2435;
wire n_954;
wire n_864;
wire n_2504;
wire n_2623;
wire n_1110;
wire n_2213;
wire n_1410;
wire n_2389;
wire n_1440;
wire n_2132;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_1483;
wire n_1834;
wire n_2331;
wire n_1372;
wire n_2292;
wire n_2330;
wire n_1457;
wire n_1719;
wire n_1339;
wire n_1787;
wire n_2701;
wire n_2475;
wire n_2511;
wire n_1993;
wire n_2281;
wire n_1427;
wire n_2416;
wire n_2617;
wire n_1466;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_1141;
wire n_1268;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_2323;
wire n_1893;
wire n_2209;
wire n_2301;
wire n_2387;
wire n_1755;
wire n_1602;
wire n_2421;
wire n_1136;
wire n_2618;
wire n_2025;
wire n_2357;
wire n_2464;
wire n_1125;
wire n_970;
wire n_2488;
wire n_2224;
wire n_1980;
wire n_642;
wire n_995;
wire n_1159;
wire n_2329;
wire n_1092;
wire n_2237;
wire n_1060;
wire n_1951;
wire n_2250;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_2115;
wire n_2410;
wire n_2552;
wire n_1053;
wire n_2374;
wire n_1681;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_2596;
wire n_2274;
wire n_775;
wire n_651;
wire n_1153;
wire n_1618;
wire n_1531;
wire n_1185;
wire n_2384;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_2585;
wire n_2621;
wire n_1653;
wire n_2352;
wire n_1679;
wire n_1625;
wire n_2601;
wire n_2160;
wire n_1453;
wire n_2146;
wire n_2226;
wire n_2131;
wire n_2502;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_2556;
wire n_2648;
wire n_1315;
wire n_1647;
wire n_2575;
wire n_1224;
wire n_2306;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_2462;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_1617;
wire n_1470;
wire n_2550;
wire n_1243;
wire n_848;
wire n_1096;
wire n_2249;
wire n_1091;
wire n_2000;
wire n_1917;
wire n_1580;
wire n_2227;
wire n_2270;
wire n_1425;
wire n_1881;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_2023;
wire n_2572;
wire n_2204;
wire n_1520;
wire n_2159;
wire n_906;
wire n_1390;
wire n_688;
wire n_2289;
wire n_1077;
wire n_1733;
wire n_2315;
wire n_1419;
wire n_1731;
wire n_2158;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_2135;
wire n_1645;
wire n_1832;
wire n_1687;
wire n_1439;
wire n_2328;
wire n_1323;
wire n_2202;
wire n_858;
wire n_2049;
wire n_1331;
wire n_736;
wire n_2627;
wire n_956;
wire n_960;
wire n_2276;
wire n_663;
wire n_856;
wire n_2100;
wire n_778;
wire n_1668;
wire n_1134;
wire n_1129;
wire n_1696;
wire n_2181;
wire n_1594;
wire n_1995;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_2379;
wire n_1905;
wire n_2016;
wire n_2343;
wire n_793;
wire n_1593;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_2515;
wire n_1744;
wire n_828;
wire n_2139;
wire n_2142;
wire n_1551;
wire n_2448;
wire n_1103;
wire n_2555;
wire n_2219;
wire n_1203;
wire n_820;
wire n_2327;
wire n_951;
wire n_2201;
wire n_725;
wire n_952;
wire n_999;
wire n_1254;
wire n_2420;
wire n_994;
wire n_2263;
wire n_2304;
wire n_1508;
wire n_2487;
wire n_732;
wire n_974;
wire n_2240;
wire n_2278;
wire n_2656;
wire n_2538;
wire n_724;
wire n_2597;
wire n_2375;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_1871;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_1549;
wire n_1510;
wire n_892;
wire n_768;
wire n_1468;
wire n_1859;
wire n_2102;
wire n_2563;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_2156;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_2598;
wire n_1270;
wire n_2549;
wire n_1187;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_2153;
wire n_2544;
wire n_2381;
wire n_1847;
wire n_2052;
wire n_2302;
wire n_1667;
wire n_667;
wire n_1206;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_923;
wire n_1409;
wire n_1841;
wire n_2637;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_2526;
wire n_2423;
wire n_1057;
wire n_2548;
wire n_991;
wire n_1657;
wire n_1126;
wire n_2412;
wire n_1997;
wire n_2636;
wire n_710;
wire n_1108;
wire n_1818;
wire n_2439;
wire n_2404;
wire n_1182;
wire n_1298;
wire n_2559;
wire n_2177;
wire n_2595;
wire n_2088;
wire n_1611;
wire n_785;
wire n_746;
wire n_1601;
wire n_1960;
wire n_2694;
wire n_2061;
wire n_1686;
wire n_2337;
wire n_2401;
wire n_1356;
wire n_1589;
wire n_2309;
wire n_2607;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_2452;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_2499;
wire n_1622;
wire n_1586;
wire n_2543;
wire n_2264;
wire n_1694;
wire n_1535;
wire n_2486;
wire n_2571;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_1983;
wire n_1938;
wire n_2498;
wire n_2220;
wire n_2577;
wire n_1262;
wire n_2472;
wire n_1891;
wire n_2171;
wire n_1213;
wire n_2235;
wire n_1350;
wire n_1673;
wire n_2232;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_2392;
wire n_2037;
wire n_2298;
wire n_782;
wire n_2326;
wire n_1539;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_2305;
wire n_2120;
wire n_1472;
wire n_2050;
wire n_2373;
wire n_2164;
wire n_2402;
wire n_2225;
wire n_1081;
wire n_1870;
wire n_1692;
wire n_1084;
wire n_800;
wire n_1171;
wire n_2169;
wire n_2371;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_2187;
wire n_662;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_2244;
wire n_2586;
wire n_1684;
wire n_921;
wire n_2446;
wire n_1346;
wire n_711;
wire n_1642;
wire n_1352;
wire n_937;
wire n_2257;
wire n_1682;
wire n_2017;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_2272;
wire n_2699;
wire n_2200;
wire n_650;
wire n_1046;
wire n_2560;
wire n_1940;
wire n_1979;
wire n_2704;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_2376;
wire n_1406;
wire n_1332;
wire n_2670;
wire n_2700;
wire n_962;
wire n_1041;
wire n_2346;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_2342;
wire n_2167;
wire n_2084;
wire n_2541;
wire n_654;
wire n_2518;
wire n_2458;
wire n_1222;
wire n_776;
wire n_1823;
wire n_2479;
wire n_1974;
wire n_2673;
wire n_2456;
wire n_1720;
wire n_2527;
wire n_934;
wire n_1637;
wire n_2635;
wire n_1407;
wire n_1795;
wire n_2688;
wire n_1341;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_2314;
wire n_942;
wire n_1524;
wire n_2229;
wire n_1964;
wire n_2288;
wire n_1920;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_2258;
wire n_1640;
wire n_804;
wire n_1846;
wire n_2406;
wire n_2390;
wire n_806;
wire n_879;
wire n_959;
wire n_2310;
wire n_2506;
wire n_2141;
wire n_2562;
wire n_2642;
wire n_1343;
wire n_1522;
wire n_1782;
wire n_2383;
wire n_2626;
wire n_1676;
wire n_833;
wire n_1830;
wire n_2351;
wire n_1567;
wire n_1319;
wire n_707;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_2536;
wire n_2196;
wire n_2629;
wire n_1633;
wire n_2195;
wire n_787;
wire n_2172;
wire n_1416;
wire n_1528;
wire n_2293;
wire n_1146;
wire n_2021;
wire n_2454;
wire n_2114;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_1282;
wire n_2561;
wire n_2567;
wire n_2322;
wire n_652;
wire n_2154;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_2533;
wire n_1758;
wire n_2283;
wire n_2422;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_2361;
wire n_1373;
wire n_1292;
wire n_2266;
wire n_2427;
wire n_1029;
wire n_1447;
wire n_2388;
wire n_2056;
wire n_790;
wire n_2611;
wire n_1706;
wire n_1498;
wire n_2653;
wire n_2417;
wire n_1210;
wire n_1248;
wire n_1556;
wire n_902;
wire n_2189;
wire n_2680;
wire n_2246;
wire n_1047;
wire n_1984;
wire n_2236;
wire n_1385;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_2668;
wire n_672;
wire n_2441;
wire n_1257;
wire n_1751;
wire n_1375;
wire n_1941;
wire n_2128;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_2398;
wire n_1872;
wire n_834;
wire n_2695;
wire n_743;
wire n_766;
wire n_1746;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1949;
wire n_2671;
wire n_1804;
wire n_1727;
wire n_2508;
wire n_1019;
wire n_636;
wire n_2054;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_2062;
wire n_2041;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_2070;
wire n_2588;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_2484;
wire n_2348;
wire n_2614;
wire n_2126;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_2253;
wire n_2366;
wire n_646;
wire n_1098;
wire n_1329;
wire n_2045;
wire n_817;
wire n_2261;
wire n_2216;
wire n_2210;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_2516;
wire n_1001;
wire n_1800;
wire n_2241;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_1191;
wire n_1826;
wire n_1023;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_2369;
wire n_1592;
wire n_855;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_1377;
wire n_1879;
wire n_853;
wire n_695;
wire n_1542;
wire n_2587;
wire n_875;
wire n_680;
wire n_1678;
wire n_2569;
wire n_661;
wire n_2400;
wire n_1716;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_1435;
wire n_969;
wire n_988;
wire n_2140;
wire n_1065;
wire n_2507;
wire n_1401;
wire n_2358;
wire n_1255;
wire n_1516;
wire n_1536;
wire n_2163;
wire n_2186;
wire n_2029;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_1074;
wire n_698;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_955;
wire n_739;
wire n_1379;
wire n_2528;
wire n_1338;
wire n_1097;
wire n_2395;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_769;
wire n_2380;
wire n_676;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_2295;
wire n_814;
wire n_1643;
wire n_2020;
wire n_2500;
wire n_2269;
wire n_1729;
wire n_669;
wire n_2290;
wire n_2048;
wire n_2005;
wire n_747;
wire n_2565;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_691;
wire n_2076;
wire n_1408;
wire n_1196;
wire n_1598;
wire n_863;
wire n_2175;
wire n_2182;
wire n_1283;
wire n_2385;
wire n_918;
wire n_748;
wire n_1848;
wire n_1114;
wire n_1785;
wire n_1147;
wire n_763;
wire n_1754;
wire n_2149;
wire n_2396;
wire n_1506;
wire n_2584;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_2450;
wire n_2485;
wire n_2284;
wire n_2566;
wire n_2287;
wire n_744;
wire n_971;
wire n_2702;
wire n_946;
wire n_761;
wire n_1303;
wire n_1205;
wire n_2492;
wire n_1258;
wire n_2438;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_2463;
wire n_1677;
wire n_1116;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_2180;
wire n_2679;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_1017;
wire n_2117;
wire n_2234;
wire n_2685;
wire n_1083;
wire n_1561;
wire n_930;
wire n_888;
wire n_2275;
wire n_1112;
wire n_2465;
wire n_2620;
wire n_2081;
wire n_2168;
wire n_2568;
wire n_2022;
wire n_2203;
wire n_1945;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_2112;
wire n_2255;
wire n_1464;
wire n_1737;
wire n_653;
wire n_2430;
wire n_1414;
wire n_908;
wire n_752;
wire n_2649;
wire n_944;
wire n_2034;
wire n_1028;
wire n_2106;
wire n_2265;
wire n_2615;
wire n_2683;
wire n_1922;
wire n_2032;
wire n_1011;
wire n_2474;
wire n_1566;
wire n_1215;
wire n_2437;
wire n_839;
wire n_2444;
wire n_708;
wire n_1973;
wire n_2267;
wire n_668;
wire n_990;
wire n_1500;
wire n_1537;
wire n_779;
wire n_1821;
wire n_2205;
wire n_1104;
wire n_1058;
wire n_854;
wire n_2312;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_1266;
wire n_709;
wire n_2242;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_2222;
wire n_712;
wire n_1276;
wire n_2015;
wire n_2118;
wire n_2111;
wire n_2466;
wire n_2530;
wire n_1148;
wire n_2188;
wire n_2505;
wire n_1989;
wire n_1161;
wire n_2609;
wire n_1085;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_771;
wire n_1584;
wire n_2425;
wire n_924;
wire n_1582;
wire n_2318;
wire n_2408;
wire n_1149;
wire n_1184;
wire n_2483;
wire n_719;
wire n_1972;
wire n_2592;
wire n_1525;
wire n_2594;
wire n_2666;
wire n_1585;
wire n_1851;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_2564;
wire n_1816;
wire n_2503;
wire n_2433;
wire n_1518;
wire n_1362;
wire n_1156;
wire n_829;
wire n_984;
wire n_2600;
wire n_1829;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_859;
wire n_2033;
wire n_735;
wire n_1789;
wire n_2531;
wire n_1770;
wire n_878;
wire n_2523;
wire n_1218;
wire n_2413;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_1144;
wire n_2071;
wire n_2429;
wire n_985;
wire n_2233;
wire n_2440;
wire n_997;
wire n_1710;
wire n_2161;
wire n_1301;
wire n_802;
wire n_980;
wire n_2681;
wire n_1306;
wire n_2010;
wire n_2282;
wire n_1651;
wire n_1198;
wire n_2360;
wire n_2047;
wire n_2651;
wire n_2095;
wire n_1609;
wire n_2174;
wire n_2334;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_2426;
wire n_2490;
wire n_756;
wire n_2303;
wire n_1619;
wire n_2478;
wire n_1981;
wire n_2285;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_2640;
wire n_1051;
wire n_1552;
wire n_1996;
wire n_2367;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_2248;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_2363;
wire n_2578;
wire n_849;
wire n_2662;
wire n_753;
wire n_1753;
wire n_2471;
wire n_2540;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_2197;
wire n_2217;
wire n_2065;
wire n_861;
wire n_857;
wire n_967;
wire n_2215;
wire n_2461;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_679;
wire n_1170;
wire n_665;
wire n_1629;
wire n_2221;
wire n_1260;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_2553;
wire n_1040;
wire n_915;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_2634;
wire n_1761;
wire n_2709;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_2477;
wire n_1888;
wire n_1557;
wire n_2280;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_2325;
wire n_670;
wire n_1850;
wire n_1898;
wire n_2443;
wire n_2697;
wire n_2308;
wire n_2162;
wire n_1868;
wire n_2333;
wire n_2079;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_2512;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_2185;
wire n_2086;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_2166;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_1958;
wire n_2077;
wire n_784;
wire n_1059;
wire n_1197;
wire n_2632;
wire n_2579;
wire n_722;
wire n_862;
wire n_2105;
wire n_2098;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_2223;
wire n_2091;
wire n_1915;
wire n_1621;
wire n_1748;
wire n_2547;
wire n_2415;
wire n_900;
wire n_1449;
wire n_827;
wire n_2659;
wire n_1025;
wire n_2419;
wire n_2116;
wire n_2320;
wire n_1885;
wire n_2677;
wire n_1013;
wire n_1259;
wire n_2183;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx2_ASAP7_75t_L g634 ( 
.A(n_159),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_520),
.Y(n_635)
);

INVx1_ASAP7_75t_SL g636 ( 
.A(n_163),
.Y(n_636)
);

BUFx10_ASAP7_75t_L g637 ( 
.A(n_298),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_442),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_359),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_35),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_377),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_124),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_74),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_229),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_591),
.Y(n_645)
);

CKINVDCx5p33_ASAP7_75t_R g646 ( 
.A(n_222),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_356),
.Y(n_647)
);

BUFx6f_ASAP7_75t_L g648 ( 
.A(n_512),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_229),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_535),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_575),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_102),
.Y(n_652)
);

CKINVDCx20_ASAP7_75t_R g653 ( 
.A(n_129),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_395),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_167),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_628),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_13),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_192),
.Y(n_658)
);

INVxp67_ASAP7_75t_SL g659 ( 
.A(n_511),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_617),
.Y(n_660)
);

BUFx10_ASAP7_75t_L g661 ( 
.A(n_457),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_557),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_66),
.Y(n_663)
);

BUFx8_ASAP7_75t_SL g664 ( 
.A(n_600),
.Y(n_664)
);

INVx2_ASAP7_75t_SL g665 ( 
.A(n_32),
.Y(n_665)
);

INVx1_ASAP7_75t_SL g666 ( 
.A(n_366),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_605),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_389),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_437),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_46),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_337),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_79),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_61),
.Y(n_673)
);

CKINVDCx20_ASAP7_75t_R g674 ( 
.A(n_216),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_560),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_286),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_263),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_521),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_419),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_3),
.Y(n_680)
);

CKINVDCx20_ASAP7_75t_R g681 ( 
.A(n_270),
.Y(n_681)
);

BUFx3_ASAP7_75t_L g682 ( 
.A(n_15),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_436),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_34),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_106),
.Y(n_685)
);

INVx1_ASAP7_75t_SL g686 ( 
.A(n_378),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_40),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_219),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_562),
.Y(n_689)
);

CKINVDCx20_ASAP7_75t_R g690 ( 
.A(n_555),
.Y(n_690)
);

INVx1_ASAP7_75t_SL g691 ( 
.A(n_254),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_393),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_581),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_580),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_387),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_384),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_380),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_438),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_162),
.Y(n_699)
);

CKINVDCx14_ASAP7_75t_R g700 ( 
.A(n_135),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_551),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_190),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_593),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_236),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_578),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_535),
.Y(n_706)
);

CKINVDCx20_ASAP7_75t_R g707 ( 
.A(n_403),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_554),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_225),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_540),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_410),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_154),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_316),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_270),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_627),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_74),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_48),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_91),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_392),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_139),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_123),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_304),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_135),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_383),
.Y(n_724)
);

BUFx10_ASAP7_75t_L g725 ( 
.A(n_12),
.Y(n_725)
);

CKINVDCx20_ASAP7_75t_R g726 ( 
.A(n_141),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_556),
.Y(n_727)
);

CKINVDCx20_ASAP7_75t_R g728 ( 
.A(n_561),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_243),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_558),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_490),
.Y(n_731)
);

CKINVDCx20_ASAP7_75t_R g732 ( 
.A(n_190),
.Y(n_732)
);

BUFx2_ASAP7_75t_L g733 ( 
.A(n_297),
.Y(n_733)
);

CKINVDCx20_ASAP7_75t_R g734 ( 
.A(n_178),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_479),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_172),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_184),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_137),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_454),
.Y(n_739)
);

INVx2_ASAP7_75t_SL g740 ( 
.A(n_251),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_386),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_488),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_403),
.Y(n_743)
);

INVx2_ASAP7_75t_SL g744 ( 
.A(n_595),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_632),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_609),
.Y(n_746)
);

BUFx3_ASAP7_75t_L g747 ( 
.A(n_589),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_52),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_121),
.Y(n_749)
);

BUFx10_ASAP7_75t_L g750 ( 
.A(n_329),
.Y(n_750)
);

CKINVDCx20_ASAP7_75t_R g751 ( 
.A(n_233),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_76),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_622),
.Y(n_753)
);

CKINVDCx20_ASAP7_75t_R g754 ( 
.A(n_613),
.Y(n_754)
);

CKINVDCx5p33_ASAP7_75t_R g755 ( 
.A(n_490),
.Y(n_755)
);

CKINVDCx5p33_ASAP7_75t_R g756 ( 
.A(n_301),
.Y(n_756)
);

BUFx6f_ASAP7_75t_L g757 ( 
.A(n_320),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_610),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_426),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_514),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_470),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_110),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_63),
.Y(n_763)
);

CKINVDCx5p33_ASAP7_75t_R g764 ( 
.A(n_264),
.Y(n_764)
);

CKINVDCx20_ASAP7_75t_R g765 ( 
.A(n_390),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_61),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_269),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_34),
.Y(n_768)
);

INVx1_ASAP7_75t_SL g769 ( 
.A(n_511),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_127),
.Y(n_770)
);

HB1xp67_ASAP7_75t_L g771 ( 
.A(n_361),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_461),
.Y(n_772)
);

BUFx6f_ASAP7_75t_L g773 ( 
.A(n_531),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_493),
.Y(n_774)
);

CKINVDCx20_ASAP7_75t_R g775 ( 
.A(n_498),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_119),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_436),
.Y(n_777)
);

CKINVDCx5p33_ASAP7_75t_R g778 ( 
.A(n_530),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_486),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_468),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_400),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_344),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_418),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_449),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_173),
.Y(n_785)
);

CKINVDCx5p33_ASAP7_75t_R g786 ( 
.A(n_485),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_332),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_435),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_39),
.Y(n_789)
);

BUFx2_ASAP7_75t_SL g790 ( 
.A(n_553),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_563),
.Y(n_791)
);

CKINVDCx5p33_ASAP7_75t_R g792 ( 
.A(n_60),
.Y(n_792)
);

CKINVDCx5p33_ASAP7_75t_R g793 ( 
.A(n_106),
.Y(n_793)
);

CKINVDCx5p33_ASAP7_75t_R g794 ( 
.A(n_319),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_332),
.Y(n_795)
);

CKINVDCx5p33_ASAP7_75t_R g796 ( 
.A(n_629),
.Y(n_796)
);

BUFx10_ASAP7_75t_L g797 ( 
.A(n_167),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_86),
.Y(n_798)
);

BUFx5_ASAP7_75t_L g799 ( 
.A(n_99),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_5),
.Y(n_800)
);

INVxp67_ASAP7_75t_L g801 ( 
.A(n_72),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_379),
.Y(n_802)
);

CKINVDCx5p33_ASAP7_75t_R g803 ( 
.A(n_291),
.Y(n_803)
);

CKINVDCx20_ASAP7_75t_R g804 ( 
.A(n_489),
.Y(n_804)
);

CKINVDCx20_ASAP7_75t_R g805 ( 
.A(n_602),
.Y(n_805)
);

CKINVDCx5p33_ASAP7_75t_R g806 ( 
.A(n_497),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_298),
.Y(n_807)
);

CKINVDCx5p33_ASAP7_75t_R g808 ( 
.A(n_163),
.Y(n_808)
);

BUFx3_ASAP7_75t_L g809 ( 
.A(n_552),
.Y(n_809)
);

CKINVDCx5p33_ASAP7_75t_R g810 ( 
.A(n_79),
.Y(n_810)
);

INVx1_ASAP7_75t_SL g811 ( 
.A(n_441),
.Y(n_811)
);

CKINVDCx5p33_ASAP7_75t_R g812 ( 
.A(n_477),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_331),
.Y(n_813)
);

CKINVDCx5p33_ASAP7_75t_R g814 ( 
.A(n_626),
.Y(n_814)
);

CKINVDCx5p33_ASAP7_75t_R g815 ( 
.A(n_255),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_250),
.Y(n_816)
);

CKINVDCx16_ASAP7_75t_R g817 ( 
.A(n_64),
.Y(n_817)
);

HB1xp67_ASAP7_75t_L g818 ( 
.A(n_458),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_216),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_215),
.Y(n_820)
);

CKINVDCx16_ASAP7_75t_R g821 ( 
.A(n_38),
.Y(n_821)
);

CKINVDCx5p33_ASAP7_75t_R g822 ( 
.A(n_206),
.Y(n_822)
);

CKINVDCx14_ASAP7_75t_R g823 ( 
.A(n_21),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_110),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_418),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_337),
.Y(n_826)
);

CKINVDCx5p33_ASAP7_75t_R g827 ( 
.A(n_437),
.Y(n_827)
);

CKINVDCx5p33_ASAP7_75t_R g828 ( 
.A(n_36),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_46),
.Y(n_829)
);

INVx1_ASAP7_75t_SL g830 ( 
.A(n_131),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_388),
.Y(n_831)
);

CKINVDCx20_ASAP7_75t_R g832 ( 
.A(n_187),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_120),
.Y(n_833)
);

INVx2_ASAP7_75t_SL g834 ( 
.A(n_300),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_508),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_379),
.Y(n_836)
);

CKINVDCx5p33_ASAP7_75t_R g837 ( 
.A(n_560),
.Y(n_837)
);

CKINVDCx5p33_ASAP7_75t_R g838 ( 
.A(n_33),
.Y(n_838)
);

CKINVDCx5p33_ASAP7_75t_R g839 ( 
.A(n_420),
.Y(n_839)
);

CKINVDCx5p33_ASAP7_75t_R g840 ( 
.A(n_559),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_397),
.Y(n_841)
);

CKINVDCx5p33_ASAP7_75t_R g842 ( 
.A(n_351),
.Y(n_842)
);

INVx2_ASAP7_75t_SL g843 ( 
.A(n_168),
.Y(n_843)
);

CKINVDCx5p33_ASAP7_75t_R g844 ( 
.A(n_514),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_518),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_10),
.Y(n_846)
);

CKINVDCx20_ASAP7_75t_R g847 ( 
.A(n_564),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_557),
.Y(n_848)
);

INVx3_ASAP7_75t_L g849 ( 
.A(n_101),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_474),
.Y(n_850)
);

CKINVDCx5p33_ASAP7_75t_R g851 ( 
.A(n_422),
.Y(n_851)
);

CKINVDCx5p33_ASAP7_75t_R g852 ( 
.A(n_235),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_273),
.Y(n_853)
);

CKINVDCx5p33_ASAP7_75t_R g854 ( 
.A(n_489),
.Y(n_854)
);

CKINVDCx5p33_ASAP7_75t_R g855 ( 
.A(n_192),
.Y(n_855)
);

BUFx2_ASAP7_75t_L g856 ( 
.A(n_3),
.Y(n_856)
);

CKINVDCx5p33_ASAP7_75t_R g857 ( 
.A(n_423),
.Y(n_857)
);

CKINVDCx5p33_ASAP7_75t_R g858 ( 
.A(n_261),
.Y(n_858)
);

BUFx3_ASAP7_75t_L g859 ( 
.A(n_552),
.Y(n_859)
);

CKINVDCx20_ASAP7_75t_R g860 ( 
.A(n_561),
.Y(n_860)
);

CKINVDCx5p33_ASAP7_75t_R g861 ( 
.A(n_433),
.Y(n_861)
);

CKINVDCx5p33_ASAP7_75t_R g862 ( 
.A(n_219),
.Y(n_862)
);

BUFx6f_ASAP7_75t_L g863 ( 
.A(n_574),
.Y(n_863)
);

CKINVDCx5p33_ASAP7_75t_R g864 ( 
.A(n_57),
.Y(n_864)
);

CKINVDCx5p33_ASAP7_75t_R g865 ( 
.A(n_407),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_799),
.Y(n_866)
);

CKINVDCx20_ASAP7_75t_R g867 ( 
.A(n_754),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_799),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_799),
.Y(n_869)
);

BUFx3_ASAP7_75t_L g870 ( 
.A(n_747),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_799),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_799),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_799),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_799),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_849),
.Y(n_875)
);

BUFx2_ASAP7_75t_L g876 ( 
.A(n_733),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_849),
.Y(n_877)
);

NOR2xp33_ASAP7_75t_L g878 ( 
.A(n_700),
.B(n_1),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_648),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_849),
.Y(n_880)
);

CKINVDCx5p33_ASAP7_75t_R g881 ( 
.A(n_823),
.Y(n_881)
);

NOR2xp67_ASAP7_75t_L g882 ( 
.A(n_801),
.B(n_0),
.Y(n_882)
);

INVxp67_ASAP7_75t_L g883 ( 
.A(n_856),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_648),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_648),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_648),
.Y(n_886)
);

CKINVDCx14_ASAP7_75t_R g887 ( 
.A(n_637),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_648),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_757),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_757),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_757),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_757),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_757),
.Y(n_893)
);

CKINVDCx20_ASAP7_75t_R g894 ( 
.A(n_754),
.Y(n_894)
);

INVxp33_ASAP7_75t_SL g895 ( 
.A(n_771),
.Y(n_895)
);

INVxp33_ASAP7_75t_L g896 ( 
.A(n_818),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_773),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_773),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_773),
.Y(n_899)
);

INVxp67_ASAP7_75t_SL g900 ( 
.A(n_747),
.Y(n_900)
);

BUFx6f_ASAP7_75t_L g901 ( 
.A(n_863),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_682),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_773),
.Y(n_903)
);

CKINVDCx5p33_ASAP7_75t_R g904 ( 
.A(n_817),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_682),
.Y(n_905)
);

CKINVDCx5p33_ASAP7_75t_R g906 ( 
.A(n_821),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_809),
.Y(n_907)
);

INVxp33_ASAP7_75t_SL g908 ( 
.A(n_635),
.Y(n_908)
);

BUFx3_ASAP7_75t_L g909 ( 
.A(n_745),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_809),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_859),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_859),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_773),
.Y(n_913)
);

CKINVDCx16_ASAP7_75t_R g914 ( 
.A(n_805),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_634),
.Y(n_915)
);

CKINVDCx5p33_ASAP7_75t_R g916 ( 
.A(n_639),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_634),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_638),
.Y(n_918)
);

NOR2xp67_ASAP7_75t_L g919 ( 
.A(n_665),
.B(n_0),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_640),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_652),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_657),
.Y(n_922)
);

INVx1_ASAP7_75t_SL g923 ( 
.A(n_637),
.Y(n_923)
);

BUFx3_ASAP7_75t_L g924 ( 
.A(n_746),
.Y(n_924)
);

INVxp67_ASAP7_75t_SL g925 ( 
.A(n_753),
.Y(n_925)
);

INVxp33_ASAP7_75t_SL g926 ( 
.A(n_635),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_669),
.Y(n_927)
);

CKINVDCx5p33_ASAP7_75t_R g928 ( 
.A(n_641),
.Y(n_928)
);

INVx1_ASAP7_75t_SL g929 ( 
.A(n_637),
.Y(n_929)
);

INVxp33_ASAP7_75t_SL g930 ( 
.A(n_658),
.Y(n_930)
);

CKINVDCx5p33_ASAP7_75t_R g931 ( 
.A(n_642),
.Y(n_931)
);

CKINVDCx16_ASAP7_75t_R g932 ( 
.A(n_805),
.Y(n_932)
);

INVxp67_ASAP7_75t_SL g933 ( 
.A(n_693),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_655),
.Y(n_934)
);

HB1xp67_ASAP7_75t_L g935 ( 
.A(n_658),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_678),
.Y(n_936)
);

HB1xp67_ASAP7_75t_L g937 ( 
.A(n_662),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_679),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_687),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_697),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_699),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_701),
.Y(n_942)
);

CKINVDCx5p33_ASAP7_75t_R g943 ( 
.A(n_643),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_704),
.Y(n_944)
);

CKINVDCx20_ASAP7_75t_R g945 ( 
.A(n_664),
.Y(n_945)
);

INVxp33_ASAP7_75t_L g946 ( 
.A(n_706),
.Y(n_946)
);

CKINVDCx16_ASAP7_75t_R g947 ( 
.A(n_661),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_712),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_713),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_655),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_696),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_696),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_748),
.Y(n_953)
);

CKINVDCx20_ASAP7_75t_R g954 ( 
.A(n_645),
.Y(n_954)
);

INVxp33_ASAP7_75t_L g955 ( 
.A(n_714),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_748),
.Y(n_956)
);

INVxp33_ASAP7_75t_L g957 ( 
.A(n_718),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_761),
.Y(n_958)
);

CKINVDCx5p33_ASAP7_75t_R g959 ( 
.A(n_644),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_761),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_762),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_762),
.Y(n_962)
);

INVxp33_ASAP7_75t_SL g963 ( 
.A(n_662),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_900),
.B(n_744),
.Y(n_964)
);

NOR2xp33_ASAP7_75t_L g965 ( 
.A(n_881),
.B(n_878),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_925),
.B(n_651),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_890),
.Y(n_967)
);

BUFx8_ASAP7_75t_SL g968 ( 
.A(n_945),
.Y(n_968)
);

BUFx3_ASAP7_75t_L g969 ( 
.A(n_870),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_870),
.B(n_694),
.Y(n_970)
);

CKINVDCx5p33_ASAP7_75t_R g971 ( 
.A(n_954),
.Y(n_971)
);

BUFx12f_ASAP7_75t_L g972 ( 
.A(n_881),
.Y(n_972)
);

AND2x4_ASAP7_75t_L g973 ( 
.A(n_933),
.B(n_863),
.Y(n_973)
);

BUFx6f_ASAP7_75t_L g974 ( 
.A(n_901),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_902),
.B(n_703),
.Y(n_975)
);

INVx2_ASAP7_75t_SL g976 ( 
.A(n_935),
.Y(n_976)
);

INVx5_ASAP7_75t_L g977 ( 
.A(n_901),
.Y(n_977)
);

AND2x2_ASAP7_75t_L g978 ( 
.A(n_905),
.B(n_665),
.Y(n_978)
);

BUFx8_ASAP7_75t_L g979 ( 
.A(n_876),
.Y(n_979)
);

INVx2_ASAP7_75t_L g980 ( 
.A(n_890),
.Y(n_980)
);

AND2x6_ASAP7_75t_L g981 ( 
.A(n_901),
.B(n_863),
.Y(n_981)
);

INVx4_ASAP7_75t_L g982 ( 
.A(n_901),
.Y(n_982)
);

BUFx8_ASAP7_75t_SL g983 ( 
.A(n_867),
.Y(n_983)
);

BUFx12f_ASAP7_75t_L g984 ( 
.A(n_904),
.Y(n_984)
);

AND2x4_ASAP7_75t_L g985 ( 
.A(n_880),
.B(n_875),
.Y(n_985)
);

BUFx6f_ASAP7_75t_L g986 ( 
.A(n_901),
.Y(n_986)
);

BUFx12f_ASAP7_75t_L g987 ( 
.A(n_904),
.Y(n_987)
);

BUFx12f_ASAP7_75t_L g988 ( 
.A(n_906),
.Y(n_988)
);

BUFx3_ASAP7_75t_L g989 ( 
.A(n_909),
.Y(n_989)
);

INVx5_ASAP7_75t_L g990 ( 
.A(n_903),
.Y(n_990)
);

INVx3_ASAP7_75t_L g991 ( 
.A(n_903),
.Y(n_991)
);

BUFx8_ASAP7_75t_L g992 ( 
.A(n_876),
.Y(n_992)
);

INVx2_ASAP7_75t_L g993 ( 
.A(n_879),
.Y(n_993)
);

AND2x4_ASAP7_75t_L g994 ( 
.A(n_880),
.B(n_863),
.Y(n_994)
);

INVx4_ASAP7_75t_L g995 ( 
.A(n_909),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_907),
.B(n_910),
.Y(n_996)
);

AND2x4_ASAP7_75t_L g997 ( 
.A(n_877),
.B(n_863),
.Y(n_997)
);

BUFx2_ASAP7_75t_L g998 ( 
.A(n_906),
.Y(n_998)
);

INVx5_ASAP7_75t_L g999 ( 
.A(n_915),
.Y(n_999)
);

AND2x4_ASAP7_75t_L g1000 ( 
.A(n_924),
.B(n_772),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_911),
.B(n_705),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_879),
.Y(n_1002)
);

HB1xp67_ASAP7_75t_L g1003 ( 
.A(n_916),
.Y(n_1003)
);

INVx3_ASAP7_75t_L g1004 ( 
.A(n_884),
.Y(n_1004)
);

NOR2xp33_ASAP7_75t_L g1005 ( 
.A(n_916),
.B(n_656),
.Y(n_1005)
);

INVx3_ASAP7_75t_L g1006 ( 
.A(n_884),
.Y(n_1006)
);

AND2x4_ASAP7_75t_L g1007 ( 
.A(n_924),
.B(n_772),
.Y(n_1007)
);

BUFx2_ASAP7_75t_L g1008 ( 
.A(n_928),
.Y(n_1008)
);

BUFx3_ASAP7_75t_L g1009 ( 
.A(n_912),
.Y(n_1009)
);

INVx5_ASAP7_75t_L g1010 ( 
.A(n_917),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_913),
.B(n_715),
.Y(n_1011)
);

CKINVDCx5p33_ASAP7_75t_R g1012 ( 
.A(n_914),
.Y(n_1012)
);

AND2x4_ASAP7_75t_L g1013 ( 
.A(n_885),
.B(n_781),
.Y(n_1013)
);

BUFx3_ASAP7_75t_L g1014 ( 
.A(n_885),
.Y(n_1014)
);

INVx3_ASAP7_75t_L g1015 ( 
.A(n_886),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_886),
.Y(n_1016)
);

BUFx2_ASAP7_75t_L g1017 ( 
.A(n_931),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_888),
.B(n_758),
.Y(n_1018)
);

NOR2x1_ASAP7_75t_L g1019 ( 
.A(n_888),
.B(n_720),
.Y(n_1019)
);

INVx2_ASAP7_75t_L g1020 ( 
.A(n_889),
.Y(n_1020)
);

AND2x2_ASAP7_75t_R g1021 ( 
.A(n_932),
.B(n_674),
.Y(n_1021)
);

NOR2x1_ASAP7_75t_L g1022 ( 
.A(n_889),
.B(n_721),
.Y(n_1022)
);

INVx3_ASAP7_75t_L g1023 ( 
.A(n_891),
.Y(n_1023)
);

INVx5_ASAP7_75t_L g1024 ( 
.A(n_917),
.Y(n_1024)
);

AND2x4_ASAP7_75t_L g1025 ( 
.A(n_891),
.B(n_781),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_892),
.B(n_796),
.Y(n_1026)
);

AND2x4_ASAP7_75t_L g1027 ( 
.A(n_969),
.B(n_989),
.Y(n_1027)
);

AND2x4_ASAP7_75t_L g1028 ( 
.A(n_969),
.B(n_934),
.Y(n_1028)
);

NOR3xp33_ASAP7_75t_L g1029 ( 
.A(n_976),
.B(n_947),
.C(n_883),
.Y(n_1029)
);

INVx2_ASAP7_75t_L g1030 ( 
.A(n_967),
.Y(n_1030)
);

AND2x2_ASAP7_75t_L g1031 ( 
.A(n_985),
.B(n_934),
.Y(n_1031)
);

INVx2_ASAP7_75t_L g1032 ( 
.A(n_967),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_1014),
.Y(n_1033)
);

NOR2xp33_ASAP7_75t_L g1034 ( 
.A(n_1005),
.B(n_908),
.Y(n_1034)
);

AND2x2_ASAP7_75t_L g1035 ( 
.A(n_985),
.B(n_950),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_1009),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_1009),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_985),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_1002),
.Y(n_1039)
);

BUFx2_ASAP7_75t_L g1040 ( 
.A(n_989),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_1002),
.Y(n_1041)
);

BUFx6f_ASAP7_75t_L g1042 ( 
.A(n_974),
.Y(n_1042)
);

INVx2_ASAP7_75t_L g1043 ( 
.A(n_980),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_1016),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_1016),
.Y(n_1045)
);

CKINVDCx20_ASAP7_75t_R g1046 ( 
.A(n_979),
.Y(n_1046)
);

BUFx6f_ASAP7_75t_L g1047 ( 
.A(n_974),
.Y(n_1047)
);

INVx2_ASAP7_75t_L g1048 ( 
.A(n_980),
.Y(n_1048)
);

BUFx3_ASAP7_75t_L g1049 ( 
.A(n_973),
.Y(n_1049)
);

BUFx3_ASAP7_75t_L g1050 ( 
.A(n_973),
.Y(n_1050)
);

BUFx6f_ASAP7_75t_L g1051 ( 
.A(n_974),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_994),
.Y(n_1052)
);

AND2x4_ASAP7_75t_L g1053 ( 
.A(n_1000),
.B(n_918),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_994),
.Y(n_1054)
);

INVx2_ASAP7_75t_L g1055 ( 
.A(n_993),
.Y(n_1055)
);

BUFx2_ASAP7_75t_L g1056 ( 
.A(n_979),
.Y(n_1056)
);

OA21x2_ASAP7_75t_L g1057 ( 
.A1(n_1018),
.A2(n_869),
.B(n_868),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_985),
.Y(n_1058)
);

BUFx2_ASAP7_75t_L g1059 ( 
.A(n_979),
.Y(n_1059)
);

INVx2_ASAP7_75t_L g1060 ( 
.A(n_993),
.Y(n_1060)
);

OR2x6_ASAP7_75t_L g1061 ( 
.A(n_984),
.B(n_790),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_994),
.Y(n_1062)
);

BUFx6f_ASAP7_75t_L g1063 ( 
.A(n_974),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_994),
.Y(n_1064)
);

BUFx2_ASAP7_75t_L g1065 ( 
.A(n_979),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_1004),
.Y(n_1066)
);

INVx2_ASAP7_75t_L g1067 ( 
.A(n_1020),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_1004),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_973),
.B(n_893),
.Y(n_1069)
);

NOR2x1_ASAP7_75t_L g1070 ( 
.A(n_995),
.B(n_919),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_1004),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_973),
.B(n_893),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_1006),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_1006),
.Y(n_1074)
);

NOR2x1_ASAP7_75t_L g1075 ( 
.A(n_995),
.B(n_871),
.Y(n_1075)
);

AND2x4_ASAP7_75t_L g1076 ( 
.A(n_1000),
.B(n_920),
.Y(n_1076)
);

INVx3_ASAP7_75t_L g1077 ( 
.A(n_974),
.Y(n_1077)
);

OAI21x1_ASAP7_75t_L g1078 ( 
.A1(n_964),
.A2(n_873),
.B(n_872),
.Y(n_1078)
);

INVx3_ASAP7_75t_L g1079 ( 
.A(n_986),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_1006),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_1015),
.Y(n_1081)
);

AND2x2_ASAP7_75t_L g1082 ( 
.A(n_978),
.B(n_950),
.Y(n_1082)
);

BUFx6f_ASAP7_75t_L g1083 ( 
.A(n_986),
.Y(n_1083)
);

INVx3_ASAP7_75t_L g1084 ( 
.A(n_986),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_1015),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_1015),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_1013),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_1013),
.Y(n_1088)
);

BUFx6f_ASAP7_75t_L g1089 ( 
.A(n_986),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_1013),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_1013),
.Y(n_1091)
);

BUFx6f_ASAP7_75t_L g1092 ( 
.A(n_986),
.Y(n_1092)
);

NAND2x1p5_ASAP7_75t_L g1093 ( 
.A(n_1019),
.B(n_866),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_1023),
.Y(n_1094)
);

AOI22xp5_ASAP7_75t_L g1095 ( 
.A1(n_965),
.A2(n_895),
.B1(n_943),
.B2(n_931),
.Y(n_1095)
);

BUFx6f_ASAP7_75t_L g1096 ( 
.A(n_977),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_1011),
.B(n_897),
.Y(n_1097)
);

AND2x2_ASAP7_75t_L g1098 ( 
.A(n_978),
.B(n_951),
.Y(n_1098)
);

OR2x2_ASAP7_75t_L g1099 ( 
.A(n_976),
.B(n_937),
.Y(n_1099)
);

INVx2_ASAP7_75t_L g1100 ( 
.A(n_1020),
.Y(n_1100)
);

AOI22xp5_ASAP7_75t_L g1101 ( 
.A1(n_966),
.A2(n_895),
.B1(n_959),
.B2(n_943),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_1025),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_1026),
.B(n_898),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_1023),
.Y(n_1104)
);

OAI22xp5_ASAP7_75t_SL g1105 ( 
.A1(n_1012),
.A2(n_653),
.B1(n_681),
.B2(n_674),
.Y(n_1105)
);

INVx2_ASAP7_75t_L g1106 ( 
.A(n_1023),
.Y(n_1106)
);

INVx2_ASAP7_75t_L g1107 ( 
.A(n_991),
.Y(n_1107)
);

INVx2_ASAP7_75t_L g1108 ( 
.A(n_991),
.Y(n_1108)
);

INVx6_ASAP7_75t_L g1109 ( 
.A(n_982),
.Y(n_1109)
);

HB1xp67_ASAP7_75t_L g1110 ( 
.A(n_970),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_SL g1111 ( 
.A(n_1034),
.B(n_1008),
.Y(n_1111)
);

AOI22xp33_ASAP7_75t_L g1112 ( 
.A1(n_1049),
.A2(n_930),
.B1(n_963),
.B2(n_926),
.Y(n_1112)
);

NAND3xp33_ASAP7_75t_L g1113 ( 
.A(n_1101),
.B(n_959),
.C(n_975),
.Y(n_1113)
);

INVx2_ASAP7_75t_L g1114 ( 
.A(n_1030),
.Y(n_1114)
);

AND2x2_ASAP7_75t_L g1115 ( 
.A(n_1082),
.B(n_1098),
.Y(n_1115)
);

INVx2_ASAP7_75t_L g1116 ( 
.A(n_1030),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_1052),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_1049),
.B(n_1001),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_SL g1119 ( 
.A(n_1027),
.B(n_1099),
.Y(n_1119)
);

INVx5_ASAP7_75t_L g1120 ( 
.A(n_1096),
.Y(n_1120)
);

AND2x6_ASAP7_75t_L g1121 ( 
.A(n_1050),
.B(n_1019),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_1052),
.Y(n_1122)
);

INVx2_ASAP7_75t_L g1123 ( 
.A(n_1032),
.Y(n_1123)
);

INVx2_ASAP7_75t_L g1124 ( 
.A(n_1032),
.Y(n_1124)
);

INVx1_ASAP7_75t_SL g1125 ( 
.A(n_1099),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_1054),
.Y(n_1126)
);

INVx2_ASAP7_75t_L g1127 ( 
.A(n_1043),
.Y(n_1127)
);

OAI22xp33_ASAP7_75t_L g1128 ( 
.A1(n_1110),
.A2(n_1017),
.B1(n_1003),
.B2(n_998),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_SL g1129 ( 
.A(n_1027),
.B(n_1017),
.Y(n_1129)
);

INVx2_ASAP7_75t_L g1130 ( 
.A(n_1043),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_1050),
.B(n_995),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_1054),
.Y(n_1132)
);

INVx3_ASAP7_75t_L g1133 ( 
.A(n_1106),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_SL g1134 ( 
.A(n_1027),
.B(n_998),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_SL g1135 ( 
.A(n_1095),
.B(n_992),
.Y(n_1135)
);

CKINVDCx5p33_ASAP7_75t_R g1136 ( 
.A(n_1046),
.Y(n_1136)
);

INVx3_ASAP7_75t_L g1137 ( 
.A(n_1106),
.Y(n_1137)
);

OR2x6_ASAP7_75t_L g1138 ( 
.A(n_1056),
.B(n_984),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_1062),
.Y(n_1139)
);

CKINVDCx5p33_ASAP7_75t_R g1140 ( 
.A(n_1046),
.Y(n_1140)
);

BUFx10_ASAP7_75t_L g1141 ( 
.A(n_1053),
.Y(n_1141)
);

INVx2_ASAP7_75t_L g1142 ( 
.A(n_1048),
.Y(n_1142)
);

INVx2_ASAP7_75t_L g1143 ( 
.A(n_1039),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_1064),
.Y(n_1144)
);

NOR2xp33_ASAP7_75t_L g1145 ( 
.A(n_1040),
.B(n_926),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_SL g1146 ( 
.A(n_1070),
.B(n_992),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_1035),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_1087),
.Y(n_1148)
);

INVx2_ASAP7_75t_L g1149 ( 
.A(n_1039),
.Y(n_1149)
);

CKINVDCx6p67_ASAP7_75t_R g1150 ( 
.A(n_1056),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_1087),
.Y(n_1151)
);

INVx2_ASAP7_75t_L g1152 ( 
.A(n_1041),
.Y(n_1152)
);

INVx2_ASAP7_75t_L g1153 ( 
.A(n_1041),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_1038),
.B(n_997),
.Y(n_1154)
);

INVx2_ASAP7_75t_L g1155 ( 
.A(n_1044),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_1058),
.B(n_997),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_1097),
.B(n_1022),
.Y(n_1157)
);

BUFx2_ASAP7_75t_L g1158 ( 
.A(n_1061),
.Y(n_1158)
);

INVx2_ASAP7_75t_L g1159 ( 
.A(n_1044),
.Y(n_1159)
);

INVx2_ASAP7_75t_L g1160 ( 
.A(n_1045),
.Y(n_1160)
);

INVx2_ASAP7_75t_L g1161 ( 
.A(n_1045),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_SL g1162 ( 
.A(n_1053),
.B(n_1076),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_1088),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_1090),
.Y(n_1164)
);

INVx2_ASAP7_75t_SL g1165 ( 
.A(n_1028),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_L g1166 ( 
.A(n_1103),
.B(n_1090),
.Y(n_1166)
);

BUFx10_ASAP7_75t_L g1167 ( 
.A(n_1053),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_1091),
.B(n_1102),
.Y(n_1168)
);

INVx1_ASAP7_75t_SL g1169 ( 
.A(n_1105),
.Y(n_1169)
);

BUFx6f_ASAP7_75t_L g1170 ( 
.A(n_1042),
.Y(n_1170)
);

INVx2_ASAP7_75t_L g1171 ( 
.A(n_1091),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_SL g1172 ( 
.A(n_1076),
.B(n_992),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_1102),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_1028),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_1028),
.Y(n_1175)
);

INVx2_ASAP7_75t_L g1176 ( 
.A(n_1055),
.Y(n_1176)
);

INVx2_ASAP7_75t_L g1177 ( 
.A(n_1055),
.Y(n_1177)
);

INVx2_ASAP7_75t_SL g1178 ( 
.A(n_1098),
.Y(n_1178)
);

BUFx6f_ASAP7_75t_L g1179 ( 
.A(n_1042),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_1060),
.Y(n_1180)
);

INVx3_ASAP7_75t_L g1181 ( 
.A(n_1060),
.Y(n_1181)
);

AND2x2_ASAP7_75t_L g1182 ( 
.A(n_1031),
.B(n_1000),
.Y(n_1182)
);

INVxp33_ASAP7_75t_L g1183 ( 
.A(n_1029),
.Y(n_1183)
);

NOR2xp33_ASAP7_75t_L g1184 ( 
.A(n_1036),
.B(n_887),
.Y(n_1184)
);

INVx2_ASAP7_75t_L g1185 ( 
.A(n_1067),
.Y(n_1185)
);

AOI21x1_ASAP7_75t_L g1186 ( 
.A1(n_1069),
.A2(n_874),
.B(n_866),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_SL g1187 ( 
.A(n_1037),
.B(n_972),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_1031),
.Y(n_1188)
);

NAND2xp33_ASAP7_75t_L g1189 ( 
.A(n_1093),
.B(n_981),
.Y(n_1189)
);

NOR2xp33_ASAP7_75t_L g1190 ( 
.A(n_1033),
.B(n_894),
.Y(n_1190)
);

INVx2_ASAP7_75t_L g1191 ( 
.A(n_1067),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_1100),
.Y(n_1192)
);

INVx2_ASAP7_75t_L g1193 ( 
.A(n_1100),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_1066),
.Y(n_1194)
);

INVx3_ASAP7_75t_L g1195 ( 
.A(n_1077),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_1068),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_1071),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_1073),
.Y(n_1198)
);

AND2x2_ASAP7_75t_L g1199 ( 
.A(n_1093),
.B(n_1007),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1074),
.Y(n_1200)
);

INVxp33_ASAP7_75t_L g1201 ( 
.A(n_1059),
.Y(n_1201)
);

INVx2_ASAP7_75t_L g1202 ( 
.A(n_1107),
.Y(n_1202)
);

INVx2_ASAP7_75t_L g1203 ( 
.A(n_1107),
.Y(n_1203)
);

INVx3_ASAP7_75t_L g1204 ( 
.A(n_1077),
.Y(n_1204)
);

CKINVDCx5p33_ASAP7_75t_R g1205 ( 
.A(n_1059),
.Y(n_1205)
);

CKINVDCx5p33_ASAP7_75t_R g1206 ( 
.A(n_1065),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_1080),
.Y(n_1207)
);

AND2x4_ASAP7_75t_L g1208 ( 
.A(n_1075),
.B(n_1007),
.Y(n_1208)
);

BUFx3_ASAP7_75t_L g1209 ( 
.A(n_1093),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_SL g1210 ( 
.A(n_1065),
.B(n_972),
.Y(n_1210)
);

INVx2_ASAP7_75t_L g1211 ( 
.A(n_1108),
.Y(n_1211)
);

INVx2_ASAP7_75t_L g1212 ( 
.A(n_1108),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1081),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_SL g1214 ( 
.A(n_1072),
.B(n_923),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_1085),
.B(n_982),
.Y(n_1215)
);

INVx3_ASAP7_75t_L g1216 ( 
.A(n_1077),
.Y(n_1216)
);

AO21x2_ASAP7_75t_L g1217 ( 
.A1(n_1078),
.A2(n_899),
.B(n_898),
.Y(n_1217)
);

AND2x2_ASAP7_75t_L g1218 ( 
.A(n_1057),
.B(n_1007),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_1086),
.B(n_982),
.Y(n_1219)
);

AOI22xp33_ASAP7_75t_L g1220 ( 
.A1(n_1057),
.A2(n_882),
.B1(n_1025),
.B2(n_659),
.Y(n_1220)
);

BUFx10_ASAP7_75t_L g1221 ( 
.A(n_1061),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_SL g1222 ( 
.A(n_1094),
.B(n_929),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1104),
.Y(n_1223)
);

AND2x2_ASAP7_75t_L g1224 ( 
.A(n_1057),
.B(n_996),
.Y(n_1224)
);

NOR2xp33_ASAP7_75t_L g1225 ( 
.A(n_1061),
.B(n_896),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1078),
.Y(n_1226)
);

BUFx6f_ASAP7_75t_SL g1227 ( 
.A(n_1061),
.Y(n_1227)
);

INVx2_ASAP7_75t_L g1228 ( 
.A(n_1079),
.Y(n_1228)
);

NOR2xp33_ASAP7_75t_L g1229 ( 
.A(n_1109),
.B(n_1012),
.Y(n_1229)
);

CKINVDCx5p33_ASAP7_75t_R g1230 ( 
.A(n_1079),
.Y(n_1230)
);

INVx2_ASAP7_75t_L g1231 ( 
.A(n_1079),
.Y(n_1231)
);

INVx8_ASAP7_75t_L g1232 ( 
.A(n_1042),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1084),
.Y(n_1233)
);

INVx2_ASAP7_75t_L g1234 ( 
.A(n_1084),
.Y(n_1234)
);

INVx2_ASAP7_75t_L g1235 ( 
.A(n_1084),
.Y(n_1235)
);

BUFx3_ASAP7_75t_L g1236 ( 
.A(n_1109),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_1042),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1117),
.Y(n_1238)
);

NOR2xp33_ASAP7_75t_L g1239 ( 
.A(n_1111),
.B(n_971),
.Y(n_1239)
);

AND2x2_ASAP7_75t_L g1240 ( 
.A(n_1115),
.B(n_971),
.Y(n_1240)
);

INVx2_ASAP7_75t_L g1241 ( 
.A(n_1171),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1117),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1132),
.Y(n_1243)
);

XOR2xp5_ASAP7_75t_L g1244 ( 
.A(n_1136),
.B(n_983),
.Y(n_1244)
);

AND2x2_ASAP7_75t_L g1245 ( 
.A(n_1115),
.B(n_987),
.Y(n_1245)
);

AND2x4_ASAP7_75t_L g1246 ( 
.A(n_1178),
.B(n_921),
.Y(n_1246)
);

NOR2xp33_ASAP7_75t_SL g1247 ( 
.A(n_1125),
.B(n_968),
.Y(n_1247)
);

HB1xp67_ASAP7_75t_L g1248 ( 
.A(n_1182),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1171),
.Y(n_1249)
);

XNOR2x1_ASAP7_75t_L g1250 ( 
.A(n_1169),
.B(n_1021),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1163),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1163),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1164),
.Y(n_1253)
);

CKINVDCx20_ASAP7_75t_R g1254 ( 
.A(n_1150),
.Y(n_1254)
);

INVxp33_ASAP7_75t_L g1255 ( 
.A(n_1145),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1164),
.Y(n_1256)
);

CKINVDCx20_ASAP7_75t_R g1257 ( 
.A(n_1150),
.Y(n_1257)
);

AND2x2_ASAP7_75t_L g1258 ( 
.A(n_1178),
.B(n_987),
.Y(n_1258)
);

BUFx6f_ASAP7_75t_L g1259 ( 
.A(n_1170),
.Y(n_1259)
);

CKINVDCx20_ASAP7_75t_R g1260 ( 
.A(n_1136),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1173),
.Y(n_1261)
);

INVx2_ASAP7_75t_L g1262 ( 
.A(n_1143),
.Y(n_1262)
);

CKINVDCx20_ASAP7_75t_R g1263 ( 
.A(n_1140),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1173),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1122),
.Y(n_1265)
);

CKINVDCx20_ASAP7_75t_R g1266 ( 
.A(n_1140),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1126),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1139),
.Y(n_1268)
);

XOR2xp5_ASAP7_75t_L g1269 ( 
.A(n_1113),
.B(n_653),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_L g1270 ( 
.A(n_1182),
.B(n_1042),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1139),
.Y(n_1271)
);

NOR2xp33_ASAP7_75t_L g1272 ( 
.A(n_1183),
.B(n_988),
.Y(n_1272)
);

INVx2_ASAP7_75t_L g1273 ( 
.A(n_1143),
.Y(n_1273)
);

XOR2xp5_ASAP7_75t_L g1274 ( 
.A(n_1205),
.B(n_681),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1144),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1144),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1148),
.Y(n_1277)
);

INVx2_ASAP7_75t_L g1278 ( 
.A(n_1149),
.Y(n_1278)
);

BUFx3_ASAP7_75t_L g1279 ( 
.A(n_1158),
.Y(n_1279)
);

NOR2xp33_ASAP7_75t_L g1280 ( 
.A(n_1119),
.B(n_690),
.Y(n_1280)
);

AND2x4_ASAP7_75t_L g1281 ( 
.A(n_1147),
.B(n_1188),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1151),
.Y(n_1282)
);

AND2x2_ASAP7_75t_L g1283 ( 
.A(n_1112),
.B(n_946),
.Y(n_1283)
);

NOR2xp33_ASAP7_75t_SL g1284 ( 
.A(n_1205),
.B(n_690),
.Y(n_1284)
);

AND2x4_ASAP7_75t_L g1285 ( 
.A(n_1165),
.B(n_922),
.Y(n_1285)
);

INVx4_ASAP7_75t_L g1286 ( 
.A(n_1232),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1174),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1175),
.Y(n_1288)
);

INVx4_ASAP7_75t_L g1289 ( 
.A(n_1232),
.Y(n_1289)
);

AND2x2_ASAP7_75t_L g1290 ( 
.A(n_1214),
.B(n_955),
.Y(n_1290)
);

NOR2xp33_ASAP7_75t_L g1291 ( 
.A(n_1128),
.B(n_707),
.Y(n_1291)
);

INVx2_ASAP7_75t_SL g1292 ( 
.A(n_1134),
.Y(n_1292)
);

INVx2_ASAP7_75t_L g1293 ( 
.A(n_1149),
.Y(n_1293)
);

NOR2xp33_ASAP7_75t_L g1294 ( 
.A(n_1190),
.B(n_707),
.Y(n_1294)
);

CKINVDCx20_ASAP7_75t_R g1295 ( 
.A(n_1206),
.Y(n_1295)
);

NOR2xp33_ASAP7_75t_L g1296 ( 
.A(n_1129),
.B(n_726),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1152),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1152),
.Y(n_1298)
);

XNOR2x2_ASAP7_75t_L g1299 ( 
.A(n_1135),
.B(n_636),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1153),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1153),
.Y(n_1301)
);

BUFx2_ASAP7_75t_L g1302 ( 
.A(n_1158),
.Y(n_1302)
);

NOR2xp33_ASAP7_75t_L g1303 ( 
.A(n_1118),
.B(n_1166),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1155),
.Y(n_1304)
);

CKINVDCx5p33_ASAP7_75t_R g1305 ( 
.A(n_1227),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1155),
.Y(n_1306)
);

XOR2x2_ASAP7_75t_L g1307 ( 
.A(n_1187),
.B(n_666),
.Y(n_1307)
);

XOR2x2_ASAP7_75t_L g1308 ( 
.A(n_1210),
.B(n_686),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_1159),
.B(n_1047),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_SL g1310 ( 
.A(n_1209),
.B(n_1047),
.Y(n_1310)
);

XNOR2x2_ASAP7_75t_L g1311 ( 
.A(n_1225),
.B(n_691),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1159),
.Y(n_1312)
);

BUFx3_ASAP7_75t_L g1313 ( 
.A(n_1138),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1160),
.Y(n_1314)
);

NOR2xp33_ASAP7_75t_L g1315 ( 
.A(n_1229),
.B(n_726),
.Y(n_1315)
);

NOR2xp33_ASAP7_75t_L g1316 ( 
.A(n_1157),
.B(n_728),
.Y(n_1316)
);

CKINVDCx5p33_ASAP7_75t_R g1317 ( 
.A(n_1138),
.Y(n_1317)
);

NOR2xp33_ASAP7_75t_L g1318 ( 
.A(n_1194),
.B(n_728),
.Y(n_1318)
);

INVxp33_ASAP7_75t_SL g1319 ( 
.A(n_1206),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1160),
.Y(n_1320)
);

AND2x2_ASAP7_75t_L g1321 ( 
.A(n_1184),
.B(n_957),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_SL g1322 ( 
.A(n_1209),
.B(n_1047),
.Y(n_1322)
);

OR2x2_ASAP7_75t_L g1323 ( 
.A(n_1222),
.B(n_769),
.Y(n_1323)
);

NOR2xp33_ASAP7_75t_L g1324 ( 
.A(n_1194),
.B(n_732),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1161),
.Y(n_1325)
);

BUFx2_ASAP7_75t_L g1326 ( 
.A(n_1138),
.Y(n_1326)
);

NOR2xp33_ASAP7_75t_L g1327 ( 
.A(n_1196),
.B(n_732),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1196),
.Y(n_1328)
);

NOR2xp33_ASAP7_75t_L g1329 ( 
.A(n_1197),
.B(n_734),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1197),
.Y(n_1330)
);

NAND2xp5_ASAP7_75t_SL g1331 ( 
.A(n_1199),
.B(n_1047),
.Y(n_1331)
);

NOR2xp33_ASAP7_75t_L g1332 ( 
.A(n_1198),
.B(n_734),
.Y(n_1332)
);

NOR2xp33_ASAP7_75t_L g1333 ( 
.A(n_1198),
.B(n_751),
.Y(n_1333)
);

INVxp33_ASAP7_75t_SL g1334 ( 
.A(n_1146),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1200),
.Y(n_1335)
);

NOR2xp33_ASAP7_75t_L g1336 ( 
.A(n_1200),
.B(n_751),
.Y(n_1336)
);

INVx3_ASAP7_75t_R g1337 ( 
.A(n_1208),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1207),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1207),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1213),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1213),
.Y(n_1341)
);

CKINVDCx14_ASAP7_75t_R g1342 ( 
.A(n_1138),
.Y(n_1342)
);

XOR2xp5_ASAP7_75t_L g1343 ( 
.A(n_1201),
.B(n_765),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1223),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1223),
.Y(n_1345)
);

BUFx6f_ASAP7_75t_L g1346 ( 
.A(n_1170),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1180),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1180),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1192),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1168),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1165),
.Y(n_1351)
);

OR2x6_ASAP7_75t_L g1352 ( 
.A(n_1172),
.B(n_740),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1202),
.Y(n_1353)
);

XOR2xp5_ASAP7_75t_L g1354 ( 
.A(n_1208),
.B(n_765),
.Y(n_1354)
);

NOR2xp33_ASAP7_75t_L g1355 ( 
.A(n_1162),
.B(n_775),
.Y(n_1355)
);

BUFx3_ASAP7_75t_L g1356 ( 
.A(n_1221),
.Y(n_1356)
);

CKINVDCx20_ASAP7_75t_R g1357 ( 
.A(n_1221),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1203),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1203),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1211),
.Y(n_1360)
);

AND2x2_ASAP7_75t_L g1361 ( 
.A(n_1199),
.B(n_661),
.Y(n_1361)
);

OR2x2_ASAP7_75t_L g1362 ( 
.A(n_1220),
.B(n_811),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1212),
.Y(n_1363)
);

CKINVDCx5p33_ASAP7_75t_R g1364 ( 
.A(n_1221),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1212),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1176),
.Y(n_1366)
);

INVxp33_ASAP7_75t_L g1367 ( 
.A(n_1224),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1176),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1177),
.Y(n_1369)
);

NOR2xp33_ASAP7_75t_L g1370 ( 
.A(n_1131),
.B(n_775),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1177),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1185),
.Y(n_1372)
);

NOR2xp33_ASAP7_75t_L g1373 ( 
.A(n_1224),
.B(n_804),
.Y(n_1373)
);

XOR2xp5_ASAP7_75t_L g1374 ( 
.A(n_1208),
.B(n_804),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1185),
.Y(n_1375)
);

INVx1_ASAP7_75t_SL g1376 ( 
.A(n_1141),
.Y(n_1376)
);

XOR2xp5_ASAP7_75t_L g1377 ( 
.A(n_1230),
.B(n_1154),
.Y(n_1377)
);

NAND2xp33_ASAP7_75t_R g1378 ( 
.A(n_1218),
.B(n_663),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1191),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1193),
.Y(n_1380)
);

NOR2xp33_ASAP7_75t_L g1381 ( 
.A(n_1156),
.B(n_832),
.Y(n_1381)
);

INVx2_ASAP7_75t_L g1382 ( 
.A(n_1114),
.Y(n_1382)
);

NOR2xp33_ASAP7_75t_SL g1383 ( 
.A(n_1141),
.B(n_832),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1116),
.Y(n_1384)
);

INVx2_ASAP7_75t_L g1385 ( 
.A(n_1116),
.Y(n_1385)
);

XNOR2xp5_ASAP7_75t_L g1386 ( 
.A(n_1186),
.B(n_847),
.Y(n_1386)
);

NOR2xp33_ASAP7_75t_L g1387 ( 
.A(n_1181),
.B(n_847),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1123),
.Y(n_1388)
);

INVx2_ASAP7_75t_L g1389 ( 
.A(n_1123),
.Y(n_1389)
);

OR2x2_ASAP7_75t_SL g1390 ( 
.A(n_1226),
.B(n_791),
.Y(n_1390)
);

CKINVDCx20_ASAP7_75t_R g1391 ( 
.A(n_1167),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1124),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1127),
.Y(n_1393)
);

NOR2xp33_ASAP7_75t_L g1394 ( 
.A(n_1181),
.B(n_1133),
.Y(n_1394)
);

CKINVDCx5p33_ASAP7_75t_R g1395 ( 
.A(n_1167),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1127),
.Y(n_1396)
);

AND2x2_ASAP7_75t_SL g1397 ( 
.A(n_1189),
.B(n_791),
.Y(n_1397)
);

AOI21xp5_ASAP7_75t_L g1398 ( 
.A1(n_1189),
.A2(n_1063),
.B(n_1051),
.Y(n_1398)
);

INVx1_ASAP7_75t_SL g1399 ( 
.A(n_1121),
.Y(n_1399)
);

INVx2_ASAP7_75t_L g1400 ( 
.A(n_1130),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_L g1401 ( 
.A(n_1236),
.B(n_1051),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1130),
.Y(n_1402)
);

INVx2_ASAP7_75t_SL g1403 ( 
.A(n_1228),
.Y(n_1403)
);

BUFx3_ASAP7_75t_L g1404 ( 
.A(n_1121),
.Y(n_1404)
);

XOR2x2_ASAP7_75t_L g1405 ( 
.A(n_1217),
.B(n_830),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1142),
.Y(n_1406)
);

CKINVDCx20_ASAP7_75t_R g1407 ( 
.A(n_1217),
.Y(n_1407)
);

NOR2xp33_ASAP7_75t_SL g1408 ( 
.A(n_1121),
.B(n_860),
.Y(n_1408)
);

INVxp33_ASAP7_75t_L g1409 ( 
.A(n_1228),
.Y(n_1409)
);

NAND2xp5_ASAP7_75t_L g1410 ( 
.A(n_1121),
.B(n_1051),
.Y(n_1410)
);

AND2x2_ASAP7_75t_SL g1411 ( 
.A(n_1226),
.B(n_798),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1133),
.Y(n_1412)
);

BUFx6f_ASAP7_75t_L g1413 ( 
.A(n_1259),
.Y(n_1413)
);

AND2x2_ASAP7_75t_L g1414 ( 
.A(n_1316),
.B(n_725),
.Y(n_1414)
);

AND2x2_ASAP7_75t_L g1415 ( 
.A(n_1316),
.B(n_1381),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_L g1416 ( 
.A(n_1303),
.B(n_1121),
.Y(n_1416)
);

NOR2xp33_ASAP7_75t_L g1417 ( 
.A(n_1255),
.B(n_1233),
.Y(n_1417)
);

NAND2x1p5_ASAP7_75t_L g1418 ( 
.A(n_1286),
.B(n_1289),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1249),
.Y(n_1419)
);

INVx2_ASAP7_75t_L g1420 ( 
.A(n_1241),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1303),
.B(n_1181),
.Y(n_1421)
);

OAI22xp5_ASAP7_75t_L g1422 ( 
.A1(n_1373),
.A2(n_860),
.B1(n_1204),
.B2(n_1195),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1238),
.Y(n_1423)
);

NOR2xp33_ASAP7_75t_L g1424 ( 
.A(n_1255),
.B(n_1233),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_SL g1425 ( 
.A(n_1408),
.B(n_1179),
.Y(n_1425)
);

NAND2xp33_ASAP7_75t_L g1426 ( 
.A(n_1350),
.B(n_1170),
.Y(n_1426)
);

AOI22xp5_ASAP7_75t_L g1427 ( 
.A1(n_1373),
.A2(n_1217),
.B1(n_1137),
.B2(n_1133),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1242),
.Y(n_1428)
);

NAND2xp5_ASAP7_75t_L g1429 ( 
.A(n_1248),
.B(n_1137),
.Y(n_1429)
);

NAND2xp5_ASAP7_75t_L g1430 ( 
.A(n_1248),
.B(n_1137),
.Y(n_1430)
);

OR2x2_ASAP7_75t_L g1431 ( 
.A(n_1240),
.B(n_1231),
.Y(n_1431)
);

OR2x2_ASAP7_75t_L g1432 ( 
.A(n_1315),
.B(n_1294),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1243),
.Y(n_1433)
);

AND2x2_ASAP7_75t_L g1434 ( 
.A(n_1381),
.B(n_750),
.Y(n_1434)
);

BUFx6f_ASAP7_75t_SL g1435 ( 
.A(n_1313),
.Y(n_1435)
);

INVx2_ASAP7_75t_L g1436 ( 
.A(n_1262),
.Y(n_1436)
);

OAI21xp5_ASAP7_75t_L g1437 ( 
.A1(n_1367),
.A2(n_1186),
.B(n_1215),
.Y(n_1437)
);

INVxp67_ASAP7_75t_L g1438 ( 
.A(n_1302),
.Y(n_1438)
);

BUFx6f_ASAP7_75t_L g1439 ( 
.A(n_1259),
.Y(n_1439)
);

AOI22xp5_ASAP7_75t_L g1440 ( 
.A1(n_1407),
.A2(n_1219),
.B1(n_1234),
.B2(n_1231),
.Y(n_1440)
);

AOI221xp5_ASAP7_75t_L g1441 ( 
.A1(n_1294),
.A2(n_759),
.B1(n_858),
.B2(n_749),
.C(n_663),
.Y(n_1441)
);

AOI22xp5_ASAP7_75t_L g1442 ( 
.A1(n_1411),
.A2(n_1235),
.B1(n_1234),
.B2(n_1025),
.Y(n_1442)
);

AOI22xp5_ASAP7_75t_L g1443 ( 
.A1(n_1411),
.A2(n_1370),
.B1(n_1281),
.B2(n_1378),
.Y(n_1443)
);

INVx2_ASAP7_75t_L g1444 ( 
.A(n_1273),
.Y(n_1444)
);

NAND2xp5_ASAP7_75t_L g1445 ( 
.A(n_1268),
.B(n_1204),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_SL g1446 ( 
.A(n_1383),
.B(n_1179),
.Y(n_1446)
);

NAND2xp5_ASAP7_75t_L g1447 ( 
.A(n_1271),
.B(n_1216),
.Y(n_1447)
);

AOI22xp33_ASAP7_75t_L g1448 ( 
.A1(n_1281),
.A2(n_1362),
.B1(n_1280),
.B2(n_1355),
.Y(n_1448)
);

INVx2_ASAP7_75t_L g1449 ( 
.A(n_1278),
.Y(n_1449)
);

BUFx2_ASAP7_75t_L g1450 ( 
.A(n_1295),
.Y(n_1450)
);

NAND2xp5_ASAP7_75t_L g1451 ( 
.A(n_1275),
.B(n_1216),
.Y(n_1451)
);

INVx2_ASAP7_75t_L g1452 ( 
.A(n_1293),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_L g1453 ( 
.A(n_1276),
.B(n_1216),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1251),
.Y(n_1454)
);

NOR2xp33_ASAP7_75t_L g1455 ( 
.A(n_1280),
.B(n_1235),
.Y(n_1455)
);

BUFx5_ASAP7_75t_L g1456 ( 
.A(n_1404),
.Y(n_1456)
);

NAND2xp5_ASAP7_75t_SL g1457 ( 
.A(n_1245),
.B(n_1179),
.Y(n_1457)
);

OR2x6_ASAP7_75t_L g1458 ( 
.A(n_1326),
.B(n_1232),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1252),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_L g1460 ( 
.A(n_1265),
.B(n_1237),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_L g1461 ( 
.A(n_1267),
.B(n_1237),
.Y(n_1461)
);

NAND2xp5_ASAP7_75t_SL g1462 ( 
.A(n_1292),
.B(n_1179),
.Y(n_1462)
);

AOI22xp5_ASAP7_75t_L g1463 ( 
.A1(n_1378),
.A2(n_814),
.B1(n_667),
.B2(n_660),
.Y(n_1463)
);

NAND2xp5_ASAP7_75t_SL g1464 ( 
.A(n_1258),
.B(n_1232),
.Y(n_1464)
);

AOI22xp5_ASAP7_75t_L g1465 ( 
.A1(n_1277),
.A2(n_1282),
.B1(n_1256),
.B2(n_1261),
.Y(n_1465)
);

AND2x2_ASAP7_75t_L g1466 ( 
.A(n_1321),
.B(n_750),
.Y(n_1466)
);

NAND2xp5_ASAP7_75t_L g1467 ( 
.A(n_1328),
.B(n_991),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_L g1468 ( 
.A(n_1330),
.B(n_646),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1253),
.Y(n_1469)
);

NAND2xp33_ASAP7_75t_L g1470 ( 
.A(n_1346),
.B(n_1051),
.Y(n_1470)
);

INVx2_ASAP7_75t_SL g1471 ( 
.A(n_1279),
.Y(n_1471)
);

INVx2_ASAP7_75t_L g1472 ( 
.A(n_1382),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1264),
.Y(n_1473)
);

BUFx6f_ASAP7_75t_L g1474 ( 
.A(n_1346),
.Y(n_1474)
);

INVx2_ASAP7_75t_L g1475 ( 
.A(n_1385),
.Y(n_1475)
);

AND2x6_ASAP7_75t_L g1476 ( 
.A(n_1399),
.B(n_798),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1318),
.B(n_1324),
.Y(n_1477)
);

BUFx3_ASAP7_75t_L g1478 ( 
.A(n_1356),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1297),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_L g1480 ( 
.A(n_1335),
.B(n_647),
.Y(n_1480)
);

BUFx3_ASAP7_75t_L g1481 ( 
.A(n_1260),
.Y(n_1481)
);

NOR2xp33_ASAP7_75t_L g1482 ( 
.A(n_1296),
.B(n_649),
.Y(n_1482)
);

AOI22xp5_ASAP7_75t_L g1483 ( 
.A1(n_1387),
.A2(n_899),
.B1(n_843),
.B2(n_834),
.Y(n_1483)
);

NAND2xp5_ASAP7_75t_L g1484 ( 
.A(n_1338),
.B(n_650),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1298),
.Y(n_1485)
);

CKINVDCx5p33_ASAP7_75t_R g1486 ( 
.A(n_1263),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1300),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_L g1488 ( 
.A(n_1339),
.B(n_654),
.Y(n_1488)
);

INVx3_ASAP7_75t_L g1489 ( 
.A(n_1286),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_L g1490 ( 
.A(n_1340),
.B(n_668),
.Y(n_1490)
);

OAI22xp33_ASAP7_75t_L g1491 ( 
.A1(n_1284),
.A2(n_843),
.B1(n_834),
.B2(n_759),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_L g1492 ( 
.A(n_1341),
.B(n_670),
.Y(n_1492)
);

NOR2xp67_ASAP7_75t_L g1493 ( 
.A(n_1272),
.B(n_571),
.Y(n_1493)
);

NOR2xp33_ASAP7_75t_L g1494 ( 
.A(n_1296),
.B(n_671),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_1344),
.B(n_672),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1301),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_L g1497 ( 
.A(n_1345),
.B(n_673),
.Y(n_1497)
);

INVx8_ASAP7_75t_L g1498 ( 
.A(n_1346),
.Y(n_1498)
);

NOR2xp33_ASAP7_75t_L g1499 ( 
.A(n_1355),
.B(n_675),
.Y(n_1499)
);

NOR2xp67_ASAP7_75t_L g1500 ( 
.A(n_1272),
.B(n_572),
.Y(n_1500)
);

NAND2xp5_ASAP7_75t_L g1501 ( 
.A(n_1361),
.B(n_676),
.Y(n_1501)
);

OA22x2_ASAP7_75t_L g1502 ( 
.A1(n_1269),
.A2(n_864),
.B1(n_858),
.B2(n_861),
.Y(n_1502)
);

INVx2_ASAP7_75t_L g1503 ( 
.A(n_1389),
.Y(n_1503)
);

NAND2xp5_ASAP7_75t_L g1504 ( 
.A(n_1246),
.B(n_677),
.Y(n_1504)
);

INVxp67_ASAP7_75t_L g1505 ( 
.A(n_1290),
.Y(n_1505)
);

OR2x2_ASAP7_75t_L g1506 ( 
.A(n_1323),
.B(n_927),
.Y(n_1506)
);

NAND2xp5_ASAP7_75t_L g1507 ( 
.A(n_1246),
.B(n_680),
.Y(n_1507)
);

INVx8_ASAP7_75t_L g1508 ( 
.A(n_1391),
.Y(n_1508)
);

NOR2xp33_ASAP7_75t_L g1509 ( 
.A(n_1239),
.B(n_683),
.Y(n_1509)
);

INVx2_ASAP7_75t_L g1510 ( 
.A(n_1400),
.Y(n_1510)
);

INVx2_ASAP7_75t_L g1511 ( 
.A(n_1304),
.Y(n_1511)
);

NOR2xp33_ASAP7_75t_L g1512 ( 
.A(n_1239),
.B(n_1377),
.Y(n_1512)
);

OAI221xp5_ASAP7_75t_L g1513 ( 
.A1(n_1291),
.A2(n_862),
.B1(n_864),
.B2(n_861),
.C(n_749),
.Y(n_1513)
);

INVx3_ASAP7_75t_L g1514 ( 
.A(n_1351),
.Y(n_1514)
);

INVx2_ASAP7_75t_L g1515 ( 
.A(n_1306),
.Y(n_1515)
);

NAND2xp5_ASAP7_75t_L g1516 ( 
.A(n_1285),
.B(n_684),
.Y(n_1516)
);

INVxp67_ASAP7_75t_L g1517 ( 
.A(n_1354),
.Y(n_1517)
);

NOR2xp33_ASAP7_75t_L g1518 ( 
.A(n_1291),
.B(n_685),
.Y(n_1518)
);

NAND2xp5_ASAP7_75t_SL g1519 ( 
.A(n_1334),
.B(n_1063),
.Y(n_1519)
);

NOR2xp33_ASAP7_75t_L g1520 ( 
.A(n_1324),
.B(n_1327),
.Y(n_1520)
);

NAND2xp5_ASAP7_75t_SL g1521 ( 
.A(n_1327),
.B(n_1063),
.Y(n_1521)
);

NOR2xp33_ASAP7_75t_L g1522 ( 
.A(n_1329),
.B(n_688),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_L g1523 ( 
.A(n_1285),
.B(n_689),
.Y(n_1523)
);

BUFx2_ASAP7_75t_L g1524 ( 
.A(n_1266),
.Y(n_1524)
);

OAI22xp5_ASAP7_75t_SL g1525 ( 
.A1(n_1274),
.A2(n_1374),
.B1(n_1343),
.B2(n_1319),
.Y(n_1525)
);

OAI22xp33_ASAP7_75t_L g1526 ( 
.A1(n_1352),
.A2(n_862),
.B1(n_833),
.B2(n_816),
.Y(n_1526)
);

INVxp67_ASAP7_75t_L g1527 ( 
.A(n_1329),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1287),
.B(n_692),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_L g1529 ( 
.A(n_1288),
.B(n_695),
.Y(n_1529)
);

AOI22xp5_ASAP7_75t_L g1530 ( 
.A1(n_1397),
.A2(n_702),
.B1(n_708),
.B2(n_698),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_L g1531 ( 
.A(n_1367),
.B(n_709),
.Y(n_1531)
);

NOR2xp33_ASAP7_75t_L g1532 ( 
.A(n_1332),
.B(n_710),
.Y(n_1532)
);

INVxp67_ASAP7_75t_L g1533 ( 
.A(n_1332),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_L g1534 ( 
.A(n_1333),
.B(n_711),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_L g1535 ( 
.A(n_1333),
.B(n_716),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1312),
.Y(n_1536)
);

BUFx6f_ASAP7_75t_L g1537 ( 
.A(n_1395),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1314),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1320),
.Y(n_1539)
);

NAND2xp5_ASAP7_75t_SL g1540 ( 
.A(n_1336),
.B(n_1376),
.Y(n_1540)
);

AND2x2_ASAP7_75t_L g1541 ( 
.A(n_1336),
.B(n_750),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1325),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_L g1543 ( 
.A(n_1347),
.B(n_717),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1348),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_L g1545 ( 
.A(n_1349),
.B(n_719),
.Y(n_1545)
);

NOR2xp33_ASAP7_75t_L g1546 ( 
.A(n_1283),
.B(n_722),
.Y(n_1546)
);

INVx4_ASAP7_75t_L g1547 ( 
.A(n_1364),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_L g1548 ( 
.A(n_1270),
.B(n_723),
.Y(n_1548)
);

INVx2_ASAP7_75t_L g1549 ( 
.A(n_1353),
.Y(n_1549)
);

INVx2_ASAP7_75t_L g1550 ( 
.A(n_1358),
.Y(n_1550)
);

INVx2_ASAP7_75t_L g1551 ( 
.A(n_1359),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_L g1552 ( 
.A(n_1409),
.B(n_727),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_L g1553 ( 
.A(n_1409),
.B(n_729),
.Y(n_1553)
);

NOR2xp33_ASAP7_75t_L g1554 ( 
.A(n_1386),
.B(n_731),
.Y(n_1554)
);

INVx2_ASAP7_75t_L g1555 ( 
.A(n_1360),
.Y(n_1555)
);

AOI22xp5_ASAP7_75t_L g1556 ( 
.A1(n_1405),
.A2(n_737),
.B1(n_738),
.B2(n_736),
.Y(n_1556)
);

NAND2xp33_ASAP7_75t_L g1557 ( 
.A(n_1410),
.B(n_1083),
.Y(n_1557)
);

CKINVDCx6p67_ASAP7_75t_R g1558 ( 
.A(n_1254),
.Y(n_1558)
);

INVx2_ASAP7_75t_L g1559 ( 
.A(n_1363),
.Y(n_1559)
);

INVx2_ASAP7_75t_L g1560 ( 
.A(n_1365),
.Y(n_1560)
);

INVx2_ASAP7_75t_L g1561 ( 
.A(n_1366),
.Y(n_1561)
);

NOR2xp33_ASAP7_75t_L g1562 ( 
.A(n_1250),
.B(n_739),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1307),
.B(n_797),
.Y(n_1563)
);

INVxp67_ASAP7_75t_L g1564 ( 
.A(n_1311),
.Y(n_1564)
);

BUFx3_ASAP7_75t_L g1565 ( 
.A(n_1257),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_L g1566 ( 
.A(n_1368),
.B(n_741),
.Y(n_1566)
);

NAND2xp5_ASAP7_75t_L g1567 ( 
.A(n_1369),
.B(n_742),
.Y(n_1567)
);

NOR2xp33_ASAP7_75t_L g1568 ( 
.A(n_1352),
.B(n_743),
.Y(n_1568)
);

NOR2xp33_ASAP7_75t_L g1569 ( 
.A(n_1352),
.B(n_752),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1308),
.B(n_797),
.Y(n_1570)
);

OR2x6_ASAP7_75t_L g1571 ( 
.A(n_1337),
.B(n_816),
.Y(n_1571)
);

INVx2_ASAP7_75t_SL g1572 ( 
.A(n_1299),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1371),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_L g1574 ( 
.A(n_1372),
.B(n_755),
.Y(n_1574)
);

AND2x6_ASAP7_75t_L g1575 ( 
.A(n_1375),
.B(n_833),
.Y(n_1575)
);

BUFx3_ASAP7_75t_L g1576 ( 
.A(n_1357),
.Y(n_1576)
);

CKINVDCx20_ASAP7_75t_R g1577 ( 
.A(n_1244),
.Y(n_1577)
);

NOR2xp33_ASAP7_75t_L g1578 ( 
.A(n_1390),
.B(n_756),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_L g1579 ( 
.A(n_1379),
.B(n_760),
.Y(n_1579)
);

INVx3_ASAP7_75t_L g1580 ( 
.A(n_1412),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1380),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1384),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1388),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1392),
.Y(n_1584)
);

OAI22xp5_ASAP7_75t_L g1585 ( 
.A1(n_1394),
.A2(n_730),
.B1(n_735),
.B2(n_724),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_SL g1586 ( 
.A(n_1247),
.B(n_1083),
.Y(n_1586)
);

NAND2xp33_ASAP7_75t_L g1587 ( 
.A(n_1403),
.B(n_1089),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1393),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_SL g1589 ( 
.A(n_1305),
.B(n_1089),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1406),
.B(n_1092),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_SL g1591 ( 
.A(n_1520),
.B(n_1317),
.Y(n_1591)
);

AOI21xp5_ASAP7_75t_L g1592 ( 
.A1(n_1426),
.A2(n_1398),
.B(n_1401),
.Y(n_1592)
);

BUFx2_ASAP7_75t_L g1593 ( 
.A(n_1438),
.Y(n_1593)
);

NOR2xp33_ASAP7_75t_L g1594 ( 
.A(n_1432),
.B(n_1342),
.Y(n_1594)
);

OAI22xp5_ASAP7_75t_L g1595 ( 
.A1(n_1443),
.A2(n_1310),
.B1(n_1322),
.B2(n_1394),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_SL g1596 ( 
.A(n_1477),
.B(n_1310),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_L g1597 ( 
.A(n_1415),
.B(n_1396),
.Y(n_1597)
);

AOI21xp5_ASAP7_75t_L g1598 ( 
.A1(n_1470),
.A2(n_1331),
.B(n_1322),
.Y(n_1598)
);

AOI22xp5_ASAP7_75t_L g1599 ( 
.A1(n_1509),
.A2(n_1342),
.B1(n_1402),
.B2(n_1309),
.Y(n_1599)
);

BUFx4f_ASAP7_75t_L g1600 ( 
.A(n_1537),
.Y(n_1600)
);

INVx4_ASAP7_75t_L g1601 ( 
.A(n_1498),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_L g1602 ( 
.A(n_1455),
.B(n_1092),
.Y(n_1602)
);

AOI21xp5_ASAP7_75t_L g1603 ( 
.A1(n_1421),
.A2(n_1120),
.B(n_1092),
.Y(n_1603)
);

AOI21xp5_ASAP7_75t_L g1604 ( 
.A1(n_1416),
.A2(n_1120),
.B(n_1092),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_SL g1605 ( 
.A(n_1443),
.B(n_797),
.Y(n_1605)
);

OAI21xp5_ASAP7_75t_L g1606 ( 
.A1(n_1427),
.A2(n_938),
.B(n_936),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1423),
.Y(n_1607)
);

NAND2xp33_ASAP7_75t_L g1608 ( 
.A(n_1456),
.B(n_1092),
.Y(n_1608)
);

INVx1_ASAP7_75t_SL g1609 ( 
.A(n_1486),
.Y(n_1609)
);

AOI33xp33_ASAP7_75t_L g1610 ( 
.A1(n_1563),
.A2(n_1570),
.A3(n_1556),
.B1(n_1441),
.B2(n_1491),
.B3(n_1541),
.Y(n_1610)
);

NOR2xp33_ASAP7_75t_L g1611 ( 
.A(n_1518),
.B(n_1527),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1448),
.B(n_1533),
.Y(n_1612)
);

INVx3_ASAP7_75t_L g1613 ( 
.A(n_1489),
.Y(n_1613)
);

BUFx4f_ASAP7_75t_L g1614 ( 
.A(n_1537),
.Y(n_1614)
);

OAI21xp33_ASAP7_75t_L g1615 ( 
.A1(n_1522),
.A2(n_764),
.B(n_763),
.Y(n_1615)
);

AOI21xp5_ASAP7_75t_L g1616 ( 
.A1(n_1587),
.A2(n_977),
.B(n_999),
.Y(n_1616)
);

NAND2xp5_ASAP7_75t_L g1617 ( 
.A(n_1499),
.B(n_767),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_SL g1618 ( 
.A(n_1512),
.B(n_766),
.Y(n_1618)
);

AOI21xp5_ASAP7_75t_L g1619 ( 
.A1(n_1557),
.A2(n_977),
.B(n_999),
.Y(n_1619)
);

O2A1O1Ixp5_ASAP7_75t_L g1620 ( 
.A1(n_1532),
.A2(n_1494),
.B(n_1482),
.C(n_1521),
.Y(n_1620)
);

AND2x4_ASAP7_75t_L g1621 ( 
.A(n_1458),
.B(n_939),
.Y(n_1621)
);

OAI22xp5_ASAP7_75t_L g1622 ( 
.A1(n_1465),
.A2(n_768),
.B1(n_779),
.B2(n_774),
.Y(n_1622)
);

O2A1O1Ixp5_ASAP7_75t_L g1623 ( 
.A1(n_1425),
.A2(n_787),
.B(n_788),
.C(n_785),
.Y(n_1623)
);

HB1xp67_ASAP7_75t_L g1624 ( 
.A(n_1505),
.Y(n_1624)
);

BUFx2_ASAP7_75t_L g1625 ( 
.A(n_1471),
.Y(n_1625)
);

INVx2_ASAP7_75t_L g1626 ( 
.A(n_1549),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1428),
.Y(n_1627)
);

A2O1A1Ixp33_ASAP7_75t_L g1628 ( 
.A1(n_1546),
.A2(n_1572),
.B(n_1535),
.C(n_1534),
.Y(n_1628)
);

NOR2xp33_ASAP7_75t_L g1629 ( 
.A(n_1564),
.B(n_1562),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_L g1630 ( 
.A(n_1417),
.B(n_789),
.Y(n_1630)
);

INVx2_ASAP7_75t_L g1631 ( 
.A(n_1550),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1433),
.Y(n_1632)
);

OR2x2_ASAP7_75t_L g1633 ( 
.A(n_1506),
.B(n_940),
.Y(n_1633)
);

BUFx4f_ASAP7_75t_L g1634 ( 
.A(n_1537),
.Y(n_1634)
);

NOR2xp33_ASAP7_75t_L g1635 ( 
.A(n_1540),
.B(n_770),
.Y(n_1635)
);

OAI21xp5_ASAP7_75t_L g1636 ( 
.A1(n_1427),
.A2(n_942),
.B(n_941),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1454),
.Y(n_1637)
);

INVxp33_ASAP7_75t_SL g1638 ( 
.A(n_1525),
.Y(n_1638)
);

AOI22xp5_ASAP7_75t_L g1639 ( 
.A1(n_1554),
.A2(n_777),
.B1(n_778),
.B2(n_776),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_L g1640 ( 
.A(n_1424),
.B(n_813),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_L g1641 ( 
.A(n_1434),
.B(n_819),
.Y(n_1641)
);

OAI21xp33_ASAP7_75t_SL g1642 ( 
.A1(n_1465),
.A2(n_825),
.B(n_820),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1459),
.Y(n_1643)
);

A2O1A1Ixp33_ASAP7_75t_L g1644 ( 
.A1(n_1483),
.A2(n_831),
.B(n_835),
.C(n_829),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_L g1645 ( 
.A(n_1414),
.B(n_836),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_SL g1646 ( 
.A(n_1431),
.B(n_780),
.Y(n_1646)
);

OAI21xp5_ASAP7_75t_L g1647 ( 
.A1(n_1437),
.A2(n_948),
.B(n_944),
.Y(n_1647)
);

BUFx2_ASAP7_75t_L g1648 ( 
.A(n_1450),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_SL g1649 ( 
.A(n_1466),
.B(n_782),
.Y(n_1649)
);

AOI21xp33_ASAP7_75t_L g1650 ( 
.A1(n_1422),
.A2(n_949),
.B(n_850),
.Y(n_1650)
);

AO21x2_ASAP7_75t_L g1651 ( 
.A1(n_1437),
.A2(n_953),
.B(n_952),
.Y(n_1651)
);

INVx4_ASAP7_75t_L g1652 ( 
.A(n_1498),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_L g1653 ( 
.A(n_1531),
.B(n_841),
.Y(n_1653)
);

INVx2_ASAP7_75t_L g1654 ( 
.A(n_1551),
.Y(n_1654)
);

BUFx6f_ASAP7_75t_L g1655 ( 
.A(n_1413),
.Y(n_1655)
);

INVx3_ASAP7_75t_L g1656 ( 
.A(n_1489),
.Y(n_1656)
);

INVx4_ASAP7_75t_L g1657 ( 
.A(n_1498),
.Y(n_1657)
);

INVx2_ASAP7_75t_L g1658 ( 
.A(n_1555),
.Y(n_1658)
);

NOR2xp33_ASAP7_75t_SL g1659 ( 
.A(n_1547),
.B(n_783),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_L g1660 ( 
.A(n_1422),
.B(n_845),
.Y(n_1660)
);

A2O1A1Ixp33_ASAP7_75t_L g1661 ( 
.A1(n_1483),
.A2(n_848),
.B(n_853),
.C(n_846),
.Y(n_1661)
);

NOR2xp33_ASAP7_75t_L g1662 ( 
.A(n_1556),
.B(n_784),
.Y(n_1662)
);

A2O1A1Ixp33_ASAP7_75t_L g1663 ( 
.A1(n_1578),
.A2(n_792),
.B(n_793),
.C(n_786),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_L g1664 ( 
.A(n_1548),
.B(n_794),
.Y(n_1664)
);

AND2x4_ASAP7_75t_SL g1665 ( 
.A(n_1547),
.B(n_956),
.Y(n_1665)
);

CKINVDCx10_ASAP7_75t_R g1666 ( 
.A(n_1435),
.Y(n_1666)
);

O2A1O1Ixp5_ASAP7_75t_L g1667 ( 
.A1(n_1446),
.A2(n_960),
.B(n_961),
.C(n_958),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_L g1668 ( 
.A(n_1552),
.B(n_795),
.Y(n_1668)
);

BUFx12f_ASAP7_75t_L g1669 ( 
.A(n_1524),
.Y(n_1669)
);

NOR2xp33_ASAP7_75t_L g1670 ( 
.A(n_1517),
.B(n_800),
.Y(n_1670)
);

BUFx3_ASAP7_75t_L g1671 ( 
.A(n_1478),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1553),
.B(n_802),
.Y(n_1672)
);

AOI22xp33_ASAP7_75t_L g1673 ( 
.A1(n_1513),
.A2(n_806),
.B1(n_807),
.B2(n_803),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_L g1674 ( 
.A(n_1501),
.B(n_808),
.Y(n_1674)
);

OAI21xp5_ASAP7_75t_L g1675 ( 
.A1(n_1440),
.A2(n_960),
.B(n_958),
.Y(n_1675)
);

BUFx12f_ASAP7_75t_L g1676 ( 
.A(n_1481),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1469),
.B(n_810),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_1473),
.B(n_812),
.Y(n_1678)
);

AND2x2_ASAP7_75t_L g1679 ( 
.A(n_1502),
.B(n_961),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_L g1680 ( 
.A(n_1544),
.B(n_815),
.Y(n_1680)
);

INVxp67_ASAP7_75t_L g1681 ( 
.A(n_1435),
.Y(n_1681)
);

AOI21xp5_ASAP7_75t_L g1682 ( 
.A1(n_1464),
.A2(n_1447),
.B(n_1445),
.Y(n_1682)
);

AOI21xp5_ASAP7_75t_L g1683 ( 
.A1(n_1451),
.A2(n_1453),
.B(n_1457),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_SL g1684 ( 
.A(n_1493),
.B(n_822),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_L g1685 ( 
.A(n_1468),
.B(n_824),
.Y(n_1685)
);

AOI21xp33_ASAP7_75t_L g1686 ( 
.A1(n_1440),
.A2(n_962),
.B(n_827),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_L g1687 ( 
.A(n_1480),
.B(n_826),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_L g1688 ( 
.A(n_1484),
.B(n_828),
.Y(n_1688)
);

AOI22xp5_ASAP7_75t_L g1689 ( 
.A1(n_1525),
.A2(n_838),
.B1(n_839),
.B2(n_837),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1488),
.B(n_840),
.Y(n_1690)
);

INVx2_ASAP7_75t_L g1691 ( 
.A(n_1559),
.Y(n_1691)
);

INVxp67_ASAP7_75t_L g1692 ( 
.A(n_1565),
.Y(n_1692)
);

AOI22xp33_ASAP7_75t_L g1693 ( 
.A1(n_1568),
.A2(n_844),
.B1(n_851),
.B2(n_842),
.Y(n_1693)
);

AOI21xp5_ASAP7_75t_L g1694 ( 
.A1(n_1460),
.A2(n_1024),
.B(n_1010),
.Y(n_1694)
);

OAI321xp33_ASAP7_75t_L g1695 ( 
.A1(n_1526),
.A2(n_857),
.A3(n_854),
.B1(n_865),
.B2(n_855),
.C(n_852),
.Y(n_1695)
);

AND2x2_ASAP7_75t_L g1696 ( 
.A(n_1463),
.B(n_1504),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_L g1697 ( 
.A(n_1490),
.B(n_1),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1573),
.Y(n_1698)
);

AOI21xp5_ASAP7_75t_L g1699 ( 
.A1(n_1461),
.A2(n_1024),
.B(n_1096),
.Y(n_1699)
);

AND2x2_ASAP7_75t_L g1700 ( 
.A(n_1463),
.B(n_2),
.Y(n_1700)
);

OAI21xp5_ASAP7_75t_L g1701 ( 
.A1(n_1442),
.A2(n_981),
.B(n_1024),
.Y(n_1701)
);

OAI21xp5_ASAP7_75t_L g1702 ( 
.A1(n_1442),
.A2(n_981),
.B(n_1024),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_L g1703 ( 
.A(n_1492),
.B(n_4),
.Y(n_1703)
);

INVx2_ASAP7_75t_SL g1704 ( 
.A(n_1508),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_L g1705 ( 
.A(n_1495),
.B(n_6),
.Y(n_1705)
);

NAND2xp5_ASAP7_75t_L g1706 ( 
.A(n_1497),
.B(n_1543),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_SL g1707 ( 
.A(n_1500),
.B(n_1024),
.Y(n_1707)
);

CKINVDCx5p33_ASAP7_75t_R g1708 ( 
.A(n_1558),
.Y(n_1708)
);

NAND2x1p5_ASAP7_75t_L g1709 ( 
.A(n_1413),
.B(n_1024),
.Y(n_1709)
);

NAND2xp5_ASAP7_75t_L g1710 ( 
.A(n_1545),
.B(n_7),
.Y(n_1710)
);

A2O1A1Ixp33_ASAP7_75t_L g1711 ( 
.A1(n_1569),
.A2(n_9),
.B(n_7),
.C(n_8),
.Y(n_1711)
);

NAND2xp5_ASAP7_75t_L g1712 ( 
.A(n_1566),
.B(n_8),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_L g1713 ( 
.A(n_1567),
.B(n_9),
.Y(n_1713)
);

AOI22xp33_ASAP7_75t_L g1714 ( 
.A1(n_1507),
.A2(n_981),
.B1(n_990),
.B2(n_12),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_1574),
.B(n_10),
.Y(n_1715)
);

INVx2_ASAP7_75t_L g1716 ( 
.A(n_1560),
.Y(n_1716)
);

BUFx6f_ASAP7_75t_L g1717 ( 
.A(n_1439),
.Y(n_1717)
);

BUFx12f_ASAP7_75t_L g1718 ( 
.A(n_1571),
.Y(n_1718)
);

CKINVDCx5p33_ASAP7_75t_R g1719 ( 
.A(n_1577),
.Y(n_1719)
);

NOR3xp33_ASAP7_75t_L g1720 ( 
.A(n_1586),
.B(n_1523),
.C(n_1516),
.Y(n_1720)
);

AOI21xp5_ASAP7_75t_L g1721 ( 
.A1(n_1429),
.A2(n_1096),
.B(n_990),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_L g1722 ( 
.A(n_1579),
.B(n_11),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1581),
.Y(n_1723)
);

INVx2_ASAP7_75t_L g1724 ( 
.A(n_1561),
.Y(n_1724)
);

HB1xp67_ASAP7_75t_L g1725 ( 
.A(n_1514),
.Y(n_1725)
);

AOI22xp5_ASAP7_75t_L g1726 ( 
.A1(n_1519),
.A2(n_990),
.B1(n_1096),
.B2(n_14),
.Y(n_1726)
);

HB1xp67_ASAP7_75t_L g1727 ( 
.A(n_1571),
.Y(n_1727)
);

NOR2xp33_ASAP7_75t_L g1728 ( 
.A(n_1528),
.B(n_11),
.Y(n_1728)
);

NOR2xp33_ASAP7_75t_L g1729 ( 
.A(n_1529),
.B(n_1530),
.Y(n_1729)
);

AOI21xp33_ASAP7_75t_L g1730 ( 
.A1(n_1585),
.A2(n_13),
.B(n_14),
.Y(n_1730)
);

O2A1O1Ixp33_ASAP7_75t_L g1731 ( 
.A1(n_1585),
.A2(n_17),
.B(n_15),
.C(n_16),
.Y(n_1731)
);

O2A1O1Ixp33_ASAP7_75t_SL g1732 ( 
.A1(n_1462),
.A2(n_576),
.B(n_577),
.C(n_573),
.Y(n_1732)
);

OAI21xp5_ASAP7_75t_L g1733 ( 
.A1(n_1590),
.A2(n_1430),
.B(n_1467),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1582),
.Y(n_1734)
);

NAND2xp5_ASAP7_75t_L g1735 ( 
.A(n_1530),
.B(n_16),
.Y(n_1735)
);

NAND2xp5_ASAP7_75t_L g1736 ( 
.A(n_1511),
.B(n_18),
.Y(n_1736)
);

CKINVDCx5p33_ASAP7_75t_R g1737 ( 
.A(n_1508),
.Y(n_1737)
);

AOI21xp5_ASAP7_75t_L g1738 ( 
.A1(n_1590),
.A2(n_990),
.B(n_582),
.Y(n_1738)
);

INVx2_ASAP7_75t_L g1739 ( 
.A(n_1515),
.Y(n_1739)
);

OAI21xp5_ASAP7_75t_L g1740 ( 
.A1(n_1419),
.A2(n_583),
.B(n_579),
.Y(n_1740)
);

NAND2xp5_ASAP7_75t_L g1741 ( 
.A(n_1479),
.B(n_18),
.Y(n_1741)
);

NAND2xp5_ASAP7_75t_L g1742 ( 
.A(n_1485),
.B(n_19),
.Y(n_1742)
);

AOI21xp33_ASAP7_75t_L g1743 ( 
.A1(n_1487),
.A2(n_19),
.B(n_20),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_SL g1744 ( 
.A(n_1576),
.B(n_20),
.Y(n_1744)
);

CKINVDCx5p33_ASAP7_75t_R g1745 ( 
.A(n_1508),
.Y(n_1745)
);

AOI21x1_ASAP7_75t_L g1746 ( 
.A1(n_1496),
.A2(n_585),
.B(n_584),
.Y(n_1746)
);

NAND2x1p5_ASAP7_75t_L g1747 ( 
.A(n_1439),
.B(n_586),
.Y(n_1747)
);

AND2x2_ASAP7_75t_SL g1748 ( 
.A(n_1536),
.B(n_21),
.Y(n_1748)
);

HB1xp67_ASAP7_75t_L g1749 ( 
.A(n_1571),
.Y(n_1749)
);

AOI21xp5_ASAP7_75t_L g1750 ( 
.A1(n_1418),
.A2(n_1539),
.B(n_1538),
.Y(n_1750)
);

NAND2xp5_ASAP7_75t_L g1751 ( 
.A(n_1542),
.B(n_22),
.Y(n_1751)
);

AND2x2_ASAP7_75t_L g1752 ( 
.A(n_1420),
.B(n_22),
.Y(n_1752)
);

AOI22xp33_ASAP7_75t_L g1753 ( 
.A1(n_1476),
.A2(n_25),
.B1(n_23),
.B2(n_24),
.Y(n_1753)
);

O2A1O1Ixp33_ASAP7_75t_L g1754 ( 
.A1(n_1589),
.A2(n_25),
.B(n_23),
.C(n_24),
.Y(n_1754)
);

AOI21x1_ASAP7_75t_L g1755 ( 
.A1(n_1583),
.A2(n_588),
.B(n_587),
.Y(n_1755)
);

NAND2xp5_ASAP7_75t_L g1756 ( 
.A(n_1584),
.B(n_1588),
.Y(n_1756)
);

NAND2xp5_ASAP7_75t_L g1757 ( 
.A(n_1436),
.B(n_26),
.Y(n_1757)
);

NOR2xp33_ASAP7_75t_SL g1758 ( 
.A(n_1600),
.B(n_1458),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1607),
.Y(n_1759)
);

NAND2xp5_ASAP7_75t_L g1760 ( 
.A(n_1611),
.B(n_1444),
.Y(n_1760)
);

NAND2xp5_ASAP7_75t_L g1761 ( 
.A(n_1729),
.B(n_1449),
.Y(n_1761)
);

AOI21xp5_ASAP7_75t_L g1762 ( 
.A1(n_1608),
.A2(n_1418),
.B(n_1458),
.Y(n_1762)
);

BUFx12f_ASAP7_75t_L g1763 ( 
.A(n_1708),
.Y(n_1763)
);

NAND2xp5_ASAP7_75t_L g1764 ( 
.A(n_1706),
.B(n_1452),
.Y(n_1764)
);

OAI21xp5_ASAP7_75t_L g1765 ( 
.A1(n_1620),
.A2(n_1575),
.B(n_1476),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_SL g1766 ( 
.A(n_1629),
.B(n_1456),
.Y(n_1766)
);

OAI22x1_ASAP7_75t_L g1767 ( 
.A1(n_1599),
.A2(n_1472),
.B1(n_1503),
.B2(n_1475),
.Y(n_1767)
);

OAI22xp5_ASAP7_75t_L g1768 ( 
.A1(n_1628),
.A2(n_1510),
.B1(n_1580),
.B2(n_1474),
.Y(n_1768)
);

NOR2xp33_ASAP7_75t_L g1769 ( 
.A(n_1638),
.B(n_1580),
.Y(n_1769)
);

NAND2x1p5_ASAP7_75t_L g1770 ( 
.A(n_1600),
.B(n_1474),
.Y(n_1770)
);

NAND2xp5_ASAP7_75t_SL g1771 ( 
.A(n_1610),
.B(n_1456),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1627),
.Y(n_1772)
);

OAI22xp5_ASAP7_75t_L g1773 ( 
.A1(n_1612),
.A2(n_1456),
.B1(n_1575),
.B2(n_1476),
.Y(n_1773)
);

AOI21xp5_ASAP7_75t_L g1774 ( 
.A1(n_1592),
.A2(n_1456),
.B(n_1575),
.Y(n_1774)
);

A2O1A1Ixp33_ASAP7_75t_L g1775 ( 
.A1(n_1728),
.A2(n_1575),
.B(n_1476),
.C(n_28),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1632),
.Y(n_1776)
);

NOR2xp33_ASAP7_75t_L g1777 ( 
.A(n_1594),
.B(n_590),
.Y(n_1777)
);

A2O1A1Ixp33_ASAP7_75t_L g1778 ( 
.A1(n_1617),
.A2(n_28),
.B(n_26),
.C(n_27),
.Y(n_1778)
);

INVxp67_ASAP7_75t_L g1779 ( 
.A(n_1593),
.Y(n_1779)
);

NAND2xp5_ASAP7_75t_L g1780 ( 
.A(n_1696),
.B(n_27),
.Y(n_1780)
);

OR2x4_ASAP7_75t_L g1781 ( 
.A(n_1662),
.B(n_29),
.Y(n_1781)
);

AOI22xp33_ASAP7_75t_L g1782 ( 
.A1(n_1735),
.A2(n_31),
.B1(n_29),
.B2(n_30),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_SL g1783 ( 
.A(n_1720),
.B(n_30),
.Y(n_1783)
);

OR2x2_ASAP7_75t_L g1784 ( 
.A(n_1648),
.B(n_31),
.Y(n_1784)
);

OAI22x1_ASAP7_75t_L g1785 ( 
.A1(n_1605),
.A2(n_1700),
.B1(n_1591),
.B2(n_1660),
.Y(n_1785)
);

NOR2xp33_ASAP7_75t_L g1786 ( 
.A(n_1618),
.B(n_592),
.Y(n_1786)
);

NAND2xp5_ASAP7_75t_SL g1787 ( 
.A(n_1748),
.B(n_33),
.Y(n_1787)
);

NAND2xp5_ASAP7_75t_L g1788 ( 
.A(n_1597),
.B(n_35),
.Y(n_1788)
);

OAI22xp5_ASAP7_75t_L g1789 ( 
.A1(n_1624),
.A2(n_38),
.B1(n_36),
.B2(n_37),
.Y(n_1789)
);

INVx3_ASAP7_75t_L g1790 ( 
.A(n_1601),
.Y(n_1790)
);

NAND2xp5_ASAP7_75t_L g1791 ( 
.A(n_1633),
.B(n_37),
.Y(n_1791)
);

AO21x1_ASAP7_75t_L g1792 ( 
.A1(n_1740),
.A2(n_39),
.B(n_40),
.Y(n_1792)
);

NAND2xp5_ASAP7_75t_L g1793 ( 
.A(n_1630),
.B(n_41),
.Y(n_1793)
);

NAND2xp5_ASAP7_75t_L g1794 ( 
.A(n_1640),
.B(n_41),
.Y(n_1794)
);

NOR2xp33_ASAP7_75t_L g1795 ( 
.A(n_1670),
.B(n_594),
.Y(n_1795)
);

AOI21xp5_ASAP7_75t_L g1796 ( 
.A1(n_1598),
.A2(n_633),
.B(n_631),
.Y(n_1796)
);

NAND2xp5_ASAP7_75t_SL g1797 ( 
.A(n_1635),
.B(n_42),
.Y(n_1797)
);

OAI22xp5_ASAP7_75t_L g1798 ( 
.A1(n_1674),
.A2(n_1685),
.B1(n_1688),
.B2(n_1687),
.Y(n_1798)
);

AOI21xp5_ASAP7_75t_L g1799 ( 
.A1(n_1707),
.A2(n_612),
.B(n_611),
.Y(n_1799)
);

AOI22xp5_ASAP7_75t_L g1800 ( 
.A1(n_1642),
.A2(n_45),
.B1(n_43),
.B2(n_44),
.Y(n_1800)
);

OAI22xp5_ASAP7_75t_L g1801 ( 
.A1(n_1690),
.A2(n_48),
.B1(n_45),
.B2(n_47),
.Y(n_1801)
);

NAND2xp5_ASAP7_75t_SL g1802 ( 
.A(n_1621),
.B(n_47),
.Y(n_1802)
);

INVxp67_ASAP7_75t_L g1803 ( 
.A(n_1625),
.Y(n_1803)
);

INVx2_ASAP7_75t_L g1804 ( 
.A(n_1626),
.Y(n_1804)
);

AO32x1_ASAP7_75t_L g1805 ( 
.A1(n_1595),
.A2(n_51),
.A3(n_49),
.B1(n_50),
.B2(n_52),
.Y(n_1805)
);

NAND2xp5_ASAP7_75t_SL g1806 ( 
.A(n_1621),
.B(n_49),
.Y(n_1806)
);

CKINVDCx8_ASAP7_75t_R g1807 ( 
.A(n_1666),
.Y(n_1807)
);

NAND2xp5_ASAP7_75t_L g1808 ( 
.A(n_1641),
.B(n_50),
.Y(n_1808)
);

AOI22xp5_ASAP7_75t_L g1809 ( 
.A1(n_1615),
.A2(n_54),
.B1(n_51),
.B2(n_53),
.Y(n_1809)
);

OR2x2_ASAP7_75t_L g1810 ( 
.A(n_1645),
.B(n_53),
.Y(n_1810)
);

NAND2xp5_ASAP7_75t_L g1811 ( 
.A(n_1664),
.B(n_54),
.Y(n_1811)
);

NAND2xp5_ASAP7_75t_L g1812 ( 
.A(n_1697),
.B(n_55),
.Y(n_1812)
);

O2A1O1Ixp33_ASAP7_75t_L g1813 ( 
.A1(n_1711),
.A2(n_57),
.B(n_55),
.C(n_56),
.Y(n_1813)
);

NAND2xp5_ASAP7_75t_L g1814 ( 
.A(n_1703),
.B(n_56),
.Y(n_1814)
);

O2A1O1Ixp33_ASAP7_75t_L g1815 ( 
.A1(n_1650),
.A2(n_60),
.B(n_58),
.C(n_59),
.Y(n_1815)
);

OAI21xp5_ASAP7_75t_L g1816 ( 
.A1(n_1668),
.A2(n_1672),
.B(n_1682),
.Y(n_1816)
);

BUFx6f_ASAP7_75t_L g1817 ( 
.A(n_1614),
.Y(n_1817)
);

NAND2xp5_ASAP7_75t_L g1818 ( 
.A(n_1705),
.B(n_58),
.Y(n_1818)
);

AOI21xp5_ASAP7_75t_L g1819 ( 
.A1(n_1595),
.A2(n_615),
.B(n_614),
.Y(n_1819)
);

NAND2xp5_ASAP7_75t_L g1820 ( 
.A(n_1710),
.B(n_62),
.Y(n_1820)
);

BUFx6f_ASAP7_75t_SL g1821 ( 
.A(n_1671),
.Y(n_1821)
);

INVx3_ASAP7_75t_L g1822 ( 
.A(n_1601),
.Y(n_1822)
);

NAND2xp5_ASAP7_75t_L g1823 ( 
.A(n_1653),
.B(n_63),
.Y(n_1823)
);

BUFx8_ASAP7_75t_L g1824 ( 
.A(n_1718),
.Y(n_1824)
);

NAND2xp5_ASAP7_75t_L g1825 ( 
.A(n_1712),
.B(n_64),
.Y(n_1825)
);

AOI21xp5_ASAP7_75t_L g1826 ( 
.A1(n_1683),
.A2(n_625),
.B(n_624),
.Y(n_1826)
);

NOR2xp33_ASAP7_75t_L g1827 ( 
.A(n_1609),
.B(n_596),
.Y(n_1827)
);

AOI21xp5_ASAP7_75t_L g1828 ( 
.A1(n_1750),
.A2(n_598),
.B(n_597),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1637),
.Y(n_1829)
);

NOR2xp33_ASAP7_75t_L g1830 ( 
.A(n_1692),
.B(n_599),
.Y(n_1830)
);

NOR2xp33_ASAP7_75t_L g1831 ( 
.A(n_1719),
.B(n_601),
.Y(n_1831)
);

NAND2xp5_ASAP7_75t_L g1832 ( 
.A(n_1713),
.B(n_65),
.Y(n_1832)
);

AND2x2_ASAP7_75t_L g1833 ( 
.A(n_1679),
.B(n_67),
.Y(n_1833)
);

AND2x2_ASAP7_75t_L g1834 ( 
.A(n_1752),
.B(n_68),
.Y(n_1834)
);

AOI21xp5_ASAP7_75t_L g1835 ( 
.A1(n_1602),
.A2(n_630),
.B(n_604),
.Y(n_1835)
);

NAND2xp5_ASAP7_75t_L g1836 ( 
.A(n_1715),
.B(n_68),
.Y(n_1836)
);

NOR2xp33_ASAP7_75t_L g1837 ( 
.A(n_1649),
.B(n_603),
.Y(n_1837)
);

NOR2xp33_ASAP7_75t_L g1838 ( 
.A(n_1722),
.B(n_606),
.Y(n_1838)
);

NAND2xp5_ASAP7_75t_SL g1839 ( 
.A(n_1695),
.B(n_69),
.Y(n_1839)
);

AOI221xp5_ASAP7_75t_L g1840 ( 
.A1(n_1650),
.A2(n_1730),
.B1(n_1622),
.B2(n_1673),
.C(n_1693),
.Y(n_1840)
);

INVx2_ASAP7_75t_L g1841 ( 
.A(n_1631),
.Y(n_1841)
);

OAI22xp33_ASAP7_75t_L g1842 ( 
.A1(n_1659),
.A2(n_71),
.B1(n_69),
.B2(n_70),
.Y(n_1842)
);

INVx4_ASAP7_75t_L g1843 ( 
.A(n_1614),
.Y(n_1843)
);

O2A1O1Ixp33_ASAP7_75t_L g1844 ( 
.A1(n_1730),
.A2(n_72),
.B(n_70),
.C(n_71),
.Y(n_1844)
);

OAI21xp5_ASAP7_75t_L g1845 ( 
.A1(n_1623),
.A2(n_73),
.B(n_75),
.Y(n_1845)
);

AOI22x1_ASAP7_75t_L g1846 ( 
.A1(n_1606),
.A2(n_76),
.B1(n_73),
.B2(n_75),
.Y(n_1846)
);

NAND2xp5_ASAP7_75t_L g1847 ( 
.A(n_1756),
.B(n_77),
.Y(n_1847)
);

NAND2xp5_ASAP7_75t_SL g1848 ( 
.A(n_1634),
.B(n_77),
.Y(n_1848)
);

INVx5_ASAP7_75t_L g1849 ( 
.A(n_1655),
.Y(n_1849)
);

NOR2xp33_ASAP7_75t_L g1850 ( 
.A(n_1689),
.B(n_607),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1643),
.Y(n_1851)
);

NOR2x1p5_ASAP7_75t_L g1852 ( 
.A(n_1669),
.B(n_608),
.Y(n_1852)
);

INVx2_ASAP7_75t_L g1853 ( 
.A(n_1654),
.Y(n_1853)
);

O2A1O1Ixp33_ASAP7_75t_L g1854 ( 
.A1(n_1744),
.A2(n_81),
.B(n_78),
.C(n_80),
.Y(n_1854)
);

CKINVDCx20_ASAP7_75t_R g1855 ( 
.A(n_1737),
.Y(n_1855)
);

NAND2xp5_ASAP7_75t_L g1856 ( 
.A(n_1596),
.B(n_80),
.Y(n_1856)
);

NOR2xp33_ASAP7_75t_R g1857 ( 
.A(n_1745),
.B(n_616),
.Y(n_1857)
);

AOI21xp5_ASAP7_75t_L g1858 ( 
.A1(n_1602),
.A2(n_623),
.B(n_619),
.Y(n_1858)
);

O2A1O1Ixp33_ASAP7_75t_L g1859 ( 
.A1(n_1663),
.A2(n_83),
.B(n_81),
.C(n_82),
.Y(n_1859)
);

BUFx2_ASAP7_75t_SL g1860 ( 
.A(n_1652),
.Y(n_1860)
);

O2A1O1Ixp33_ASAP7_75t_SL g1861 ( 
.A1(n_1740),
.A2(n_1684),
.B(n_1661),
.C(n_1644),
.Y(n_1861)
);

NAND2xp5_ASAP7_75t_L g1862 ( 
.A(n_1658),
.B(n_82),
.Y(n_1862)
);

NAND2xp5_ASAP7_75t_SL g1863 ( 
.A(n_1634),
.B(n_83),
.Y(n_1863)
);

NOR2xp33_ASAP7_75t_L g1864 ( 
.A(n_1646),
.B(n_618),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1698),
.Y(n_1865)
);

OA22x2_ASAP7_75t_L g1866 ( 
.A1(n_1639),
.A2(n_86),
.B1(n_84),
.B2(n_85),
.Y(n_1866)
);

OAI321xp33_ASAP7_75t_L g1867 ( 
.A1(n_1753),
.A2(n_87),
.A3(n_89),
.B1(n_84),
.B2(n_85),
.C(n_88),
.Y(n_1867)
);

NOR2xp33_ASAP7_75t_L g1868 ( 
.A(n_1727),
.B(n_620),
.Y(n_1868)
);

OAI22xp5_ASAP7_75t_L g1869 ( 
.A1(n_1704),
.A2(n_90),
.B1(n_88),
.B2(n_89),
.Y(n_1869)
);

NOR2xp33_ASAP7_75t_L g1870 ( 
.A(n_1749),
.B(n_1676),
.Y(n_1870)
);

AOI21xp5_ASAP7_75t_L g1871 ( 
.A1(n_1651),
.A2(n_621),
.B(n_90),
.Y(n_1871)
);

NAND2x1p5_ASAP7_75t_L g1872 ( 
.A(n_1652),
.B(n_91),
.Y(n_1872)
);

AND2x2_ASAP7_75t_L g1873 ( 
.A(n_1691),
.B(n_92),
.Y(n_1873)
);

AOI22xp5_ASAP7_75t_L g1874 ( 
.A1(n_1622),
.A2(n_94),
.B1(n_92),
.B2(n_93),
.Y(n_1874)
);

AOI21xp5_ASAP7_75t_L g1875 ( 
.A1(n_1651),
.A2(n_93),
.B(n_94),
.Y(n_1875)
);

AO22x1_ASAP7_75t_L g1876 ( 
.A1(n_1681),
.A2(n_97),
.B1(n_95),
.B2(n_96),
.Y(n_1876)
);

AOI21xp5_ASAP7_75t_L g1877 ( 
.A1(n_1603),
.A2(n_95),
.B(n_96),
.Y(n_1877)
);

BUFx6f_ASAP7_75t_L g1878 ( 
.A(n_1655),
.Y(n_1878)
);

AOI21x1_ASAP7_75t_L g1879 ( 
.A1(n_1604),
.A2(n_97),
.B(n_98),
.Y(n_1879)
);

AOI21xp5_ASAP7_75t_L g1880 ( 
.A1(n_1701),
.A2(n_570),
.B(n_98),
.Y(n_1880)
);

OAI22xp5_ASAP7_75t_L g1881 ( 
.A1(n_1723),
.A2(n_101),
.B1(n_99),
.B2(n_100),
.Y(n_1881)
);

OAI321xp33_ASAP7_75t_L g1882 ( 
.A1(n_1731),
.A2(n_103),
.A3(n_105),
.B1(n_100),
.B2(n_102),
.C(n_104),
.Y(n_1882)
);

AO32x1_ASAP7_75t_L g1883 ( 
.A1(n_1734),
.A2(n_107),
.A3(n_104),
.B1(n_105),
.B2(n_108),
.Y(n_1883)
);

NAND2xp5_ASAP7_75t_L g1884 ( 
.A(n_1716),
.B(n_107),
.Y(n_1884)
);

NAND2xp5_ASAP7_75t_L g1885 ( 
.A(n_1724),
.B(n_108),
.Y(n_1885)
);

NAND2xp5_ASAP7_75t_L g1886 ( 
.A(n_1739),
.B(n_109),
.Y(n_1886)
);

AOI21xp5_ASAP7_75t_L g1887 ( 
.A1(n_1701),
.A2(n_111),
.B(n_112),
.Y(n_1887)
);

NAND2xp5_ASAP7_75t_L g1888 ( 
.A(n_1677),
.B(n_111),
.Y(n_1888)
);

INVx1_ASAP7_75t_SL g1889 ( 
.A(n_1725),
.Y(n_1889)
);

OAI22xp5_ASAP7_75t_L g1890 ( 
.A1(n_1677),
.A2(n_114),
.B1(n_112),
.B2(n_113),
.Y(n_1890)
);

NAND2xp5_ASAP7_75t_L g1891 ( 
.A(n_1678),
.B(n_113),
.Y(n_1891)
);

NOR2xp33_ASAP7_75t_L g1892 ( 
.A(n_1665),
.B(n_114),
.Y(n_1892)
);

AND2x2_ASAP7_75t_L g1893 ( 
.A(n_1680),
.B(n_115),
.Y(n_1893)
);

OAI21xp5_ASAP7_75t_L g1894 ( 
.A1(n_1647),
.A2(n_116),
.B(n_117),
.Y(n_1894)
);

AOI21xp5_ASAP7_75t_L g1895 ( 
.A1(n_1702),
.A2(n_570),
.B(n_118),
.Y(n_1895)
);

BUFx12f_ASAP7_75t_L g1896 ( 
.A(n_1657),
.Y(n_1896)
);

AOI21xp5_ASAP7_75t_L g1897 ( 
.A1(n_1702),
.A2(n_569),
.B(n_119),
.Y(n_1897)
);

O2A1O1Ixp5_ASAP7_75t_SL g1898 ( 
.A1(n_1686),
.A2(n_122),
.B(n_120),
.C(n_121),
.Y(n_1898)
);

NAND2xp5_ASAP7_75t_SL g1899 ( 
.A(n_1741),
.B(n_122),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1757),
.Y(n_1900)
);

AOI21xp5_ASAP7_75t_L g1901 ( 
.A1(n_1733),
.A2(n_569),
.B(n_124),
.Y(n_1901)
);

NOR2xp33_ASAP7_75t_L g1902 ( 
.A(n_1742),
.B(n_125),
.Y(n_1902)
);

AOI21xp5_ASAP7_75t_L g1903 ( 
.A1(n_1738),
.A2(n_1647),
.B(n_1636),
.Y(n_1903)
);

OAI22xp5_ASAP7_75t_L g1904 ( 
.A1(n_1751),
.A2(n_128),
.B1(n_126),
.B2(n_127),
.Y(n_1904)
);

OAI22xp5_ASAP7_75t_L g1905 ( 
.A1(n_1736),
.A2(n_129),
.B1(n_126),
.B2(n_128),
.Y(n_1905)
);

NAND2xp5_ASAP7_75t_L g1906 ( 
.A(n_1636),
.B(n_130),
.Y(n_1906)
);

NAND2xp5_ASAP7_75t_L g1907 ( 
.A(n_1686),
.B(n_130),
.Y(n_1907)
);

OAI21xp33_ASAP7_75t_L g1908 ( 
.A1(n_1743),
.A2(n_131),
.B(n_132),
.Y(n_1908)
);

INVx1_ASAP7_75t_L g1909 ( 
.A(n_1667),
.Y(n_1909)
);

INVx2_ASAP7_75t_SL g1910 ( 
.A(n_1655),
.Y(n_1910)
);

NOR2xp67_ASAP7_75t_SL g1911 ( 
.A(n_1657),
.B(n_133),
.Y(n_1911)
);

NAND2xp5_ASAP7_75t_L g1912 ( 
.A(n_1675),
.B(n_133),
.Y(n_1912)
);

NAND2xp5_ASAP7_75t_L g1913 ( 
.A(n_1613),
.B(n_134),
.Y(n_1913)
);

OAI21xp5_ASAP7_75t_L g1914 ( 
.A1(n_1726),
.A2(n_134),
.B(n_136),
.Y(n_1914)
);

AOI22xp5_ASAP7_75t_L g1915 ( 
.A1(n_1840),
.A2(n_1743),
.B1(n_1714),
.B2(n_1747),
.Y(n_1915)
);

NAND2x1p5_ASAP7_75t_L g1916 ( 
.A(n_1849),
.B(n_1613),
.Y(n_1916)
);

CKINVDCx20_ASAP7_75t_R g1917 ( 
.A(n_1855),
.Y(n_1917)
);

AND2x2_ASAP7_75t_L g1918 ( 
.A(n_1834),
.B(n_1747),
.Y(n_1918)
);

OAI21x1_ASAP7_75t_L g1919 ( 
.A1(n_1774),
.A2(n_1755),
.B(n_1746),
.Y(n_1919)
);

NAND2xp5_ASAP7_75t_L g1920 ( 
.A(n_1761),
.B(n_1754),
.Y(n_1920)
);

NAND2xp5_ASAP7_75t_L g1921 ( 
.A(n_1764),
.B(n_1656),
.Y(n_1921)
);

AND2x4_ASAP7_75t_L g1922 ( 
.A(n_1843),
.B(n_1889),
.Y(n_1922)
);

AOI21xp5_ASAP7_75t_L g1923 ( 
.A1(n_1903),
.A2(n_1619),
.B(n_1732),
.Y(n_1923)
);

NAND2x1p5_ASAP7_75t_L g1924 ( 
.A(n_1849),
.B(n_1717),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1759),
.Y(n_1925)
);

AND2x2_ASAP7_75t_L g1926 ( 
.A(n_1833),
.B(n_1717),
.Y(n_1926)
);

NAND2x1_ASAP7_75t_L g1927 ( 
.A(n_1762),
.B(n_1717),
.Y(n_1927)
);

AOI21xp5_ASAP7_75t_L g1928 ( 
.A1(n_1816),
.A2(n_1616),
.B(n_1699),
.Y(n_1928)
);

AND2x2_ASAP7_75t_L g1929 ( 
.A(n_1780),
.B(n_136),
.Y(n_1929)
);

OAI21xp33_ASAP7_75t_L g1930 ( 
.A1(n_1894),
.A2(n_1721),
.B(n_1694),
.Y(n_1930)
);

BUFx6f_ASAP7_75t_L g1931 ( 
.A(n_1817),
.Y(n_1931)
);

AND2x2_ASAP7_75t_L g1932 ( 
.A(n_1873),
.B(n_137),
.Y(n_1932)
);

OAI21xp5_ASAP7_75t_L g1933 ( 
.A1(n_1880),
.A2(n_1709),
.B(n_138),
.Y(n_1933)
);

AO22x2_ASAP7_75t_L g1934 ( 
.A1(n_1887),
.A2(n_140),
.B1(n_138),
.B2(n_139),
.Y(n_1934)
);

O2A1O1Ixp5_ASAP7_75t_L g1935 ( 
.A1(n_1792),
.A2(n_1709),
.B(n_143),
.C(n_141),
.Y(n_1935)
);

OAI21xp5_ASAP7_75t_L g1936 ( 
.A1(n_1895),
.A2(n_142),
.B(n_143),
.Y(n_1936)
);

AOI21xp5_ASAP7_75t_L g1937 ( 
.A1(n_1819),
.A2(n_142),
.B(n_144),
.Y(n_1937)
);

INVx5_ASAP7_75t_L g1938 ( 
.A(n_1817),
.Y(n_1938)
);

AOI21xp5_ASAP7_75t_L g1939 ( 
.A1(n_1765),
.A2(n_145),
.B(n_146),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1772),
.Y(n_1940)
);

OAI21x1_ASAP7_75t_L g1941 ( 
.A1(n_1826),
.A2(n_146),
.B(n_147),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1776),
.Y(n_1942)
);

OAI21xp5_ASAP7_75t_L g1943 ( 
.A1(n_1897),
.A2(n_147),
.B(n_148),
.Y(n_1943)
);

NAND2xp5_ASAP7_75t_L g1944 ( 
.A(n_1900),
.B(n_568),
.Y(n_1944)
);

NAND2xp33_ASAP7_75t_SL g1945 ( 
.A(n_1817),
.B(n_1857),
.Y(n_1945)
);

NOR2xp33_ASAP7_75t_L g1946 ( 
.A(n_1798),
.B(n_149),
.Y(n_1946)
);

OAI21x1_ASAP7_75t_L g1947 ( 
.A1(n_1879),
.A2(n_150),
.B(n_151),
.Y(n_1947)
);

OAI21x1_ASAP7_75t_L g1948 ( 
.A1(n_1796),
.A2(n_152),
.B(n_153),
.Y(n_1948)
);

INVx1_ASAP7_75t_SL g1949 ( 
.A(n_1766),
.Y(n_1949)
);

A2O1A1Ixp33_ASAP7_75t_L g1950 ( 
.A1(n_1850),
.A2(n_154),
.B(n_152),
.C(n_153),
.Y(n_1950)
);

AOI21xp5_ASAP7_75t_L g1951 ( 
.A1(n_1861),
.A2(n_155),
.B(n_156),
.Y(n_1951)
);

AO31x2_ASAP7_75t_L g1952 ( 
.A1(n_1773),
.A2(n_157),
.A3(n_155),
.B(n_156),
.Y(n_1952)
);

CKINVDCx5p33_ASAP7_75t_R g1953 ( 
.A(n_1807),
.Y(n_1953)
);

NAND2xp5_ASAP7_75t_L g1954 ( 
.A(n_1907),
.B(n_157),
.Y(n_1954)
);

OAI21x1_ASAP7_75t_L g1955 ( 
.A1(n_1828),
.A2(n_158),
.B(n_159),
.Y(n_1955)
);

NAND2xp5_ASAP7_75t_L g1956 ( 
.A(n_1847),
.B(n_158),
.Y(n_1956)
);

INVx1_ASAP7_75t_L g1957 ( 
.A(n_1829),
.Y(n_1957)
);

INVx1_ASAP7_75t_SL g1958 ( 
.A(n_1760),
.Y(n_1958)
);

OAI21x1_ASAP7_75t_L g1959 ( 
.A1(n_1871),
.A2(n_160),
.B(n_161),
.Y(n_1959)
);

NAND2xp5_ASAP7_75t_L g1960 ( 
.A(n_1788),
.B(n_568),
.Y(n_1960)
);

NAND2xp5_ASAP7_75t_SL g1961 ( 
.A(n_1838),
.B(n_160),
.Y(n_1961)
);

NAND2xp5_ASAP7_75t_L g1962 ( 
.A(n_1902),
.B(n_567),
.Y(n_1962)
);

NAND2xp5_ASAP7_75t_SL g1963 ( 
.A(n_1777),
.B(n_161),
.Y(n_1963)
);

OAI21x1_ASAP7_75t_L g1964 ( 
.A1(n_1877),
.A2(n_162),
.B(n_164),
.Y(n_1964)
);

AOI21xp5_ASAP7_75t_L g1965 ( 
.A1(n_1906),
.A2(n_164),
.B(n_165),
.Y(n_1965)
);

INVx4_ASAP7_75t_L g1966 ( 
.A(n_1849),
.Y(n_1966)
);

OAI21xp5_ASAP7_75t_L g1967 ( 
.A1(n_1901),
.A2(n_165),
.B(n_166),
.Y(n_1967)
);

CKINVDCx5p33_ASAP7_75t_R g1968 ( 
.A(n_1763),
.Y(n_1968)
);

A2O1A1Ixp33_ASAP7_75t_L g1969 ( 
.A1(n_1813),
.A2(n_1914),
.B(n_1795),
.C(n_1859),
.Y(n_1969)
);

OAI21x1_ASAP7_75t_L g1970 ( 
.A1(n_1835),
.A2(n_166),
.B(n_168),
.Y(n_1970)
);

NOR2xp33_ASAP7_75t_L g1971 ( 
.A(n_1769),
.B(n_169),
.Y(n_1971)
);

OAI21xp33_ASAP7_75t_L g1972 ( 
.A1(n_1908),
.A2(n_567),
.B(n_169),
.Y(n_1972)
);

AOI21xp5_ASAP7_75t_L g1973 ( 
.A1(n_1768),
.A2(n_170),
.B(n_171),
.Y(n_1973)
);

INVx4_ASAP7_75t_L g1974 ( 
.A(n_1843),
.Y(n_1974)
);

NAND2xp5_ASAP7_75t_L g1975 ( 
.A(n_1804),
.B(n_566),
.Y(n_1975)
);

AOI21xp5_ASAP7_75t_L g1976 ( 
.A1(n_1771),
.A2(n_170),
.B(n_171),
.Y(n_1976)
);

AND2x2_ASAP7_75t_L g1977 ( 
.A(n_1893),
.B(n_174),
.Y(n_1977)
);

AND2x2_ASAP7_75t_L g1978 ( 
.A(n_1841),
.B(n_174),
.Y(n_1978)
);

NAND2xp5_ASAP7_75t_SL g1979 ( 
.A(n_1785),
.B(n_175),
.Y(n_1979)
);

NAND2xp5_ASAP7_75t_L g1980 ( 
.A(n_1853),
.B(n_175),
.Y(n_1980)
);

AOI22xp5_ASAP7_75t_L g1981 ( 
.A1(n_1787),
.A2(n_178),
.B1(n_176),
.B2(n_177),
.Y(n_1981)
);

AOI21xp5_ASAP7_75t_L g1982 ( 
.A1(n_1805),
.A2(n_176),
.B(n_177),
.Y(n_1982)
);

NAND2xp5_ASAP7_75t_L g1983 ( 
.A(n_1793),
.B(n_179),
.Y(n_1983)
);

AOI21xp5_ASAP7_75t_L g1984 ( 
.A1(n_1805),
.A2(n_179),
.B(n_180),
.Y(n_1984)
);

INVx1_ASAP7_75t_L g1985 ( 
.A(n_1851),
.Y(n_1985)
);

BUFx6f_ASAP7_75t_L g1986 ( 
.A(n_1878),
.Y(n_1986)
);

BUFx6f_ASAP7_75t_L g1987 ( 
.A(n_1878),
.Y(n_1987)
);

OAI21x1_ASAP7_75t_L g1988 ( 
.A1(n_1858),
.A2(n_180),
.B(n_181),
.Y(n_1988)
);

O2A1O1Ixp5_ASAP7_75t_L g1989 ( 
.A1(n_1783),
.A2(n_183),
.B(n_181),
.C(n_182),
.Y(n_1989)
);

NOR2xp67_ASAP7_75t_L g1990 ( 
.A(n_1767),
.B(n_182),
.Y(n_1990)
);

NAND2xp5_ASAP7_75t_L g1991 ( 
.A(n_1794),
.B(n_183),
.Y(n_1991)
);

OAI21x1_ASAP7_75t_L g1992 ( 
.A1(n_1875),
.A2(n_185),
.B(n_186),
.Y(n_1992)
);

OAI22xp5_ASAP7_75t_L g1993 ( 
.A1(n_1809),
.A2(n_1912),
.B1(n_1781),
.B2(n_1779),
.Y(n_1993)
);

NAND2x1_ASAP7_75t_L g1994 ( 
.A(n_1790),
.B(n_185),
.Y(n_1994)
);

OAI21x1_ASAP7_75t_L g1995 ( 
.A1(n_1909),
.A2(n_186),
.B(n_187),
.Y(n_1995)
);

OAI21x1_ASAP7_75t_SL g1996 ( 
.A1(n_1846),
.A2(n_188),
.B(n_189),
.Y(n_1996)
);

INVx1_ASAP7_75t_L g1997 ( 
.A(n_1865),
.Y(n_1997)
);

CKINVDCx20_ASAP7_75t_R g1998 ( 
.A(n_1824),
.Y(n_1998)
);

NAND2xp5_ASAP7_75t_L g1999 ( 
.A(n_1856),
.B(n_188),
.Y(n_1999)
);

NAND2xp33_ASAP7_75t_L g2000 ( 
.A(n_1809),
.B(n_189),
.Y(n_2000)
);

OAI21x1_ASAP7_75t_L g2001 ( 
.A1(n_1799),
.A2(n_191),
.B(n_193),
.Y(n_2001)
);

NAND2xp5_ASAP7_75t_L g2002 ( 
.A(n_1888),
.B(n_191),
.Y(n_2002)
);

INVx4_ASAP7_75t_L g2003 ( 
.A(n_1821),
.Y(n_2003)
);

A2O1A1Ixp33_ASAP7_75t_L g2004 ( 
.A1(n_1775),
.A2(n_195),
.B(n_193),
.C(n_194),
.Y(n_2004)
);

OAI21x1_ASAP7_75t_L g2005 ( 
.A1(n_1898),
.A2(n_194),
.B(n_195),
.Y(n_2005)
);

NAND2xp5_ASAP7_75t_L g2006 ( 
.A(n_1812),
.B(n_196),
.Y(n_2006)
);

NAND2xp5_ASAP7_75t_L g2007 ( 
.A(n_1814),
.B(n_196),
.Y(n_2007)
);

AND2x2_ASAP7_75t_SL g2008 ( 
.A(n_1758),
.B(n_566),
.Y(n_2008)
);

OAI21x1_ASAP7_75t_L g2009 ( 
.A1(n_1845),
.A2(n_197),
.B(n_198),
.Y(n_2009)
);

OAI21x1_ASAP7_75t_SL g2010 ( 
.A1(n_1844),
.A2(n_199),
.B(n_200),
.Y(n_2010)
);

OAI21x1_ASAP7_75t_L g2011 ( 
.A1(n_1913),
.A2(n_199),
.B(n_201),
.Y(n_2011)
);

NAND2x1p5_ASAP7_75t_L g2012 ( 
.A(n_1790),
.B(n_201),
.Y(n_2012)
);

NAND2xp5_ASAP7_75t_L g2013 ( 
.A(n_1818),
.B(n_565),
.Y(n_2013)
);

INVx2_ASAP7_75t_L g2014 ( 
.A(n_1862),
.Y(n_2014)
);

NAND2xp5_ASAP7_75t_L g2015 ( 
.A(n_1820),
.B(n_565),
.Y(n_2015)
);

NAND2xp5_ASAP7_75t_L g2016 ( 
.A(n_1825),
.B(n_202),
.Y(n_2016)
);

INVx2_ASAP7_75t_L g2017 ( 
.A(n_1884),
.Y(n_2017)
);

AOI21x1_ASAP7_75t_L g2018 ( 
.A1(n_1911),
.A2(n_202),
.B(n_203),
.Y(n_2018)
);

AOI31xp67_ASAP7_75t_L g2019 ( 
.A1(n_1800),
.A2(n_205),
.A3(n_203),
.B(n_204),
.Y(n_2019)
);

AOI21xp5_ASAP7_75t_L g2020 ( 
.A1(n_2000),
.A2(n_1805),
.B(n_1883),
.Y(n_2020)
);

BUFx6f_ASAP7_75t_L g2021 ( 
.A(n_1931),
.Y(n_2021)
);

INVx3_ASAP7_75t_L g2022 ( 
.A(n_1986),
.Y(n_2022)
);

NAND2xp5_ASAP7_75t_L g2023 ( 
.A(n_1958),
.B(n_1832),
.Y(n_2023)
);

BUFx3_ASAP7_75t_L g2024 ( 
.A(n_1922),
.Y(n_2024)
);

AND2x2_ASAP7_75t_L g2025 ( 
.A(n_1926),
.B(n_1831),
.Y(n_2025)
);

AND2x4_ASAP7_75t_L g2026 ( 
.A(n_1925),
.B(n_1870),
.Y(n_2026)
);

INVx3_ASAP7_75t_L g2027 ( 
.A(n_1986),
.Y(n_2027)
);

NOR2x1_ASAP7_75t_SL g2028 ( 
.A(n_1966),
.B(n_1860),
.Y(n_2028)
);

INVx1_ASAP7_75t_SL g2029 ( 
.A(n_1958),
.Y(n_2029)
);

AND2x4_ASAP7_75t_L g2030 ( 
.A(n_1940),
.B(n_1822),
.Y(n_2030)
);

NAND2xp5_ASAP7_75t_L g2031 ( 
.A(n_2014),
.B(n_1836),
.Y(n_2031)
);

HB1xp67_ASAP7_75t_L g2032 ( 
.A(n_1942),
.Y(n_2032)
);

BUFx3_ASAP7_75t_L g2033 ( 
.A(n_1917),
.Y(n_2033)
);

INVx1_ASAP7_75t_L g2034 ( 
.A(n_1957),
.Y(n_2034)
);

CKINVDCx11_ASAP7_75t_R g2035 ( 
.A(n_1998),
.Y(n_2035)
);

HB1xp67_ASAP7_75t_L g2036 ( 
.A(n_1985),
.Y(n_2036)
);

NOR2xp33_ASAP7_75t_SL g2037 ( 
.A(n_1968),
.B(n_1821),
.Y(n_2037)
);

BUFx2_ASAP7_75t_L g2038 ( 
.A(n_1922),
.Y(n_2038)
);

INVx3_ASAP7_75t_L g2039 ( 
.A(n_1986),
.Y(n_2039)
);

OR2x6_ASAP7_75t_L g2040 ( 
.A(n_1927),
.B(n_1951),
.Y(n_2040)
);

CKINVDCx5p33_ASAP7_75t_R g2041 ( 
.A(n_1953),
.Y(n_2041)
);

AOI22xp5_ASAP7_75t_L g2042 ( 
.A1(n_1946),
.A2(n_1797),
.B1(n_1786),
.B2(n_1801),
.Y(n_2042)
);

NAND2xp5_ASAP7_75t_L g2043 ( 
.A(n_2017),
.B(n_1811),
.Y(n_2043)
);

NAND2xp5_ASAP7_75t_L g2044 ( 
.A(n_1921),
.B(n_1791),
.Y(n_2044)
);

AOI21xp5_ASAP7_75t_L g2045 ( 
.A1(n_1923),
.A2(n_1883),
.B(n_1882),
.Y(n_2045)
);

CKINVDCx5p33_ASAP7_75t_R g2046 ( 
.A(n_2003),
.Y(n_2046)
);

AOI21xp5_ASAP7_75t_L g2047 ( 
.A1(n_1928),
.A2(n_1883),
.B(n_1867),
.Y(n_2047)
);

OR2x6_ASAP7_75t_L g2048 ( 
.A(n_1933),
.B(n_1896),
.Y(n_2048)
);

AOI21xp5_ASAP7_75t_L g2049 ( 
.A1(n_1933),
.A2(n_1864),
.B(n_1839),
.Y(n_2049)
);

AND2x2_ASAP7_75t_L g2050 ( 
.A(n_1918),
.B(n_1949),
.Y(n_2050)
);

INVx2_ASAP7_75t_L g2051 ( 
.A(n_1997),
.Y(n_2051)
);

O2A1O1Ixp33_ASAP7_75t_L g2052 ( 
.A1(n_1969),
.A2(n_1778),
.B(n_1854),
.C(n_1842),
.Y(n_2052)
);

AOI21xp5_ASAP7_75t_L g2053 ( 
.A1(n_1936),
.A2(n_1815),
.B(n_1837),
.Y(n_2053)
);

NAND2x1p5_ASAP7_75t_L g2054 ( 
.A(n_1949),
.B(n_1800),
.Y(n_2054)
);

AOI21xp5_ASAP7_75t_L g2055 ( 
.A1(n_1936),
.A2(n_1874),
.B(n_1866),
.Y(n_2055)
);

INVx2_ASAP7_75t_SL g2056 ( 
.A(n_1987),
.Y(n_2056)
);

NOR2xp33_ASAP7_75t_L g2057 ( 
.A(n_1993),
.B(n_1899),
.Y(n_2057)
);

AND2x6_ASAP7_75t_L g2058 ( 
.A(n_1915),
.B(n_1868),
.Y(n_2058)
);

AOI21xp5_ASAP7_75t_L g2059 ( 
.A1(n_1943),
.A2(n_1823),
.B(n_1891),
.Y(n_2059)
);

BUFx3_ASAP7_75t_L g2060 ( 
.A(n_1931),
.Y(n_2060)
);

NAND2xp5_ASAP7_75t_L g2061 ( 
.A(n_1920),
.B(n_1810),
.Y(n_2061)
);

AND2x4_ASAP7_75t_L g2062 ( 
.A(n_2003),
.B(n_1910),
.Y(n_2062)
);

AND2x2_ASAP7_75t_L g2063 ( 
.A(n_1929),
.B(n_1932),
.Y(n_2063)
);

INVxp67_ASAP7_75t_SL g2064 ( 
.A(n_1919),
.Y(n_2064)
);

AOI21x1_ASAP7_75t_L g2065 ( 
.A1(n_1979),
.A2(n_1890),
.B(n_1905),
.Y(n_2065)
);

INVx3_ASAP7_75t_L g2066 ( 
.A(n_1987),
.Y(n_2066)
);

NAND3xp33_ASAP7_75t_L g2067 ( 
.A(n_1967),
.B(n_1782),
.C(n_1904),
.Y(n_2067)
);

INVx1_ASAP7_75t_L g2068 ( 
.A(n_1952),
.Y(n_2068)
);

AND2x2_ASAP7_75t_L g2069 ( 
.A(n_1977),
.B(n_1827),
.Y(n_2069)
);

INVx2_ASAP7_75t_L g2070 ( 
.A(n_1978),
.Y(n_2070)
);

INVx2_ASAP7_75t_SL g2071 ( 
.A(n_1987),
.Y(n_2071)
);

NAND2x1p5_ASAP7_75t_L g2072 ( 
.A(n_1966),
.B(n_1848),
.Y(n_2072)
);

INVx2_ASAP7_75t_SL g2073 ( 
.A(n_1931),
.Y(n_2073)
);

INVx1_ASAP7_75t_L g2074 ( 
.A(n_1952),
.Y(n_2074)
);

NOR3xp33_ASAP7_75t_SL g2075 ( 
.A(n_1950),
.B(n_1789),
.C(n_1881),
.Y(n_2075)
);

A2O1A1Ixp33_ASAP7_75t_L g2076 ( 
.A1(n_1972),
.A2(n_1863),
.B(n_1892),
.C(n_1808),
.Y(n_2076)
);

BUFx3_ASAP7_75t_L g2077 ( 
.A(n_1938),
.Y(n_2077)
);

AO21x1_ASAP7_75t_L g2078 ( 
.A1(n_1967),
.A2(n_1943),
.B(n_1939),
.Y(n_2078)
);

INVx3_ASAP7_75t_SL g2079 ( 
.A(n_1938),
.Y(n_2079)
);

INVx2_ASAP7_75t_L g2080 ( 
.A(n_1975),
.Y(n_2080)
);

INVx3_ASAP7_75t_L g2081 ( 
.A(n_1974),
.Y(n_2081)
);

NAND2xp5_ASAP7_75t_L g2082 ( 
.A(n_1954),
.B(n_1885),
.Y(n_2082)
);

O2A1O1Ixp33_ASAP7_75t_L g2083 ( 
.A1(n_2004),
.A2(n_1806),
.B(n_1802),
.C(n_1869),
.Y(n_2083)
);

INVx1_ASAP7_75t_L g2084 ( 
.A(n_2032),
.Y(n_2084)
);

OAI22xp5_ASAP7_75t_L g2085 ( 
.A1(n_2042),
.A2(n_1981),
.B1(n_2008),
.B2(n_1934),
.Y(n_2085)
);

AND2x4_ASAP7_75t_L g2086 ( 
.A(n_2024),
.B(n_1990),
.Y(n_2086)
);

CKINVDCx5p33_ASAP7_75t_R g2087 ( 
.A(n_2035),
.Y(n_2087)
);

BUFx3_ASAP7_75t_L g2088 ( 
.A(n_2024),
.Y(n_2088)
);

CKINVDCx5p33_ASAP7_75t_R g2089 ( 
.A(n_2035),
.Y(n_2089)
);

OAI22xp33_ASAP7_75t_L g2090 ( 
.A1(n_2048),
.A2(n_1981),
.B1(n_1915),
.B2(n_1937),
.Y(n_2090)
);

AOI22xp33_ASAP7_75t_L g2091 ( 
.A1(n_2058),
.A2(n_1972),
.B1(n_1934),
.B2(n_1963),
.Y(n_2091)
);

INVx3_ASAP7_75t_L g2092 ( 
.A(n_2051),
.Y(n_2092)
);

INVx1_ASAP7_75t_L g2093 ( 
.A(n_2032),
.Y(n_2093)
);

INVx2_ASAP7_75t_SL g2094 ( 
.A(n_2038),
.Y(n_2094)
);

INVx6_ASAP7_75t_L g2095 ( 
.A(n_2077),
.Y(n_2095)
);

INVx4_ASAP7_75t_L g2096 ( 
.A(n_2079),
.Y(n_2096)
);

INVx1_ASAP7_75t_L g2097 ( 
.A(n_2036),
.Y(n_2097)
);

INVx1_ASAP7_75t_L g2098 ( 
.A(n_2036),
.Y(n_2098)
);

AOI22xp33_ASAP7_75t_L g2099 ( 
.A1(n_2058),
.A2(n_1961),
.B1(n_1965),
.B2(n_1971),
.Y(n_2099)
);

OAI22xp33_ASAP7_75t_L g2100 ( 
.A1(n_2048),
.A2(n_1973),
.B1(n_1990),
.B2(n_1976),
.Y(n_2100)
);

BUFx3_ASAP7_75t_L g2101 ( 
.A(n_2062),
.Y(n_2101)
);

BUFx6f_ASAP7_75t_L g2102 ( 
.A(n_2077),
.Y(n_2102)
);

BUFx12f_ASAP7_75t_L g2103 ( 
.A(n_2041),
.Y(n_2103)
);

BUFx10_ASAP7_75t_L g2104 ( 
.A(n_2046),
.Y(n_2104)
);

AOI22xp33_ASAP7_75t_L g2105 ( 
.A1(n_2058),
.A2(n_1962),
.B1(n_2010),
.B2(n_1996),
.Y(n_2105)
);

INVx3_ASAP7_75t_L g2106 ( 
.A(n_2030),
.Y(n_2106)
);

BUFx4f_ASAP7_75t_SL g2107 ( 
.A(n_2033),
.Y(n_2107)
);

BUFx6f_ASAP7_75t_L g2108 ( 
.A(n_2079),
.Y(n_2108)
);

INVx2_ASAP7_75t_L g2109 ( 
.A(n_2034),
.Y(n_2109)
);

INVx1_ASAP7_75t_L g2110 ( 
.A(n_2068),
.Y(n_2110)
);

OAI22xp5_ASAP7_75t_L g2111 ( 
.A1(n_2067),
.A2(n_2012),
.B1(n_1956),
.B2(n_2002),
.Y(n_2111)
);

INVx1_ASAP7_75t_L g2112 ( 
.A(n_2074),
.Y(n_2112)
);

BUFx2_ASAP7_75t_L g2113 ( 
.A(n_2030),
.Y(n_2113)
);

INVx1_ASAP7_75t_L g2114 ( 
.A(n_2029),
.Y(n_2114)
);

OAI22xp5_ASAP7_75t_L g2115 ( 
.A1(n_2055),
.A2(n_1960),
.B1(n_1991),
.B2(n_1983),
.Y(n_2115)
);

NAND2xp5_ASAP7_75t_L g2116 ( 
.A(n_2044),
.B(n_2006),
.Y(n_2116)
);

NAND2xp5_ASAP7_75t_L g2117 ( 
.A(n_2023),
.B(n_2007),
.Y(n_2117)
);

BUFx3_ASAP7_75t_L g2118 ( 
.A(n_2062),
.Y(n_2118)
);

AOI22xp33_ASAP7_75t_L g2119 ( 
.A1(n_2058),
.A2(n_2009),
.B1(n_1930),
.B2(n_1999),
.Y(n_2119)
);

CKINVDCx20_ASAP7_75t_R g2120 ( 
.A(n_2063),
.Y(n_2120)
);

OAI21xp5_ASAP7_75t_SL g2121 ( 
.A1(n_2057),
.A2(n_1872),
.B(n_2013),
.Y(n_2121)
);

AOI22xp33_ASAP7_75t_SL g2122 ( 
.A1(n_2058),
.A2(n_1959),
.B1(n_1992),
.B2(n_1988),
.Y(n_2122)
);

INVx4_ASAP7_75t_L g2123 ( 
.A(n_2081),
.Y(n_2123)
);

AOI22xp33_ASAP7_75t_SL g2124 ( 
.A1(n_2057),
.A2(n_1970),
.B1(n_1948),
.B2(n_1941),
.Y(n_2124)
);

CKINVDCx11_ASAP7_75t_R g2125 ( 
.A(n_2021),
.Y(n_2125)
);

BUFx6f_ASAP7_75t_L g2126 ( 
.A(n_2021),
.Y(n_2126)
);

OR2x2_ASAP7_75t_L g2127 ( 
.A(n_2093),
.B(n_2064),
.Y(n_2127)
);

OAI22xp5_ASAP7_75t_L g2128 ( 
.A1(n_2091),
.A2(n_2055),
.B1(n_2053),
.B2(n_2049),
.Y(n_2128)
);

INVx2_ASAP7_75t_L g2129 ( 
.A(n_2110),
.Y(n_2129)
);

AND2x2_ASAP7_75t_L g2130 ( 
.A(n_2113),
.B(n_2050),
.Y(n_2130)
);

AND2x2_ASAP7_75t_L g2131 ( 
.A(n_2113),
.B(n_2064),
.Y(n_2131)
);

AND2x2_ASAP7_75t_L g2132 ( 
.A(n_2094),
.B(n_2026),
.Y(n_2132)
);

INVx1_ASAP7_75t_L g2133 ( 
.A(n_2093),
.Y(n_2133)
);

INVx2_ASAP7_75t_L g2134 ( 
.A(n_2112),
.Y(n_2134)
);

INVx1_ASAP7_75t_L g2135 ( 
.A(n_2084),
.Y(n_2135)
);

NOR2xp33_ASAP7_75t_L g2136 ( 
.A(n_2087),
.B(n_2061),
.Y(n_2136)
);

INVx1_ASAP7_75t_L g2137 ( 
.A(n_2097),
.Y(n_2137)
);

AND2x2_ASAP7_75t_L g2138 ( 
.A(n_2094),
.B(n_2106),
.Y(n_2138)
);

NOR2xp67_ASAP7_75t_L g2139 ( 
.A(n_2096),
.B(n_2081),
.Y(n_2139)
);

INVx2_ASAP7_75t_L g2140 ( 
.A(n_2109),
.Y(n_2140)
);

AOI21xp5_ASAP7_75t_SL g2141 ( 
.A1(n_2085),
.A2(n_2048),
.B(n_2053),
.Y(n_2141)
);

AND2x2_ASAP7_75t_L g2142 ( 
.A(n_2106),
.B(n_2026),
.Y(n_2142)
);

OAI22xp5_ASAP7_75t_L g2143 ( 
.A1(n_2099),
.A2(n_2049),
.B1(n_2076),
.B2(n_2054),
.Y(n_2143)
);

O2A1O1Ixp5_ASAP7_75t_L g2144 ( 
.A1(n_2090),
.A2(n_2078),
.B(n_2059),
.C(n_2020),
.Y(n_2144)
);

OAI22xp5_ASAP7_75t_L g2145 ( 
.A1(n_2105),
.A2(n_2076),
.B1(n_2054),
.B2(n_2075),
.Y(n_2145)
);

OAI22xp5_ASAP7_75t_L g2146 ( 
.A1(n_2120),
.A2(n_2075),
.B1(n_2059),
.B2(n_2052),
.Y(n_2146)
);

INVx2_ASAP7_75t_L g2147 ( 
.A(n_2109),
.Y(n_2147)
);

AND2x2_ASAP7_75t_L g2148 ( 
.A(n_2106),
.B(n_2025),
.Y(n_2148)
);

INVx2_ASAP7_75t_L g2149 ( 
.A(n_2092),
.Y(n_2149)
);

OAI31xp33_ASAP7_75t_L g2150 ( 
.A1(n_2100),
.A2(n_2052),
.A3(n_2083),
.B(n_2045),
.Y(n_2150)
);

INVx2_ASAP7_75t_L g2151 ( 
.A(n_2140),
.Y(n_2151)
);

AND2x4_ASAP7_75t_SL g2152 ( 
.A(n_2132),
.B(n_2104),
.Y(n_2152)
);

NAND2xp33_ASAP7_75t_R g2153 ( 
.A(n_2136),
.B(n_2087),
.Y(n_2153)
);

AND2x4_ASAP7_75t_L g2154 ( 
.A(n_2139),
.B(n_2096),
.Y(n_2154)
);

NAND2xp5_ASAP7_75t_L g2155 ( 
.A(n_2128),
.B(n_2114),
.Y(n_2155)
);

NAND2xp5_ASAP7_75t_L g2156 ( 
.A(n_2128),
.B(n_2092),
.Y(n_2156)
);

AND2x2_ASAP7_75t_L g2157 ( 
.A(n_2142),
.B(n_2132),
.Y(n_2157)
);

AND2x2_ASAP7_75t_L g2158 ( 
.A(n_2142),
.B(n_2088),
.Y(n_2158)
);

INVx2_ASAP7_75t_L g2159 ( 
.A(n_2140),
.Y(n_2159)
);

CKINVDCx5p33_ASAP7_75t_R g2160 ( 
.A(n_2146),
.Y(n_2160)
);

INVx2_ASAP7_75t_L g2161 ( 
.A(n_2151),
.Y(n_2161)
);

BUFx6f_ASAP7_75t_L g2162 ( 
.A(n_2154),
.Y(n_2162)
);

INVx1_ASAP7_75t_L g2163 ( 
.A(n_2151),
.Y(n_2163)
);

AND2x2_ASAP7_75t_L g2164 ( 
.A(n_2154),
.B(n_2138),
.Y(n_2164)
);

AND2x2_ASAP7_75t_L g2165 ( 
.A(n_2154),
.B(n_2138),
.Y(n_2165)
);

OA21x2_ASAP7_75t_L g2166 ( 
.A1(n_2159),
.A2(n_2144),
.B(n_2134),
.Y(n_2166)
);

INVx1_ASAP7_75t_L g2167 ( 
.A(n_2159),
.Y(n_2167)
);

NAND4xp25_ASAP7_75t_L g2168 ( 
.A(n_2155),
.B(n_2150),
.C(n_2141),
.D(n_2146),
.Y(n_2168)
);

INVx1_ASAP7_75t_L g2169 ( 
.A(n_2163),
.Y(n_2169)
);

INVx2_ASAP7_75t_L g2170 ( 
.A(n_2166),
.Y(n_2170)
);

NAND2x1_ASAP7_75t_L g2171 ( 
.A(n_2162),
.B(n_2141),
.Y(n_2171)
);

AND2x2_ASAP7_75t_L g2172 ( 
.A(n_2164),
.B(n_2152),
.Y(n_2172)
);

NAND2xp5_ASAP7_75t_L g2173 ( 
.A(n_2168),
.B(n_2160),
.Y(n_2173)
);

AND2x2_ASAP7_75t_L g2174 ( 
.A(n_2164),
.B(n_2152),
.Y(n_2174)
);

INVxp67_ASAP7_75t_SL g2175 ( 
.A(n_2162),
.Y(n_2175)
);

INVx1_ASAP7_75t_L g2176 ( 
.A(n_2163),
.Y(n_2176)
);

AND2x2_ASAP7_75t_L g2177 ( 
.A(n_2165),
.B(n_2157),
.Y(n_2177)
);

INVx2_ASAP7_75t_L g2178 ( 
.A(n_2166),
.Y(n_2178)
);

NAND2xp5_ASAP7_75t_L g2179 ( 
.A(n_2175),
.B(n_2160),
.Y(n_2179)
);

INVx2_ASAP7_75t_L g2180 ( 
.A(n_2177),
.Y(n_2180)
);

INVx2_ASAP7_75t_L g2181 ( 
.A(n_2177),
.Y(n_2181)
);

AND2x2_ASAP7_75t_L g2182 ( 
.A(n_2172),
.B(n_2174),
.Y(n_2182)
);

AOI22xp5_ASAP7_75t_L g2183 ( 
.A1(n_2173),
.A2(n_2143),
.B1(n_2145),
.B2(n_2115),
.Y(n_2183)
);

NAND2xp5_ASAP7_75t_L g2184 ( 
.A(n_2172),
.B(n_2156),
.Y(n_2184)
);

AOI22xp33_ASAP7_75t_L g2185 ( 
.A1(n_2171),
.A2(n_2143),
.B1(n_2150),
.B2(n_2145),
.Y(n_2185)
);

NAND3xp33_ASAP7_75t_L g2186 ( 
.A(n_2169),
.B(n_2162),
.C(n_2119),
.Y(n_2186)
);

NOR2xp33_ASAP7_75t_L g2187 ( 
.A(n_2174),
.B(n_2089),
.Y(n_2187)
);

INVx2_ASAP7_75t_L g2188 ( 
.A(n_2178),
.Y(n_2188)
);

AOI221xp5_ASAP7_75t_L g2189 ( 
.A1(n_2176),
.A2(n_2111),
.B1(n_2162),
.B2(n_1876),
.C(n_2121),
.Y(n_2189)
);

INVx2_ASAP7_75t_L g2190 ( 
.A(n_2180),
.Y(n_2190)
);

NAND2xp5_ASAP7_75t_L g2191 ( 
.A(n_2179),
.B(n_2165),
.Y(n_2191)
);

INVx2_ASAP7_75t_SL g2192 ( 
.A(n_2182),
.Y(n_2192)
);

AND2x2_ASAP7_75t_L g2193 ( 
.A(n_2181),
.B(n_2162),
.Y(n_2193)
);

AND2x2_ASAP7_75t_L g2194 ( 
.A(n_2187),
.B(n_2170),
.Y(n_2194)
);

INVx1_ASAP7_75t_L g2195 ( 
.A(n_2188),
.Y(n_2195)
);

INVx1_ASAP7_75t_L g2196 ( 
.A(n_2186),
.Y(n_2196)
);

AND2x4_ASAP7_75t_L g2197 ( 
.A(n_2184),
.B(n_2170),
.Y(n_2197)
);

AND2x2_ASAP7_75t_L g2198 ( 
.A(n_2185),
.B(n_2178),
.Y(n_2198)
);

INVx1_ASAP7_75t_L g2199 ( 
.A(n_2190),
.Y(n_2199)
);

BUFx2_ASAP7_75t_L g2200 ( 
.A(n_2192),
.Y(n_2200)
);

NOR2xp33_ASAP7_75t_L g2201 ( 
.A(n_2192),
.B(n_2089),
.Y(n_2201)
);

INVx1_ASAP7_75t_L g2202 ( 
.A(n_2190),
.Y(n_2202)
);

O2A1O1Ixp33_ASAP7_75t_SL g2203 ( 
.A1(n_2201),
.A2(n_2196),
.B(n_2189),
.C(n_2195),
.Y(n_2203)
);

AND2x4_ASAP7_75t_L g2204 ( 
.A(n_2200),
.B(n_2193),
.Y(n_2204)
);

INVx1_ASAP7_75t_L g2205 ( 
.A(n_2199),
.Y(n_2205)
);

INVx1_ASAP7_75t_SL g2206 ( 
.A(n_2201),
.Y(n_2206)
);

A2O1A1Ixp33_ASAP7_75t_L g2207 ( 
.A1(n_2204),
.A2(n_2198),
.B(n_2183),
.C(n_2197),
.Y(n_2207)
);

OAI21xp33_ASAP7_75t_L g2208 ( 
.A1(n_2206),
.A2(n_2198),
.B(n_2191),
.Y(n_2208)
);

BUFx2_ASAP7_75t_SL g2209 ( 
.A(n_2204),
.Y(n_2209)
);

AND2x4_ASAP7_75t_L g2210 ( 
.A(n_2205),
.B(n_2202),
.Y(n_2210)
);

OA22x2_ASAP7_75t_L g2211 ( 
.A1(n_2203),
.A2(n_2183),
.B1(n_2195),
.B2(n_2194),
.Y(n_2211)
);

AOI21xp5_ASAP7_75t_L g2212 ( 
.A1(n_2203),
.A2(n_2194),
.B(n_2197),
.Y(n_2212)
);

INVx1_ASAP7_75t_L g2213 ( 
.A(n_2209),
.Y(n_2213)
);

OR2x2_ASAP7_75t_L g2214 ( 
.A(n_2207),
.B(n_2197),
.Y(n_2214)
);

AND2x2_ASAP7_75t_L g2215 ( 
.A(n_2208),
.B(n_2193),
.Y(n_2215)
);

HB1xp67_ASAP7_75t_L g2216 ( 
.A(n_2210),
.Y(n_2216)
);

AND2x4_ASAP7_75t_L g2217 ( 
.A(n_2212),
.B(n_2161),
.Y(n_2217)
);

INVx1_ASAP7_75t_SL g2218 ( 
.A(n_2211),
.Y(n_2218)
);

OR2x6_ASAP7_75t_L g2219 ( 
.A(n_2209),
.B(n_2103),
.Y(n_2219)
);

HB1xp67_ASAP7_75t_L g2220 ( 
.A(n_2209),
.Y(n_2220)
);

AND2x2_ASAP7_75t_L g2221 ( 
.A(n_2209),
.B(n_2103),
.Y(n_2221)
);

AND2x4_ASAP7_75t_L g2222 ( 
.A(n_2210),
.B(n_2161),
.Y(n_2222)
);

NAND3xp33_ASAP7_75t_L g2223 ( 
.A(n_2220),
.B(n_1824),
.C(n_2037),
.Y(n_2223)
);

INVxp67_ASAP7_75t_SL g2224 ( 
.A(n_2216),
.Y(n_2224)
);

INVx2_ASAP7_75t_L g2225 ( 
.A(n_2221),
.Y(n_2225)
);

INVx1_ASAP7_75t_L g2226 ( 
.A(n_2213),
.Y(n_2226)
);

AND2x2_ASAP7_75t_L g2227 ( 
.A(n_2219),
.B(n_2104),
.Y(n_2227)
);

NAND2xp5_ASAP7_75t_L g2228 ( 
.A(n_2213),
.B(n_2166),
.Y(n_2228)
);

AOI21xp33_ASAP7_75t_L g2229 ( 
.A1(n_2219),
.A2(n_2153),
.B(n_2016),
.Y(n_2229)
);

INVx1_ASAP7_75t_L g2230 ( 
.A(n_2215),
.Y(n_2230)
);

OAI22xp33_ASAP7_75t_SL g2231 ( 
.A1(n_2214),
.A2(n_2167),
.B1(n_2096),
.B2(n_2095),
.Y(n_2231)
);

NOR2xp33_ASAP7_75t_L g2232 ( 
.A(n_2218),
.B(n_2107),
.Y(n_2232)
);

NAND3xp33_ASAP7_75t_L g2233 ( 
.A(n_2217),
.B(n_2015),
.C(n_1944),
.Y(n_2233)
);

AOI21xp33_ASAP7_75t_L g2234 ( 
.A1(n_2217),
.A2(n_2166),
.B(n_2082),
.Y(n_2234)
);

OAI22xp5_ASAP7_75t_L g2235 ( 
.A1(n_2222),
.A2(n_2167),
.B1(n_2120),
.B2(n_2139),
.Y(n_2235)
);

INVx2_ASAP7_75t_L g2236 ( 
.A(n_2227),
.Y(n_2236)
);

OAI21xp5_ASAP7_75t_L g2237 ( 
.A1(n_2224),
.A2(n_2222),
.B(n_1803),
.Y(n_2237)
);

AND2x2_ASAP7_75t_L g2238 ( 
.A(n_2232),
.B(n_2104),
.Y(n_2238)
);

OR2x2_ASAP7_75t_L g2239 ( 
.A(n_2230),
.B(n_2116),
.Y(n_2239)
);

INVx2_ASAP7_75t_SL g2240 ( 
.A(n_2226),
.Y(n_2240)
);

NAND2xp5_ASAP7_75t_L g2241 ( 
.A(n_2225),
.B(n_2117),
.Y(n_2241)
);

NAND2xp5_ASAP7_75t_L g2242 ( 
.A(n_2229),
.B(n_2069),
.Y(n_2242)
);

AO21x1_ASAP7_75t_L g2243 ( 
.A1(n_2228),
.A2(n_1784),
.B(n_1830),
.Y(n_2243)
);

OAI22xp5_ASAP7_75t_L g2244 ( 
.A1(n_2223),
.A2(n_2095),
.B1(n_2108),
.B2(n_2102),
.Y(n_2244)
);

INVx1_ASAP7_75t_SL g2245 ( 
.A(n_2233),
.Y(n_2245)
);

AOI22xp33_ASAP7_75t_SL g2246 ( 
.A1(n_2231),
.A2(n_2108),
.B1(n_2095),
.B2(n_1938),
.Y(n_2246)
);

AO22x1_ASAP7_75t_L g2247 ( 
.A1(n_2235),
.A2(n_1974),
.B1(n_1852),
.B2(n_2108),
.Y(n_2247)
);

OAI22xp5_ASAP7_75t_L g2248 ( 
.A1(n_2234),
.A2(n_2095),
.B1(n_2108),
.B2(n_2102),
.Y(n_2248)
);

NAND5xp2_ASAP7_75t_SL g2249 ( 
.A(n_2227),
.B(n_2158),
.C(n_2083),
.D(n_1984),
.E(n_1982),
.Y(n_2249)
);

INVx2_ASAP7_75t_L g2250 ( 
.A(n_2227),
.Y(n_2250)
);

AND2x2_ASAP7_75t_L g2251 ( 
.A(n_2238),
.B(n_2158),
.Y(n_2251)
);

OR2x2_ASAP7_75t_L g2252 ( 
.A(n_2240),
.B(n_2135),
.Y(n_2252)
);

NAND2x1_ASAP7_75t_L g2253 ( 
.A(n_2237),
.B(n_2108),
.Y(n_2253)
);

INVx1_ASAP7_75t_L g2254 ( 
.A(n_2242),
.Y(n_2254)
);

AND2x2_ASAP7_75t_L g2255 ( 
.A(n_2236),
.B(n_2148),
.Y(n_2255)
);

NAND2xp5_ASAP7_75t_L g2256 ( 
.A(n_2245),
.B(n_2135),
.Y(n_2256)
);

INVx1_ASAP7_75t_L g2257 ( 
.A(n_2239),
.Y(n_2257)
);

AND2x2_ASAP7_75t_L g2258 ( 
.A(n_2250),
.B(n_2148),
.Y(n_2258)
);

AND2x2_ASAP7_75t_L g2259 ( 
.A(n_2241),
.B(n_2130),
.Y(n_2259)
);

AND2x2_ASAP7_75t_L g2260 ( 
.A(n_2246),
.B(n_2130),
.Y(n_2260)
);

NOR2xp33_ASAP7_75t_L g2261 ( 
.A(n_2243),
.B(n_2043),
.Y(n_2261)
);

OR2x2_ASAP7_75t_L g2262 ( 
.A(n_2248),
.B(n_2137),
.Y(n_2262)
);

AND2x2_ASAP7_75t_L g2263 ( 
.A(n_2244),
.B(n_2131),
.Y(n_2263)
);

INVx1_ASAP7_75t_L g2264 ( 
.A(n_2247),
.Y(n_2264)
);

NAND2xp5_ASAP7_75t_SL g2265 ( 
.A(n_2257),
.B(n_2249),
.Y(n_2265)
);

NOR2xp33_ASAP7_75t_SL g2266 ( 
.A(n_2264),
.B(n_1770),
.Y(n_2266)
);

AOI211xp5_ASAP7_75t_SL g2267 ( 
.A1(n_2264),
.A2(n_1886),
.B(n_1980),
.C(n_2031),
.Y(n_2267)
);

NOR3xp33_ASAP7_75t_L g2268 ( 
.A(n_2254),
.B(n_2253),
.C(n_2256),
.Y(n_2268)
);

NAND3xp33_ASAP7_75t_SL g2269 ( 
.A(n_2252),
.B(n_1945),
.C(n_1994),
.Y(n_2269)
);

AOI222xp33_ASAP7_75t_L g2270 ( 
.A1(n_2260),
.A2(n_2263),
.B1(n_2258),
.B2(n_2255),
.C1(n_2251),
.C2(n_2261),
.Y(n_2270)
);

NAND2xp5_ASAP7_75t_L g2271 ( 
.A(n_2259),
.B(n_2262),
.Y(n_2271)
);

AOI21xp5_ASAP7_75t_L g2272 ( 
.A1(n_2253),
.A2(n_2011),
.B(n_1989),
.Y(n_2272)
);

NAND3xp33_ASAP7_75t_SL g2273 ( 
.A(n_2257),
.B(n_2072),
.C(n_1935),
.Y(n_2273)
);

AOI221xp5_ASAP7_75t_L g2274 ( 
.A1(n_2264),
.A2(n_2137),
.B1(n_2080),
.B2(n_2045),
.C(n_2102),
.Y(n_2274)
);

NAND2xp5_ASAP7_75t_L g2275 ( 
.A(n_2251),
.B(n_2133),
.Y(n_2275)
);

OAI211xp5_ASAP7_75t_L g2276 ( 
.A1(n_2264),
.A2(n_2018),
.B(n_2125),
.C(n_206),
.Y(n_2276)
);

INVx2_ASAP7_75t_L g2277 ( 
.A(n_2251),
.Y(n_2277)
);

NOR2xp33_ASAP7_75t_L g2278 ( 
.A(n_2251),
.B(n_204),
.Y(n_2278)
);

NOR3x1_ASAP7_75t_L g2279 ( 
.A(n_2253),
.B(n_1995),
.C(n_1964),
.Y(n_2279)
);

OR2x2_ASAP7_75t_L g2280 ( 
.A(n_2257),
.B(n_2133),
.Y(n_2280)
);

INVx1_ASAP7_75t_L g2281 ( 
.A(n_2255),
.Y(n_2281)
);

NOR3x1_ASAP7_75t_L g2282 ( 
.A(n_2253),
.B(n_2001),
.C(n_205),
.Y(n_2282)
);

OAI211xp5_ASAP7_75t_L g2283 ( 
.A1(n_2264),
.A2(n_2125),
.B(n_209),
.C(n_207),
.Y(n_2283)
);

AOI221xp5_ASAP7_75t_L g2284 ( 
.A1(n_2264),
.A2(n_2102),
.B1(n_2047),
.B2(n_2086),
.C(n_209),
.Y(n_2284)
);

NOR3xp33_ASAP7_75t_SL g2285 ( 
.A(n_2264),
.B(n_207),
.C(n_208),
.Y(n_2285)
);

AND4x1_ASAP7_75t_L g2286 ( 
.A(n_2257),
.B(n_211),
.C(n_208),
.D(n_210),
.Y(n_2286)
);

NAND3xp33_ASAP7_75t_L g2287 ( 
.A(n_2285),
.B(n_210),
.C(n_211),
.Y(n_2287)
);

OAI211xp5_ASAP7_75t_L g2288 ( 
.A1(n_2283),
.A2(n_214),
.B(n_212),
.C(n_213),
.Y(n_2288)
);

INVx1_ASAP7_75t_SL g2289 ( 
.A(n_2277),
.Y(n_2289)
);

NAND2xp5_ASAP7_75t_L g2290 ( 
.A(n_2286),
.B(n_2278),
.Y(n_2290)
);

NAND2xp5_ASAP7_75t_L g2291 ( 
.A(n_2270),
.B(n_212),
.Y(n_2291)
);

NAND2xp5_ASAP7_75t_L g2292 ( 
.A(n_2281),
.B(n_213),
.Y(n_2292)
);

NOR2x1_ASAP7_75t_L g2293 ( 
.A(n_2271),
.B(n_214),
.Y(n_2293)
);

INVx1_ASAP7_75t_L g2294 ( 
.A(n_2280),
.Y(n_2294)
);

NAND2x1_ASAP7_75t_L g2295 ( 
.A(n_2268),
.B(n_1878),
.Y(n_2295)
);

INVx1_ASAP7_75t_L g2296 ( 
.A(n_2266),
.Y(n_2296)
);

NOR3xp33_ASAP7_75t_L g2297 ( 
.A(n_2265),
.B(n_2065),
.C(n_217),
.Y(n_2297)
);

NAND2xp5_ASAP7_75t_SL g2298 ( 
.A(n_2284),
.B(n_2102),
.Y(n_2298)
);

NAND4xp25_ASAP7_75t_L g2299 ( 
.A(n_2282),
.B(n_220),
.C(n_217),
.D(n_218),
.Y(n_2299)
);

INVx1_ASAP7_75t_L g2300 ( 
.A(n_2275),
.Y(n_2300)
);

O2A1O1Ixp33_ASAP7_75t_SL g2301 ( 
.A1(n_2276),
.A2(n_221),
.B(n_218),
.C(n_220),
.Y(n_2301)
);

INVx1_ASAP7_75t_L g2302 ( 
.A(n_2269),
.Y(n_2302)
);

NAND2xp5_ASAP7_75t_L g2303 ( 
.A(n_2267),
.B(n_221),
.Y(n_2303)
);

NAND3xp33_ASAP7_75t_L g2304 ( 
.A(n_2274),
.B(n_222),
.C(n_223),
.Y(n_2304)
);

INVx1_ASAP7_75t_L g2305 ( 
.A(n_2273),
.Y(n_2305)
);

NAND2xp5_ASAP7_75t_L g2306 ( 
.A(n_2272),
.B(n_223),
.Y(n_2306)
);

HB1xp67_ASAP7_75t_L g2307 ( 
.A(n_2279),
.Y(n_2307)
);

AND2x2_ASAP7_75t_L g2308 ( 
.A(n_2277),
.B(n_2131),
.Y(n_2308)
);

NOR2xp67_ASAP7_75t_L g2309 ( 
.A(n_2283),
.B(n_224),
.Y(n_2309)
);

NOR2x1_ASAP7_75t_L g2310 ( 
.A(n_2283),
.B(n_224),
.Y(n_2310)
);

OAI322xp33_ASAP7_75t_L g2311 ( 
.A1(n_2266),
.A2(n_2072),
.A3(n_231),
.B1(n_227),
.B2(n_230),
.C1(n_225),
.C2(n_226),
.Y(n_2311)
);

NAND4xp25_ASAP7_75t_SL g2312 ( 
.A(n_2270),
.B(n_2122),
.C(n_2124),
.D(n_2127),
.Y(n_2312)
);

NOR3xp33_ASAP7_75t_L g2313 ( 
.A(n_2277),
.B(n_226),
.C(n_227),
.Y(n_2313)
);

OAI22xp5_ASAP7_75t_L g2314 ( 
.A1(n_2277),
.A2(n_2127),
.B1(n_2126),
.B2(n_2123),
.Y(n_2314)
);

NAND3xp33_ASAP7_75t_SL g2315 ( 
.A(n_2283),
.B(n_1924),
.C(n_228),
.Y(n_2315)
);

NOR3xp33_ASAP7_75t_SL g2316 ( 
.A(n_2283),
.B(n_228),
.C(n_230),
.Y(n_2316)
);

AOI221xp5_ASAP7_75t_L g2317 ( 
.A1(n_2283),
.A2(n_233),
.B1(n_231),
.B2(n_232),
.C(n_234),
.Y(n_2317)
);

NAND2xp5_ASAP7_75t_L g2318 ( 
.A(n_2286),
.B(n_232),
.Y(n_2318)
);

NAND2xp5_ASAP7_75t_L g2319 ( 
.A(n_2286),
.B(n_234),
.Y(n_2319)
);

INVx1_ASAP7_75t_L g2320 ( 
.A(n_2286),
.Y(n_2320)
);

NOR2xp33_ASAP7_75t_L g2321 ( 
.A(n_2286),
.B(n_235),
.Y(n_2321)
);

AOI22x1_ASAP7_75t_L g2322 ( 
.A1(n_2277),
.A2(n_238),
.B1(n_236),
.B2(n_237),
.Y(n_2322)
);

INVx1_ASAP7_75t_L g2323 ( 
.A(n_2286),
.Y(n_2323)
);

INVx1_ASAP7_75t_L g2324 ( 
.A(n_2293),
.Y(n_2324)
);

NOR2x1_ASAP7_75t_L g2325 ( 
.A(n_2287),
.B(n_237),
.Y(n_2325)
);

NAND2xp5_ASAP7_75t_L g2326 ( 
.A(n_2289),
.B(n_238),
.Y(n_2326)
);

INVx2_ASAP7_75t_SL g2327 ( 
.A(n_2295),
.Y(n_2327)
);

NOR2xp67_ASAP7_75t_L g2328 ( 
.A(n_2299),
.B(n_239),
.Y(n_2328)
);

O2A1O1Ixp33_ASAP7_75t_L g2329 ( 
.A1(n_2301),
.A2(n_241),
.B(n_239),
.C(n_240),
.Y(n_2329)
);

OAI221xp5_ASAP7_75t_L g2330 ( 
.A1(n_2317),
.A2(n_2040),
.B1(n_2070),
.B2(n_242),
.C(n_240),
.Y(n_2330)
);

NOR3xp33_ASAP7_75t_L g2331 ( 
.A(n_2291),
.B(n_241),
.C(n_242),
.Y(n_2331)
);

AOI21xp5_ASAP7_75t_L g2332 ( 
.A1(n_2290),
.A2(n_2028),
.B(n_243),
.Y(n_2332)
);

NAND2xp5_ASAP7_75t_L g2333 ( 
.A(n_2289),
.B(n_244),
.Y(n_2333)
);

NAND2xp5_ASAP7_75t_L g2334 ( 
.A(n_2321),
.B(n_244),
.Y(n_2334)
);

NAND2xp5_ASAP7_75t_L g2335 ( 
.A(n_2308),
.B(n_245),
.Y(n_2335)
);

NAND3xp33_ASAP7_75t_SL g2336 ( 
.A(n_2288),
.B(n_245),
.C(n_246),
.Y(n_2336)
);

NAND3xp33_ASAP7_75t_L g2337 ( 
.A(n_2316),
.B(n_246),
.C(n_247),
.Y(n_2337)
);

INVx1_ASAP7_75t_L g2338 ( 
.A(n_2318),
.Y(n_2338)
);

NOR2xp33_ASAP7_75t_L g2339 ( 
.A(n_2319),
.B(n_2320),
.Y(n_2339)
);

NAND2xp5_ASAP7_75t_L g2340 ( 
.A(n_2309),
.B(n_247),
.Y(n_2340)
);

OAI21xp5_ASAP7_75t_L g2341 ( 
.A1(n_2310),
.A2(n_1955),
.B(n_2005),
.Y(n_2341)
);

INVx1_ASAP7_75t_L g2342 ( 
.A(n_2292),
.Y(n_2342)
);

AND4x1_ASAP7_75t_L g2343 ( 
.A(n_2313),
.B(n_250),
.C(n_248),
.D(n_249),
.Y(n_2343)
);

AND4x1_ASAP7_75t_L g2344 ( 
.A(n_2323),
.B(n_251),
.C(n_248),
.D(n_249),
.Y(n_2344)
);

NAND4xp25_ASAP7_75t_L g2345 ( 
.A(n_2304),
.B(n_254),
.C(n_252),
.D(n_253),
.Y(n_2345)
);

NOR3x1_ASAP7_75t_L g2346 ( 
.A(n_2315),
.B(n_252),
.C(n_253),
.Y(n_2346)
);

NOR2xp33_ASAP7_75t_SL g2347 ( 
.A(n_2322),
.B(n_2060),
.Y(n_2347)
);

INVx1_ASAP7_75t_L g2348 ( 
.A(n_2303),
.Y(n_2348)
);

NOR2xp33_ASAP7_75t_L g2349 ( 
.A(n_2298),
.B(n_255),
.Y(n_2349)
);

NOR3x1_ASAP7_75t_L g2350 ( 
.A(n_2296),
.B(n_256),
.C(n_257),
.Y(n_2350)
);

AOI22xp5_ASAP7_75t_L g2351 ( 
.A1(n_2297),
.A2(n_2086),
.B1(n_2126),
.B2(n_2073),
.Y(n_2351)
);

AOI21xp5_ASAP7_75t_L g2352 ( 
.A1(n_2306),
.A2(n_256),
.B(n_257),
.Y(n_2352)
);

NAND3xp33_ASAP7_75t_L g2353 ( 
.A(n_2302),
.B(n_258),
.C(n_259),
.Y(n_2353)
);

NAND2xp5_ASAP7_75t_L g2354 ( 
.A(n_2294),
.B(n_258),
.Y(n_2354)
);

NAND2xp5_ASAP7_75t_L g2355 ( 
.A(n_2307),
.B(n_2300),
.Y(n_2355)
);

NAND2xp5_ASAP7_75t_L g2356 ( 
.A(n_2305),
.B(n_259),
.Y(n_2356)
);

NAND2xp5_ASAP7_75t_L g2357 ( 
.A(n_2314),
.B(n_260),
.Y(n_2357)
);

A2O1A1Ixp33_ASAP7_75t_L g2358 ( 
.A1(n_2311),
.A2(n_262),
.B(n_260),
.C(n_261),
.Y(n_2358)
);

NOR2x1p5_ASAP7_75t_SL g2359 ( 
.A(n_2312),
.B(n_262),
.Y(n_2359)
);

OAI21xp5_ASAP7_75t_L g2360 ( 
.A1(n_2287),
.A2(n_2019),
.B(n_1947),
.Y(n_2360)
);

NOR3xp33_ASAP7_75t_SL g2361 ( 
.A(n_2315),
.B(n_263),
.C(n_264),
.Y(n_2361)
);

NAND4xp25_ASAP7_75t_L g2362 ( 
.A(n_2346),
.B(n_267),
.C(n_265),
.D(n_266),
.Y(n_2362)
);

NOR2xp33_ASAP7_75t_L g2363 ( 
.A(n_2343),
.B(n_265),
.Y(n_2363)
);

NOR2xp67_ASAP7_75t_L g2364 ( 
.A(n_2324),
.B(n_266),
.Y(n_2364)
);

OAI211xp5_ASAP7_75t_L g2365 ( 
.A1(n_2329),
.A2(n_269),
.B(n_267),
.C(n_268),
.Y(n_2365)
);

OAI211xp5_ASAP7_75t_L g2366 ( 
.A1(n_2326),
.A2(n_272),
.B(n_268),
.C(n_271),
.Y(n_2366)
);

NOR3xp33_ASAP7_75t_L g2367 ( 
.A(n_2355),
.B(n_271),
.C(n_272),
.Y(n_2367)
);

NAND2xp5_ASAP7_75t_L g2368 ( 
.A(n_2344),
.B(n_273),
.Y(n_2368)
);

NOR2xp33_ASAP7_75t_L g2369 ( 
.A(n_2337),
.B(n_274),
.Y(n_2369)
);

NAND4xp75_ASAP7_75t_L g2370 ( 
.A(n_2350),
.B(n_276),
.C(n_274),
.D(n_275),
.Y(n_2370)
);

INVx1_ASAP7_75t_L g2371 ( 
.A(n_2333),
.Y(n_2371)
);

O2A1O1Ixp33_ASAP7_75t_L g2372 ( 
.A1(n_2327),
.A2(n_277),
.B(n_275),
.C(n_276),
.Y(n_2372)
);

NAND3xp33_ASAP7_75t_SL g2373 ( 
.A(n_2331),
.B(n_277),
.C(n_278),
.Y(n_2373)
);

NOR3xp33_ASAP7_75t_L g2374 ( 
.A(n_2334),
.B(n_278),
.C(n_279),
.Y(n_2374)
);

NOR4xp25_ASAP7_75t_L g2375 ( 
.A(n_2336),
.B(n_281),
.C(n_279),
.D(n_280),
.Y(n_2375)
);

NOR3xp33_ASAP7_75t_SL g2376 ( 
.A(n_2349),
.B(n_280),
.C(n_281),
.Y(n_2376)
);

NAND2xp5_ASAP7_75t_L g2377 ( 
.A(n_2328),
.B(n_282),
.Y(n_2377)
);

AOI211xp5_ASAP7_75t_SL g2378 ( 
.A1(n_2356),
.A2(n_284),
.B(n_282),
.C(n_283),
.Y(n_2378)
);

AND2x2_ASAP7_75t_L g2379 ( 
.A(n_2361),
.B(n_2101),
.Y(n_2379)
);

AO221x1_ASAP7_75t_L g2380 ( 
.A1(n_2338),
.A2(n_2126),
.B1(n_2021),
.B2(n_2027),
.C(n_2039),
.Y(n_2380)
);

NAND2xp5_ASAP7_75t_L g2381 ( 
.A(n_2358),
.B(n_284),
.Y(n_2381)
);

NAND3xp33_ASAP7_75t_L g2382 ( 
.A(n_2353),
.B(n_285),
.C(n_286),
.Y(n_2382)
);

NAND2xp5_ASAP7_75t_L g2383 ( 
.A(n_2352),
.B(n_285),
.Y(n_2383)
);

NOR3xp33_ASAP7_75t_L g2384 ( 
.A(n_2340),
.B(n_287),
.C(n_288),
.Y(n_2384)
);

NOR3xp33_ASAP7_75t_L g2385 ( 
.A(n_2339),
.B(n_2348),
.C(n_2342),
.Y(n_2385)
);

AO221x1_ASAP7_75t_L g2386 ( 
.A1(n_2359),
.A2(n_2126),
.B1(n_2021),
.B2(n_2027),
.C(n_2039),
.Y(n_2386)
);

NAND4xp25_ASAP7_75t_SL g2387 ( 
.A(n_2332),
.B(n_289),
.C(n_287),
.D(n_288),
.Y(n_2387)
);

NAND2xp5_ASAP7_75t_L g2388 ( 
.A(n_2354),
.B(n_289),
.Y(n_2388)
);

INVx1_ASAP7_75t_L g2389 ( 
.A(n_2335),
.Y(n_2389)
);

INVx1_ASAP7_75t_L g2390 ( 
.A(n_2325),
.Y(n_2390)
);

OAI211xp5_ASAP7_75t_L g2391 ( 
.A1(n_2345),
.A2(n_292),
.B(n_290),
.C(n_291),
.Y(n_2391)
);

AOI211x1_ASAP7_75t_L g2392 ( 
.A1(n_2330),
.A2(n_2357),
.B(n_2360),
.C(n_2341),
.Y(n_2392)
);

NAND4xp25_ASAP7_75t_L g2393 ( 
.A(n_2347),
.B(n_293),
.C(n_290),
.D(n_292),
.Y(n_2393)
);

OA211x2_ASAP7_75t_L g2394 ( 
.A1(n_2351),
.A2(n_295),
.B(n_293),
.C(n_294),
.Y(n_2394)
);

NAND4xp25_ASAP7_75t_L g2395 ( 
.A(n_2346),
.B(n_296),
.C(n_294),
.D(n_295),
.Y(n_2395)
);

AOI221x1_ASAP7_75t_L g2396 ( 
.A1(n_2331),
.A2(n_299),
.B1(n_296),
.B2(n_297),
.C(n_300),
.Y(n_2396)
);

NOR2xp33_ASAP7_75t_L g2397 ( 
.A(n_2343),
.B(n_299),
.Y(n_2397)
);

NAND3xp33_ASAP7_75t_L g2398 ( 
.A(n_2353),
.B(n_301),
.C(n_302),
.Y(n_2398)
);

AOI211xp5_ASAP7_75t_L g2399 ( 
.A1(n_2337),
.A2(n_304),
.B(n_302),
.C(n_303),
.Y(n_2399)
);

NAND3xp33_ASAP7_75t_L g2400 ( 
.A(n_2353),
.B(n_303),
.C(n_305),
.Y(n_2400)
);

NOR4xp25_ASAP7_75t_SL g2401 ( 
.A(n_2324),
.B(n_307),
.C(n_305),
.D(n_306),
.Y(n_2401)
);

NOR2xp67_ASAP7_75t_SL g2402 ( 
.A(n_2324),
.B(n_306),
.Y(n_2402)
);

NOR3xp33_ASAP7_75t_L g2403 ( 
.A(n_2355),
.B(n_307),
.C(n_308),
.Y(n_2403)
);

OAI321xp33_ASAP7_75t_L g2404 ( 
.A1(n_2355),
.A2(n_308),
.A3(n_309),
.B1(n_310),
.B2(n_311),
.C(n_312),
.Y(n_2404)
);

AOI22xp5_ASAP7_75t_L g2405 ( 
.A1(n_2347),
.A2(n_2126),
.B1(n_2123),
.B2(n_2071),
.Y(n_2405)
);

NAND3xp33_ASAP7_75t_L g2406 ( 
.A(n_2353),
.B(n_309),
.C(n_310),
.Y(n_2406)
);

NOR3xp33_ASAP7_75t_L g2407 ( 
.A(n_2355),
.B(n_311),
.C(n_312),
.Y(n_2407)
);

NOR2x1p5_ASAP7_75t_L g2408 ( 
.A(n_2337),
.B(n_313),
.Y(n_2408)
);

NAND5xp2_ASAP7_75t_L g2409 ( 
.A(n_2339),
.B(n_315),
.C(n_313),
.D(n_314),
.E(n_316),
.Y(n_2409)
);

AOI221xp5_ASAP7_75t_L g2410 ( 
.A1(n_2329),
.A2(n_317),
.B1(n_314),
.B2(n_315),
.C(n_318),
.Y(n_2410)
);

AOI221xp5_ASAP7_75t_L g2411 ( 
.A1(n_2329),
.A2(n_319),
.B1(n_317),
.B2(n_318),
.C(n_320),
.Y(n_2411)
);

OR2x2_ASAP7_75t_L g2412 ( 
.A(n_2326),
.B(n_321),
.Y(n_2412)
);

NOR2xp33_ASAP7_75t_L g2413 ( 
.A(n_2343),
.B(n_321),
.Y(n_2413)
);

NOR3xp33_ASAP7_75t_L g2414 ( 
.A(n_2355),
.B(n_322),
.C(n_323),
.Y(n_2414)
);

NOR2xp67_ASAP7_75t_L g2415 ( 
.A(n_2324),
.B(n_322),
.Y(n_2415)
);

NOR3xp33_ASAP7_75t_SL g2416 ( 
.A(n_2336),
.B(n_323),
.C(n_324),
.Y(n_2416)
);

NOR3xp33_ASAP7_75t_L g2417 ( 
.A(n_2355),
.B(n_324),
.C(n_325),
.Y(n_2417)
);

OAI211xp5_ASAP7_75t_L g2418 ( 
.A1(n_2329),
.A2(n_327),
.B(n_325),
.C(n_326),
.Y(n_2418)
);

NAND3xp33_ASAP7_75t_SL g2419 ( 
.A(n_2329),
.B(n_326),
.C(n_327),
.Y(n_2419)
);

OAI211xp5_ASAP7_75t_L g2420 ( 
.A1(n_2329),
.A2(n_330),
.B(n_328),
.C(n_329),
.Y(n_2420)
);

NOR3xp33_ASAP7_75t_L g2421 ( 
.A(n_2355),
.B(n_328),
.C(n_330),
.Y(n_2421)
);

NAND2xp5_ASAP7_75t_SL g2422 ( 
.A(n_2324),
.B(n_2123),
.Y(n_2422)
);

NAND5xp2_ASAP7_75t_L g2423 ( 
.A(n_2339),
.B(n_334),
.C(n_331),
.D(n_333),
.E(n_335),
.Y(n_2423)
);

OAI211xp5_ASAP7_75t_SL g2424 ( 
.A1(n_2416),
.A2(n_335),
.B(n_333),
.C(n_334),
.Y(n_2424)
);

BUFx6f_ASAP7_75t_L g2425 ( 
.A(n_2390),
.Y(n_2425)
);

INVx1_ASAP7_75t_L g2426 ( 
.A(n_2402),
.Y(n_2426)
);

INVx1_ASAP7_75t_L g2427 ( 
.A(n_2364),
.Y(n_2427)
);

INVx1_ASAP7_75t_L g2428 ( 
.A(n_2415),
.Y(n_2428)
);

NAND2xp5_ASAP7_75t_L g2429 ( 
.A(n_2378),
.B(n_336),
.Y(n_2429)
);

NOR3xp33_ASAP7_75t_L g2430 ( 
.A(n_2377),
.B(n_336),
.C(n_338),
.Y(n_2430)
);

NAND2xp33_ASAP7_75t_SL g2431 ( 
.A(n_2401),
.B(n_338),
.Y(n_2431)
);

NOR2xp33_ASAP7_75t_R g2432 ( 
.A(n_2419),
.B(n_339),
.Y(n_2432)
);

XOR2x2_ASAP7_75t_L g2433 ( 
.A(n_2370),
.B(n_339),
.Y(n_2433)
);

AOI211xp5_ASAP7_75t_SL g2434 ( 
.A1(n_2369),
.A2(n_342),
.B(n_340),
.C(n_341),
.Y(n_2434)
);

AOI22xp5_ASAP7_75t_L g2435 ( 
.A1(n_2363),
.A2(n_2056),
.B1(n_2149),
.B2(n_2066),
.Y(n_2435)
);

INVx2_ASAP7_75t_SL g2436 ( 
.A(n_2386),
.Y(n_2436)
);

HB1xp67_ASAP7_75t_L g2437 ( 
.A(n_2394),
.Y(n_2437)
);

AOI211xp5_ASAP7_75t_SL g2438 ( 
.A1(n_2365),
.A2(n_342),
.B(n_340),
.C(n_341),
.Y(n_2438)
);

NOR2xp33_ASAP7_75t_R g2439 ( 
.A(n_2373),
.B(n_343),
.Y(n_2439)
);

NAND2xp5_ASAP7_75t_L g2440 ( 
.A(n_2397),
.B(n_343),
.Y(n_2440)
);

INVx1_ASAP7_75t_L g2441 ( 
.A(n_2368),
.Y(n_2441)
);

NAND2xp5_ASAP7_75t_L g2442 ( 
.A(n_2413),
.B(n_344),
.Y(n_2442)
);

OAI211xp5_ASAP7_75t_L g2443 ( 
.A1(n_2410),
.A2(n_347),
.B(n_345),
.C(n_346),
.Y(n_2443)
);

AOI21xp33_ASAP7_75t_SL g2444 ( 
.A1(n_2372),
.A2(n_345),
.B(n_346),
.Y(n_2444)
);

OAI221xp5_ASAP7_75t_SL g2445 ( 
.A1(n_2375),
.A2(n_2040),
.B1(n_349),
.B2(n_347),
.C(n_348),
.Y(n_2445)
);

NAND2xp33_ASAP7_75t_R g2446 ( 
.A(n_2376),
.B(n_348),
.Y(n_2446)
);

OAI211xp5_ASAP7_75t_L g2447 ( 
.A1(n_2411),
.A2(n_351),
.B(n_349),
.C(n_350),
.Y(n_2447)
);

INVx1_ASAP7_75t_SL g2448 ( 
.A(n_2412),
.Y(n_2448)
);

INVx1_ASAP7_75t_SL g2449 ( 
.A(n_2381),
.Y(n_2449)
);

AOI21xp5_ASAP7_75t_L g2450 ( 
.A1(n_2383),
.A2(n_350),
.B(n_352),
.Y(n_2450)
);

NAND2xp5_ASAP7_75t_SL g2451 ( 
.A(n_2399),
.B(n_2149),
.Y(n_2451)
);

NAND4xp75_ASAP7_75t_L g2452 ( 
.A(n_2396),
.B(n_354),
.C(n_352),
.D(n_353),
.Y(n_2452)
);

INVx1_ASAP7_75t_SL g2453 ( 
.A(n_2388),
.Y(n_2453)
);

O2A1O1Ixp33_ASAP7_75t_L g2454 ( 
.A1(n_2367),
.A2(n_2403),
.B(n_2414),
.C(n_2407),
.Y(n_2454)
);

HB1xp67_ASAP7_75t_L g2455 ( 
.A(n_2387),
.Y(n_2455)
);

NOR2xp33_ASAP7_75t_L g2456 ( 
.A(n_2409),
.B(n_353),
.Y(n_2456)
);

AOI22xp5_ASAP7_75t_L g2457 ( 
.A1(n_2379),
.A2(n_2149),
.B1(n_2066),
.B2(n_2022),
.Y(n_2457)
);

NAND2xp5_ASAP7_75t_L g2458 ( 
.A(n_2417),
.B(n_354),
.Y(n_2458)
);

NAND2xp33_ASAP7_75t_SL g2459 ( 
.A(n_2408),
.B(n_355),
.Y(n_2459)
);

AOI221xp5_ASAP7_75t_L g2460 ( 
.A1(n_2362),
.A2(n_355),
.B1(n_356),
.B2(n_357),
.C(n_358),
.Y(n_2460)
);

INVx1_ASAP7_75t_SL g2461 ( 
.A(n_2422),
.Y(n_2461)
);

CKINVDCx16_ASAP7_75t_R g2462 ( 
.A(n_2389),
.Y(n_2462)
);

A2O1A1Ixp33_ASAP7_75t_SL g2463 ( 
.A1(n_2385),
.A2(n_359),
.B(n_357),
.C(n_358),
.Y(n_2463)
);

OAI322xp33_ASAP7_75t_L g2464 ( 
.A1(n_2371),
.A2(n_360),
.A3(n_361),
.B1(n_362),
.B2(n_363),
.C1(n_364),
.C2(n_365),
.Y(n_2464)
);

INVx1_ASAP7_75t_L g2465 ( 
.A(n_2423),
.Y(n_2465)
);

XNOR2xp5_ASAP7_75t_L g2466 ( 
.A(n_2395),
.B(n_360),
.Y(n_2466)
);

INVx1_ASAP7_75t_SL g2467 ( 
.A(n_2382),
.Y(n_2467)
);

AOI21xp5_ASAP7_75t_L g2468 ( 
.A1(n_2418),
.A2(n_2420),
.B(n_2391),
.Y(n_2468)
);

AO22x2_ASAP7_75t_L g2469 ( 
.A1(n_2384),
.A2(n_2398),
.B1(n_2406),
.B2(n_2400),
.Y(n_2469)
);

AOI21xp5_ASAP7_75t_L g2470 ( 
.A1(n_2393),
.A2(n_362),
.B(n_363),
.Y(n_2470)
);

INVx1_ASAP7_75t_L g2471 ( 
.A(n_2366),
.Y(n_2471)
);

AOI221xp5_ASAP7_75t_L g2472 ( 
.A1(n_2392),
.A2(n_364),
.B1(n_365),
.B2(n_366),
.C(n_367),
.Y(n_2472)
);

NAND2xp33_ASAP7_75t_SL g2473 ( 
.A(n_2404),
.B(n_367),
.Y(n_2473)
);

A2O1A1Ixp33_ASAP7_75t_SL g2474 ( 
.A1(n_2421),
.A2(n_370),
.B(n_368),
.C(n_369),
.Y(n_2474)
);

BUFx2_ASAP7_75t_L g2475 ( 
.A(n_2405),
.Y(n_2475)
);

NAND2xp5_ASAP7_75t_SL g2476 ( 
.A(n_2374),
.B(n_368),
.Y(n_2476)
);

OR2x2_ASAP7_75t_L g2477 ( 
.A(n_2380),
.B(n_369),
.Y(n_2477)
);

INVx2_ASAP7_75t_SL g2478 ( 
.A(n_2404),
.Y(n_2478)
);

NAND2xp33_ASAP7_75t_R g2479 ( 
.A(n_2401),
.B(n_370),
.Y(n_2479)
);

INVx1_ASAP7_75t_L g2480 ( 
.A(n_2402),
.Y(n_2480)
);

OAI22xp5_ASAP7_75t_L g2481 ( 
.A1(n_2405),
.A2(n_2040),
.B1(n_2022),
.B2(n_2129),
.Y(n_2481)
);

NOR4xp25_ASAP7_75t_L g2482 ( 
.A(n_2419),
.B(n_373),
.C(n_371),
.D(n_372),
.Y(n_2482)
);

XOR2x2_ASAP7_75t_L g2483 ( 
.A(n_2370),
.B(n_371),
.Y(n_2483)
);

INVx1_ASAP7_75t_L g2484 ( 
.A(n_2402),
.Y(n_2484)
);

AOI221xp5_ASAP7_75t_L g2485 ( 
.A1(n_2375),
.A2(n_372),
.B1(n_373),
.B2(n_374),
.C(n_375),
.Y(n_2485)
);

OAI221xp5_ASAP7_75t_L g2486 ( 
.A1(n_2410),
.A2(n_375),
.B1(n_376),
.B2(n_377),
.C(n_378),
.Y(n_2486)
);

BUFx6f_ASAP7_75t_L g2487 ( 
.A(n_2390),
.Y(n_2487)
);

OAI221xp5_ASAP7_75t_L g2488 ( 
.A1(n_2410),
.A2(n_376),
.B1(n_381),
.B2(n_382),
.C(n_383),
.Y(n_2488)
);

INVx1_ASAP7_75t_SL g2489 ( 
.A(n_2370),
.Y(n_2489)
);

AOI22xp5_ASAP7_75t_L g2490 ( 
.A1(n_2363),
.A2(n_2101),
.B1(n_2118),
.B2(n_2129),
.Y(n_2490)
);

NAND2xp5_ASAP7_75t_SL g2491 ( 
.A(n_2425),
.B(n_381),
.Y(n_2491)
);

INVx1_ASAP7_75t_L g2492 ( 
.A(n_2433),
.Y(n_2492)
);

INVx1_ASAP7_75t_L g2493 ( 
.A(n_2483),
.Y(n_2493)
);

INVx1_ASAP7_75t_L g2494 ( 
.A(n_2452),
.Y(n_2494)
);

NAND2xp5_ASAP7_75t_L g2495 ( 
.A(n_2438),
.B(n_382),
.Y(n_2495)
);

NAND3xp33_ASAP7_75t_L g2496 ( 
.A(n_2434),
.B(n_384),
.C(n_385),
.Y(n_2496)
);

INVx1_ASAP7_75t_L g2497 ( 
.A(n_2437),
.Y(n_2497)
);

NAND2xp5_ASAP7_75t_L g2498 ( 
.A(n_2456),
.B(n_385),
.Y(n_2498)
);

NOR2xp67_ASAP7_75t_L g2499 ( 
.A(n_2444),
.B(n_386),
.Y(n_2499)
);

CKINVDCx14_ASAP7_75t_R g2500 ( 
.A(n_2431),
.Y(n_2500)
);

INVx2_ASAP7_75t_L g2501 ( 
.A(n_2477),
.Y(n_2501)
);

INVxp67_ASAP7_75t_L g2502 ( 
.A(n_2479),
.Y(n_2502)
);

BUFx12f_ASAP7_75t_L g2503 ( 
.A(n_2425),
.Y(n_2503)
);

NAND4xp75_ASAP7_75t_L g2504 ( 
.A(n_2440),
.B(n_390),
.C(n_387),
.D(n_388),
.Y(n_2504)
);

INVxp67_ASAP7_75t_L g2505 ( 
.A(n_2429),
.Y(n_2505)
);

AND2x4_ASAP7_75t_L g2506 ( 
.A(n_2427),
.B(n_391),
.Y(n_2506)
);

O2A1O1Ixp33_ASAP7_75t_L g2507 ( 
.A1(n_2463),
.A2(n_2474),
.B(n_2478),
.C(n_2442),
.Y(n_2507)
);

INVx1_ASAP7_75t_L g2508 ( 
.A(n_2466),
.Y(n_2508)
);

NAND4xp75_ASAP7_75t_L g2509 ( 
.A(n_2426),
.B(n_393),
.C(n_391),
.D(n_392),
.Y(n_2509)
);

AO22x2_ASAP7_75t_L g2510 ( 
.A1(n_2489),
.A2(n_396),
.B1(n_394),
.B2(n_395),
.Y(n_2510)
);

NAND4xp75_ASAP7_75t_L g2511 ( 
.A(n_2480),
.B(n_397),
.C(n_394),
.D(n_396),
.Y(n_2511)
);

AOI22xp5_ASAP7_75t_L g2512 ( 
.A1(n_2446),
.A2(n_2118),
.B1(n_2134),
.B2(n_2129),
.Y(n_2512)
);

NOR2x1_ASAP7_75t_L g2513 ( 
.A(n_2428),
.B(n_398),
.Y(n_2513)
);

NAND2xp5_ASAP7_75t_L g2514 ( 
.A(n_2482),
.B(n_398),
.Y(n_2514)
);

HB1xp67_ASAP7_75t_L g2515 ( 
.A(n_2425),
.Y(n_2515)
);

INVx1_ASAP7_75t_L g2516 ( 
.A(n_2455),
.Y(n_2516)
);

NOR4xp75_ASAP7_75t_L g2517 ( 
.A(n_2476),
.B(n_401),
.C(n_399),
.D(n_400),
.Y(n_2517)
);

XOR2xp5_ASAP7_75t_L g2518 ( 
.A(n_2465),
.B(n_399),
.Y(n_2518)
);

INVx1_ASAP7_75t_L g2519 ( 
.A(n_2458),
.Y(n_2519)
);

HB1xp67_ASAP7_75t_L g2520 ( 
.A(n_2487),
.Y(n_2520)
);

NOR2x1_ASAP7_75t_L g2521 ( 
.A(n_2484),
.B(n_401),
.Y(n_2521)
);

INVx1_ASAP7_75t_L g2522 ( 
.A(n_2487),
.Y(n_2522)
);

NOR2x1_ASAP7_75t_L g2523 ( 
.A(n_2464),
.B(n_402),
.Y(n_2523)
);

OR2x2_ASAP7_75t_L g2524 ( 
.A(n_2445),
.B(n_402),
.Y(n_2524)
);

NOR2x1_ASAP7_75t_L g2525 ( 
.A(n_2471),
.B(n_404),
.Y(n_2525)
);

INVxp67_ASAP7_75t_L g2526 ( 
.A(n_2473),
.Y(n_2526)
);

INVx2_ASAP7_75t_L g2527 ( 
.A(n_2487),
.Y(n_2527)
);

INVx1_ASAP7_75t_L g2528 ( 
.A(n_2469),
.Y(n_2528)
);

A2O1A1Ixp33_ASAP7_75t_L g2529 ( 
.A1(n_2470),
.A2(n_406),
.B(n_404),
.C(n_405),
.Y(n_2529)
);

NOR2x1_ASAP7_75t_L g2530 ( 
.A(n_2424),
.B(n_2450),
.Y(n_2530)
);

OR2x2_ASAP7_75t_L g2531 ( 
.A(n_2461),
.B(n_405),
.Y(n_2531)
);

INVx1_ASAP7_75t_L g2532 ( 
.A(n_2469),
.Y(n_2532)
);

OAI221xp5_ASAP7_75t_L g2533 ( 
.A1(n_2485),
.A2(n_406),
.B1(n_407),
.B2(n_408),
.C(n_409),
.Y(n_2533)
);

AOI22xp33_ASAP7_75t_L g2534 ( 
.A1(n_2436),
.A2(n_2134),
.B1(n_2098),
.B2(n_2088),
.Y(n_2534)
);

NOR2x1_ASAP7_75t_L g2535 ( 
.A(n_2443),
.B(n_408),
.Y(n_2535)
);

INVx2_ASAP7_75t_L g2536 ( 
.A(n_2441),
.Y(n_2536)
);

INVx1_ASAP7_75t_L g2537 ( 
.A(n_2430),
.Y(n_2537)
);

INVx1_ASAP7_75t_L g2538 ( 
.A(n_2447),
.Y(n_2538)
);

INVxp67_ASAP7_75t_L g2539 ( 
.A(n_2459),
.Y(n_2539)
);

NOR2xp33_ASAP7_75t_L g2540 ( 
.A(n_2486),
.B(n_409),
.Y(n_2540)
);

INVxp67_ASAP7_75t_SL g2541 ( 
.A(n_2454),
.Y(n_2541)
);

NOR2x1_ASAP7_75t_L g2542 ( 
.A(n_2448),
.B(n_410),
.Y(n_2542)
);

AOI22xp33_ASAP7_75t_SL g2543 ( 
.A1(n_2462),
.A2(n_411),
.B1(n_412),
.B2(n_413),
.Y(n_2543)
);

NAND2xp5_ASAP7_75t_L g2544 ( 
.A(n_2472),
.B(n_411),
.Y(n_2544)
);

INVx1_ASAP7_75t_L g2545 ( 
.A(n_2475),
.Y(n_2545)
);

INVx2_ASAP7_75t_L g2546 ( 
.A(n_2453),
.Y(n_2546)
);

NAND2x1p5_ASAP7_75t_L g2547 ( 
.A(n_2467),
.B(n_412),
.Y(n_2547)
);

AND2x2_ASAP7_75t_L g2548 ( 
.A(n_2460),
.B(n_2140),
.Y(n_2548)
);

INVx2_ASAP7_75t_L g2549 ( 
.A(n_2449),
.Y(n_2549)
);

NAND4xp75_ASAP7_75t_L g2550 ( 
.A(n_2468),
.B(n_413),
.C(n_414),
.D(n_415),
.Y(n_2550)
);

AND2x4_ASAP7_75t_L g2551 ( 
.A(n_2490),
.B(n_414),
.Y(n_2551)
);

AND2x2_ASAP7_75t_L g2552 ( 
.A(n_2432),
.B(n_2147),
.Y(n_2552)
);

OR2x2_ASAP7_75t_L g2553 ( 
.A(n_2451),
.B(n_415),
.Y(n_2553)
);

NOR3xp33_ASAP7_75t_L g2554 ( 
.A(n_2497),
.B(n_2488),
.C(n_2439),
.Y(n_2554)
);

AND2x2_ASAP7_75t_L g2555 ( 
.A(n_2502),
.B(n_2435),
.Y(n_2555)
);

XNOR2xp5_ASAP7_75t_L g2556 ( 
.A(n_2518),
.B(n_2457),
.Y(n_2556)
);

AND3x4_ASAP7_75t_L g2557 ( 
.A(n_2517),
.B(n_2481),
.C(n_416),
.Y(n_2557)
);

INVx2_ASAP7_75t_L g2558 ( 
.A(n_2510),
.Y(n_2558)
);

NOR4xp25_ASAP7_75t_L g2559 ( 
.A(n_2507),
.B(n_416),
.C(n_417),
.D(n_419),
.Y(n_2559)
);

NOR2xp33_ASAP7_75t_L g2560 ( 
.A(n_2531),
.B(n_417),
.Y(n_2560)
);

NOR3xp33_ASAP7_75t_SL g2561 ( 
.A(n_2498),
.B(n_420),
.C(n_421),
.Y(n_2561)
);

INVx1_ASAP7_75t_L g2562 ( 
.A(n_2542),
.Y(n_2562)
);

NAND4xp75_ASAP7_75t_L g2563 ( 
.A(n_2525),
.B(n_421),
.C(n_422),
.D(n_423),
.Y(n_2563)
);

NAND3xp33_ASAP7_75t_SL g2564 ( 
.A(n_2547),
.B(n_424),
.C(n_425),
.Y(n_2564)
);

OR2x2_ASAP7_75t_L g2565 ( 
.A(n_2514),
.B(n_425),
.Y(n_2565)
);

INVx3_ASAP7_75t_L g2566 ( 
.A(n_2503),
.Y(n_2566)
);

NOR3xp33_ASAP7_75t_SL g2567 ( 
.A(n_2545),
.B(n_426),
.C(n_427),
.Y(n_2567)
);

NOR3xp33_ASAP7_75t_L g2568 ( 
.A(n_2500),
.B(n_427),
.C(n_428),
.Y(n_2568)
);

NOR4xp25_ASAP7_75t_L g2569 ( 
.A(n_2522),
.B(n_428),
.C(n_429),
.D(n_430),
.Y(n_2569)
);

NOR4xp75_ASAP7_75t_L g2570 ( 
.A(n_2495),
.B(n_429),
.C(n_430),
.D(n_431),
.Y(n_2570)
);

INVx1_ASAP7_75t_L g2571 ( 
.A(n_2521),
.Y(n_2571)
);

AO22x2_ASAP7_75t_L g2572 ( 
.A1(n_2494),
.A2(n_431),
.B1(n_432),
.B2(n_433),
.Y(n_2572)
);

AOI21xp5_ASAP7_75t_L g2573 ( 
.A1(n_2515),
.A2(n_432),
.B(n_434),
.Y(n_2573)
);

NOR3xp33_ASAP7_75t_SL g2574 ( 
.A(n_2496),
.B(n_2516),
.C(n_2528),
.Y(n_2574)
);

NAND2xp5_ASAP7_75t_L g2575 ( 
.A(n_2513),
.B(n_434),
.Y(n_2575)
);

INVx1_ASAP7_75t_L g2576 ( 
.A(n_2520),
.Y(n_2576)
);

OAI22xp5_ASAP7_75t_L g2577 ( 
.A1(n_2526),
.A2(n_2147),
.B1(n_1916),
.B2(n_2092),
.Y(n_2577)
);

NAND4xp75_ASAP7_75t_L g2578 ( 
.A(n_2532),
.B(n_435),
.C(n_439),
.D(n_440),
.Y(n_2578)
);

NOR3xp33_ASAP7_75t_L g2579 ( 
.A(n_2527),
.B(n_439),
.C(n_440),
.Y(n_2579)
);

NAND2xp5_ASAP7_75t_L g2580 ( 
.A(n_2499),
.B(n_441),
.Y(n_2580)
);

NOR3xp33_ASAP7_75t_L g2581 ( 
.A(n_2539),
.B(n_442),
.C(n_443),
.Y(n_2581)
);

NAND4xp75_ASAP7_75t_L g2582 ( 
.A(n_2523),
.B(n_443),
.C(n_444),
.D(n_445),
.Y(n_2582)
);

NAND4xp25_ASAP7_75t_L g2583 ( 
.A(n_2540),
.B(n_445),
.C(n_446),
.D(n_447),
.Y(n_2583)
);

INVx2_ASAP7_75t_SL g2584 ( 
.A(n_2506),
.Y(n_2584)
);

OR2x2_ASAP7_75t_L g2585 ( 
.A(n_2524),
.B(n_446),
.Y(n_2585)
);

NOR3xp33_ASAP7_75t_L g2586 ( 
.A(n_2541),
.B(n_447),
.C(n_448),
.Y(n_2586)
);

NOR3xp33_ASAP7_75t_SL g2587 ( 
.A(n_2538),
.B(n_448),
.C(n_449),
.Y(n_2587)
);

AND4x1_ASAP7_75t_L g2588 ( 
.A(n_2530),
.B(n_450),
.C(n_451),
.D(n_452),
.Y(n_2588)
);

NOR2x1_ASAP7_75t_L g2589 ( 
.A(n_2550),
.B(n_450),
.Y(n_2589)
);

NAND4xp25_ASAP7_75t_L g2590 ( 
.A(n_2544),
.B(n_451),
.C(n_452),
.D(n_453),
.Y(n_2590)
);

NOR3xp33_ASAP7_75t_L g2591 ( 
.A(n_2546),
.B(n_453),
.C(n_454),
.Y(n_2591)
);

NAND3xp33_ASAP7_75t_SL g2592 ( 
.A(n_2529),
.B(n_455),
.C(n_456),
.Y(n_2592)
);

NAND2xp5_ASAP7_75t_L g2593 ( 
.A(n_2543),
.B(n_455),
.Y(n_2593)
);

OR2x2_ASAP7_75t_L g2594 ( 
.A(n_2553),
.B(n_456),
.Y(n_2594)
);

AND2x2_ASAP7_75t_L g2595 ( 
.A(n_2501),
.B(n_2147),
.Y(n_2595)
);

NOR3xp33_ASAP7_75t_SL g2596 ( 
.A(n_2533),
.B(n_457),
.C(n_458),
.Y(n_2596)
);

BUFx4f_ASAP7_75t_SL g2597 ( 
.A(n_2549),
.Y(n_2597)
);

NOR3xp33_ASAP7_75t_L g2598 ( 
.A(n_2536),
.B(n_459),
.C(n_460),
.Y(n_2598)
);

CKINVDCx16_ASAP7_75t_R g2599 ( 
.A(n_2585),
.Y(n_2599)
);

HB1xp67_ASAP7_75t_L g2600 ( 
.A(n_2588),
.Y(n_2600)
);

BUFx2_ASAP7_75t_L g2601 ( 
.A(n_2567),
.Y(n_2601)
);

BUFx6f_ASAP7_75t_L g2602 ( 
.A(n_2584),
.Y(n_2602)
);

CKINVDCx5p33_ASAP7_75t_R g2603 ( 
.A(n_2574),
.Y(n_2603)
);

INVx1_ASAP7_75t_L g2604 ( 
.A(n_2575),
.Y(n_2604)
);

INVx1_ASAP7_75t_SL g2605 ( 
.A(n_2570),
.Y(n_2605)
);

BUFx6f_ASAP7_75t_L g2606 ( 
.A(n_2566),
.Y(n_2606)
);

AOI21xp5_ASAP7_75t_L g2607 ( 
.A1(n_2580),
.A2(n_2535),
.B(n_2505),
.Y(n_2607)
);

HB1xp67_ASAP7_75t_L g2608 ( 
.A(n_2578),
.Y(n_2608)
);

HB1xp67_ASAP7_75t_L g2609 ( 
.A(n_2563),
.Y(n_2609)
);

BUFx2_ASAP7_75t_L g2610 ( 
.A(n_2561),
.Y(n_2610)
);

XOR2xp5_ASAP7_75t_L g2611 ( 
.A(n_2582),
.B(n_2504),
.Y(n_2611)
);

HB1xp67_ASAP7_75t_L g2612 ( 
.A(n_2558),
.Y(n_2612)
);

NOR2xp33_ASAP7_75t_R g2613 ( 
.A(n_2564),
.B(n_2537),
.Y(n_2613)
);

AOI22xp5_ASAP7_75t_L g2614 ( 
.A1(n_2576),
.A2(n_2492),
.B1(n_2493),
.B2(n_2551),
.Y(n_2614)
);

INVx1_ASAP7_75t_L g2615 ( 
.A(n_2594),
.Y(n_2615)
);

AOI22xp5_ASAP7_75t_L g2616 ( 
.A1(n_2597),
.A2(n_2551),
.B1(n_2508),
.B2(n_2552),
.Y(n_2616)
);

INVx2_ASAP7_75t_L g2617 ( 
.A(n_2572),
.Y(n_2617)
);

INVxp67_ASAP7_75t_SL g2618 ( 
.A(n_2589),
.Y(n_2618)
);

CKINVDCx20_ASAP7_75t_R g2619 ( 
.A(n_2556),
.Y(n_2619)
);

INVx1_ASAP7_75t_SL g2620 ( 
.A(n_2565),
.Y(n_2620)
);

NAND2xp5_ASAP7_75t_L g2621 ( 
.A(n_2568),
.B(n_2491),
.Y(n_2621)
);

OAI21xp33_ASAP7_75t_L g2622 ( 
.A1(n_2566),
.A2(n_2519),
.B(n_2548),
.Y(n_2622)
);

CKINVDCx5p33_ASAP7_75t_R g2623 ( 
.A(n_2562),
.Y(n_2623)
);

BUFx6f_ASAP7_75t_L g2624 ( 
.A(n_2571),
.Y(n_2624)
);

NOR2xp33_ASAP7_75t_R g2625 ( 
.A(n_2592),
.B(n_2506),
.Y(n_2625)
);

HB1xp67_ASAP7_75t_L g2626 ( 
.A(n_2569),
.Y(n_2626)
);

INVx1_ASAP7_75t_L g2627 ( 
.A(n_2593),
.Y(n_2627)
);

NOR2xp33_ASAP7_75t_R g2628 ( 
.A(n_2560),
.B(n_2509),
.Y(n_2628)
);

CKINVDCx5p33_ASAP7_75t_R g2629 ( 
.A(n_2555),
.Y(n_2629)
);

INVx1_ASAP7_75t_SL g2630 ( 
.A(n_2572),
.Y(n_2630)
);

NAND2xp33_ASAP7_75t_SL g2631 ( 
.A(n_2587),
.B(n_2510),
.Y(n_2631)
);

NAND2xp5_ASAP7_75t_L g2632 ( 
.A(n_2559),
.B(n_2586),
.Y(n_2632)
);

CKINVDCx5p33_ASAP7_75t_R g2633 ( 
.A(n_2596),
.Y(n_2633)
);

INVxp67_ASAP7_75t_L g2634 ( 
.A(n_2626),
.Y(n_2634)
);

OAI32xp33_ASAP7_75t_L g2635 ( 
.A1(n_2612),
.A2(n_2554),
.A3(n_2590),
.B1(n_2583),
.B2(n_2591),
.Y(n_2635)
);

AOI322xp5_ASAP7_75t_L g2636 ( 
.A1(n_2631),
.A2(n_2605),
.A3(n_2618),
.B1(n_2622),
.B2(n_2608),
.C1(n_2609),
.C2(n_2619),
.Y(n_2636)
);

NAND3xp33_ASAP7_75t_L g2637 ( 
.A(n_2606),
.B(n_2598),
.C(n_2579),
.Y(n_2637)
);

AOI322xp5_ASAP7_75t_L g2638 ( 
.A1(n_2600),
.A2(n_2595),
.A3(n_2581),
.B1(n_2534),
.B2(n_2557),
.C1(n_2512),
.C2(n_2573),
.Y(n_2638)
);

AOI322xp5_ASAP7_75t_L g2639 ( 
.A1(n_2630),
.A2(n_2511),
.A3(n_2577),
.B1(n_461),
.B2(n_462),
.C1(n_463),
.C2(n_464),
.Y(n_2639)
);

OAI221xp5_ASAP7_75t_L g2640 ( 
.A1(n_2614),
.A2(n_459),
.B1(n_460),
.B2(n_462),
.C(n_463),
.Y(n_2640)
);

NOR2xp33_ASAP7_75t_L g2641 ( 
.A(n_2602),
.B(n_464),
.Y(n_2641)
);

NAND2xp5_ASAP7_75t_L g2642 ( 
.A(n_2617),
.B(n_465),
.Y(n_2642)
);

AOI322xp5_ASAP7_75t_L g2643 ( 
.A1(n_2603),
.A2(n_465),
.A3(n_466),
.B1(n_467),
.B2(n_468),
.C1(n_469),
.C2(n_470),
.Y(n_2643)
);

AOI322xp5_ASAP7_75t_L g2644 ( 
.A1(n_2620),
.A2(n_466),
.A3(n_467),
.B1(n_469),
.B2(n_471),
.C1(n_472),
.C2(n_473),
.Y(n_2644)
);

AOI221xp5_ASAP7_75t_L g2645 ( 
.A1(n_2606),
.A2(n_471),
.B1(n_472),
.B2(n_473),
.C(n_474),
.Y(n_2645)
);

AOI22x1_ASAP7_75t_L g2646 ( 
.A1(n_2629),
.A2(n_475),
.B1(n_476),
.B2(n_477),
.Y(n_2646)
);

AOI322xp5_ASAP7_75t_L g2647 ( 
.A1(n_2632),
.A2(n_475),
.A3(n_476),
.B1(n_478),
.B2(n_479),
.C1(n_480),
.C2(n_481),
.Y(n_2647)
);

INVx1_ASAP7_75t_L g2648 ( 
.A(n_2611),
.Y(n_2648)
);

OAI22xp5_ASAP7_75t_L g2649 ( 
.A1(n_2623),
.A2(n_478),
.B1(n_480),
.B2(n_481),
.Y(n_2649)
);

A2O1A1Ixp33_ASAP7_75t_L g2650 ( 
.A1(n_2607),
.A2(n_482),
.B(n_483),
.C(n_484),
.Y(n_2650)
);

AO22x2_ASAP7_75t_L g2651 ( 
.A1(n_2615),
.A2(n_2627),
.B1(n_2604),
.B2(n_2621),
.Y(n_2651)
);

AOI221xp5_ASAP7_75t_L g2652 ( 
.A1(n_2602),
.A2(n_482),
.B1(n_483),
.B2(n_484),
.C(n_485),
.Y(n_2652)
);

INVx2_ASAP7_75t_L g2653 ( 
.A(n_2624),
.Y(n_2653)
);

AOI322xp5_ASAP7_75t_L g2654 ( 
.A1(n_2601),
.A2(n_2610),
.A3(n_2599),
.B1(n_2616),
.B2(n_2633),
.C1(n_2624),
.C2(n_2613),
.Y(n_2654)
);

OR2x2_ASAP7_75t_L g2655 ( 
.A(n_2624),
.B(n_486),
.Y(n_2655)
);

AOI22xp5_ASAP7_75t_L g2656 ( 
.A1(n_2628),
.A2(n_2625),
.B1(n_488),
.B2(n_491),
.Y(n_2656)
);

NOR2xp67_ASAP7_75t_L g2657 ( 
.A(n_2617),
.B(n_487),
.Y(n_2657)
);

OAI322xp33_ASAP7_75t_L g2658 ( 
.A1(n_2630),
.A2(n_487),
.A3(n_491),
.B1(n_492),
.B2(n_493),
.C1(n_494),
.C2(n_495),
.Y(n_2658)
);

INVx1_ASAP7_75t_L g2659 ( 
.A(n_2626),
.Y(n_2659)
);

AOI22xp5_ASAP7_75t_L g2660 ( 
.A1(n_2634),
.A2(n_492),
.B1(n_494),
.B2(n_495),
.Y(n_2660)
);

OAI22xp5_ASAP7_75t_L g2661 ( 
.A1(n_2659),
.A2(n_496),
.B1(n_497),
.B2(n_498),
.Y(n_2661)
);

INVx1_ASAP7_75t_L g2662 ( 
.A(n_2657),
.Y(n_2662)
);

OAI22xp5_ASAP7_75t_L g2663 ( 
.A1(n_2653),
.A2(n_496),
.B1(n_499),
.B2(n_500),
.Y(n_2663)
);

INVx1_ASAP7_75t_L g2664 ( 
.A(n_2655),
.Y(n_2664)
);

OAI22xp5_ASAP7_75t_L g2665 ( 
.A1(n_2637),
.A2(n_499),
.B1(n_500),
.B2(n_501),
.Y(n_2665)
);

OAI22xp5_ASAP7_75t_L g2666 ( 
.A1(n_2656),
.A2(n_501),
.B1(n_502),
.B2(n_503),
.Y(n_2666)
);

OAI22x1_ASAP7_75t_L g2667 ( 
.A1(n_2646),
.A2(n_502),
.B1(n_503),
.B2(n_504),
.Y(n_2667)
);

AOI221xp5_ASAP7_75t_SL g2668 ( 
.A1(n_2635),
.A2(n_2648),
.B1(n_2640),
.B2(n_2658),
.C(n_2650),
.Y(n_2668)
);

AOI22xp5_ASAP7_75t_L g2669 ( 
.A1(n_2651),
.A2(n_504),
.B1(n_505),
.B2(n_506),
.Y(n_2669)
);

AOI22xp5_ASAP7_75t_L g2670 ( 
.A1(n_2651),
.A2(n_505),
.B1(n_506),
.B2(n_507),
.Y(n_2670)
);

AO22x2_ASAP7_75t_L g2671 ( 
.A1(n_2636),
.A2(n_507),
.B1(n_508),
.B2(n_509),
.Y(n_2671)
);

OAI22xp5_ASAP7_75t_SL g2672 ( 
.A1(n_2641),
.A2(n_509),
.B1(n_510),
.B2(n_512),
.Y(n_2672)
);

INVx1_ASAP7_75t_L g2673 ( 
.A(n_2642),
.Y(n_2673)
);

INVx1_ASAP7_75t_L g2674 ( 
.A(n_2649),
.Y(n_2674)
);

INVx1_ASAP7_75t_L g2675 ( 
.A(n_2652),
.Y(n_2675)
);

INVx1_ASAP7_75t_L g2676 ( 
.A(n_2645),
.Y(n_2676)
);

INVxp33_ASAP7_75t_SL g2677 ( 
.A(n_2664),
.Y(n_2677)
);

NAND5xp2_ASAP7_75t_L g2678 ( 
.A(n_2668),
.B(n_2654),
.C(n_2638),
.D(n_2639),
.E(n_2643),
.Y(n_2678)
);

OAI322xp33_ASAP7_75t_L g2679 ( 
.A1(n_2674),
.A2(n_2644),
.A3(n_2647),
.B1(n_515),
.B2(n_516),
.C1(n_517),
.C2(n_518),
.Y(n_2679)
);

NAND4xp25_ASAP7_75t_SL g2680 ( 
.A(n_2662),
.B(n_510),
.C(n_513),
.D(n_515),
.Y(n_2680)
);

OAI221xp5_ASAP7_75t_L g2681 ( 
.A1(n_2666),
.A2(n_2669),
.B1(n_2670),
.B2(n_2675),
.C(n_2676),
.Y(n_2681)
);

OAI221xp5_ASAP7_75t_L g2682 ( 
.A1(n_2673),
.A2(n_513),
.B1(n_516),
.B2(n_517),
.C(n_519),
.Y(n_2682)
);

INVx1_ASAP7_75t_L g2683 ( 
.A(n_2671),
.Y(n_2683)
);

NOR3xp33_ASAP7_75t_L g2684 ( 
.A(n_2672),
.B(n_519),
.C(n_520),
.Y(n_2684)
);

AOI221x1_ASAP7_75t_L g2685 ( 
.A1(n_2671),
.A2(n_521),
.B1(n_522),
.B2(n_523),
.C(n_524),
.Y(n_2685)
);

NAND3xp33_ASAP7_75t_L g2686 ( 
.A(n_2660),
.B(n_522),
.C(n_523),
.Y(n_2686)
);

XNOR2x1_ASAP7_75t_L g2687 ( 
.A(n_2667),
.B(n_524),
.Y(n_2687)
);

AOI221xp5_ASAP7_75t_L g2688 ( 
.A1(n_2665),
.A2(n_525),
.B1(n_526),
.B2(n_527),
.C(n_528),
.Y(n_2688)
);

INVx1_ASAP7_75t_L g2689 ( 
.A(n_2687),
.Y(n_2689)
);

INVx1_ASAP7_75t_L g2690 ( 
.A(n_2679),
.Y(n_2690)
);

NAND2xp5_ASAP7_75t_L g2691 ( 
.A(n_2684),
.B(n_2661),
.Y(n_2691)
);

OA21x2_ASAP7_75t_L g2692 ( 
.A1(n_2683),
.A2(n_2663),
.B(n_526),
.Y(n_2692)
);

AOI22xp33_ASAP7_75t_L g2693 ( 
.A1(n_2677),
.A2(n_525),
.B1(n_527),
.B2(n_528),
.Y(n_2693)
);

NAND2xp5_ASAP7_75t_L g2694 ( 
.A(n_2685),
.B(n_529),
.Y(n_2694)
);

AND2x2_ASAP7_75t_L g2695 ( 
.A(n_2686),
.B(n_529),
.Y(n_2695)
);

INVx1_ASAP7_75t_L g2696 ( 
.A(n_2694),
.Y(n_2696)
);

AOI21xp5_ASAP7_75t_L g2697 ( 
.A1(n_2691),
.A2(n_2678),
.B(n_2681),
.Y(n_2697)
);

OA22x2_ASAP7_75t_L g2698 ( 
.A1(n_2695),
.A2(n_2688),
.B1(n_2680),
.B2(n_2682),
.Y(n_2698)
);

OAI22xp5_ASAP7_75t_SL g2699 ( 
.A1(n_2692),
.A2(n_530),
.B1(n_531),
.B2(n_532),
.Y(n_2699)
);

OAI22x1_ASAP7_75t_L g2700 ( 
.A1(n_2690),
.A2(n_532),
.B1(n_533),
.B2(n_534),
.Y(n_2700)
);

OAI21xp33_ASAP7_75t_L g2701 ( 
.A1(n_2689),
.A2(n_533),
.B(n_534),
.Y(n_2701)
);

AO21x1_ASAP7_75t_L g2702 ( 
.A1(n_2697),
.A2(n_2693),
.B(n_537),
.Y(n_2702)
);

OAI21xp5_ASAP7_75t_L g2703 ( 
.A1(n_2698),
.A2(n_536),
.B(n_537),
.Y(n_2703)
);

OAI21xp5_ASAP7_75t_L g2704 ( 
.A1(n_2696),
.A2(n_536),
.B(n_538),
.Y(n_2704)
);

NAND2xp5_ASAP7_75t_SL g2705 ( 
.A(n_2702),
.B(n_2699),
.Y(n_2705)
);

OAI21xp5_ASAP7_75t_L g2706 ( 
.A1(n_2703),
.A2(n_2701),
.B(n_2700),
.Y(n_2706)
);

AOI22xp5_ASAP7_75t_L g2707 ( 
.A1(n_2704),
.A2(n_538),
.B1(n_539),
.B2(n_540),
.Y(n_2707)
);

OAI22xp33_ASAP7_75t_L g2708 ( 
.A1(n_2707),
.A2(n_539),
.B1(n_541),
.B2(n_542),
.Y(n_2708)
);

OAI22xp33_ASAP7_75t_L g2709 ( 
.A1(n_2706),
.A2(n_541),
.B1(n_542),
.B2(n_543),
.Y(n_2709)
);

AO21x2_ASAP7_75t_L g2710 ( 
.A1(n_2708),
.A2(n_2705),
.B(n_544),
.Y(n_2710)
);

AO21x1_ASAP7_75t_L g2711 ( 
.A1(n_2710),
.A2(n_2709),
.B(n_544),
.Y(n_2711)
);

AOI221xp5_ASAP7_75t_L g2712 ( 
.A1(n_2711),
.A2(n_543),
.B1(n_545),
.B2(n_546),
.C(n_547),
.Y(n_2712)
);

AOI221xp5_ASAP7_75t_L g2713 ( 
.A1(n_2712),
.A2(n_545),
.B1(n_546),
.B2(n_547),
.C(n_548),
.Y(n_2713)
);

AOI211xp5_ASAP7_75t_L g2714 ( 
.A1(n_2713),
.A2(n_548),
.B(n_549),
.C(n_550),
.Y(n_2714)
);


endmodule