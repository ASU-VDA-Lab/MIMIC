module fake_netlist_6_2620_n_83 (n_16, n_1, n_9, n_8, n_18, n_10, n_21, n_6, n_15, n_3, n_14, n_0, n_4, n_22, n_13, n_11, n_17, n_12, n_20, n_7, n_2, n_5, n_19, n_83);

input n_16;
input n_1;
input n_9;
input n_8;
input n_18;
input n_10;
input n_21;
input n_6;
input n_15;
input n_3;
input n_14;
input n_0;
input n_4;
input n_22;
input n_13;
input n_11;
input n_17;
input n_12;
input n_20;
input n_7;
input n_2;
input n_5;
input n_19;

output n_83;

wire n_52;
wire n_46;
wire n_39;
wire n_63;
wire n_73;
wire n_68;
wire n_28;
wire n_50;
wire n_49;
wire n_77;
wire n_42;
wire n_24;
wire n_54;
wire n_32;
wire n_66;
wire n_78;
wire n_23;
wire n_47;
wire n_62;
wire n_29;
wire n_75;
wire n_45;
wire n_34;
wire n_70;
wire n_37;
wire n_67;
wire n_33;
wire n_82;
wire n_27;
wire n_38;
wire n_61;
wire n_81;
wire n_59;
wire n_76;
wire n_36;
wire n_26;
wire n_55;
wire n_58;
wire n_64;
wire n_48;
wire n_65;
wire n_25;
wire n_40;
wire n_80;
wire n_41;
wire n_71;
wire n_74;
wire n_72;
wire n_60;
wire n_35;
wire n_69;
wire n_30;
wire n_79;
wire n_43;
wire n_31;
wire n_57;
wire n_53;
wire n_51;
wire n_44;
wire n_56;

INVx2_ASAP7_75t_L g23 ( 
.A(n_18),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_19),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

AND2x4_ASAP7_75t_L g27 ( 
.A(n_1),
.B(n_2),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_4),
.B(n_7),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_21),
.B(n_14),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_22),
.A2(n_11),
.B1(n_0),
.B2(n_2),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

BUFx2_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

OA21x2_ASAP7_75t_L g39 ( 
.A1(n_6),
.A2(n_13),
.B(n_20),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g40 ( 
.A(n_38),
.B(n_3),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx2_ASAP7_75t_SL g42 ( 
.A(n_26),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_27),
.A2(n_15),
.B1(n_33),
.B2(n_36),
.Y(n_43)
);

NAND3xp33_ASAP7_75t_L g44 ( 
.A(n_27),
.B(n_30),
.C(n_26),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_27),
.B(n_30),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_34),
.B(n_25),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_26),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

NAND2x1p5_ASAP7_75t_L g49 ( 
.A(n_39),
.B(n_37),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_30),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_48),
.B(n_42),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_48),
.B(n_24),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_45),
.B(n_41),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_43),
.A2(n_37),
.B1(n_25),
.B2(n_34),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_51),
.Y(n_55)
);

HB1xp67_ASAP7_75t_L g56 ( 
.A(n_52),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_53),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_54),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_53),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_53),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_57),
.B(n_49),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_59),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_60),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_56),
.B(n_58),
.Y(n_64)
);

INVxp67_ASAP7_75t_SL g65 ( 
.A(n_56),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_55),
.B(n_49),
.Y(n_66)
);

NAND2x1_ASAP7_75t_L g67 ( 
.A(n_62),
.B(n_39),
.Y(n_67)
);

INVx2_ASAP7_75t_SL g68 ( 
.A(n_63),
.Y(n_68)
);

AOI211xp5_ASAP7_75t_L g69 ( 
.A1(n_64),
.A2(n_40),
.B(n_45),
.C(n_46),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_65),
.B(n_24),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_68),
.A2(n_62),
.B1(n_66),
.B2(n_61),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_SL g72 ( 
.A1(n_70),
.A2(n_28),
.B(n_34),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_71),
.Y(n_73)
);

INVx1_ASAP7_75t_SL g74 ( 
.A(n_72),
.Y(n_74)
);

AND4x2_ASAP7_75t_L g75 ( 
.A(n_74),
.B(n_69),
.C(n_67),
.D(n_39),
.Y(n_75)
);

NOR3xp33_ASAP7_75t_L g76 ( 
.A(n_73),
.B(n_69),
.C(n_32),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_76),
.A2(n_31),
.B1(n_23),
.B2(n_29),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_L g78 ( 
.A1(n_75),
.A2(n_44),
.B(n_29),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_78),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_77),
.B(n_23),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_79),
.B(n_47),
.Y(n_81)
);

OAI22xp33_ASAP7_75t_L g82 ( 
.A1(n_80),
.A2(n_35),
.B1(n_50),
.B2(n_41),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_82),
.A2(n_35),
.B(n_81),
.Y(n_83)
);


endmodule