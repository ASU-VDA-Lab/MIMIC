module fake_jpeg_30896_n_521 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_521);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_521;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_518;
wire n_378;
wire n_133;
wire n_419;
wire n_132;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_1),
.B(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_6),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_9),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_3),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

BUFx12_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

INVx1_ASAP7_75t_SL g42 ( 
.A(n_12),
.Y(n_42)
);

CKINVDCx14_ASAP7_75t_R g43 ( 
.A(n_8),
.Y(n_43)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

OR2x2_ASAP7_75t_L g46 ( 
.A(n_10),
.B(n_11),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_6),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_7),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_1),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_15),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_0),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_5),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_13),
.Y(n_53)
);

INVx2_ASAP7_75t_SL g54 ( 
.A(n_17),
.Y(n_54)
);

CKINVDCx14_ASAP7_75t_R g153 ( 
.A(n_54),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_28),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_55),
.Y(n_126)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_56),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_28),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_57),
.Y(n_150)
);

BUFx12_ASAP7_75t_L g58 ( 
.A(n_52),
.Y(n_58)
);

INVx13_ASAP7_75t_L g130 ( 
.A(n_58),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_28),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_59),
.Y(n_159)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_60),
.Y(n_116)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_61),
.Y(n_117)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_62),
.Y(n_127)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_63),
.Y(n_123)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_64),
.Y(n_125)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_24),
.Y(n_65)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_65),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_46),
.B(n_15),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_66),
.B(n_67),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_46),
.B(n_14),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_31),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_68),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_31),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_69),
.Y(n_169)
);

BUFx16f_ASAP7_75t_L g70 ( 
.A(n_52),
.Y(n_70)
);

INVx13_ASAP7_75t_L g149 ( 
.A(n_70),
.Y(n_149)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_21),
.Y(n_71)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_71),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_17),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_72),
.B(n_93),
.Y(n_134)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_16),
.Y(n_73)
);

INVx11_ASAP7_75t_L g111 ( 
.A(n_73),
.Y(n_111)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_21),
.Y(n_74)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_74),
.Y(n_162)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_31),
.Y(n_75)
);

BUFx5_ASAP7_75t_L g132 ( 
.A(n_75),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_46),
.B(n_14),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_76),
.B(n_83),
.Y(n_133)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_16),
.Y(n_77)
);

INVx8_ASAP7_75t_L g114 ( 
.A(n_77),
.Y(n_114)
);

BUFx5_ASAP7_75t_L g78 ( 
.A(n_24),
.Y(n_78)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_78),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_38),
.Y(n_79)
);

INVx6_ASAP7_75t_L g131 ( 
.A(n_79),
.Y(n_131)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_24),
.Y(n_80)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_80),
.Y(n_146)
);

BUFx5_ASAP7_75t_L g81 ( 
.A(n_24),
.Y(n_81)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_81),
.Y(n_135)
);

INVx11_ASAP7_75t_L g82 ( 
.A(n_44),
.Y(n_82)
);

INVx5_ASAP7_75t_L g158 ( 
.A(n_82),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_18),
.B(n_0),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_19),
.B(n_0),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_84),
.B(n_87),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_38),
.Y(n_85)
);

INVx6_ASAP7_75t_L g140 ( 
.A(n_85),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_45),
.Y(n_86)
);

INVx5_ASAP7_75t_L g165 ( 
.A(n_86),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_19),
.B(n_2),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_45),
.Y(n_88)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_88),
.Y(n_110)
);

BUFx5_ASAP7_75t_L g89 ( 
.A(n_44),
.Y(n_89)
);

BUFx2_ASAP7_75t_L g115 ( 
.A(n_89),
.Y(n_115)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_20),
.Y(n_90)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_90),
.Y(n_128)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_20),
.Y(n_91)
);

INVx8_ASAP7_75t_L g161 ( 
.A(n_91),
.Y(n_161)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_38),
.Y(n_92)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_92),
.Y(n_154)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_26),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_40),
.Y(n_94)
);

INVx6_ASAP7_75t_L g144 ( 
.A(n_94),
.Y(n_144)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_25),
.Y(n_95)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_95),
.Y(n_141)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_25),
.Y(n_96)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_96),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_40),
.Y(n_97)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_97),
.Y(n_170)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_29),
.Y(n_98)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_98),
.Y(n_148)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_29),
.Y(n_99)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_99),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_41),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_100),
.B(n_102),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_22),
.B(n_2),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_101),
.B(n_33),
.Y(n_137)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_26),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_41),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_103),
.B(n_107),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_40),
.Y(n_104)
);

BUFx12f_ASAP7_75t_L g124 ( 
.A(n_104),
.Y(n_124)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_27),
.Y(n_105)
);

BUFx12f_ASAP7_75t_L g164 ( 
.A(n_105),
.Y(n_164)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_27),
.Y(n_106)
);

INVx2_ASAP7_75t_SL g168 ( 
.A(n_106),
.Y(n_168)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_35),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_30),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_108),
.Y(n_136)
);

BUFx4f_ASAP7_75t_SL g113 ( 
.A(n_70),
.Y(n_113)
);

INVx6_ASAP7_75t_SL g196 ( 
.A(n_113),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_105),
.A2(n_42),
.B1(n_32),
.B2(n_30),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_118),
.A2(n_42),
.B1(n_77),
.B2(n_75),
.Y(n_179)
);

INVx6_ASAP7_75t_SL g119 ( 
.A(n_58),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_119),
.B(n_137),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_86),
.B(n_88),
.C(n_80),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_121),
.B(n_50),
.C(n_27),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_92),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_138),
.B(n_142),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_65),
.B(n_33),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_78),
.B(n_53),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_147),
.B(n_151),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_108),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_54),
.B(n_53),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_152),
.B(n_155),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_58),
.B(n_43),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_91),
.B(n_36),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_157),
.B(n_23),
.Y(n_204)
);

BUFx2_ASAP7_75t_R g160 ( 
.A(n_73),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_160),
.B(n_32),
.Y(n_183)
);

HB1xp67_ASAP7_75t_L g166 ( 
.A(n_89),
.Y(n_166)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_166),
.Y(n_177)
);

OAI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_129),
.A2(n_106),
.B1(n_104),
.B2(n_97),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_171),
.A2(n_198),
.B1(n_212),
.B2(n_168),
.Y(n_243)
);

INVx11_ASAP7_75t_L g172 ( 
.A(n_158),
.Y(n_172)
);

INVx11_ASAP7_75t_L g231 ( 
.A(n_172),
.Y(n_231)
);

BUFx2_ASAP7_75t_L g173 ( 
.A(n_165),
.Y(n_173)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_173),
.Y(n_228)
);

BUFx12f_ASAP7_75t_L g174 ( 
.A(n_149),
.Y(n_174)
);

INVx3_ASAP7_75t_L g253 ( 
.A(n_174),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_126),
.Y(n_175)
);

INVx8_ASAP7_75t_L g224 ( 
.A(n_175),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_L g176 ( 
.A1(n_117),
.A2(n_85),
.B1(n_57),
.B2(n_59),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_176),
.A2(n_168),
.B1(n_144),
.B2(n_140),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_126),
.Y(n_178)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_178),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_179),
.A2(n_211),
.B1(n_120),
.B2(n_135),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_150),
.Y(n_180)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_180),
.Y(n_234)
);

BUFx2_ASAP7_75t_L g181 ( 
.A(n_165),
.Y(n_181)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_181),
.Y(n_242)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_124),
.Y(n_182)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_182),
.Y(n_246)
);

AND2x2_ASAP7_75t_L g236 ( 
.A(n_183),
.B(n_191),
.Y(n_236)
);

BUFx2_ASAP7_75t_L g184 ( 
.A(n_110),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_184),
.Y(n_227)
);

INVx2_ASAP7_75t_SL g186 ( 
.A(n_160),
.Y(n_186)
);

INVx2_ASAP7_75t_SL g233 ( 
.A(n_186),
.Y(n_233)
);

HB1xp67_ASAP7_75t_L g187 ( 
.A(n_122),
.Y(n_187)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_187),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_156),
.B(n_162),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_188),
.B(n_203),
.Y(n_222)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_127),
.Y(n_189)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_189),
.Y(n_256)
);

OA22x2_ASAP7_75t_L g190 ( 
.A1(n_109),
.A2(n_75),
.B1(n_55),
.B2(n_79),
.Y(n_190)
);

AO22x1_ASAP7_75t_L g247 ( 
.A1(n_190),
.A2(n_211),
.B1(n_183),
.B2(n_212),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_166),
.A2(n_39),
.B1(n_35),
.B2(n_51),
.Y(n_191)
);

HAxp5_ASAP7_75t_SL g192 ( 
.A(n_133),
.B(n_34),
.CON(n_192),
.SN(n_192)
);

AND2x2_ASAP7_75t_L g240 ( 
.A(n_192),
.B(n_198),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_153),
.A2(n_39),
.B1(n_49),
.B2(n_51),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_194),
.Y(n_226)
);

AND2x2_ASAP7_75t_L g198 ( 
.A(n_116),
.B(n_94),
.Y(n_198)
);

INVx11_ASAP7_75t_L g199 ( 
.A(n_158),
.Y(n_199)
);

BUFx24_ASAP7_75t_L g251 ( 
.A(n_199),
.Y(n_251)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_134),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_200),
.B(n_201),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_139),
.Y(n_201)
);

BUFx2_ASAP7_75t_L g202 ( 
.A(n_110),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_202),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_145),
.B(n_49),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_204),
.B(n_206),
.Y(n_244)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_128),
.Y(n_205)
);

AND2x2_ASAP7_75t_L g259 ( 
.A(n_205),
.B(n_212),
.Y(n_259)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_141),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_123),
.B(n_23),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_207),
.B(n_215),
.Y(n_230)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_143),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_208),
.B(n_209),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_115),
.Y(n_209)
);

INVx5_ASAP7_75t_L g210 ( 
.A(n_111),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_210),
.B(n_213),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_125),
.A2(n_69),
.B1(n_68),
.B2(n_82),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g212 ( 
.A(n_148),
.B(n_50),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_146),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_170),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_214),
.B(n_216),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_163),
.B(n_36),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_154),
.Y(n_216)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_112),
.B(n_50),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_217),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_113),
.B(n_34),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_218),
.Y(n_258)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_161),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_219),
.B(n_220),
.Y(n_241)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_131),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_221),
.B(n_115),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_L g225 ( 
.A1(n_190),
.A2(n_140),
.B1(n_131),
.B2(n_144),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_225),
.A2(n_238),
.B1(n_239),
.B2(n_252),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_229),
.B(n_183),
.C(n_190),
.Y(n_265)
);

OAI32xp33_ASAP7_75t_L g237 ( 
.A1(n_188),
.A2(n_153),
.A3(n_136),
.B1(n_118),
.B2(n_164),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_237),
.B(n_191),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_L g239 ( 
.A1(n_190),
.A2(n_150),
.B1(n_159),
.B2(n_167),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g274 ( 
.A(n_243),
.B(n_247),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_221),
.A2(n_169),
.B1(n_167),
.B2(n_159),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_254),
.A2(n_198),
.B1(n_193),
.B2(n_114),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_186),
.A2(n_120),
.B(n_135),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_255),
.A2(n_254),
.B(n_233),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_245),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_260),
.B(n_266),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_230),
.B(n_207),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_262),
.B(n_264),
.Y(n_295)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_256),
.Y(n_263)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_263),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_230),
.B(n_215),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_265),
.B(n_267),
.C(n_272),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_245),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_226),
.A2(n_217),
.B1(n_186),
.B2(n_189),
.Y(n_267)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_267),
.Y(n_314)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_256),
.Y(n_268)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_268),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_222),
.B(n_217),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_269),
.B(n_285),
.Y(n_308)
);

OAI32xp33_ASAP7_75t_L g301 ( 
.A1(n_270),
.A2(n_240),
.A3(n_250),
.B1(n_255),
.B2(n_248),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_241),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_271),
.B(n_287),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_272),
.A2(n_273),
.B1(n_283),
.B2(n_233),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_247),
.A2(n_195),
.B1(n_205),
.B2(n_197),
.Y(n_273)
);

AND2x6_ASAP7_75t_L g275 ( 
.A(n_237),
.B(n_192),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_SL g311 ( 
.A(n_275),
.B(n_278),
.C(n_282),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_L g292 ( 
.A1(n_276),
.A2(n_282),
.B(n_236),
.Y(n_292)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_223),
.Y(n_277)
);

CKINVDCx14_ASAP7_75t_R g304 ( 
.A(n_277),
.Y(n_304)
);

AND2x6_ASAP7_75t_L g278 ( 
.A(n_229),
.B(n_130),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_223),
.Y(n_279)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_279),
.Y(n_302)
);

INVx3_ASAP7_75t_L g280 ( 
.A(n_253),
.Y(n_280)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_280),
.Y(n_309)
);

INVx13_ASAP7_75t_L g281 ( 
.A(n_253),
.Y(n_281)
);

BUFx2_ASAP7_75t_SL g307 ( 
.A(n_281),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_L g282 ( 
.A1(n_236),
.A2(n_185),
.B(n_203),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_247),
.A2(n_216),
.B1(n_169),
.B2(n_220),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_241),
.Y(n_284)
);

CKINVDCx16_ASAP7_75t_R g310 ( 
.A(n_284),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_244),
.B(n_177),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_222),
.B(n_177),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_286),
.B(n_291),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_244),
.B(n_213),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_235),
.B(n_174),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_288),
.B(n_290),
.Y(n_320)
);

AND2x2_ASAP7_75t_L g289 ( 
.A(n_259),
.B(n_214),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_289),
.Y(n_315)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_250),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_258),
.B(n_22),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g328 ( 
.A(n_292),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_274),
.A2(n_232),
.B1(n_236),
.B2(n_252),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_294),
.A2(n_321),
.B1(n_261),
.B2(n_265),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_276),
.A2(n_243),
.B1(n_240),
.B2(n_259),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_296),
.A2(n_300),
.B1(n_303),
.B2(n_289),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_274),
.A2(n_240),
.B1(n_259),
.B2(n_233),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g338 ( 
.A(n_297),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_299),
.B(n_278),
.C(n_263),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_301),
.B(n_317),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_271),
.A2(n_238),
.B1(n_248),
.B2(n_178),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_262),
.B(n_235),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_306),
.B(n_264),
.Y(n_336)
);

INVx13_ASAP7_75t_L g333 ( 
.A(n_311),
.Y(n_333)
);

MAJx2_ASAP7_75t_L g312 ( 
.A(n_269),
.B(n_249),
.C(n_196),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_312),
.B(n_313),
.Y(n_324)
);

XNOR2x1_ASAP7_75t_SL g313 ( 
.A(n_274),
.B(n_249),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g317 ( 
.A(n_288),
.Y(n_317)
);

OA21x2_ASAP7_75t_L g319 ( 
.A1(n_270),
.A2(n_251),
.B(n_257),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_L g326 ( 
.A1(n_319),
.A2(n_283),
.B(n_289),
.Y(n_326)
);

AOI22xp33_ASAP7_75t_L g321 ( 
.A1(n_266),
.A2(n_175),
.B1(n_180),
.B2(n_228),
.Y(n_321)
);

XOR2x2_ASAP7_75t_L g322 ( 
.A(n_313),
.B(n_311),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_322),
.B(n_312),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_323),
.A2(n_314),
.B1(n_310),
.B2(n_308),
.Y(n_355)
);

AOI21xp5_ASAP7_75t_L g367 ( 
.A1(n_326),
.A2(n_341),
.B(n_350),
.Y(n_367)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_293),
.Y(n_327)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_327),
.Y(n_364)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_293),
.Y(n_329)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_329),
.Y(n_375)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_298),
.Y(n_330)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_330),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_316),
.B(n_285),
.Y(n_331)
);

INVxp33_ASAP7_75t_L g366 ( 
.A(n_331),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_316),
.B(n_320),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_332),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_334),
.A2(n_335),
.B1(n_349),
.B2(n_350),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_294),
.A2(n_261),
.B1(n_284),
.B2(n_275),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_336),
.B(n_342),
.Y(n_352)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_298),
.Y(n_337)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_337),
.Y(n_378)
);

OR2x2_ASAP7_75t_L g339 ( 
.A(n_318),
.B(n_290),
.Y(n_339)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_339),
.Y(n_382)
);

INVx13_ASAP7_75t_L g340 ( 
.A(n_307),
.Y(n_340)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_340),
.Y(n_353)
);

OAI21xp5_ASAP7_75t_L g341 ( 
.A1(n_319),
.A2(n_292),
.B(n_297),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_306),
.B(n_295),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_308),
.B(n_286),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_343),
.B(n_345),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_SL g344 ( 
.A(n_305),
.B(n_273),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_SL g359 ( 
.A(n_344),
.B(n_300),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_295),
.B(n_287),
.Y(n_345)
);

INVx13_ASAP7_75t_L g346 ( 
.A(n_304),
.Y(n_346)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_346),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_347),
.B(n_312),
.C(n_315),
.Y(n_363)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_318),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_348),
.B(n_351),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_299),
.A2(n_268),
.B1(n_234),
.B2(n_224),
.Y(n_349)
);

AOI21xp5_ASAP7_75t_L g350 ( 
.A1(n_296),
.A2(n_280),
.B(n_227),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_305),
.B(n_291),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_355),
.A2(n_357),
.B1(n_334),
.B2(n_325),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_SL g385 ( 
.A(n_356),
.B(n_324),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_L g357 ( 
.A1(n_344),
.A2(n_310),
.B1(n_320),
.B2(n_303),
.Y(n_357)
);

BUFx3_ASAP7_75t_L g358 ( 
.A(n_349),
.Y(n_358)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_358),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_359),
.B(n_360),
.Y(n_383)
);

HB1xp67_ASAP7_75t_L g360 ( 
.A(n_348),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_SL g361 ( 
.A(n_351),
.B(n_309),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_361),
.B(n_368),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_339),
.B(n_281),
.Y(n_362)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_362),
.Y(n_390)
);

XOR2xp5_ASAP7_75t_L g391 ( 
.A(n_363),
.B(n_324),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_365),
.B(n_323),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_SL g368 ( 
.A(n_339),
.B(n_309),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_331),
.B(n_281),
.Y(n_372)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_372),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_332),
.B(n_319),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_373),
.B(n_374),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_345),
.B(n_319),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_342),
.B(n_302),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_376),
.B(n_379),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_336),
.B(n_257),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_322),
.B(n_301),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_380),
.B(n_335),
.Y(n_400)
);

INVxp67_ASAP7_75t_L g381 ( 
.A(n_326),
.Y(n_381)
);

AOI21xp5_ASAP7_75t_L g389 ( 
.A1(n_381),
.A2(n_326),
.B(n_341),
.Y(n_389)
);

OAI21xp5_ASAP7_75t_L g384 ( 
.A1(n_367),
.A2(n_381),
.B(n_373),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g430 ( 
.A(n_384),
.B(n_392),
.Y(n_430)
);

XOR2xp5_ASAP7_75t_L g429 ( 
.A(n_385),
.B(n_391),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_363),
.B(n_347),
.C(n_322),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_386),
.B(n_396),
.C(n_403),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_SL g414 ( 
.A1(n_387),
.A2(n_394),
.B1(n_382),
.B2(n_370),
.Y(n_414)
);

CKINVDCx14_ASAP7_75t_R g419 ( 
.A(n_389),
.Y(n_419)
);

OAI21xp5_ASAP7_75t_L g392 ( 
.A1(n_367),
.A2(n_325),
.B(n_341),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_SL g393 ( 
.A(n_356),
.B(n_324),
.Y(n_393)
);

XOR2xp5_ASAP7_75t_SL g417 ( 
.A(n_393),
.B(n_399),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_380),
.B(n_347),
.C(n_328),
.Y(n_396)
);

AND2x2_ASAP7_75t_L g398 ( 
.A(n_371),
.B(n_365),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_398),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_SL g399 ( 
.A(n_371),
.B(n_343),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_400),
.B(n_406),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_L g402 ( 
.A1(n_358),
.A2(n_338),
.B1(n_327),
.B2(n_337),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_SL g418 ( 
.A(n_402),
.B(n_405),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_376),
.B(n_333),
.C(n_330),
.Y(n_403)
);

XOR2xp5_ASAP7_75t_L g404 ( 
.A(n_355),
.B(n_333),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_404),
.B(n_411),
.C(n_279),
.Y(n_433)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_369),
.A2(n_329),
.B1(n_302),
.B2(n_333),
.Y(n_405)
);

INVxp67_ASAP7_75t_L g406 ( 
.A(n_374),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_SL g407 ( 
.A(n_352),
.B(n_227),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_407),
.B(n_408),
.Y(n_422)
);

INVxp67_ASAP7_75t_L g408 ( 
.A(n_364),
.Y(n_408)
);

AND2x2_ASAP7_75t_L g410 ( 
.A(n_382),
.B(n_346),
.Y(n_410)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_410),
.Y(n_415)
);

XOR2xp5_ASAP7_75t_L g411 ( 
.A(n_352),
.B(n_346),
.Y(n_411)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_414),
.A2(n_423),
.B1(n_426),
.B2(n_427),
.Y(n_446)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_409),
.Y(n_416)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_416),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_398),
.A2(n_378),
.B1(n_377),
.B2(n_375),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_SL g454 ( 
.A1(n_420),
.A2(n_425),
.B1(n_340),
.B2(n_231),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_SL g421 ( 
.A(n_395),
.B(n_366),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_421),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_SL g423 ( 
.A1(n_406),
.A2(n_370),
.B1(n_377),
.B2(n_375),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_390),
.Y(n_424)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_424),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_404),
.A2(n_378),
.B1(n_364),
.B2(n_354),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_SL g426 ( 
.A1(n_397),
.A2(n_354),
.B1(n_353),
.B2(n_224),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_SL g427 ( 
.A1(n_392),
.A2(n_353),
.B1(n_224),
.B2(n_234),
.Y(n_427)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_410),
.Y(n_431)
);

CKINVDCx16_ASAP7_75t_R g447 ( 
.A(n_431),
.Y(n_447)
);

INVxp67_ASAP7_75t_SL g432 ( 
.A(n_383),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_432),
.B(n_401),
.Y(n_435)
);

XOR2xp5_ASAP7_75t_L g440 ( 
.A(n_433),
.B(n_400),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_403),
.B(n_246),
.C(n_242),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_434),
.B(n_433),
.C(n_428),
.Y(n_441)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_435),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_412),
.B(n_399),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_SL g457 ( 
.A(n_437),
.B(n_450),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_422),
.B(n_408),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_L g459 ( 
.A(n_439),
.B(n_440),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_441),
.B(n_443),
.C(n_451),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_428),
.B(n_396),
.C(n_386),
.Y(n_443)
);

OR2x2_ASAP7_75t_L g444 ( 
.A(n_415),
.B(n_384),
.Y(n_444)
);

OAI21xp5_ASAP7_75t_L g464 ( 
.A1(n_444),
.A2(n_446),
.B(n_439),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_416),
.B(n_411),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g471 ( 
.A(n_445),
.B(n_449),
.Y(n_471)
);

AOI22xp5_ASAP7_75t_L g448 ( 
.A1(n_414),
.A2(n_388),
.B1(n_391),
.B2(n_393),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_SL g462 ( 
.A1(n_448),
.A2(n_446),
.B1(n_445),
.B2(n_417),
.Y(n_462)
);

XOR2xp5_ASAP7_75t_L g449 ( 
.A(n_429),
.B(n_385),
.Y(n_449)
);

CKINVDCx16_ASAP7_75t_R g450 ( 
.A(n_420),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_434),
.B(n_246),
.C(n_277),
.Y(n_451)
);

HB1xp67_ASAP7_75t_L g452 ( 
.A(n_415),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_SL g470 ( 
.A(n_452),
.B(n_202),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_425),
.B(n_242),
.C(n_228),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_453),
.B(n_427),
.C(n_426),
.Y(n_463)
);

AOI22xp5_ASAP7_75t_L g465 ( 
.A1(n_454),
.A2(n_417),
.B1(n_210),
.B2(n_231),
.Y(n_465)
);

AOI21xp5_ASAP7_75t_L g455 ( 
.A1(n_444),
.A2(n_430),
.B(n_413),
.Y(n_455)
);

OAI21xp5_ASAP7_75t_SL g476 ( 
.A1(n_455),
.A2(n_440),
.B(n_449),
.Y(n_476)
);

OAI22xp5_ASAP7_75t_L g458 ( 
.A1(n_442),
.A2(n_419),
.B1(n_418),
.B2(n_423),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_458),
.B(n_463),
.Y(n_480)
);

NOR2xp67_ASAP7_75t_L g460 ( 
.A(n_447),
.B(n_430),
.Y(n_460)
);

OAI21x1_ASAP7_75t_L g485 ( 
.A1(n_460),
.A2(n_149),
.B(n_130),
.Y(n_485)
);

XNOR2xp5_ASAP7_75t_L g472 ( 
.A(n_462),
.B(n_470),
.Y(n_472)
);

AOI21xp5_ASAP7_75t_SL g473 ( 
.A1(n_464),
.A2(n_454),
.B(n_448),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_465),
.B(n_467),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_441),
.B(n_429),
.C(n_182),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_466),
.B(n_469),
.C(n_451),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_SL g467 ( 
.A1(n_436),
.A2(n_114),
.B1(n_340),
.B2(n_173),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_L g468 ( 
.A1(n_438),
.A2(n_196),
.B1(n_181),
.B2(n_184),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_468),
.B(n_453),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_443),
.B(n_251),
.C(n_161),
.Y(n_469)
);

CKINVDCx14_ASAP7_75t_R g493 ( 
.A(n_473),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_474),
.B(n_477),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_SL g497 ( 
.A(n_475),
.B(n_484),
.Y(n_497)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_476),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_459),
.B(n_461),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_461),
.B(n_251),
.C(n_199),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_478),
.B(n_479),
.C(n_471),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_459),
.B(n_251),
.C(n_172),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_SL g482 ( 
.A(n_456),
.B(n_124),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_482),
.B(n_486),
.Y(n_489)
);

OAI22xp5_ASAP7_75t_L g483 ( 
.A1(n_464),
.A2(n_111),
.B1(n_132),
.B2(n_124),
.Y(n_483)
);

AOI22xp5_ASAP7_75t_L g491 ( 
.A1(n_483),
.A2(n_485),
.B1(n_467),
.B2(n_3),
.Y(n_491)
);

AOI21xp5_ASAP7_75t_L g484 ( 
.A1(n_469),
.A2(n_174),
.B(n_3),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_SL g486 ( 
.A(n_466),
.B(n_164),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_SL g488 ( 
.A(n_472),
.B(n_457),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_488),
.B(n_490),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_480),
.B(n_475),
.C(n_478),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_491),
.B(n_492),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_473),
.B(n_463),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_495),
.B(n_498),
.C(n_41),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_479),
.B(n_462),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_SL g501 ( 
.A(n_496),
.B(n_499),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_481),
.B(n_471),
.C(n_465),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_477),
.B(n_164),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_500),
.B(n_506),
.Y(n_511)
);

A2O1A1Ixp33_ASAP7_75t_SL g503 ( 
.A1(n_493),
.A2(n_2),
.B(n_3),
.C(n_5),
.Y(n_503)
);

AOI21xp5_ASAP7_75t_L g509 ( 
.A1(n_503),
.A2(n_7),
.B(n_8),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_487),
.B(n_41),
.C(n_6),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_SL g508 ( 
.A(n_504),
.B(n_505),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_494),
.B(n_5),
.C(n_6),
.Y(n_505)
);

AND2x2_ASAP7_75t_L g506 ( 
.A(n_495),
.B(n_7),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_SL g513 ( 
.A(n_509),
.B(n_510),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_SL g510 ( 
.A(n_502),
.B(n_489),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_SL g512 ( 
.A(n_507),
.B(n_493),
.Y(n_512)
);

AOI21xp5_ASAP7_75t_L g514 ( 
.A1(n_512),
.A2(n_501),
.B(n_497),
.Y(n_514)
);

INVxp67_ASAP7_75t_L g516 ( 
.A(n_514),
.Y(n_516)
);

A2O1A1Ixp33_ASAP7_75t_SL g515 ( 
.A1(n_511),
.A2(n_503),
.B(n_498),
.C(n_13),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_515),
.B(n_508),
.C(n_8),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_SL g518 ( 
.A(n_517),
.B(n_513),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_518),
.Y(n_519)
);

OAI21xp5_ASAP7_75t_SL g520 ( 
.A1(n_519),
.A2(n_516),
.B(n_11),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_520),
.Y(n_521)
);


endmodule