module fake_jpeg_5032_n_98 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_98);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_98;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;
wire n_96;

INVx4_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

INVx3_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

OR2x2_ASAP7_75t_L g22 ( 
.A(n_7),
.B(n_9),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_22),
.B(n_0),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_25),
.B(n_31),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_13),
.B(n_1),
.Y(n_27)
);

OAI21xp33_ASAP7_75t_L g49 ( 
.A1(n_27),
.A2(n_2),
.B(n_4),
.Y(n_49)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_21),
.Y(n_29)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_30),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_13),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_32),
.B(n_24),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_21),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_33),
.A2(n_18),
.B1(n_4),
.B2(n_5),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_20),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_34),
.B(n_19),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g35 ( 
.A1(n_30),
.A2(n_23),
.B1(n_14),
.B2(n_18),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_35),
.A2(n_39),
.B1(n_45),
.B2(n_6),
.Y(n_58)
);

INVx13_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_36),
.B(n_41),
.Y(n_59)
);

OA22x2_ASAP7_75t_L g39 ( 
.A1(n_29),
.A2(n_23),
.B1(n_14),
.B2(n_17),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_34),
.Y(n_41)
);

XNOR2xp5_ASAP7_75t_L g42 ( 
.A(n_25),
.B(n_15),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_42),
.B(n_49),
.Y(n_61)
);

OAI22xp33_ASAP7_75t_L g45 ( 
.A1(n_29),
.A2(n_19),
.B1(n_15),
.B2(n_12),
.Y(n_45)
);

INVx13_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

INVx13_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

A2O1A1Ixp33_ASAP7_75t_L g47 ( 
.A1(n_31),
.A2(n_12),
.B(n_10),
.C(n_11),
.Y(n_47)
);

AOI21xp5_ASAP7_75t_SL g55 ( 
.A1(n_47),
.A2(n_51),
.B(n_39),
.Y(n_55)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_24),
.Y(n_48)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_L g65 ( 
.A1(n_50),
.A2(n_54),
.B(n_38),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_L g62 ( 
.A1(n_52),
.A2(n_8),
.B(n_47),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

OR2x2_ASAP7_75t_L g66 ( 
.A(n_53),
.B(n_45),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_55),
.Y(n_71)
);

OAI32xp33_ASAP7_75t_L g57 ( 
.A1(n_39),
.A2(n_32),
.A3(n_27),
.B1(n_26),
.B2(n_2),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_57),
.B(n_36),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_58),
.B(n_65),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_53),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_60),
.A2(n_67),
.B1(n_68),
.B2(n_46),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_62),
.Y(n_74)
);

OAI21xp33_ASAP7_75t_SL g63 ( 
.A1(n_39),
.A2(n_42),
.B(n_35),
.Y(n_63)
);

OAI21x1_ASAP7_75t_L g79 ( 
.A1(n_63),
.A2(n_66),
.B(n_57),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_50),
.A2(n_44),
.B1(n_48),
.B2(n_43),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_44),
.A2(n_43),
.B1(n_40),
.B2(n_37),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_69),
.A2(n_73),
.B1(n_79),
.B2(n_60),
.Y(n_80)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_67),
.Y(n_70)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_70),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_59),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_SL g82 ( 
.A1(n_72),
.A2(n_64),
.B(n_62),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_56),
.Y(n_75)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_75),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_61),
.B(n_65),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_77),
.B(n_78),
.C(n_61),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_61),
.B(n_55),
.Y(n_78)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_80),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_82),
.B(n_74),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_83),
.B(n_84),
.C(n_85),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_77),
.B(n_64),
.C(n_68),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_78),
.B(n_58),
.C(n_66),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_SL g93 ( 
.A1(n_89),
.A2(n_71),
.B(n_76),
.Y(n_93)
);

BUFx24_ASAP7_75t_SL g90 ( 
.A(n_86),
.Y(n_90)
);

NAND2xp33_ASAP7_75t_L g92 ( 
.A(n_90),
.B(n_79),
.Y(n_92)
);

INVxp33_ASAP7_75t_L g91 ( 
.A(n_81),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_91),
.A2(n_73),
.B1(n_72),
.B2(n_70),
.Y(n_94)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_92),
.Y(n_96)
);

AOI322xp5_ASAP7_75t_L g95 ( 
.A1(n_93),
.A2(n_94),
.A3(n_71),
.B1(n_88),
.B2(n_83),
.C1(n_69),
.C2(n_87),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_95),
.B(n_66),
.C(n_56),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_97),
.A2(n_75),
.B1(n_96),
.B2(n_71),
.Y(n_98)
);


endmodule