module fake_jpeg_24156_n_253 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_253);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_253;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_122;
wire n_75;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx12_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_15),
.Y(n_22)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_9),
.Y(n_29)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_35),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_30),
.B(n_0),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_36),
.B(n_41),
.Y(n_48)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_37),
.B(n_30),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_22),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_38),
.B(n_40),
.Y(n_52)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_19),
.B(n_0),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_22),
.Y(n_41)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

HB1xp67_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_45),
.B(n_46),
.Y(n_75)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_47),
.B(n_58),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_39),
.A2(n_32),
.B1(n_34),
.B2(n_20),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_50),
.A2(n_54),
.B1(n_33),
.B2(n_21),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_37),
.A2(n_34),
.B1(n_20),
.B2(n_31),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_53),
.A2(n_42),
.B1(n_31),
.B2(n_17),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_39),
.A2(n_34),
.B1(n_17),
.B2(n_33),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_36),
.B(n_28),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_57),
.B(n_25),
.Y(n_70)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_59),
.B(n_63),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_39),
.A2(n_24),
.B1(n_27),
.B2(n_21),
.Y(n_60)
);

OAI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_60),
.A2(n_18),
.B1(n_27),
.B2(n_41),
.Y(n_94)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_61),
.Y(n_66)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_64),
.Y(n_67)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_65),
.B(n_33),
.Y(n_88)
);

OAI22xp33_ASAP7_75t_L g68 ( 
.A1(n_51),
.A2(n_42),
.B1(n_37),
.B2(n_36),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_68),
.A2(n_72),
.B1(n_76),
.B2(n_90),
.Y(n_104)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_62),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_69),
.B(n_71),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_70),
.B(n_79),
.Y(n_106)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_62),
.Y(n_71)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_53),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_73),
.B(n_77),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_48),
.A2(n_24),
.B1(n_40),
.B2(n_17),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_74),
.A2(n_80),
.B(n_86),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_51),
.A2(n_18),
.B1(n_27),
.B2(n_21),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_61),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_52),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_78),
.B(n_81),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_48),
.B(n_30),
.Y(n_79)
);

AO22x1_ASAP7_75t_L g80 ( 
.A1(n_49),
.A2(n_44),
.B1(n_30),
.B2(n_25),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_52),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_57),
.B(n_24),
.C(n_44),
.Y(n_82)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_82),
.B(n_83),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_56),
.B(n_44),
.C(n_30),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_63),
.B(n_41),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_85),
.B(n_93),
.Y(n_101)
);

AO21x1_ASAP7_75t_L g86 ( 
.A1(n_49),
.A2(n_65),
.B(n_31),
.Y(n_86)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_88),
.Y(n_112)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_55),
.Y(n_89)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_89),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_46),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_91),
.Y(n_118)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_55),
.Y(n_92)
);

HB1xp67_ASAP7_75t_L g102 ( 
.A(n_92),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_55),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_94),
.B(n_99),
.Y(n_113)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_64),
.Y(n_95)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_95),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_47),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_96),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g97 ( 
.A(n_45),
.B(n_28),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_97),
.B(n_98),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_56),
.B(n_25),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_58),
.B(n_38),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_73),
.A2(n_59),
.B1(n_38),
.B2(n_25),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_100),
.A2(n_119),
.B1(n_92),
.B2(n_95),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_70),
.B(n_23),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_109),
.B(n_120),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_81),
.A2(n_26),
.B1(n_29),
.B2(n_18),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_110),
.A2(n_115),
.B1(n_116),
.B2(n_120),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_78),
.A2(n_72),
.B1(n_79),
.B2(n_82),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_86),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_116),
.B(n_125),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_66),
.A2(n_29),
.B1(n_26),
.B2(n_23),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_74),
.B(n_66),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_77),
.B(n_23),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_122),
.B(n_124),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_85),
.B(n_97),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_87),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_126),
.B(n_127),
.Y(n_158)
);

CKINVDCx14_ASAP7_75t_R g127 ( 
.A(n_121),
.Y(n_127)
);

MAJx2_ASAP7_75t_L g128 ( 
.A(n_124),
.B(n_68),
.C(n_80),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_128),
.B(n_115),
.C(n_104),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_111),
.B(n_83),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_129),
.B(n_122),
.Y(n_160)
);

INVx13_ASAP7_75t_L g130 ( 
.A(n_102),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_130),
.B(n_131),
.Y(n_153)
);

INVx11_ASAP7_75t_L g131 ( 
.A(n_114),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_121),
.A2(n_80),
.B1(n_98),
.B2(n_69),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_132),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_111),
.B(n_96),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_133),
.A2(n_139),
.B(n_141),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_118),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_134),
.Y(n_156)
);

OAI211xp5_ASAP7_75t_L g136 ( 
.A1(n_105),
.A2(n_91),
.B(n_75),
.C(n_23),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_136),
.B(n_123),
.Y(n_155)
);

AO21x1_ASAP7_75t_L g139 ( 
.A1(n_105),
.A2(n_71),
.B(n_67),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_118),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_140),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_108),
.A2(n_67),
.B(n_84),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_SL g142 ( 
.A(n_108),
.B(n_23),
.C(n_19),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_142),
.A2(n_147),
.B(n_150),
.Y(n_173)
);

CKINVDCx14_ASAP7_75t_R g143 ( 
.A(n_100),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_143),
.B(n_145),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_144),
.A2(n_149),
.B1(n_113),
.B2(n_112),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_123),
.B(n_117),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_106),
.B(n_89),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_146),
.B(n_148),
.Y(n_170)
);

NOR2x1_ASAP7_75t_L g147 ( 
.A(n_110),
.B(n_19),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_106),
.B(n_109),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_107),
.A2(n_19),
.B1(n_2),
.B2(n_3),
.Y(n_149)
);

AOI21xp33_ASAP7_75t_L g150 ( 
.A1(n_107),
.A2(n_1),
.B(n_2),
.Y(n_150)
);

CKINVDCx10_ASAP7_75t_R g151 ( 
.A(n_102),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_151),
.B(n_1),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_101),
.B(n_19),
.Y(n_152)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_152),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_154),
.B(n_160),
.Y(n_179)
);

AOI221xp5_ASAP7_75t_L g181 ( 
.A1(n_155),
.A2(n_135),
.B1(n_152),
.B2(n_148),
.C(n_137),
.Y(n_181)
);

OR2x2_ASAP7_75t_L g157 ( 
.A(n_147),
.B(n_103),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_157),
.B(n_138),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_L g161 ( 
.A1(n_147),
.A2(n_104),
.B1(n_103),
.B2(n_112),
.Y(n_161)
);

CKINVDCx14_ASAP7_75t_R g178 ( 
.A(n_161),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_133),
.B(n_101),
.C(n_125),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_162),
.B(n_174),
.C(n_138),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_163),
.B(n_171),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_142),
.A2(n_113),
.B1(n_114),
.B2(n_119),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_167),
.A2(n_169),
.B(n_6),
.Y(n_194)
);

AO22x1_ASAP7_75t_L g169 ( 
.A1(n_139),
.A2(n_117),
.B1(n_2),
.B2(n_4),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_134),
.B(n_4),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_172),
.B(n_175),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_129),
.B(n_5),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_146),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_140),
.B(n_5),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_176),
.Y(n_180)
);

AOI221xp5_ASAP7_75t_SL g177 ( 
.A1(n_154),
.A2(n_128),
.B1(n_139),
.B2(n_126),
.C(n_141),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_177),
.A2(n_193),
.B1(n_194),
.B2(n_159),
.Y(n_203)
);

BUFx24_ASAP7_75t_SL g199 ( 
.A(n_181),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_183),
.B(n_164),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_184),
.B(n_192),
.C(n_173),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_170),
.B(n_135),
.Y(n_185)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_185),
.Y(n_207)
);

INVxp67_ASAP7_75t_SL g186 ( 
.A(n_169),
.Y(n_186)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_186),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_165),
.B(n_160),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_187),
.B(n_188),
.Y(n_208)
);

MAJx2_ASAP7_75t_L g188 ( 
.A(n_165),
.B(n_133),
.C(n_137),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_174),
.B(n_151),
.C(n_132),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_189),
.B(n_190),
.C(n_191),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_162),
.B(n_144),
.C(n_149),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_170),
.B(n_130),
.C(n_131),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_175),
.B(n_5),
.C(n_6),
.Y(n_192)
);

XOR2x2_ASAP7_75t_L g193 ( 
.A(n_159),
.B(n_6),
.Y(n_193)
);

HB1xp67_ASAP7_75t_L g196 ( 
.A(n_169),
.Y(n_196)
);

BUFx2_ASAP7_75t_L g204 ( 
.A(n_196),
.Y(n_204)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_197),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_198),
.B(n_200),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_195),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_180),
.B(n_156),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_201),
.B(n_166),
.Y(n_218)
);

BUFx12_ASAP7_75t_L g202 ( 
.A(n_193),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_202),
.B(n_210),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_203),
.A2(n_167),
.B1(n_155),
.B2(n_178),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_191),
.B(n_156),
.Y(n_205)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_205),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_179),
.B(n_168),
.C(n_158),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_206),
.B(n_184),
.Y(n_222)
);

BUFx12_ASAP7_75t_L g210 ( 
.A(n_179),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_212),
.B(n_222),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_209),
.A2(n_183),
.B1(n_190),
.B2(n_189),
.Y(n_216)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_216),
.Y(n_225)
);

NOR3xp33_ASAP7_75t_L g217 ( 
.A(n_202),
.B(n_166),
.C(n_173),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_217),
.B(n_218),
.Y(n_228)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_204),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_219),
.B(n_223),
.Y(n_229)
);

OA21x2_ASAP7_75t_L g221 ( 
.A1(n_204),
.A2(n_157),
.B(n_194),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_221),
.A2(n_157),
.B(n_168),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_207),
.A2(n_185),
.B1(n_182),
.B2(n_188),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_221),
.A2(n_206),
.B(n_202),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_226),
.A2(n_227),
.B(n_230),
.Y(n_236)
);

MAJx2_ASAP7_75t_L g227 ( 
.A(n_215),
.B(n_208),
.C(n_187),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_214),
.B(n_153),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_231),
.B(n_233),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_SL g232 ( 
.A1(n_221),
.A2(n_208),
.B1(n_210),
.B2(n_192),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_232),
.A2(n_211),
.B(n_198),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_213),
.B(n_163),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_228),
.B(n_220),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_234),
.B(n_229),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_224),
.B(n_211),
.C(n_216),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_235),
.B(n_236),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_238),
.B(n_240),
.Y(n_241)
);

AOI21xp33_ASAP7_75t_L g239 ( 
.A1(n_225),
.A2(n_210),
.B(n_199),
.Y(n_239)
);

NOR2xp67_ASAP7_75t_SL g243 ( 
.A(n_239),
.B(n_232),
.Y(n_243)
);

AOI322xp5_ASAP7_75t_L g240 ( 
.A1(n_226),
.A2(n_222),
.A3(n_223),
.B1(n_10),
.B2(n_11),
.C1(n_12),
.C2(n_8),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_242),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_247)
);

AOI31xp33_ASAP7_75t_L g248 ( 
.A1(n_243),
.A2(n_15),
.A3(n_10),
.B(n_11),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_237),
.B(n_224),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_244),
.B(n_245),
.C(n_8),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_241),
.B(n_235),
.C(n_227),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_246),
.A2(n_248),
.B(n_12),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_247),
.B(n_249),
.Y(n_250)
);

OAI321xp33_ASAP7_75t_L g252 ( 
.A1(n_251),
.A2(n_12),
.A3(n_13),
.B1(n_14),
.B2(n_15),
.C(n_246),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_252),
.B(n_250),
.Y(n_253)
);


endmodule