module fake_jpeg_12179_n_647 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_647);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_647;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_384;
wire n_296;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_18),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx8_ASAP7_75t_SL g29 ( 
.A(n_5),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_11),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

OR2x2_ASAP7_75t_L g38 ( 
.A(n_15),
.B(n_2),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_17),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_4),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_0),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_15),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_12),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_1),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_9),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_7),
.Y(n_49)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_17),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_2),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_12),
.Y(n_52)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_1),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_16),
.B(n_10),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_8),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_3),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_16),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_18),
.Y(n_58)
);

BUFx12_ASAP7_75t_L g59 ( 
.A(n_15),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_4),
.Y(n_60)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_52),
.Y(n_61)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_61),
.Y(n_136)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_28),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_62),
.Y(n_131)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_29),
.Y(n_63)
);

INVx11_ASAP7_75t_L g133 ( 
.A(n_63),
.Y(n_133)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

INVx5_ASAP7_75t_L g199 ( 
.A(n_64),
.Y(n_199)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_19),
.Y(n_65)
);

HB1xp67_ASAP7_75t_L g149 ( 
.A(n_65),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_22),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_66),
.Y(n_139)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_19),
.Y(n_67)
);

HB1xp67_ASAP7_75t_L g162 ( 
.A(n_67),
.Y(n_162)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_29),
.Y(n_68)
);

INVx11_ASAP7_75t_L g177 ( 
.A(n_68),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_54),
.B(n_18),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_69),
.B(n_75),
.Y(n_174)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_70),
.Y(n_127)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_71),
.Y(n_170)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

BUFx2_ASAP7_75t_L g138 ( 
.A(n_72),
.Y(n_138)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_73),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_54),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_74),
.B(n_88),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_23),
.B(n_18),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_22),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_76),
.Y(n_155)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_40),
.Y(n_77)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_77),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_22),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_78),
.Y(n_161)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_24),
.Y(n_79)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_79),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_22),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_80),
.Y(n_164)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_19),
.Y(n_81)
);

BUFx2_ASAP7_75t_L g163 ( 
.A(n_81),
.Y(n_163)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_40),
.Y(n_82)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_82),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_23),
.B(n_17),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_83),
.B(n_104),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_38),
.B(n_17),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_84),
.B(n_114),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_31),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_85),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_31),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_86),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_31),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_87),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_39),
.B(n_14),
.Y(n_88)
);

BUFx5_ASAP7_75t_L g89 ( 
.A(n_28),
.Y(n_89)
);

BUFx2_ASAP7_75t_L g179 ( 
.A(n_89),
.Y(n_179)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_24),
.Y(n_90)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_90),
.Y(n_143)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_36),
.Y(n_91)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_91),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_31),
.Y(n_92)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_92),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_59),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_93),
.B(n_109),
.Y(n_150)
);

NAND2x1_ASAP7_75t_L g94 ( 
.A(n_36),
.B(n_14),
.Y(n_94)
);

OR2x2_ASAP7_75t_L g167 ( 
.A(n_94),
.B(n_38),
.Y(n_167)
);

BUFx12f_ASAP7_75t_L g95 ( 
.A(n_52),
.Y(n_95)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_95),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_28),
.Y(n_96)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_96),
.Y(n_135)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_50),
.Y(n_97)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_97),
.Y(n_141)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_28),
.Y(n_98)
);

INVx6_ASAP7_75t_L g137 ( 
.A(n_98),
.Y(n_137)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_36),
.Y(n_99)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_99),
.Y(n_185)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_50),
.Y(n_100)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_100),
.Y(n_156)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_34),
.Y(n_101)
);

INVx6_ASAP7_75t_L g140 ( 
.A(n_101),
.Y(n_140)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_53),
.Y(n_102)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_102),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_34),
.Y(n_103)
);

INVx6_ASAP7_75t_L g147 ( 
.A(n_103),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_39),
.B(n_14),
.Y(n_104)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_53),
.Y(n_105)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_105),
.Y(n_188)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_44),
.Y(n_106)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_106),
.Y(n_157)
);

INVx11_ASAP7_75t_L g107 ( 
.A(n_20),
.Y(n_107)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_107),
.Y(n_165)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_19),
.Y(n_108)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_108),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_58),
.B(n_14),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_45),
.Y(n_110)
);

INVx4_ASAP7_75t_L g205 ( 
.A(n_110),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_34),
.Y(n_111)
);

INVx6_ASAP7_75t_L g151 ( 
.A(n_111),
.Y(n_151)
);

INVx11_ASAP7_75t_L g112 ( 
.A(n_20),
.Y(n_112)
);

INVx4_ASAP7_75t_L g206 ( 
.A(n_112),
.Y(n_206)
);

OR2x2_ASAP7_75t_L g113 ( 
.A(n_44),
.B(n_13),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_113),
.B(n_124),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_38),
.B(n_13),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_34),
.Y(n_115)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_115),
.Y(n_195)
);

AND2x4_ASAP7_75t_SL g116 ( 
.A(n_38),
.B(n_0),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_116),
.B(n_0),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_46),
.Y(n_117)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_117),
.Y(n_189)
);

BUFx2_ASAP7_75t_L g118 ( 
.A(n_50),
.Y(n_118)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_118),
.Y(n_197)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_45),
.Y(n_119)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_119),
.Y(n_200)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_45),
.Y(n_120)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_120),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_46),
.Y(n_121)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_121),
.Y(n_176)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_19),
.Y(n_122)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_122),
.Y(n_190)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_55),
.Y(n_123)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_123),
.Y(n_198)
);

BUFx12f_ASAP7_75t_L g124 ( 
.A(n_48),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_46),
.Y(n_125)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_125),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_62),
.A2(n_53),
.B1(n_46),
.B2(n_30),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_129),
.A2(n_158),
.B1(n_159),
.B2(n_192),
.Y(n_277)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_64),
.A2(n_21),
.B1(n_20),
.B2(n_30),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g258 ( 
.A1(n_130),
.A2(n_142),
.B1(n_145),
.B2(n_148),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_72),
.A2(n_21),
.B1(n_30),
.B2(n_33),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_63),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_144),
.B(n_175),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_118),
.A2(n_21),
.B1(n_33),
.B2(n_48),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_70),
.A2(n_33),
.B1(n_60),
.B2(n_48),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_70),
.A2(n_60),
.B1(n_49),
.B2(n_55),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g275 ( 
.A1(n_152),
.A2(n_171),
.B1(n_178),
.B2(n_180),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_L g158 ( 
.A1(n_98),
.A2(n_58),
.B1(n_43),
.B2(n_26),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_101),
.A2(n_57),
.B1(n_60),
.B2(n_47),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_167),
.B(n_81),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_113),
.B(n_57),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_169),
.B(n_196),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_97),
.A2(n_55),
.B1(n_45),
.B2(n_56),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_116),
.B(n_42),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_172),
.B(n_194),
.Y(n_217)
);

OAI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_66),
.A2(n_25),
.B1(n_56),
.B2(n_37),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_173),
.A2(n_191),
.B1(n_125),
.B2(n_121),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_116),
.B(n_42),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_100),
.A2(n_55),
.B1(n_45),
.B2(n_51),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_107),
.A2(n_55),
.B1(n_37),
.B2(n_51),
.Y(n_180)
);

NAND2x1_ASAP7_75t_L g220 ( 
.A(n_183),
.B(n_35),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_96),
.A2(n_32),
.B1(n_47),
.B2(n_43),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_112),
.A2(n_61),
.B1(n_108),
.B2(n_123),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_65),
.A2(n_35),
.B1(n_27),
.B2(n_25),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_193),
.A2(n_85),
.B1(n_76),
.B2(n_78),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_94),
.B(n_32),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_124),
.B(n_26),
.Y(n_196)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_120),
.Y(n_202)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_202),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_124),
.B(n_73),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_203),
.B(n_117),
.Y(n_261)
);

INVx11_ASAP7_75t_L g209 ( 
.A(n_133),
.Y(n_209)
);

INVx4_ASAP7_75t_L g313 ( 
.A(n_209),
.Y(n_313)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_197),
.Y(n_210)
);

INVx3_ASAP7_75t_L g340 ( 
.A(n_210),
.Y(n_340)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_189),
.Y(n_211)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_211),
.Y(n_285)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_136),
.Y(n_212)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_212),
.Y(n_305)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_132),
.Y(n_213)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_213),
.Y(n_316)
);

BUFx3_ASAP7_75t_L g215 ( 
.A(n_179),
.Y(n_215)
);

INVx5_ASAP7_75t_L g287 ( 
.A(n_215),
.Y(n_287)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_146),
.Y(n_216)
);

INVx1_ASAP7_75t_SL g296 ( 
.A(n_216),
.Y(n_296)
);

INVx4_ASAP7_75t_L g218 ( 
.A(n_146),
.Y(n_218)
);

INVx6_ASAP7_75t_L g284 ( 
.A(n_218),
.Y(n_284)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_136),
.Y(n_219)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_219),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_220),
.B(n_230),
.C(n_5),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_174),
.B(n_27),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_221),
.B(n_229),
.Y(n_299)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_143),
.Y(n_222)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_222),
.Y(n_328)
);

OAI21xp33_ASAP7_75t_L g224 ( 
.A1(n_183),
.A2(n_68),
.B(n_13),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_224),
.B(n_226),
.Y(n_310)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_170),
.Y(n_225)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_225),
.Y(n_333)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_139),
.Y(n_227)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_227),
.Y(n_335)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_157),
.Y(n_228)
);

INVx1_ASAP7_75t_SL g308 ( 
.A(n_228),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_149),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_134),
.B(n_122),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_181),
.Y(n_231)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_231),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_128),
.B(n_67),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_232),
.B(n_236),
.Y(n_309)
);

O2A1O1Ixp33_ASAP7_75t_L g233 ( 
.A1(n_154),
.A2(n_73),
.B(n_95),
.C(n_110),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g292 ( 
.A1(n_233),
.A2(n_152),
.B(n_192),
.Y(n_292)
);

INVx3_ASAP7_75t_L g234 ( 
.A(n_160),
.Y(n_234)
);

INVx1_ASAP7_75t_SL g329 ( 
.A(n_234),
.Y(n_329)
);

OAI22xp33_ASAP7_75t_SL g293 ( 
.A1(n_235),
.A2(n_195),
.B1(n_207),
.B2(n_204),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_162),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_166),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_237),
.B(n_239),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_139),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_SL g289 ( 
.A1(n_238),
.A2(n_246),
.B1(n_248),
.B2(n_251),
.Y(n_289)
);

INVx5_ASAP7_75t_L g239 ( 
.A(n_160),
.Y(n_239)
);

INVx2_ASAP7_75t_SL g240 ( 
.A(n_133),
.Y(n_240)
);

AND2x2_ASAP7_75t_L g338 ( 
.A(n_240),
.B(n_249),
.Y(n_338)
);

BUFx3_ASAP7_75t_L g241 ( 
.A(n_179),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_241),
.B(n_243),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_150),
.B(n_95),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g295 ( 
.A(n_242),
.Y(n_295)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_168),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_176),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_244),
.Y(n_301)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_201),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_245),
.Y(n_321)
);

INVx6_ASAP7_75t_L g246 ( 
.A(n_155),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_153),
.B(n_119),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g334 ( 
.A(n_247),
.Y(n_334)
);

INVx6_ASAP7_75t_L g248 ( 
.A(n_155),
.Y(n_248)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_168),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_186),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_250),
.Y(n_306)
);

BUFx3_ASAP7_75t_L g251 ( 
.A(n_163),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_188),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_252),
.Y(n_315)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_161),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_SL g294 ( 
.A1(n_253),
.A2(n_256),
.B1(n_257),
.B2(n_259),
.Y(n_294)
);

INVx3_ASAP7_75t_L g254 ( 
.A(n_205),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_254),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_177),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_255),
.B(n_260),
.Y(n_290)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_182),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_190),
.Y(n_257)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_198),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_167),
.B(n_13),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_261),
.B(n_263),
.Y(n_297)
);

INVx4_ASAP7_75t_L g262 ( 
.A(n_205),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_SL g320 ( 
.A1(n_262),
.A2(n_264),
.B1(n_266),
.B2(n_269),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_184),
.B(n_86),
.Y(n_263)
);

INVx3_ASAP7_75t_L g264 ( 
.A(n_199),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_185),
.B(n_87),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_265),
.B(n_270),
.Y(n_302)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_161),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_SL g342 ( 
.A1(n_267),
.A2(n_11),
.B(n_8),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_145),
.A2(n_92),
.B1(n_80),
.B2(n_103),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_268),
.A2(n_126),
.B1(n_151),
.B2(n_147),
.Y(n_300)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_163),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_141),
.Y(n_270)
);

INVx3_ASAP7_75t_L g271 ( 
.A(n_199),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_271),
.B(n_273),
.Y(n_304)
);

OAI22xp33_ASAP7_75t_SL g272 ( 
.A1(n_130),
.A2(n_115),
.B1(n_111),
.B2(n_59),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_272),
.A2(n_274),
.B1(n_138),
.B2(n_151),
.Y(n_291)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_141),
.Y(n_273)
);

CKINVDCx14_ASAP7_75t_R g274 ( 
.A(n_177),
.Y(n_274)
);

INVx3_ASAP7_75t_L g276 ( 
.A(n_200),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_276),
.B(n_278),
.Y(n_311)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_156),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_127),
.B(n_0),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_279),
.B(n_280),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_173),
.B(n_0),
.Y(n_280)
);

HB1xp67_ASAP7_75t_L g281 ( 
.A(n_156),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_281),
.B(n_282),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_127),
.B(n_1),
.Y(n_282)
);

AOI22xp33_ASAP7_75t_L g283 ( 
.A1(n_195),
.A2(n_59),
.B1(n_2),
.B2(n_3),
.Y(n_283)
);

OAI22xp33_ASAP7_75t_L g286 ( 
.A1(n_283),
.A2(n_180),
.B1(n_142),
.B2(n_193),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_286),
.A2(n_288),
.B1(n_293),
.B2(n_298),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_258),
.A2(n_148),
.B1(n_171),
.B2(n_178),
.Y(n_288)
);

OAI21xp33_ASAP7_75t_SL g348 ( 
.A1(n_291),
.A2(n_209),
.B(n_240),
.Y(n_348)
);

AND2x2_ASAP7_75t_L g375 ( 
.A(n_292),
.B(n_342),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_258),
.A2(n_140),
.B1(n_137),
.B2(n_131),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g386 ( 
.A1(n_300),
.A2(n_314),
.B1(n_324),
.B2(n_302),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_235),
.A2(n_140),
.B1(n_137),
.B2(n_131),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_303),
.A2(n_307),
.B1(n_319),
.B2(n_322),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_275),
.A2(n_126),
.B1(n_135),
.B2(n_147),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_L g312 ( 
.A1(n_208),
.A2(n_138),
.B(n_204),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_L g361 ( 
.A1(n_312),
.A2(n_215),
.B(n_241),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_277),
.A2(n_135),
.B1(n_187),
.B2(n_164),
.Y(n_314)
);

AOI32xp33_ASAP7_75t_L g317 ( 
.A1(n_217),
.A2(n_206),
.A3(n_165),
.B1(n_187),
.B2(n_207),
.Y(n_317)
);

A2O1A1Ixp33_ASAP7_75t_L g365 ( 
.A1(n_317),
.A2(n_262),
.B(n_227),
.C(n_276),
.Y(n_365)
);

OAI22xp33_ASAP7_75t_L g319 ( 
.A1(n_267),
.A2(n_165),
.B1(n_206),
.B2(n_164),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_275),
.A2(n_59),
.B1(n_2),
.B2(n_3),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_SL g323 ( 
.A(n_230),
.B(n_59),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_323),
.B(n_341),
.C(n_254),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_268),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_L g330 ( 
.A1(n_246),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_330),
.A2(n_337),
.B1(n_216),
.B2(n_234),
.Y(n_371)
);

AOI21xp5_ASAP7_75t_L g332 ( 
.A1(n_226),
.A2(n_5),
.B(n_6),
.Y(n_332)
);

AOI21xp5_ASAP7_75t_L g356 ( 
.A1(n_332),
.A2(n_271),
.B(n_264),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_223),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_339),
.B(n_341),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_220),
.B(n_6),
.C(n_7),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_225),
.B(n_7),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_344),
.B(n_345),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_231),
.B(n_9),
.Y(n_345)
);

OR2x4_ASAP7_75t_L g346 ( 
.A(n_224),
.B(n_9),
.Y(n_346)
);

AO21x1_ASAP7_75t_L g347 ( 
.A1(n_346),
.A2(n_233),
.B(n_10),
.Y(n_347)
);

INVxp67_ASAP7_75t_L g417 ( 
.A(n_347),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_348),
.A2(n_352),
.B1(n_364),
.B2(n_386),
.Y(n_411)
);

INVxp67_ASAP7_75t_L g349 ( 
.A(n_318),
.Y(n_349)
);

INVxp67_ASAP7_75t_L g429 ( 
.A(n_349),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_290),
.B(n_214),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_SL g409 ( 
.A(n_351),
.B(n_368),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_314),
.A2(n_256),
.B1(n_211),
.B2(n_248),
.Y(n_352)
);

INVxp67_ASAP7_75t_L g353 ( 
.A(n_318),
.Y(n_353)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_353),
.Y(n_401)
);

AOI22xp33_ASAP7_75t_L g354 ( 
.A1(n_303),
.A2(n_212),
.B1(n_219),
.B2(n_270),
.Y(n_354)
);

CKINVDCx16_ASAP7_75t_R g402 ( 
.A(n_354),
.Y(n_402)
);

INVxp33_ASAP7_75t_L g355 ( 
.A(n_325),
.Y(n_355)
);

CKINVDCx16_ASAP7_75t_R g420 ( 
.A(n_355),
.Y(n_420)
);

OAI21xp5_ASAP7_75t_L g434 ( 
.A1(n_356),
.A2(n_361),
.B(n_390),
.Y(n_434)
);

XNOR2xp5_ASAP7_75t_L g399 ( 
.A(n_357),
.B(n_344),
.Y(n_399)
);

INVx1_ASAP7_75t_SL g358 ( 
.A(n_338),
.Y(n_358)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_358),
.Y(n_407)
);

INVx5_ASAP7_75t_L g359 ( 
.A(n_284),
.Y(n_359)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_359),
.Y(n_410)
);

BUFx2_ASAP7_75t_L g360 ( 
.A(n_335),
.Y(n_360)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_360),
.Y(n_418)
);

NOR2x1_ASAP7_75t_L g362 ( 
.A(n_310),
.B(n_273),
.Y(n_362)
);

AOI21xp5_ASAP7_75t_SL g398 ( 
.A1(n_362),
.A2(n_376),
.B(n_346),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_300),
.A2(n_238),
.B1(n_266),
.B2(n_253),
.Y(n_364)
);

AOI21xp5_ASAP7_75t_L g433 ( 
.A1(n_365),
.A2(n_393),
.B(n_287),
.Y(n_433)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_304),
.Y(n_367)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_367),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_290),
.B(n_269),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_309),
.B(n_218),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_SL g413 ( 
.A(n_369),
.B(n_378),
.Y(n_413)
);

INVx3_ASAP7_75t_L g370 ( 
.A(n_284),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_370),
.B(n_371),
.Y(n_416)
);

AO21x2_ASAP7_75t_L g372 ( 
.A1(n_292),
.A2(n_251),
.B(n_239),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_L g408 ( 
.A1(n_372),
.A2(n_374),
.B1(n_379),
.B2(n_388),
.Y(n_408)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_305),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_373),
.B(n_381),
.Y(n_424)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_298),
.A2(n_11),
.B1(n_9),
.B2(n_10),
.Y(n_374)
);

O2A1O1Ixp33_ASAP7_75t_L g376 ( 
.A1(n_342),
.A2(n_317),
.B(n_291),
.C(n_338),
.Y(n_376)
);

XOR2xp5_ASAP7_75t_L g377 ( 
.A(n_323),
.B(n_339),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_377),
.B(n_321),
.C(n_301),
.Y(n_404)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_304),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_288),
.A2(n_307),
.B1(n_322),
.B2(n_326),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_309),
.B(n_299),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_380),
.B(n_383),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_336),
.B(n_323),
.Y(n_381)
);

XOR2xp5_ASAP7_75t_L g396 ( 
.A(n_382),
.B(n_345),
.Y(n_396)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_311),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_311),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_384),
.B(n_387),
.Y(n_432)
);

BUFx2_ASAP7_75t_L g385 ( 
.A(n_335),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_385),
.Y(n_405)
);

INVxp67_ASAP7_75t_L g387 ( 
.A(n_325),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_326),
.A2(n_336),
.B1(n_310),
.B2(n_297),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_338),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_389),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_299),
.B(n_308),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_310),
.A2(n_297),
.B1(n_302),
.B2(n_312),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_L g422 ( 
.A1(n_391),
.A2(n_327),
.B1(n_296),
.B2(n_329),
.Y(n_422)
);

INVxp67_ASAP7_75t_L g392 ( 
.A(n_332),
.Y(n_392)
);

HAxp5_ASAP7_75t_SL g421 ( 
.A(n_392),
.B(n_331),
.CON(n_421),
.SN(n_421)
);

AOI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_334),
.A2(n_295),
.B1(n_346),
.B2(n_337),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_305),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_394),
.A2(n_296),
.B1(n_329),
.B2(n_313),
.Y(n_400)
);

CKINVDCx16_ASAP7_75t_R g395 ( 
.A(n_294),
.Y(n_395)
);

AOI22xp33_ASAP7_75t_L g397 ( 
.A1(n_395),
.A2(n_329),
.B1(n_296),
.B2(n_313),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_396),
.B(n_399),
.C(n_404),
.Y(n_441)
);

OAI21xp5_ASAP7_75t_SL g443 ( 
.A1(n_397),
.A2(n_398),
.B(n_400),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_SL g403 ( 
.A1(n_379),
.A2(n_324),
.B1(n_289),
.B2(n_308),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g462 ( 
.A1(n_403),
.A2(n_406),
.B1(n_419),
.B2(n_422),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_350),
.A2(n_308),
.B1(n_320),
.B2(n_315),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_SL g412 ( 
.A1(n_375),
.A2(n_330),
.B1(n_306),
.B2(n_315),
.Y(n_412)
);

INVxp67_ASAP7_75t_L g456 ( 
.A(n_412),
.Y(n_456)
);

A2O1A1O1Ixp25_ASAP7_75t_L g414 ( 
.A1(n_381),
.A2(n_327),
.B(n_343),
.C(n_333),
.D(n_285),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_SL g464 ( 
.A(n_414),
.B(n_389),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_377),
.B(n_343),
.C(n_333),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_415),
.B(n_427),
.C(n_404),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_350),
.A2(n_306),
.B1(n_331),
.B2(n_285),
.Y(n_419)
);

CKINVDCx14_ASAP7_75t_R g457 ( 
.A(n_421),
.Y(n_457)
);

AOI22xp33_ASAP7_75t_L g423 ( 
.A1(n_367),
.A2(n_313),
.B1(n_284),
.B2(n_340),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_L g446 ( 
.A1(n_423),
.A2(n_372),
.B1(n_360),
.B2(n_385),
.Y(n_446)
);

XOR2xp5_ASAP7_75t_L g427 ( 
.A(n_357),
.B(n_382),
.Y(n_427)
);

AOI21xp5_ASAP7_75t_SL g430 ( 
.A1(n_375),
.A2(n_316),
.B(n_328),
.Y(n_430)
);

A2O1A1Ixp33_ASAP7_75t_L g472 ( 
.A1(n_430),
.A2(n_347),
.B(n_358),
.C(n_356),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_SL g431 ( 
.A1(n_366),
.A2(n_316),
.B1(n_328),
.B2(n_340),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_431),
.B(n_435),
.Y(n_445)
);

AOI21xp5_ASAP7_75t_L g474 ( 
.A1(n_433),
.A2(n_395),
.B(n_359),
.Y(n_474)
);

OAI22xp5_ASAP7_75t_SL g435 ( 
.A1(n_366),
.A2(n_372),
.B1(n_391),
.B2(n_384),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_L g436 ( 
.A(n_388),
.B(n_363),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_SL g471 ( 
.A(n_436),
.B(n_376),
.Y(n_471)
);

OAI22xp5_ASAP7_75t_SL g437 ( 
.A1(n_372),
.A2(n_287),
.B1(n_383),
.B2(n_378),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_437),
.B(n_386),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_433),
.A2(n_372),
.B1(n_393),
.B2(n_365),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_L g488 ( 
.A1(n_438),
.A2(n_439),
.B1(n_460),
.B2(n_466),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_412),
.A2(n_411),
.B1(n_398),
.B2(n_372),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_432),
.Y(n_440)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_440),
.Y(n_480)
);

XOR2xp5_ASAP7_75t_L g442 ( 
.A(n_427),
.B(n_369),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_442),
.B(n_452),
.C(n_453),
.Y(n_479)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_432),
.Y(n_444)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_444),
.Y(n_484)
);

AND2x2_ASAP7_75t_L g507 ( 
.A(n_446),
.B(n_448),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_426),
.B(n_390),
.Y(n_447)
);

CKINVDCx14_ASAP7_75t_R g492 ( 
.A(n_447),
.Y(n_492)
);

AND2x2_ASAP7_75t_L g448 ( 
.A(n_407),
.B(n_361),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_425),
.Y(n_449)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_449),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_SL g450 ( 
.A(n_428),
.B(n_380),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_SL g477 ( 
.A(n_450),
.B(n_459),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_426),
.B(n_368),
.Y(n_451)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_451),
.Y(n_504)
);

XOR2xp5_ASAP7_75t_L g452 ( 
.A(n_399),
.B(n_375),
.Y(n_452)
);

XOR2xp5_ASAP7_75t_L g453 ( 
.A(n_436),
.B(n_362),
.Y(n_453)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_413),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_454),
.B(n_464),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_455),
.B(n_458),
.C(n_401),
.Y(n_483)
);

XOR2xp5_ASAP7_75t_L g458 ( 
.A(n_396),
.B(n_362),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_SL g459 ( 
.A(n_428),
.B(n_351),
.Y(n_459)
);

OAI22xp5_ASAP7_75t_L g460 ( 
.A1(n_411),
.A2(n_365),
.B1(n_374),
.B2(n_371),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_425),
.Y(n_461)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_461),
.Y(n_485)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_463),
.Y(n_491)
);

XNOR2x1_ASAP7_75t_L g465 ( 
.A(n_424),
.B(n_363),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_SL g482 ( 
.A(n_465),
.B(n_471),
.Y(n_482)
);

OAI22xp33_ASAP7_75t_SL g466 ( 
.A1(n_417),
.A2(n_376),
.B1(n_358),
.B2(n_347),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_413),
.B(n_373),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_467),
.B(n_468),
.Y(n_508)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_423),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_409),
.B(n_401),
.Y(n_469)
);

CKINVDCx20_ASAP7_75t_R g497 ( 
.A(n_469),
.Y(n_497)
);

CKINVDCx16_ASAP7_75t_R g470 ( 
.A(n_422),
.Y(n_470)
);

BUFx10_ASAP7_75t_L g481 ( 
.A(n_470),
.Y(n_481)
);

AOI21xp5_ASAP7_75t_L g510 ( 
.A1(n_472),
.A2(n_474),
.B(n_418),
.Y(n_510)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_419),
.Y(n_473)
);

OAI22xp5_ASAP7_75t_L g499 ( 
.A1(n_473),
.A2(n_420),
.B1(n_434),
.B2(n_416),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_409),
.B(n_394),
.Y(n_475)
);

CKINVDCx16_ASAP7_75t_R g486 ( 
.A(n_475),
.Y(n_486)
);

AOI22x1_ASAP7_75t_SL g476 ( 
.A1(n_438),
.A2(n_435),
.B1(n_437),
.B2(n_406),
.Y(n_476)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_476),
.Y(n_523)
);

XNOR2xp5_ASAP7_75t_L g478 ( 
.A(n_455),
.B(n_415),
.Y(n_478)
);

XOR2xp5_ASAP7_75t_L g517 ( 
.A(n_478),
.B(n_493),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_483),
.B(n_487),
.C(n_496),
.Y(n_511)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_442),
.B(n_424),
.C(n_407),
.Y(n_487)
);

XNOR2xp5_ASAP7_75t_SL g489 ( 
.A(n_452),
.B(n_408),
.Y(n_489)
);

XNOR2xp5_ASAP7_75t_SL g518 ( 
.A(n_489),
.B(n_471),
.Y(n_518)
);

XNOR2xp5_ASAP7_75t_L g493 ( 
.A(n_441),
.B(n_430),
.Y(n_493)
);

XOR2xp5_ASAP7_75t_L g494 ( 
.A(n_441),
.B(n_458),
.Y(n_494)
);

XOR2xp5_ASAP7_75t_L g524 ( 
.A(n_494),
.B(n_501),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_453),
.B(n_430),
.C(n_398),
.Y(n_496)
);

AOI22xp5_ASAP7_75t_L g498 ( 
.A1(n_470),
.A2(n_408),
.B1(n_403),
.B2(n_434),
.Y(n_498)
);

OAI22xp5_ASAP7_75t_SL g516 ( 
.A1(n_498),
.A2(n_502),
.B1(n_503),
.B2(n_445),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_499),
.B(n_456),
.Y(n_522)
);

OAI22xp5_ASAP7_75t_L g500 ( 
.A1(n_462),
.A2(n_429),
.B1(n_420),
.B2(n_416),
.Y(n_500)
);

CKINVDCx16_ASAP7_75t_R g512 ( 
.A(n_500),
.Y(n_512)
);

XNOR2xp5_ASAP7_75t_L g501 ( 
.A(n_471),
.B(n_414),
.Y(n_501)
);

AOI22xp5_ASAP7_75t_L g502 ( 
.A1(n_460),
.A2(n_431),
.B1(n_402),
.B2(n_352),
.Y(n_502)
);

AOI22xp5_ASAP7_75t_L g503 ( 
.A1(n_463),
.A2(n_402),
.B1(n_364),
.B2(n_405),
.Y(n_503)
);

CKINVDCx16_ASAP7_75t_R g505 ( 
.A(n_447),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_SL g514 ( 
.A(n_505),
.B(n_454),
.Y(n_514)
);

OAI22xp5_ASAP7_75t_SL g506 ( 
.A1(n_462),
.A2(n_397),
.B1(n_414),
.B2(n_400),
.Y(n_506)
);

AOI22xp5_ASAP7_75t_L g520 ( 
.A1(n_506),
.A2(n_509),
.B1(n_446),
.B2(n_439),
.Y(n_520)
);

OAI22xp5_ASAP7_75t_SL g509 ( 
.A1(n_473),
.A2(n_405),
.B1(n_418),
.B2(n_410),
.Y(n_509)
);

OAI21xp5_ASAP7_75t_L g526 ( 
.A1(n_510),
.A2(n_474),
.B(n_443),
.Y(n_526)
);

CKINVDCx16_ASAP7_75t_R g513 ( 
.A(n_495),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_513),
.B(n_522),
.Y(n_558)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_514),
.Y(n_548)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_478),
.B(n_483),
.C(n_494),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g562 ( 
.A(n_515),
.B(n_519),
.C(n_521),
.Y(n_562)
);

AOI22xp5_ASAP7_75t_SL g555 ( 
.A1(n_516),
.A2(n_481),
.B1(n_507),
.B2(n_476),
.Y(n_555)
);

XNOR2xp5_ASAP7_75t_SL g547 ( 
.A(n_518),
.B(n_482),
.Y(n_547)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_479),
.B(n_448),
.C(n_465),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_520),
.B(n_527),
.Y(n_546)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_479),
.B(n_448),
.C(n_465),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_SL g525 ( 
.A(n_477),
.B(n_450),
.Y(n_525)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_525),
.Y(n_551)
);

AOI21xp5_ASAP7_75t_L g564 ( 
.A1(n_526),
.A2(n_541),
.B(n_410),
.Y(n_564)
);

AOI22xp5_ASAP7_75t_L g527 ( 
.A1(n_506),
.A2(n_445),
.B1(n_444),
.B2(n_440),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_485),
.Y(n_528)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_528),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_SL g529 ( 
.A(n_504),
.B(n_459),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_SL g550 ( 
.A(n_529),
.B(n_480),
.Y(n_550)
);

AOI22xp5_ASAP7_75t_L g530 ( 
.A1(n_491),
.A2(n_507),
.B1(n_481),
.B2(n_492),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_530),
.B(n_533),
.Y(n_554)
);

OAI22xp5_ASAP7_75t_SL g531 ( 
.A1(n_488),
.A2(n_464),
.B1(n_451),
.B2(n_469),
.Y(n_531)
);

AOI22xp5_ASAP7_75t_L g542 ( 
.A1(n_531),
.A2(n_486),
.B1(n_481),
.B2(n_484),
.Y(n_542)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_485),
.Y(n_532)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_532),
.Y(n_559)
);

AOI22xp5_ASAP7_75t_L g533 ( 
.A1(n_491),
.A2(n_448),
.B1(n_468),
.B2(n_457),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_497),
.B(n_461),
.Y(n_534)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_534),
.Y(n_567)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_508),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g553 ( 
.A(n_535),
.B(n_537),
.Y(n_553)
);

MAJIxp5_ASAP7_75t_L g536 ( 
.A(n_493),
.B(n_475),
.C(n_467),
.Y(n_536)
);

MAJIxp5_ASAP7_75t_L g565 ( 
.A(n_536),
.B(n_538),
.C(n_370),
.Y(n_565)
);

FAx1_ASAP7_75t_SL g537 ( 
.A(n_496),
.B(n_472),
.CI(n_457),
.CON(n_537),
.SN(n_537)
);

MAJIxp5_ASAP7_75t_L g538 ( 
.A(n_487),
.B(n_443),
.C(n_449),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_508),
.Y(n_539)
);

CKINVDCx20_ASAP7_75t_R g566 ( 
.A(n_539),
.Y(n_566)
);

XOR2xp5_ASAP7_75t_L g540 ( 
.A(n_489),
.B(n_472),
.Y(n_540)
);

XOR2xp5_ASAP7_75t_L g552 ( 
.A(n_540),
.B(n_482),
.Y(n_552)
);

CKINVDCx20_ASAP7_75t_R g541 ( 
.A(n_507),
.Y(n_541)
);

OAI22xp5_ASAP7_75t_L g588 ( 
.A1(n_542),
.A2(n_555),
.B1(n_527),
.B2(n_532),
.Y(n_588)
);

XNOR2xp5_ASAP7_75t_L g543 ( 
.A(n_511),
.B(n_498),
.Y(n_543)
);

XNOR2xp5_ASAP7_75t_L g572 ( 
.A(n_543),
.B(n_544),
.Y(n_572)
);

XNOR2xp5_ASAP7_75t_L g544 ( 
.A(n_511),
.B(n_501),
.Y(n_544)
);

XNOR2xp5_ASAP7_75t_L g545 ( 
.A(n_515),
.B(n_488),
.Y(n_545)
);

XNOR2xp5_ASAP7_75t_L g577 ( 
.A(n_545),
.B(n_549),
.Y(n_577)
);

XNOR2xp5_ASAP7_75t_SL g576 ( 
.A(n_547),
.B(n_552),
.Y(n_576)
);

XNOR2xp5_ASAP7_75t_L g549 ( 
.A(n_519),
.B(n_495),
.Y(n_549)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_550),
.Y(n_571)
);

XOR2xp5_ASAP7_75t_L g556 ( 
.A(n_524),
.B(n_510),
.Y(n_556)
);

XNOR2xp5_ASAP7_75t_SL g579 ( 
.A(n_556),
.B(n_540),
.Y(n_579)
);

XNOR2xp5_ASAP7_75t_L g560 ( 
.A(n_521),
.B(n_481),
.Y(n_560)
);

XOR2xp5_ASAP7_75t_L g569 ( 
.A(n_560),
.B(n_561),
.Y(n_569)
);

XNOR2xp5_ASAP7_75t_L g561 ( 
.A(n_538),
.B(n_509),
.Y(n_561)
);

AOI22xp5_ASAP7_75t_SL g563 ( 
.A1(n_523),
.A2(n_490),
.B1(n_502),
.B2(n_503),
.Y(n_563)
);

XOR2xp5_ASAP7_75t_L g578 ( 
.A(n_563),
.B(n_530),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_564),
.B(n_541),
.Y(n_573)
);

MAJIxp5_ASAP7_75t_L g582 ( 
.A(n_565),
.B(n_517),
.C(n_524),
.Y(n_582)
);

FAx1_ASAP7_75t_L g568 ( 
.A(n_553),
.B(n_526),
.CI(n_537),
.CON(n_568),
.SN(n_568)
);

AOI21x1_ASAP7_75t_SL g603 ( 
.A1(n_568),
.A2(n_573),
.B(n_537),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_SL g570 ( 
.A(n_551),
.B(n_525),
.Y(n_570)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_570),
.Y(n_598)
);

NOR2xp33_ASAP7_75t_L g574 ( 
.A(n_548),
.B(n_512),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_574),
.B(n_580),
.Y(n_590)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_557),
.Y(n_575)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_575),
.Y(n_601)
);

XNOR2xp5_ASAP7_75t_L g593 ( 
.A(n_578),
.B(n_579),
.Y(n_593)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_559),
.Y(n_580)
);

AOI22xp5_ASAP7_75t_L g581 ( 
.A1(n_567),
.A2(n_516),
.B1(n_531),
.B2(n_523),
.Y(n_581)
);

OAI22xp5_ASAP7_75t_SL g596 ( 
.A1(n_581),
.A2(n_583),
.B1(n_586),
.B2(n_563),
.Y(n_596)
);

MAJIxp5_ASAP7_75t_L g592 ( 
.A(n_582),
.B(n_587),
.C(n_562),
.Y(n_592)
);

AOI22xp5_ASAP7_75t_L g583 ( 
.A1(n_546),
.A2(n_535),
.B1(n_539),
.B2(n_522),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_558),
.Y(n_584)
);

CKINVDCx20_ASAP7_75t_R g589 ( 
.A(n_584),
.Y(n_589)
);

AOI22xp5_ASAP7_75t_L g585 ( 
.A1(n_546),
.A2(n_534),
.B1(n_536),
.B2(n_520),
.Y(n_585)
);

OAI22xp5_ASAP7_75t_SL g606 ( 
.A1(n_585),
.A2(n_518),
.B1(n_528),
.B2(n_360),
.Y(n_606)
);

CKINVDCx20_ASAP7_75t_R g586 ( 
.A(n_566),
.Y(n_586)
);

MAJIxp5_ASAP7_75t_L g587 ( 
.A(n_543),
.B(n_517),
.C(n_533),
.Y(n_587)
);

AOI22xp5_ASAP7_75t_SL g594 ( 
.A1(n_588),
.A2(n_554),
.B1(n_555),
.B2(n_542),
.Y(n_594)
);

OAI21xp5_ASAP7_75t_L g591 ( 
.A1(n_573),
.A2(n_554),
.B(n_564),
.Y(n_591)
);

AOI21xp5_ASAP7_75t_SL g617 ( 
.A1(n_591),
.A2(n_578),
.B(n_568),
.Y(n_617)
);

XNOR2xp5_ASAP7_75t_L g611 ( 
.A(n_592),
.B(n_600),
.Y(n_611)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_594),
.Y(n_619)
);

AND2x2_ASAP7_75t_L g595 ( 
.A(n_569),
.B(n_549),
.Y(n_595)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_595),
.Y(n_620)
);

OR2x2_ASAP7_75t_L g614 ( 
.A(n_596),
.B(n_603),
.Y(n_614)
);

XNOR2xp5_ASAP7_75t_L g597 ( 
.A(n_577),
.B(n_545),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_597),
.B(n_599),
.Y(n_616)
);

MAJIxp5_ASAP7_75t_L g599 ( 
.A(n_577),
.B(n_565),
.C(n_562),
.Y(n_599)
);

XNOR2xp5_ASAP7_75t_L g600 ( 
.A(n_569),
.B(n_572),
.Y(n_600)
);

MAJIxp5_ASAP7_75t_L g602 ( 
.A(n_572),
.B(n_561),
.C(n_560),
.Y(n_602)
);

MAJIxp5_ASAP7_75t_L g613 ( 
.A(n_602),
.B(n_604),
.C(n_605),
.Y(n_613)
);

MAJIxp5_ASAP7_75t_L g604 ( 
.A(n_582),
.B(n_544),
.C(n_556),
.Y(n_604)
);

MAJIxp5_ASAP7_75t_L g605 ( 
.A(n_587),
.B(n_552),
.C(n_547),
.Y(n_605)
);

INVxp67_ASAP7_75t_L g607 ( 
.A(n_606),
.Y(n_607)
);

XOR2xp5_ASAP7_75t_L g608 ( 
.A(n_597),
.B(n_585),
.Y(n_608)
);

XNOR2xp5_ASAP7_75t_L g623 ( 
.A(n_608),
.B(n_594),
.Y(n_623)
);

CKINVDCx20_ASAP7_75t_R g609 ( 
.A(n_590),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_609),
.B(n_610),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_L g610 ( 
.A(n_589),
.B(n_571),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_L g612 ( 
.A(n_598),
.B(n_599),
.Y(n_612)
);

NOR2xp33_ASAP7_75t_SL g629 ( 
.A(n_612),
.B(n_615),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_SL g615 ( 
.A(n_592),
.B(n_568),
.Y(n_615)
);

XOR2xp5_ASAP7_75t_L g622 ( 
.A(n_617),
.B(n_591),
.Y(n_622)
);

O2A1O1Ixp33_ASAP7_75t_SL g618 ( 
.A1(n_603),
.A2(n_583),
.B(n_581),
.C(n_579),
.Y(n_618)
);

INVxp67_ASAP7_75t_L g625 ( 
.A(n_618),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_SL g621 ( 
.A(n_611),
.B(n_604),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_621),
.B(n_622),
.Y(n_635)
);

XOR2xp5_ASAP7_75t_L g634 ( 
.A(n_623),
.B(n_614),
.Y(n_634)
);

OAI22xp5_ASAP7_75t_SL g624 ( 
.A1(n_619),
.A2(n_601),
.B1(n_602),
.B2(n_605),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_624),
.B(n_626),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_SL g626 ( 
.A(n_616),
.B(n_595),
.Y(n_626)
);

MAJIxp5_ASAP7_75t_L g627 ( 
.A(n_608),
.B(n_600),
.C(n_593),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_SL g637 ( 
.A(n_627),
.B(n_613),
.Y(n_637)
);

NOR2xp67_ASAP7_75t_L g628 ( 
.A(n_620),
.B(n_593),
.Y(n_628)
);

OAI21xp5_ASAP7_75t_SL g632 ( 
.A1(n_628),
.A2(n_625),
.B(n_630),
.Y(n_632)
);

OAI21xp33_ASAP7_75t_L g631 ( 
.A1(n_625),
.A2(n_617),
.B(n_618),
.Y(n_631)
);

OAI31xp33_ASAP7_75t_SL g640 ( 
.A1(n_631),
.A2(n_614),
.A3(n_622),
.B(n_607),
.Y(n_640)
);

AOI21xp5_ASAP7_75t_L g639 ( 
.A1(n_632),
.A2(n_633),
.B(n_627),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_SL g633 ( 
.A(n_629),
.B(n_613),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_634),
.B(n_637),
.Y(n_638)
);

OAI21xp5_ASAP7_75t_L g643 ( 
.A1(n_639),
.A2(n_640),
.B(n_641),
.Y(n_643)
);

MAJIxp5_ASAP7_75t_L g641 ( 
.A(n_635),
.B(n_636),
.C(n_623),
.Y(n_641)
);

INVxp67_ASAP7_75t_L g642 ( 
.A(n_638),
.Y(n_642)
);

MAJIxp5_ASAP7_75t_L g644 ( 
.A(n_642),
.B(n_607),
.C(n_631),
.Y(n_644)
);

BUFx24_ASAP7_75t_SL g645 ( 
.A(n_644),
.Y(n_645)
);

OAI22xp5_ASAP7_75t_L g646 ( 
.A1(n_645),
.A2(n_643),
.B1(n_385),
.B2(n_359),
.Y(n_646)
);

AOI22xp5_ASAP7_75t_L g647 ( 
.A1(n_646),
.A2(n_287),
.B1(n_576),
.B2(n_586),
.Y(n_647)
);


endmodule