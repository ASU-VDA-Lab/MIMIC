module fake_ariane_2105_n_1740 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_148, n_52, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_127, n_35, n_54, n_25, n_1740);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_52;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1740;

wire n_913;
wire n_1681;
wire n_1507;
wire n_1486;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_1682;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_829;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_167;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_645;
wire n_242;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_365;
wire n_238;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1597;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1594;
wire n_680;
wire n_287;
wire n_1716;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_1083;
wire n_967;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_824;
wire n_428;
wire n_159;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_155;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_162;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1163;
wire n_186;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_158;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1304;
wire n_1608;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_1726;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_163;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_321;
wire n_221;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_888;
wire n_845;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_534;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1572;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_157;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_1475;
wire n_642;
wire n_211;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_169;
wire n_1201;
wire n_1288;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_166;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_168;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_683;
wire n_601;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_820;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_161;
wire n_532;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_164;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_1536;
wire n_1471;
wire n_160;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_908;
wire n_788;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1735;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_898;
wire n_857;
wire n_363;
wire n_1067;
wire n_968;
wire n_1323;
wire n_1235;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1727;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1732;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_156;
wire n_174;
wire n_275;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_165;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1233;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_154),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_16),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_34),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_89),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_85),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_98),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_68),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_56),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_129),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_49),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_80),
.Y(n_165)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_126),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_119),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_152),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_100),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_18),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_26),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_137),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_59),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_141),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_95),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_14),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_83),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_84),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_90),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_107),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_91),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_22),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_49),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_53),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_40),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_117),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_103),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_45),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_127),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_48),
.Y(n_190)
);

BUFx10_ASAP7_75t_L g191 ( 
.A(n_144),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_55),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_150),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_112),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_108),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_33),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_21),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_21),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_5),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_149),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_148),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_62),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_114),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_69),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_53),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_63),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_60),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_37),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_29),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_1),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_118),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_18),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_78),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_143),
.Y(n_214)
);

INVx2_ASAP7_75t_SL g215 ( 
.A(n_134),
.Y(n_215)
);

CKINVDCx14_ASAP7_75t_R g216 ( 
.A(n_86),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_4),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_151),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_146),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_111),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_120),
.Y(n_221)
);

INVx2_ASAP7_75t_SL g222 ( 
.A(n_70),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_99),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_123),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_109),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_7),
.Y(n_226)
);

BUFx2_ASAP7_75t_L g227 ( 
.A(n_1),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_122),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_66),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_67),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_5),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_72),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_73),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_14),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_47),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_27),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_128),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_33),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_82),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_71),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_97),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_57),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_136),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_133),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_145),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_92),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_8),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_44),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_23),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_88),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_76),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_24),
.Y(n_252)
);

BUFx10_ASAP7_75t_L g253 ( 
.A(n_3),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_47),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_87),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_102),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_105),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_20),
.Y(n_258)
);

CKINVDCx14_ASAP7_75t_R g259 ( 
.A(n_25),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_110),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_37),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_96),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_74),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_124),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_54),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_16),
.Y(n_266)
);

HB1xp67_ASAP7_75t_L g267 ( 
.A(n_46),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_48),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_44),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_32),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_77),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_6),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_138),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_75),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_64),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_125),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_153),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_20),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_43),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_52),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_23),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_11),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_132),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_131),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_4),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_25),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_106),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_50),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_42),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_8),
.Y(n_290)
);

BUFx10_ASAP7_75t_L g291 ( 
.A(n_24),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_65),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_12),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_6),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_36),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_139),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_42),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_140),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_130),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_28),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_45),
.Y(n_301)
);

BUFx10_ASAP7_75t_L g302 ( 
.A(n_116),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_22),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_35),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_12),
.Y(n_305)
);

BUFx2_ASAP7_75t_L g306 ( 
.A(n_51),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_121),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_147),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_159),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_159),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_161),
.Y(n_311)
);

NOR2xp67_ASAP7_75t_L g312 ( 
.A(n_166),
.B(n_0),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_172),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_259),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_161),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_R g316 ( 
.A(n_216),
.B(n_142),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_203),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_162),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_162),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_219),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_165),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_246),
.Y(n_322)
);

CKINVDCx16_ASAP7_75t_R g323 ( 
.A(n_191),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_250),
.Y(n_324)
);

CKINVDCx16_ASAP7_75t_R g325 ( 
.A(n_191),
.Y(n_325)
);

BUFx3_ASAP7_75t_L g326 ( 
.A(n_166),
.Y(n_326)
);

NOR2xp67_ASAP7_75t_L g327 ( 
.A(n_166),
.B(n_0),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g328 ( 
.A(n_227),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_255),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_275),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_165),
.B(n_167),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_157),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_167),
.B(n_2),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_168),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_168),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_170),
.Y(n_336)
);

INVxp67_ASAP7_75t_SL g337 ( 
.A(n_156),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_175),
.B(n_2),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_175),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_181),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_171),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_181),
.B(n_3),
.Y(n_342)
);

INVxp67_ASAP7_75t_SL g343 ( 
.A(n_156),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_176),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_182),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_192),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_192),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_214),
.B(n_7),
.Y(n_348)
);

AND2x2_ASAP7_75t_L g349 ( 
.A(n_227),
.B(n_9),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_164),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_214),
.Y(n_351)
);

NOR2xp67_ASAP7_75t_L g352 ( 
.A(n_267),
.B(n_9),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_185),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_220),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_220),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_272),
.Y(n_356)
);

HB1xp67_ASAP7_75t_L g357 ( 
.A(n_306),
.Y(n_357)
);

INVx1_ASAP7_75t_SL g358 ( 
.A(n_306),
.Y(n_358)
);

INVx3_ASAP7_75t_L g359 ( 
.A(n_191),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_188),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_290),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_224),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_295),
.Y(n_363)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_224),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_228),
.Y(n_365)
);

AND2x2_ASAP7_75t_L g366 ( 
.A(n_253),
.B(n_10),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_198),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_199),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_297),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_210),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_228),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_237),
.B(n_10),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_237),
.Y(n_373)
);

HB1xp67_ASAP7_75t_L g374 ( 
.A(n_183),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_244),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_226),
.Y(n_376)
);

INVxp67_ASAP7_75t_SL g377 ( 
.A(n_183),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_231),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_244),
.Y(n_379)
);

BUFx6f_ASAP7_75t_L g380 ( 
.A(n_326),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_326),
.B(n_359),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_359),
.B(n_260),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_311),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_311),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_311),
.Y(n_385)
);

HB1xp67_ASAP7_75t_L g386 ( 
.A(n_358),
.Y(n_386)
);

INVxp67_ASAP7_75t_L g387 ( 
.A(n_358),
.Y(n_387)
);

BUFx6f_ASAP7_75t_L g388 ( 
.A(n_326),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_315),
.Y(n_389)
);

BUFx6f_ASAP7_75t_L g390 ( 
.A(n_315),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_359),
.B(n_260),
.Y(n_391)
);

INVx3_ASAP7_75t_L g392 ( 
.A(n_315),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_359),
.B(n_273),
.Y(n_393)
);

NAND2xp33_ASAP7_75t_SL g394 ( 
.A(n_366),
.B(n_197),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_364),
.Y(n_395)
);

INVx2_ASAP7_75t_SL g396 ( 
.A(n_364),
.Y(n_396)
);

BUFx6f_ASAP7_75t_L g397 ( 
.A(n_364),
.Y(n_397)
);

INVx3_ASAP7_75t_L g398 ( 
.A(n_375),
.Y(n_398)
);

INVx3_ASAP7_75t_L g399 ( 
.A(n_375),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_375),
.Y(n_400)
);

AND2x2_ASAP7_75t_L g401 ( 
.A(n_309),
.B(n_197),
.Y(n_401)
);

INVx3_ASAP7_75t_L g402 ( 
.A(n_309),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_310),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_310),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_331),
.B(n_273),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_318),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_318),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_319),
.B(n_274),
.Y(n_408)
);

NOR3xp33_ASAP7_75t_L g409 ( 
.A(n_342),
.B(n_190),
.C(n_184),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_319),
.B(n_274),
.Y(n_410)
);

HB1xp67_ASAP7_75t_L g411 ( 
.A(n_357),
.Y(n_411)
);

HB1xp67_ASAP7_75t_L g412 ( 
.A(n_357),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_321),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_321),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_334),
.Y(n_415)
);

AND2x2_ASAP7_75t_L g416 ( 
.A(n_334),
.B(n_212),
.Y(n_416)
);

BUFx8_ASAP7_75t_L g417 ( 
.A(n_366),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_335),
.Y(n_418)
);

INVx3_ASAP7_75t_L g419 ( 
.A(n_335),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_339),
.B(n_200),
.Y(n_420)
);

INVx3_ASAP7_75t_L g421 ( 
.A(n_339),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_340),
.B(n_202),
.Y(n_422)
);

HB1xp67_ASAP7_75t_L g423 ( 
.A(n_328),
.Y(n_423)
);

AND2x2_ASAP7_75t_L g424 ( 
.A(n_340),
.B(n_212),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_346),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_346),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_347),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_316),
.B(n_191),
.Y(n_428)
);

AND2x4_ASAP7_75t_L g429 ( 
.A(n_347),
.B(n_184),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_351),
.Y(n_430)
);

AND2x4_ASAP7_75t_L g431 ( 
.A(n_351),
.B(n_190),
.Y(n_431)
);

INVx3_ASAP7_75t_L g432 ( 
.A(n_354),
.Y(n_432)
);

AND2x2_ASAP7_75t_L g433 ( 
.A(n_354),
.B(n_302),
.Y(n_433)
);

BUFx2_ASAP7_75t_L g434 ( 
.A(n_332),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_323),
.B(n_302),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_355),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_355),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_362),
.Y(n_438)
);

BUFx6f_ASAP7_75t_L g439 ( 
.A(n_362),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_365),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_365),
.B(n_206),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_371),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_371),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_373),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_428),
.B(n_323),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_434),
.B(n_325),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_433),
.B(n_325),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_SL g448 ( 
.A(n_434),
.B(n_336),
.Y(n_448)
);

AND2x2_ASAP7_75t_L g449 ( 
.A(n_433),
.B(n_349),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_428),
.B(n_341),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_439),
.Y(n_451)
);

INVx4_ASAP7_75t_L g452 ( 
.A(n_380),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_390),
.Y(n_453)
);

BUFx3_ASAP7_75t_L g454 ( 
.A(n_380),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_390),
.Y(n_455)
);

AND2x6_ASAP7_75t_L g456 ( 
.A(n_433),
.B(n_349),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_439),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_439),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g459 ( 
.A(n_434),
.B(n_344),
.Y(n_459)
);

INVx3_ASAP7_75t_L g460 ( 
.A(n_380),
.Y(n_460)
);

NAND2xp33_ASAP7_75t_L g461 ( 
.A(n_405),
.B(n_381),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_387),
.B(n_345),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g463 ( 
.A(n_387),
.B(n_353),
.Y(n_463)
);

BUFx6f_ASAP7_75t_L g464 ( 
.A(n_390),
.Y(n_464)
);

AND2x2_ASAP7_75t_SL g465 ( 
.A(n_409),
.B(n_342),
.Y(n_465)
);

INVx3_ASAP7_75t_L g466 ( 
.A(n_380),
.Y(n_466)
);

INVx3_ASAP7_75t_L g467 ( 
.A(n_380),
.Y(n_467)
);

INVx3_ASAP7_75t_L g468 ( 
.A(n_380),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_L g469 ( 
.A1(n_405),
.A2(n_328),
.B1(n_312),
.B2(n_327),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_439),
.Y(n_470)
);

CKINVDCx20_ASAP7_75t_R g471 ( 
.A(n_386),
.Y(n_471)
);

INVx4_ASAP7_75t_L g472 ( 
.A(n_380),
.Y(n_472)
);

INVx2_ASAP7_75t_SL g473 ( 
.A(n_386),
.Y(n_473)
);

AND2x2_ASAP7_75t_L g474 ( 
.A(n_401),
.B(n_337),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_439),
.Y(n_475)
);

INVx3_ASAP7_75t_L g476 ( 
.A(n_380),
.Y(n_476)
);

BUFx3_ASAP7_75t_L g477 ( 
.A(n_380),
.Y(n_477)
);

INVx3_ASAP7_75t_L g478 ( 
.A(n_388),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_SL g479 ( 
.A(n_435),
.B(n_360),
.Y(n_479)
);

BUFx4f_ASAP7_75t_L g480 ( 
.A(n_390),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_390),
.Y(n_481)
);

XNOR2xp5_ASAP7_75t_L g482 ( 
.A(n_435),
.B(n_350),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_439),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_439),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_SL g485 ( 
.A(n_409),
.B(n_367),
.Y(n_485)
);

NAND3xp33_ASAP7_75t_L g486 ( 
.A(n_394),
.B(n_370),
.C(n_368),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_439),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_381),
.B(n_376),
.Y(n_488)
);

INVx3_ASAP7_75t_L g489 ( 
.A(n_388),
.Y(n_489)
);

INVx3_ASAP7_75t_L g490 ( 
.A(n_388),
.Y(n_490)
);

NOR2x1p5_ASAP7_75t_L g491 ( 
.A(n_408),
.B(n_337),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_390),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_439),
.Y(n_493)
);

BUFx6f_ASAP7_75t_L g494 ( 
.A(n_390),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_389),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_389),
.Y(n_496)
);

INVx1_ASAP7_75t_SL g497 ( 
.A(n_423),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_389),
.Y(n_498)
);

AOI22xp33_ASAP7_75t_L g499 ( 
.A1(n_394),
.A2(n_417),
.B1(n_338),
.B2(n_348),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_389),
.Y(n_500)
);

XNOR2xp5_ASAP7_75t_L g501 ( 
.A(n_411),
.B(n_356),
.Y(n_501)
);

INVx3_ASAP7_75t_L g502 ( 
.A(n_388),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_390),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_395),
.Y(n_504)
);

BUFx6f_ASAP7_75t_L g505 ( 
.A(n_390),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_397),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_397),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_382),
.B(n_378),
.Y(n_508)
);

INVx3_ASAP7_75t_L g509 ( 
.A(n_388),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_382),
.B(n_373),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_395),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_395),
.Y(n_512)
);

NOR2x1p5_ASAP7_75t_L g513 ( 
.A(n_408),
.B(n_343),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_SL g514 ( 
.A(n_391),
.B(n_393),
.Y(n_514)
);

INVx6_ASAP7_75t_L g515 ( 
.A(n_388),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_SL g516 ( 
.A(n_391),
.B(n_313),
.Y(n_516)
);

INVx1_ASAP7_75t_SL g517 ( 
.A(n_423),
.Y(n_517)
);

INVx1_ASAP7_75t_SL g518 ( 
.A(n_411),
.Y(n_518)
);

AND2x2_ASAP7_75t_L g519 ( 
.A(n_401),
.B(n_343),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_397),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_397),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_395),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_393),
.B(n_379),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_403),
.B(n_314),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_397),
.Y(n_525)
);

INVx3_ASAP7_75t_L g526 ( 
.A(n_388),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_383),
.Y(n_527)
);

INVx2_ASAP7_75t_SL g528 ( 
.A(n_417),
.Y(n_528)
);

AND2x2_ASAP7_75t_L g529 ( 
.A(n_401),
.B(n_377),
.Y(n_529)
);

AOI22xp33_ASAP7_75t_L g530 ( 
.A1(n_417),
.A2(n_333),
.B1(n_372),
.B2(n_352),
.Y(n_530)
);

AND2x6_ASAP7_75t_L g531 ( 
.A(n_429),
.B(n_379),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_412),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_397),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_SL g534 ( 
.A(n_429),
.B(n_317),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_397),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_383),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_384),
.Y(n_537)
);

BUFx3_ASAP7_75t_L g538 ( 
.A(n_388),
.Y(n_538)
);

INVx3_ASAP7_75t_L g539 ( 
.A(n_388),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_412),
.Y(n_540)
);

HB1xp67_ASAP7_75t_L g541 ( 
.A(n_416),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_403),
.B(n_377),
.Y(n_542)
);

AND2x2_ASAP7_75t_L g543 ( 
.A(n_416),
.B(n_374),
.Y(n_543)
);

BUFx3_ASAP7_75t_L g544 ( 
.A(n_402),
.Y(n_544)
);

INVx5_ASAP7_75t_L g545 ( 
.A(n_397),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_402),
.B(n_312),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_384),
.Y(n_547)
);

AND2x2_ASAP7_75t_L g548 ( 
.A(n_416),
.B(n_374),
.Y(n_548)
);

INVxp67_ASAP7_75t_SL g549 ( 
.A(n_417),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_402),
.B(n_327),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_397),
.Y(n_551)
);

INVx5_ASAP7_75t_L g552 ( 
.A(n_402),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_384),
.Y(n_553)
);

AOI21x1_ASAP7_75t_L g554 ( 
.A1(n_385),
.A2(n_256),
.B(n_207),
.Y(n_554)
);

BUFx4f_ASAP7_75t_L g555 ( 
.A(n_402),
.Y(n_555)
);

OAI22xp5_ASAP7_75t_L g556 ( 
.A1(n_403),
.A2(n_352),
.B1(n_249),
.B2(n_238),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_392),
.Y(n_557)
);

INVx2_ASAP7_75t_SL g558 ( 
.A(n_417),
.Y(n_558)
);

INVx4_ASAP7_75t_L g559 ( 
.A(n_402),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_385),
.Y(n_560)
);

AOI22xp33_ASAP7_75t_L g561 ( 
.A1(n_417),
.A2(n_270),
.B1(n_289),
.B2(n_235),
.Y(n_561)
);

INVxp67_ASAP7_75t_L g562 ( 
.A(n_424),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_SL g563 ( 
.A(n_424),
.B(n_320),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_392),
.Y(n_564)
);

AND2x4_ASAP7_75t_L g565 ( 
.A(n_429),
.B(n_217),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_385),
.Y(n_566)
);

INVx5_ASAP7_75t_L g567 ( 
.A(n_419),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_419),
.B(n_215),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_400),
.Y(n_569)
);

NOR2xp33_ASAP7_75t_L g570 ( 
.A(n_444),
.B(n_322),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_400),
.Y(n_571)
);

INVx3_ASAP7_75t_L g572 ( 
.A(n_419),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_419),
.B(n_215),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_419),
.B(n_222),
.Y(n_574)
);

BUFx2_ASAP7_75t_L g575 ( 
.A(n_429),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_392),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_392),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_400),
.Y(n_578)
);

INVx3_ASAP7_75t_L g579 ( 
.A(n_419),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_392),
.Y(n_580)
);

INVx3_ASAP7_75t_L g581 ( 
.A(n_421),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_421),
.Y(n_582)
);

INVx5_ASAP7_75t_L g583 ( 
.A(n_421),
.Y(n_583)
);

AND2x6_ASAP7_75t_L g584 ( 
.A(n_429),
.B(n_217),
.Y(n_584)
);

AOI22xp33_ASAP7_75t_L g585 ( 
.A1(n_429),
.A2(n_289),
.B1(n_266),
.B2(n_261),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_421),
.B(n_222),
.Y(n_586)
);

BUFx2_ASAP7_75t_L g587 ( 
.A(n_431),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_421),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_392),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_421),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_398),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_508),
.B(n_432),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_488),
.B(n_432),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_542),
.B(n_456),
.Y(n_594)
);

AND2x4_ASAP7_75t_L g595 ( 
.A(n_474),
.B(n_431),
.Y(n_595)
);

NOR2xp33_ASAP7_75t_L g596 ( 
.A(n_447),
.B(n_432),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_456),
.B(n_449),
.Y(n_597)
);

NOR2xp33_ASAP7_75t_L g598 ( 
.A(n_445),
.B(n_432),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_527),
.Y(n_599)
);

AOI22xp5_ASAP7_75t_L g600 ( 
.A1(n_456),
.A2(n_396),
.B1(n_431),
.B2(n_442),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_L g601 ( 
.A(n_516),
.B(n_432),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_456),
.B(n_432),
.Y(n_602)
);

INVx3_ASAP7_75t_L g603 ( 
.A(n_544),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_456),
.B(n_406),
.Y(n_604)
);

INVx2_ASAP7_75t_SL g605 ( 
.A(n_473),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_456),
.B(n_406),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_456),
.B(n_406),
.Y(n_607)
);

INVx4_ASAP7_75t_L g608 ( 
.A(n_531),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_527),
.Y(n_609)
);

NAND3xp33_ASAP7_75t_L g610 ( 
.A(n_570),
.B(n_324),
.C(n_413),
.Y(n_610)
);

NOR2xp67_ASAP7_75t_L g611 ( 
.A(n_473),
.B(n_396),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_495),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_495),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_496),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_449),
.B(n_413),
.Y(n_615)
);

AND2x4_ASAP7_75t_L g616 ( 
.A(n_474),
.B(n_431),
.Y(n_616)
);

NOR2xp67_ASAP7_75t_L g617 ( 
.A(n_450),
.B(n_396),
.Y(n_617)
);

AND2x6_ASAP7_75t_SL g618 ( 
.A(n_524),
.B(n_234),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_491),
.B(n_415),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_SL g620 ( 
.A(n_555),
.B(n_415),
.Y(n_620)
);

INVx1_ASAP7_75t_SL g621 ( 
.A(n_471),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_SL g622 ( 
.A(n_575),
.B(n_431),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_SL g623 ( 
.A(n_575),
.B(n_431),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_SL g624 ( 
.A(n_587),
.B(n_465),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_SL g625 ( 
.A(n_555),
.B(n_415),
.Y(n_625)
);

INVx4_ASAP7_75t_L g626 ( 
.A(n_531),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_513),
.B(n_418),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g628 ( 
.A(n_485),
.B(n_418),
.Y(n_628)
);

INVxp67_ASAP7_75t_L g629 ( 
.A(n_497),
.Y(n_629)
);

A2O1A1Ixp33_ASAP7_75t_L g630 ( 
.A1(n_465),
.A2(n_444),
.B(n_418),
.C(n_442),
.Y(n_630)
);

INVx3_ASAP7_75t_L g631 ( 
.A(n_544),
.Y(n_631)
);

INVx8_ASAP7_75t_L g632 ( 
.A(n_531),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_496),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_513),
.B(n_426),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_498),
.Y(n_635)
);

AOI22xp33_ASAP7_75t_L g636 ( 
.A1(n_465),
.A2(n_396),
.B1(n_443),
.B2(n_404),
.Y(n_636)
);

INVx3_ASAP7_75t_L g637 ( 
.A(n_544),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_587),
.B(n_426),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_498),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_510),
.B(n_426),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_536),
.Y(n_641)
);

INVx2_ASAP7_75t_SL g642 ( 
.A(n_517),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_SL g643 ( 
.A(n_555),
.B(n_430),
.Y(n_643)
);

NOR2x1_ASAP7_75t_L g644 ( 
.A(n_486),
.B(n_420),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_500),
.Y(n_645)
);

BUFx6f_ASAP7_75t_L g646 ( 
.A(n_454),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_523),
.B(n_430),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_519),
.B(n_430),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_L g649 ( 
.A(n_479),
.B(n_437),
.Y(n_649)
);

AOI22xp33_ASAP7_75t_L g650 ( 
.A1(n_561),
.A2(n_425),
.B1(n_443),
.B2(n_404),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_536),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_519),
.B(n_437),
.Y(n_652)
);

NOR2xp33_ASAP7_75t_L g653 ( 
.A(n_562),
.B(n_437),
.Y(n_653)
);

OR2x2_ASAP7_75t_L g654 ( 
.A(n_518),
.B(n_424),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_500),
.Y(n_655)
);

NOR2xp33_ASAP7_75t_L g656 ( 
.A(n_534),
.B(n_438),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_SL g657 ( 
.A(n_462),
.B(n_438),
.Y(n_657)
);

NOR2xp33_ASAP7_75t_L g658 ( 
.A(n_541),
.B(n_438),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_529),
.B(n_440),
.Y(n_659)
);

BUFx3_ASAP7_75t_L g660 ( 
.A(n_543),
.Y(n_660)
);

AOI22x1_ASAP7_75t_L g661 ( 
.A1(n_559),
.A2(n_444),
.B1(n_440),
.B2(n_442),
.Y(n_661)
);

NAND2x1_ASAP7_75t_L g662 ( 
.A(n_531),
.B(n_440),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_529),
.B(n_514),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_461),
.B(n_404),
.Y(n_664)
);

AND2x2_ASAP7_75t_L g665 ( 
.A(n_543),
.B(n_329),
.Y(n_665)
);

INVx3_ASAP7_75t_L g666 ( 
.A(n_559),
.Y(n_666)
);

BUFx4f_ASAP7_75t_L g667 ( 
.A(n_584),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_537),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_537),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_547),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_565),
.B(n_404),
.Y(n_671)
);

INVxp67_ASAP7_75t_L g672 ( 
.A(n_563),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_547),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_553),
.Y(n_674)
);

AOI22xp5_ASAP7_75t_L g675 ( 
.A1(n_499),
.A2(n_441),
.B1(n_420),
.B2(n_422),
.Y(n_675)
);

BUFx6f_ASAP7_75t_L g676 ( 
.A(n_454),
.Y(n_676)
);

AO22x2_ASAP7_75t_L g677 ( 
.A1(n_469),
.A2(n_549),
.B1(n_558),
.B2(n_528),
.Y(n_677)
);

BUFx6f_ASAP7_75t_L g678 ( 
.A(n_454),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_565),
.B(n_407),
.Y(n_679)
);

NOR2xp33_ASAP7_75t_L g680 ( 
.A(n_559),
.B(n_422),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_565),
.B(n_407),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_565),
.B(n_407),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_572),
.B(n_407),
.Y(n_683)
);

NOR2xp33_ASAP7_75t_SL g684 ( 
.A(n_532),
.B(n_330),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_SL g685 ( 
.A(n_555),
.B(n_559),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_572),
.B(n_414),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_553),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_504),
.Y(n_688)
);

BUFx6f_ASAP7_75t_L g689 ( 
.A(n_477),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_560),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_572),
.B(n_414),
.Y(n_691)
);

NOR2xp67_ASAP7_75t_L g692 ( 
.A(n_463),
.B(n_448),
.Y(n_692)
);

BUFx6f_ASAP7_75t_L g693 ( 
.A(n_477),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_504),
.Y(n_694)
);

AND2x2_ASAP7_75t_L g695 ( 
.A(n_548),
.B(n_361),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_560),
.Y(n_696)
);

INVxp67_ASAP7_75t_L g697 ( 
.A(n_501),
.Y(n_697)
);

AOI22xp5_ASAP7_75t_L g698 ( 
.A1(n_530),
.A2(n_441),
.B1(n_410),
.B2(n_436),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_572),
.B(n_414),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_511),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_579),
.B(n_414),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_SL g702 ( 
.A(n_552),
.B(n_425),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_579),
.B(n_425),
.Y(n_703)
);

INVxp33_ASAP7_75t_L g704 ( 
.A(n_501),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_566),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_566),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_569),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_569),
.Y(n_708)
);

A2O1A1Ixp33_ASAP7_75t_L g709 ( 
.A1(n_579),
.A2(n_581),
.B(n_588),
.C(n_582),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_579),
.B(n_425),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_581),
.B(n_427),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_581),
.B(n_427),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_511),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_SL g714 ( 
.A(n_552),
.B(n_427),
.Y(n_714)
);

NAND2xp33_ASAP7_75t_L g715 ( 
.A(n_531),
.B(n_427),
.Y(n_715)
);

INVx4_ASAP7_75t_L g716 ( 
.A(n_531),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_581),
.B(n_436),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_531),
.B(n_436),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_571),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_571),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_584),
.B(n_548),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_578),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_584),
.B(n_436),
.Y(n_723)
);

INVxp67_ASAP7_75t_L g724 ( 
.A(n_540),
.Y(n_724)
);

OAI22xp5_ASAP7_75t_L g725 ( 
.A1(n_582),
.A2(n_590),
.B1(n_588),
.B2(n_550),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_584),
.B(n_443),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_512),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_SL g728 ( 
.A(n_552),
.B(n_443),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_584),
.B(n_410),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_578),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_SL g731 ( 
.A(n_552),
.B(n_398),
.Y(n_731)
);

O2A1O1Ixp5_ASAP7_75t_L g732 ( 
.A1(n_546),
.A2(n_399),
.B(n_398),
.C(n_270),
.Y(n_732)
);

NOR2xp33_ASAP7_75t_L g733 ( 
.A(n_446),
.B(n_398),
.Y(n_733)
);

BUFx2_ASAP7_75t_L g734 ( 
.A(n_584),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_590),
.Y(n_735)
);

AOI22xp33_ASAP7_75t_L g736 ( 
.A1(n_584),
.A2(n_399),
.B1(n_398),
.B2(n_279),
.Y(n_736)
);

AND2x2_ASAP7_75t_L g737 ( 
.A(n_459),
.B(n_363),
.Y(n_737)
);

INVx3_ASAP7_75t_L g738 ( 
.A(n_557),
.Y(n_738)
);

O2A1O1Ixp33_ASAP7_75t_L g739 ( 
.A1(n_568),
.A2(n_235),
.B(n_279),
.C(n_266),
.Y(n_739)
);

O2A1O1Ixp33_ASAP7_75t_L g740 ( 
.A1(n_573),
.A2(n_278),
.B(n_281),
.C(n_261),
.Y(n_740)
);

AOI22xp5_ASAP7_75t_L g741 ( 
.A1(n_528),
.A2(n_179),
.B1(n_399),
.B2(n_398),
.Y(n_741)
);

OAI22xp5_ASAP7_75t_SL g742 ( 
.A1(n_482),
.A2(n_369),
.B1(n_254),
.B2(n_288),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_564),
.Y(n_743)
);

BUFx6f_ASAP7_75t_L g744 ( 
.A(n_477),
.Y(n_744)
);

BUFx6f_ASAP7_75t_L g745 ( 
.A(n_538),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_564),
.B(n_399),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_576),
.B(n_399),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_576),
.Y(n_748)
);

OR2x2_ASAP7_75t_L g749 ( 
.A(n_482),
.B(n_399),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_577),
.Y(n_750)
);

NOR2xp33_ASAP7_75t_L g751 ( 
.A(n_558),
.B(n_552),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_SL g752 ( 
.A(n_552),
.B(n_155),
.Y(n_752)
);

AO22x2_ASAP7_75t_L g753 ( 
.A1(n_556),
.A2(n_234),
.B1(n_248),
.B2(n_278),
.Y(n_753)
);

NAND2xp33_ASAP7_75t_L g754 ( 
.A(n_567),
.B(n_236),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_577),
.B(n_248),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_580),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_SL g757 ( 
.A(n_567),
.B(n_158),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_512),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_580),
.B(n_281),
.Y(n_759)
);

NOR2xp33_ASAP7_75t_L g760 ( 
.A(n_567),
.B(n_247),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_612),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_613),
.Y(n_762)
);

AOI21x1_ASAP7_75t_L g763 ( 
.A1(n_620),
.A2(n_586),
.B(n_574),
.Y(n_763)
);

OAI321xp33_ASAP7_75t_L g764 ( 
.A1(n_675),
.A2(n_585),
.A3(n_304),
.B1(n_282),
.B2(n_209),
.C(n_205),
.Y(n_764)
);

CKINVDCx10_ASAP7_75t_R g765 ( 
.A(n_684),
.Y(n_765)
);

NAND2x1p5_ASAP7_75t_L g766 ( 
.A(n_608),
.B(n_567),
.Y(n_766)
);

AOI21xp5_ASAP7_75t_L g767 ( 
.A1(n_680),
.A2(n_480),
.B(n_472),
.Y(n_767)
);

OAI21x1_ASAP7_75t_L g768 ( 
.A1(n_661),
.A2(n_455),
.B(n_453),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_595),
.B(n_522),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_614),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_595),
.B(n_522),
.Y(n_771)
);

A2O1A1Ixp33_ASAP7_75t_L g772 ( 
.A1(n_598),
.A2(n_591),
.B(n_589),
.C(n_557),
.Y(n_772)
);

AOI21xp5_ASAP7_75t_L g773 ( 
.A1(n_680),
.A2(n_593),
.B(n_592),
.Y(n_773)
);

AOI21xp5_ASAP7_75t_L g774 ( 
.A1(n_685),
.A2(n_480),
.B(n_472),
.Y(n_774)
);

AOI21xp5_ASAP7_75t_L g775 ( 
.A1(n_685),
.A2(n_480),
.B(n_472),
.Y(n_775)
);

OAI321xp33_ASAP7_75t_L g776 ( 
.A1(n_598),
.A2(n_282),
.A3(n_304),
.B1(n_258),
.B2(n_196),
.C(n_303),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_SL g777 ( 
.A(n_608),
.B(n_567),
.Y(n_777)
);

OAI21xp5_ASAP7_75t_L g778 ( 
.A1(n_709),
.A2(n_480),
.B(n_457),
.Y(n_778)
);

INVx4_ASAP7_75t_L g779 ( 
.A(n_632),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_616),
.B(n_557),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_599),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_633),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_SL g783 ( 
.A(n_626),
.B(n_567),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_609),
.Y(n_784)
);

INVx4_ASAP7_75t_L g785 ( 
.A(n_632),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_616),
.B(n_589),
.Y(n_786)
);

AOI22xp5_ASAP7_75t_L g787 ( 
.A1(n_624),
.A2(n_583),
.B1(n_589),
.B2(n_591),
.Y(n_787)
);

A2O1A1Ixp33_ASAP7_75t_L g788 ( 
.A1(n_653),
.A2(n_591),
.B(n_208),
.C(n_458),
.Y(n_788)
);

OAI21xp33_ASAP7_75t_L g789 ( 
.A1(n_628),
.A2(n_268),
.B(n_252),
.Y(n_789)
);

O2A1O1Ixp33_ASAP7_75t_L g790 ( 
.A1(n_663),
.A2(n_457),
.B(n_458),
.C(n_470),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_635),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_653),
.B(n_583),
.Y(n_792)
);

NOR3xp33_ASAP7_75t_L g793 ( 
.A(n_724),
.B(n_280),
.C(n_269),
.Y(n_793)
);

AOI21xp5_ASAP7_75t_L g794 ( 
.A1(n_620),
.A2(n_472),
.B(n_452),
.Y(n_794)
);

AOI21xp5_ASAP7_75t_L g795 ( 
.A1(n_625),
.A2(n_452),
.B(n_460),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_658),
.B(n_583),
.Y(n_796)
);

A2O1A1Ixp33_ASAP7_75t_L g797 ( 
.A1(n_628),
.A2(n_487),
.B(n_470),
.C(n_451),
.Y(n_797)
);

INVx4_ASAP7_75t_L g798 ( 
.A(n_632),
.Y(n_798)
);

AOI21xp5_ASAP7_75t_L g799 ( 
.A1(n_625),
.A2(n_452),
.B(n_460),
.Y(n_799)
);

BUFx2_ASAP7_75t_SL g800 ( 
.A(n_642),
.Y(n_800)
);

INVx1_ASAP7_75t_SL g801 ( 
.A(n_621),
.Y(n_801)
);

OAI22xp5_ASAP7_75t_L g802 ( 
.A1(n_594),
.A2(n_583),
.B1(n_451),
.B2(n_475),
.Y(n_802)
);

O2A1O1Ixp5_ASAP7_75t_L g803 ( 
.A1(n_732),
.A2(n_554),
.B(n_453),
.C(n_507),
.Y(n_803)
);

OAI22xp5_ASAP7_75t_L g804 ( 
.A1(n_626),
.A2(n_583),
.B1(n_475),
.B2(n_483),
.Y(n_804)
);

AOI22xp5_ASAP7_75t_L g805 ( 
.A1(n_721),
.A2(n_583),
.B1(n_487),
.B2(n_493),
.Y(n_805)
);

HB1xp67_ASAP7_75t_L g806 ( 
.A(n_629),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_658),
.B(n_460),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_596),
.B(n_460),
.Y(n_808)
);

OAI21xp5_ASAP7_75t_L g809 ( 
.A1(n_630),
.A2(n_484),
.B(n_483),
.Y(n_809)
);

BUFx2_ASAP7_75t_L g810 ( 
.A(n_629),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_596),
.B(n_466),
.Y(n_811)
);

O2A1O1Ixp33_ASAP7_75t_L g812 ( 
.A1(n_648),
.A2(n_493),
.B(n_484),
.C(n_539),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_652),
.B(n_466),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_659),
.B(n_466),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_605),
.B(n_466),
.Y(n_815)
);

INVx4_ASAP7_75t_L g816 ( 
.A(n_716),
.Y(n_816)
);

AOI21xp5_ASAP7_75t_L g817 ( 
.A1(n_643),
.A2(n_452),
.B(n_467),
.Y(n_817)
);

AOI21xp5_ASAP7_75t_L g818 ( 
.A1(n_643),
.A2(n_467),
.B(n_468),
.Y(n_818)
);

AOI21xp5_ASAP7_75t_L g819 ( 
.A1(n_664),
.A2(n_467),
.B(n_468),
.Y(n_819)
);

OAI22xp5_ASAP7_75t_L g820 ( 
.A1(n_716),
.A2(n_467),
.B1(n_468),
.B2(n_476),
.Y(n_820)
);

INVx3_ASAP7_75t_L g821 ( 
.A(n_603),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_656),
.B(n_468),
.Y(n_822)
);

AOI21xp33_ASAP7_75t_L g823 ( 
.A1(n_729),
.A2(n_481),
.B(n_551),
.Y(n_823)
);

OAI22xp5_ASAP7_75t_L g824 ( 
.A1(n_600),
.A2(n_502),
.B1(n_476),
.B2(n_478),
.Y(n_824)
);

AOI22xp5_ASAP7_75t_L g825 ( 
.A1(n_597),
.A2(n_507),
.B1(n_455),
.B2(n_453),
.Y(n_825)
);

A2O1A1Ixp33_ASAP7_75t_L g826 ( 
.A1(n_656),
.A2(n_502),
.B(n_478),
.C(n_489),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_639),
.Y(n_827)
);

A2O1A1Ixp33_ASAP7_75t_L g828 ( 
.A1(n_649),
.A2(n_502),
.B(n_478),
.C(n_489),
.Y(n_828)
);

AOI21xp5_ASAP7_75t_L g829 ( 
.A1(n_683),
.A2(n_476),
.B(n_478),
.Y(n_829)
);

CKINVDCx10_ASAP7_75t_R g830 ( 
.A(n_704),
.Y(n_830)
);

AOI21xp5_ASAP7_75t_L g831 ( 
.A1(n_686),
.A2(n_509),
.B(n_476),
.Y(n_831)
);

A2O1A1Ixp33_ASAP7_75t_L g832 ( 
.A1(n_649),
.A2(n_509),
.B(n_489),
.C(n_526),
.Y(n_832)
);

A2O1A1Ixp33_ASAP7_75t_L g833 ( 
.A1(n_615),
.A2(n_507),
.B(n_455),
.C(n_551),
.Y(n_833)
);

NOR2xp33_ASAP7_75t_L g834 ( 
.A(n_672),
.B(n_489),
.Y(n_834)
);

AND2x4_ASAP7_75t_L g835 ( 
.A(n_672),
.B(n_538),
.Y(n_835)
);

OAI21xp5_ASAP7_75t_L g836 ( 
.A1(n_732),
.A2(n_506),
.B(n_481),
.Y(n_836)
);

OR2x6_ASAP7_75t_SL g837 ( 
.A(n_654),
.B(n_285),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_SL g838 ( 
.A(n_667),
.B(n_464),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_641),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_638),
.B(n_490),
.Y(n_840)
);

AOI21xp5_ASAP7_75t_L g841 ( 
.A1(n_691),
.A2(n_490),
.B(n_502),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_651),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_619),
.B(n_490),
.Y(n_843)
);

A2O1A1Ixp33_ASAP7_75t_L g844 ( 
.A1(n_601),
.A2(n_509),
.B(n_526),
.C(n_539),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_627),
.B(n_509),
.Y(n_845)
);

HB1xp67_ASAP7_75t_L g846 ( 
.A(n_660),
.Y(n_846)
);

A2O1A1Ixp33_ASAP7_75t_L g847 ( 
.A1(n_698),
.A2(n_521),
.B(n_492),
.C(n_520),
.Y(n_847)
);

NOR3xp33_ASAP7_75t_L g848 ( 
.A(n_724),
.B(n_294),
.C(n_301),
.Y(n_848)
);

AOI21xp5_ASAP7_75t_L g849 ( 
.A1(n_699),
.A2(n_526),
.B(n_539),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_SL g850 ( 
.A(n_667),
.B(n_464),
.Y(n_850)
);

NAND2x1p5_ASAP7_75t_L g851 ( 
.A(n_734),
.B(n_545),
.Y(n_851)
);

OAI21xp33_ASAP7_75t_L g852 ( 
.A1(n_601),
.A2(n_679),
.B(n_671),
.Y(n_852)
);

BUFx6f_ASAP7_75t_L g853 ( 
.A(n_646),
.Y(n_853)
);

OAI21xp33_ASAP7_75t_L g854 ( 
.A1(n_681),
.A2(n_286),
.B(n_293),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_634),
.B(n_526),
.Y(n_855)
);

AOI21xp33_ASAP7_75t_L g856 ( 
.A1(n_733),
.A2(n_520),
.B(n_492),
.Y(n_856)
);

AOI21xp5_ASAP7_75t_L g857 ( 
.A1(n_701),
.A2(n_539),
.B(n_538),
.Y(n_857)
);

A2O1A1Ixp33_ASAP7_75t_L g858 ( 
.A1(n_668),
.A2(n_525),
.B(n_506),
.C(n_535),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_645),
.Y(n_859)
);

AOI21xp5_ASAP7_75t_L g860 ( 
.A1(n_703),
.A2(n_521),
.B(n_503),
.Y(n_860)
);

A2O1A1Ixp33_ASAP7_75t_L g861 ( 
.A1(n_669),
.A2(n_503),
.B(n_525),
.C(n_535),
.Y(n_861)
);

O2A1O1Ixp33_ASAP7_75t_L g862 ( 
.A1(n_682),
.A2(n_533),
.B(n_291),
.C(n_253),
.Y(n_862)
);

AOI21xp5_ASAP7_75t_L g863 ( 
.A1(n_710),
.A2(n_533),
.B(n_464),
.Y(n_863)
);

AOI21xp5_ASAP7_75t_L g864 ( 
.A1(n_711),
.A2(n_717),
.B(n_712),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_611),
.B(n_464),
.Y(n_865)
);

INVx4_ASAP7_75t_L g866 ( 
.A(n_603),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_670),
.Y(n_867)
);

BUFx6f_ASAP7_75t_L g868 ( 
.A(n_646),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_733),
.B(n_464),
.Y(n_869)
);

AOI21xp5_ASAP7_75t_L g870 ( 
.A1(n_640),
.A2(n_464),
.B(n_505),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_SL g871 ( 
.A(n_666),
.B(n_494),
.Y(n_871)
);

NOR3xp33_ASAP7_75t_L g872 ( 
.A(n_610),
.B(n_665),
.C(n_695),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_647),
.B(n_494),
.Y(n_873)
);

NOR2xp33_ASAP7_75t_L g874 ( 
.A(n_749),
.B(n_622),
.Y(n_874)
);

INVx3_ASAP7_75t_L g875 ( 
.A(n_631),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_623),
.B(n_494),
.Y(n_876)
);

AOI21x1_ASAP7_75t_L g877 ( 
.A1(n_702),
.A2(n_728),
.B(n_714),
.Y(n_877)
);

INVx2_ASAP7_75t_L g878 ( 
.A(n_655),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_673),
.B(n_494),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_674),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_687),
.B(n_494),
.Y(n_881)
);

OAI21xp33_ASAP7_75t_L g882 ( 
.A1(n_636),
.A2(n_305),
.B(n_300),
.Y(n_882)
);

CKINVDCx20_ASAP7_75t_R g883 ( 
.A(n_742),
.Y(n_883)
);

OAI321xp33_ASAP7_75t_L g884 ( 
.A1(n_736),
.A2(n_554),
.A3(n_291),
.B1(n_253),
.B2(n_302),
.C(n_505),
.Y(n_884)
);

NOR2xp33_ASAP7_75t_L g885 ( 
.A(n_657),
.B(n_515),
.Y(n_885)
);

AND2x4_ASAP7_75t_L g886 ( 
.A(n_692),
.B(n_494),
.Y(n_886)
);

HB1xp67_ASAP7_75t_L g887 ( 
.A(n_604),
.Y(n_887)
);

INVx2_ASAP7_75t_L g888 ( 
.A(n_688),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_SL g889 ( 
.A(n_666),
.B(n_505),
.Y(n_889)
);

AOI21xp5_ASAP7_75t_L g890 ( 
.A1(n_715),
.A2(n_505),
.B(n_545),
.Y(n_890)
);

AOI21x1_ASAP7_75t_L g891 ( 
.A1(n_702),
.A2(n_515),
.B(n_545),
.Y(n_891)
);

AND2x2_ASAP7_75t_L g892 ( 
.A(n_737),
.B(n_253),
.Y(n_892)
);

AND2x2_ASAP7_75t_L g893 ( 
.A(n_697),
.B(n_291),
.Y(n_893)
);

HB1xp67_ASAP7_75t_L g894 ( 
.A(n_606),
.Y(n_894)
);

HB1xp67_ASAP7_75t_L g895 ( 
.A(n_607),
.Y(n_895)
);

NOR2xp67_ASAP7_75t_L g896 ( 
.A(n_697),
.B(n_545),
.Y(n_896)
);

INVx4_ASAP7_75t_L g897 ( 
.A(n_631),
.Y(n_897)
);

O2A1O1Ixp33_ASAP7_75t_L g898 ( 
.A1(n_690),
.A2(n_291),
.B(n_13),
.C(n_15),
.Y(n_898)
);

OAI21xp5_ASAP7_75t_L g899 ( 
.A1(n_725),
.A2(n_545),
.B(n_515),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_696),
.B(n_505),
.Y(n_900)
);

AOI21xp5_ASAP7_75t_L g901 ( 
.A1(n_602),
.A2(n_505),
.B(n_545),
.Y(n_901)
);

AND2x2_ASAP7_75t_L g902 ( 
.A(n_753),
.B(n_302),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_694),
.Y(n_903)
);

INVx2_ASAP7_75t_L g904 ( 
.A(n_700),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_705),
.B(n_515),
.Y(n_905)
);

O2A1O1Ixp33_ASAP7_75t_L g906 ( 
.A1(n_706),
.A2(n_11),
.B(n_13),
.C(n_15),
.Y(n_906)
);

NOR2xp33_ASAP7_75t_SL g907 ( 
.A(n_617),
.B(n_160),
.Y(n_907)
);

AND2x2_ASAP7_75t_L g908 ( 
.A(n_753),
.B(n_17),
.Y(n_908)
);

O2A1O1Ixp33_ASAP7_75t_L g909 ( 
.A1(n_707),
.A2(n_17),
.B(n_19),
.C(n_26),
.Y(n_909)
);

INVx4_ASAP7_75t_L g910 ( 
.A(n_637),
.Y(n_910)
);

AOI21xp5_ASAP7_75t_L g911 ( 
.A1(n_746),
.A2(n_193),
.B(n_307),
.Y(n_911)
);

NOR2xp67_ASAP7_75t_L g912 ( 
.A(n_760),
.B(n_163),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_713),
.Y(n_913)
);

INVx2_ASAP7_75t_SL g914 ( 
.A(n_644),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_SL g915 ( 
.A(n_718),
.B(n_308),
.Y(n_915)
);

AOI21xp5_ASAP7_75t_L g916 ( 
.A1(n_747),
.A2(n_189),
.B(n_298),
.Y(n_916)
);

AOI21xp5_ASAP7_75t_L g917 ( 
.A1(n_735),
.A2(n_727),
.B(n_758),
.Y(n_917)
);

AOI21xp5_ASAP7_75t_L g918 ( 
.A1(n_743),
.A2(n_187),
.B(n_296),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_708),
.Y(n_919)
);

INVx2_ASAP7_75t_L g920 ( 
.A(n_738),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_719),
.B(n_169),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_720),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_722),
.B(n_173),
.Y(n_923)
);

AOI21xp5_ASAP7_75t_L g924 ( 
.A1(n_748),
.A2(n_756),
.B(n_750),
.Y(n_924)
);

AOI21xp5_ASAP7_75t_L g925 ( 
.A1(n_738),
.A2(n_194),
.B(n_292),
.Y(n_925)
);

INVx2_ASAP7_75t_L g926 ( 
.A(n_730),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_636),
.B(n_637),
.Y(n_927)
);

BUFx6f_ASAP7_75t_L g928 ( 
.A(n_646),
.Y(n_928)
);

AOI21xp5_ASAP7_75t_L g929 ( 
.A1(n_714),
.A2(n_186),
.B(n_287),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_SL g930 ( 
.A(n_646),
.B(n_174),
.Y(n_930)
);

AOI21xp5_ASAP7_75t_L g931 ( 
.A1(n_728),
.A2(n_180),
.B(n_284),
.Y(n_931)
);

AND2x2_ASAP7_75t_L g932 ( 
.A(n_753),
.B(n_736),
.Y(n_932)
);

O2A1O1Ixp33_ASAP7_75t_L g933 ( 
.A1(n_739),
.A2(n_19),
.B(n_27),
.C(n_28),
.Y(n_933)
);

AOI21xp5_ASAP7_75t_L g934 ( 
.A1(n_731),
.A2(n_201),
.B(n_283),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_650),
.B(n_195),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_650),
.B(n_178),
.Y(n_936)
);

HB1xp67_ASAP7_75t_L g937 ( 
.A(n_723),
.Y(n_937)
);

NAND3xp33_ASAP7_75t_L g938 ( 
.A(n_760),
.B(n_204),
.C(n_277),
.Y(n_938)
);

OAI21xp5_ASAP7_75t_L g939 ( 
.A1(n_726),
.A2(n_177),
.B(n_276),
.Y(n_939)
);

OAI22x1_ASAP7_75t_L g940 ( 
.A1(n_618),
.A2(n_299),
.B1(n_271),
.B2(n_265),
.Y(n_940)
);

OAI22x1_ASAP7_75t_L g941 ( 
.A1(n_741),
.A2(n_264),
.B1(n_263),
.B2(n_262),
.Y(n_941)
);

AO21x1_ASAP7_75t_L g942 ( 
.A1(n_751),
.A2(n_104),
.B(n_135),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_755),
.B(n_257),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_759),
.Y(n_944)
);

AOI21xp5_ASAP7_75t_L g945 ( 
.A1(n_731),
.A2(n_251),
.B(n_245),
.Y(n_945)
);

O2A1O1Ixp33_ASAP7_75t_L g946 ( 
.A1(n_740),
.A2(n_29),
.B(n_30),
.C(n_31),
.Y(n_946)
);

AOI21xp5_ASAP7_75t_L g947 ( 
.A1(n_773),
.A2(n_751),
.B(n_752),
.Y(n_947)
);

AOI22xp5_ASAP7_75t_L g948 ( 
.A1(n_874),
.A2(n_677),
.B1(n_662),
.B2(n_754),
.Y(n_948)
);

A2O1A1Ixp33_ASAP7_75t_L g949 ( 
.A1(n_852),
.A2(n_757),
.B(n_752),
.C(n_745),
.Y(n_949)
);

AOI21xp5_ASAP7_75t_L g950 ( 
.A1(n_873),
.A2(n_767),
.B(n_864),
.Y(n_950)
);

NOR2xp33_ASAP7_75t_L g951 ( 
.A(n_801),
.B(n_757),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_781),
.Y(n_952)
);

BUFx3_ASAP7_75t_L g953 ( 
.A(n_810),
.Y(n_953)
);

BUFx6f_ASAP7_75t_L g954 ( 
.A(n_853),
.Y(n_954)
);

BUFx6f_ASAP7_75t_L g955 ( 
.A(n_853),
.Y(n_955)
);

NOR2xp33_ASAP7_75t_L g956 ( 
.A(n_806),
.B(n_745),
.Y(n_956)
);

INVxp67_ASAP7_75t_L g957 ( 
.A(n_806),
.Y(n_957)
);

A2O1A1Ixp33_ASAP7_75t_L g958 ( 
.A1(n_834),
.A2(n_745),
.B(n_744),
.C(n_693),
.Y(n_958)
);

OAI22xp5_ASAP7_75t_L g959 ( 
.A1(n_784),
.A2(n_677),
.B1(n_744),
.B2(n_693),
.Y(n_959)
);

AOI21xp5_ASAP7_75t_L g960 ( 
.A1(n_808),
.A2(n_745),
.B(n_744),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_SL g961 ( 
.A(n_872),
.B(n_874),
.Y(n_961)
);

BUFx2_ASAP7_75t_R g962 ( 
.A(n_837),
.Y(n_962)
);

AND2x2_ASAP7_75t_L g963 ( 
.A(n_892),
.B(n_677),
.Y(n_963)
);

OAI21xp5_ASAP7_75t_L g964 ( 
.A1(n_847),
.A2(n_239),
.B(n_213),
.Y(n_964)
);

AOI21xp5_ASAP7_75t_L g965 ( 
.A1(n_811),
.A2(n_744),
.B(n_693),
.Y(n_965)
);

INVx2_ASAP7_75t_L g966 ( 
.A(n_761),
.Y(n_966)
);

INVx2_ASAP7_75t_SL g967 ( 
.A(n_765),
.Y(n_967)
);

INVxp33_ASAP7_75t_SL g968 ( 
.A(n_846),
.Y(n_968)
);

NOR2xp33_ASAP7_75t_L g969 ( 
.A(n_893),
.B(n_693),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_SL g970 ( 
.A(n_872),
.B(n_689),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_932),
.B(n_689),
.Y(n_971)
);

INVx4_ASAP7_75t_L g972 ( 
.A(n_779),
.Y(n_972)
);

NOR2xp33_ASAP7_75t_L g973 ( 
.A(n_846),
.B(n_689),
.Y(n_973)
);

HB1xp67_ASAP7_75t_L g974 ( 
.A(n_800),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_944),
.B(n_887),
.Y(n_975)
);

NAND3xp33_ASAP7_75t_SL g976 ( 
.A(n_793),
.B(n_225),
.C(n_223),
.Y(n_976)
);

AOI22xp5_ASAP7_75t_L g977 ( 
.A1(n_793),
.A2(n_848),
.B1(n_883),
.B2(n_789),
.Y(n_977)
);

A2O1A1Ixp33_ASAP7_75t_L g978 ( 
.A1(n_834),
.A2(n_689),
.B(n_678),
.C(n_676),
.Y(n_978)
);

INVx2_ASAP7_75t_L g979 ( 
.A(n_762),
.Y(n_979)
);

NOR2xp33_ASAP7_75t_L g980 ( 
.A(n_914),
.B(n_678),
.Y(n_980)
);

AO21x1_ASAP7_75t_L g981 ( 
.A1(n_927),
.A2(n_678),
.B(n_676),
.Y(n_981)
);

A2O1A1Ixp33_ASAP7_75t_SL g982 ( 
.A1(n_812),
.A2(n_678),
.B(n_676),
.C(n_32),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_SL g983 ( 
.A(n_816),
.B(n_676),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_839),
.B(n_842),
.Y(n_984)
);

OAI22xp5_ASAP7_75t_L g985 ( 
.A1(n_867),
.A2(n_243),
.B1(n_242),
.B2(n_241),
.Y(n_985)
);

AOI21xp5_ASAP7_75t_L g986 ( 
.A1(n_870),
.A2(n_899),
.B(n_775),
.Y(n_986)
);

BUFx12f_ASAP7_75t_L g987 ( 
.A(n_908),
.Y(n_987)
);

HB1xp67_ASAP7_75t_L g988 ( 
.A(n_835),
.Y(n_988)
);

NOR3xp33_ASAP7_75t_SL g989 ( 
.A(n_906),
.B(n_240),
.C(n_233),
.Y(n_989)
);

A2O1A1Ixp33_ASAP7_75t_L g990 ( 
.A1(n_776),
.A2(n_232),
.B(n_230),
.C(n_229),
.Y(n_990)
);

NOR2xp33_ASAP7_75t_L g991 ( 
.A(n_880),
.B(n_221),
.Y(n_991)
);

OAI321xp33_ASAP7_75t_L g992 ( 
.A1(n_882),
.A2(n_909),
.A3(n_946),
.B1(n_933),
.B2(n_898),
.C(n_902),
.Y(n_992)
);

AOI21xp5_ASAP7_75t_L g993 ( 
.A1(n_774),
.A2(n_863),
.B(n_792),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_919),
.B(n_30),
.Y(n_994)
);

A2O1A1Ixp33_ASAP7_75t_L g995 ( 
.A1(n_764),
.A2(n_218),
.B(n_211),
.C(n_35),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_922),
.B(n_31),
.Y(n_996)
);

A2O1A1Ixp33_ASAP7_75t_L g997 ( 
.A1(n_790),
.A2(n_34),
.B(n_36),
.C(n_38),
.Y(n_997)
);

NOR2xp33_ASAP7_75t_L g998 ( 
.A(n_926),
.B(n_38),
.Y(n_998)
);

NAND3xp33_ASAP7_75t_L g999 ( 
.A(n_848),
.B(n_39),
.C(n_40),
.Y(n_999)
);

INVx2_ASAP7_75t_L g1000 ( 
.A(n_770),
.Y(n_1000)
);

NOR2xp33_ASAP7_75t_L g1001 ( 
.A(n_821),
.B(n_39),
.Y(n_1001)
);

NOR2xp33_ASAP7_75t_L g1002 ( 
.A(n_821),
.B(n_41),
.Y(n_1002)
);

AOI22xp5_ASAP7_75t_L g1003 ( 
.A1(n_941),
.A2(n_41),
.B1(n_43),
.B2(n_46),
.Y(n_1003)
);

AOI21xp5_ASAP7_75t_L g1004 ( 
.A1(n_819),
.A2(n_81),
.B(n_113),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_887),
.B(n_894),
.Y(n_1005)
);

INVx1_ASAP7_75t_SL g1006 ( 
.A(n_830),
.Y(n_1006)
);

INVx2_ASAP7_75t_L g1007 ( 
.A(n_782),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_791),
.Y(n_1008)
);

AOI21xp5_ASAP7_75t_L g1009 ( 
.A1(n_822),
.A2(n_79),
.B(n_101),
.Y(n_1009)
);

INVx2_ASAP7_75t_L g1010 ( 
.A(n_827),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_SL g1011 ( 
.A(n_816),
.B(n_50),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_894),
.B(n_51),
.Y(n_1012)
);

AO32x1_ASAP7_75t_L g1013 ( 
.A1(n_802),
.A2(n_52),
.A3(n_58),
.B1(n_61),
.B2(n_93),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_859),
.Y(n_1014)
);

INVx3_ASAP7_75t_SL g1015 ( 
.A(n_886),
.Y(n_1015)
);

INVx2_ASAP7_75t_SL g1016 ( 
.A(n_886),
.Y(n_1016)
);

INVxp67_ASAP7_75t_L g1017 ( 
.A(n_780),
.Y(n_1017)
);

BUFx2_ASAP7_75t_L g1018 ( 
.A(n_853),
.Y(n_1018)
);

OAI22xp5_ASAP7_75t_L g1019 ( 
.A1(n_769),
.A2(n_94),
.B1(n_115),
.B2(n_771),
.Y(n_1019)
);

AOI22x1_ASAP7_75t_L g1020 ( 
.A1(n_866),
.A2(n_910),
.B1(n_897),
.B2(n_818),
.Y(n_1020)
);

NOR2xp33_ASAP7_75t_L g1021 ( 
.A(n_875),
.B(n_786),
.Y(n_1021)
);

INVx2_ASAP7_75t_L g1022 ( 
.A(n_878),
.Y(n_1022)
);

OAI22xp5_ASAP7_75t_L g1023 ( 
.A1(n_807),
.A2(n_788),
.B1(n_796),
.B2(n_814),
.Y(n_1023)
);

INVx3_ASAP7_75t_SL g1024 ( 
.A(n_930),
.Y(n_1024)
);

BUFx6f_ASAP7_75t_L g1025 ( 
.A(n_853),
.Y(n_1025)
);

INVx2_ASAP7_75t_SL g1026 ( 
.A(n_888),
.Y(n_1026)
);

AOI21x1_ASAP7_75t_L g1027 ( 
.A1(n_763),
.A2(n_869),
.B(n_891),
.Y(n_1027)
);

NOR2xp33_ASAP7_75t_R g1028 ( 
.A(n_907),
.B(n_868),
.Y(n_1028)
);

AOI21xp5_ASAP7_75t_L g1029 ( 
.A1(n_857),
.A2(n_841),
.B(n_829),
.Y(n_1029)
);

OAI22x1_ASAP7_75t_L g1030 ( 
.A1(n_930),
.A2(n_913),
.B1(n_903),
.B2(n_904),
.Y(n_1030)
);

AOI22xp5_ASAP7_75t_L g1031 ( 
.A1(n_895),
.A2(n_940),
.B1(n_854),
.B2(n_937),
.Y(n_1031)
);

AOI22xp5_ASAP7_75t_L g1032 ( 
.A1(n_895),
.A2(n_937),
.B1(n_885),
.B2(n_779),
.Y(n_1032)
);

BUFx6f_ASAP7_75t_L g1033 ( 
.A(n_868),
.Y(n_1033)
);

BUFx6f_ASAP7_75t_L g1034 ( 
.A(n_868),
.Y(n_1034)
);

NAND2x1p5_ASAP7_75t_L g1035 ( 
.A(n_785),
.B(n_798),
.Y(n_1035)
);

BUFx12f_ASAP7_75t_L g1036 ( 
.A(n_868),
.Y(n_1036)
);

NOR2xp33_ASAP7_75t_L g1037 ( 
.A(n_875),
.B(n_920),
.Y(n_1037)
);

AOI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_831),
.A2(n_849),
.B(n_879),
.Y(n_1038)
);

NOR2xp33_ASAP7_75t_SL g1039 ( 
.A(n_785),
.B(n_798),
.Y(n_1039)
);

BUFx6f_ASAP7_75t_L g1040 ( 
.A(n_928),
.Y(n_1040)
);

NAND2x1p5_ASAP7_75t_L g1041 ( 
.A(n_928),
.B(n_866),
.Y(n_1041)
);

AOI21xp5_ASAP7_75t_L g1042 ( 
.A1(n_881),
.A2(n_900),
.B(n_860),
.Y(n_1042)
);

AOI22xp33_ASAP7_75t_L g1043 ( 
.A1(n_935),
.A2(n_936),
.B1(n_923),
.B2(n_921),
.Y(n_1043)
);

NOR2xp33_ASAP7_75t_L g1044 ( 
.A(n_815),
.B(n_897),
.Y(n_1044)
);

A2O1A1Ixp33_ASAP7_75t_L g1045 ( 
.A1(n_885),
.A2(n_788),
.B(n_939),
.C(n_917),
.Y(n_1045)
);

OR2x6_ASAP7_75t_L g1046 ( 
.A(n_851),
.B(n_896),
.Y(n_1046)
);

AND2x2_ASAP7_75t_L g1047 ( 
.A(n_943),
.B(n_912),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_876),
.Y(n_1048)
);

INVx2_ASAP7_75t_L g1049 ( 
.A(n_877),
.Y(n_1049)
);

NOR2xp33_ASAP7_75t_L g1050 ( 
.A(n_910),
.B(n_928),
.Y(n_1050)
);

HB1xp67_ASAP7_75t_L g1051 ( 
.A(n_928),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_924),
.Y(n_1052)
);

A2O1A1Ixp33_ASAP7_75t_SL g1053 ( 
.A1(n_836),
.A2(n_809),
.B(n_778),
.C(n_916),
.Y(n_1053)
);

INVx2_ASAP7_75t_L g1054 ( 
.A(n_905),
.Y(n_1054)
);

OAI22xp5_ASAP7_75t_L g1055 ( 
.A1(n_813),
.A2(n_840),
.B1(n_805),
.B2(n_787),
.Y(n_1055)
);

AOI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_794),
.A2(n_889),
.B(n_871),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_SL g1057 ( 
.A(n_851),
.B(n_884),
.Y(n_1057)
);

OAI22xp5_ASAP7_75t_L g1058 ( 
.A1(n_847),
.A2(n_797),
.B1(n_772),
.B2(n_833),
.Y(n_1058)
);

BUFx3_ASAP7_75t_L g1059 ( 
.A(n_766),
.Y(n_1059)
);

OAI22xp5_ASAP7_75t_L g1060 ( 
.A1(n_833),
.A2(n_855),
.B1(n_845),
.B2(n_843),
.Y(n_1060)
);

A2O1A1Ixp33_ASAP7_75t_SL g1061 ( 
.A1(n_911),
.A2(n_795),
.B(n_817),
.C(n_799),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_SL g1062 ( 
.A(n_865),
.B(n_938),
.Y(n_1062)
);

BUFx3_ASAP7_75t_L g1063 ( 
.A(n_766),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_858),
.Y(n_1064)
);

A2O1A1Ixp33_ASAP7_75t_L g1065 ( 
.A1(n_862),
.A2(n_826),
.B(n_832),
.C(n_828),
.Y(n_1065)
);

AND2x2_ASAP7_75t_L g1066 ( 
.A(n_934),
.B(n_945),
.Y(n_1066)
);

OAI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_803),
.A2(n_858),
.B(n_861),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_871),
.B(n_889),
.Y(n_1068)
);

O2A1O1Ixp33_ASAP7_75t_L g1069 ( 
.A1(n_844),
.A2(n_861),
.B(n_824),
.C(n_918),
.Y(n_1069)
);

BUFx3_ASAP7_75t_L g1070 ( 
.A(n_942),
.Y(n_1070)
);

A2O1A1Ixp33_ASAP7_75t_L g1071 ( 
.A1(n_856),
.A2(n_838),
.B(n_850),
.C(n_915),
.Y(n_1071)
);

O2A1O1Ixp33_ASAP7_75t_L g1072 ( 
.A1(n_820),
.A2(n_915),
.B(n_804),
.C(n_783),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_825),
.B(n_850),
.Y(n_1073)
);

NOR2xp33_ASAP7_75t_L g1074 ( 
.A(n_925),
.B(n_838),
.Y(n_1074)
);

OAI21x1_ASAP7_75t_L g1075 ( 
.A1(n_768),
.A2(n_803),
.B(n_890),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_929),
.Y(n_1076)
);

AND2x2_ASAP7_75t_L g1077 ( 
.A(n_931),
.B(n_823),
.Y(n_1077)
);

O2A1O1Ixp33_ASAP7_75t_L g1078 ( 
.A1(n_777),
.A2(n_508),
.B(n_724),
.C(n_570),
.Y(n_1078)
);

CKINVDCx16_ASAP7_75t_R g1079 ( 
.A(n_777),
.Y(n_1079)
);

OAI21xp5_ASAP7_75t_L g1080 ( 
.A1(n_901),
.A2(n_847),
.B(n_773),
.Y(n_1080)
);

OAI22xp5_ASAP7_75t_L g1081 ( 
.A1(n_783),
.A2(n_594),
.B1(n_652),
.B2(n_648),
.Y(n_1081)
);

NOR2xp33_ASAP7_75t_L g1082 ( 
.A(n_801),
.B(n_313),
.Y(n_1082)
);

BUFx3_ASAP7_75t_L g1083 ( 
.A(n_810),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_781),
.Y(n_1084)
);

CKINVDCx5p33_ASAP7_75t_R g1085 ( 
.A(n_765),
.Y(n_1085)
);

A2O1A1Ixp33_ASAP7_75t_L g1086 ( 
.A1(n_852),
.A2(n_598),
.B(n_508),
.C(n_628),
.Y(n_1086)
);

NOR2xp33_ASAP7_75t_L g1087 ( 
.A(n_801),
.B(n_313),
.Y(n_1087)
);

BUFx6f_ASAP7_75t_L g1088 ( 
.A(n_853),
.Y(n_1088)
);

AOI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_773),
.A2(n_873),
.B(n_767),
.Y(n_1089)
);

NAND3xp33_ASAP7_75t_SL g1090 ( 
.A(n_793),
.B(n_434),
.C(n_532),
.Y(n_1090)
);

BUFx2_ASAP7_75t_L g1091 ( 
.A(n_953),
.Y(n_1091)
);

AO31x2_ASAP7_75t_L g1092 ( 
.A1(n_981),
.A2(n_959),
.A3(n_1030),
.B(n_1058),
.Y(n_1092)
);

A2O1A1Ixp33_ASAP7_75t_L g1093 ( 
.A1(n_1078),
.A2(n_1086),
.B(n_995),
.C(n_977),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_975),
.B(n_957),
.Y(n_1094)
);

AO31x2_ASAP7_75t_L g1095 ( 
.A1(n_959),
.A2(n_1058),
.A3(n_1060),
.B(n_1049),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_975),
.B(n_1005),
.Y(n_1096)
);

O2A1O1Ixp33_ASAP7_75t_L g1097 ( 
.A1(n_1090),
.A2(n_992),
.B(n_997),
.C(n_961),
.Y(n_1097)
);

AND2x2_ASAP7_75t_L g1098 ( 
.A(n_1083),
.B(n_967),
.Y(n_1098)
);

OAI22xp33_ASAP7_75t_L g1099 ( 
.A1(n_1003),
.A2(n_992),
.B1(n_999),
.B2(n_1024),
.Y(n_1099)
);

AOI21xp5_ASAP7_75t_L g1100 ( 
.A1(n_1089),
.A2(n_950),
.B(n_986),
.Y(n_1100)
);

A2O1A1Ixp33_ASAP7_75t_L g1101 ( 
.A1(n_1070),
.A2(n_998),
.B(n_1045),
.C(n_1047),
.Y(n_1101)
);

AOI21xp5_ASAP7_75t_SL g1102 ( 
.A1(n_1081),
.A2(n_1055),
.B(n_958),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_952),
.Y(n_1103)
);

BUFx6f_ASAP7_75t_L g1104 ( 
.A(n_1036),
.Y(n_1104)
);

A2O1A1Ixp33_ASAP7_75t_L g1105 ( 
.A1(n_1043),
.A2(n_964),
.B(n_969),
.C(n_989),
.Y(n_1105)
);

BUFx6f_ASAP7_75t_L g1106 ( 
.A(n_1015),
.Y(n_1106)
);

OR2x2_ASAP7_75t_L g1107 ( 
.A(n_1005),
.B(n_984),
.Y(n_1107)
);

AND2x2_ASAP7_75t_L g1108 ( 
.A(n_1085),
.B(n_1082),
.Y(n_1108)
);

AND2x2_ASAP7_75t_L g1109 ( 
.A(n_1087),
.B(n_988),
.Y(n_1109)
);

OAI22xp5_ASAP7_75t_L g1110 ( 
.A1(n_1081),
.A2(n_994),
.B1(n_996),
.B2(n_1084),
.Y(n_1110)
);

OA21x2_ASAP7_75t_L g1111 ( 
.A1(n_1075),
.A2(n_1080),
.B(n_1067),
.Y(n_1111)
);

CKINVDCx11_ASAP7_75t_R g1112 ( 
.A(n_1006),
.Y(n_1112)
);

AOI22xp5_ASAP7_75t_L g1113 ( 
.A1(n_1079),
.A2(n_951),
.B1(n_963),
.B2(n_968),
.Y(n_1113)
);

AO31x2_ASAP7_75t_L g1114 ( 
.A1(n_1060),
.A2(n_1071),
.A3(n_1023),
.B(n_1065),
.Y(n_1114)
);

O2A1O1Ixp33_ASAP7_75t_L g1115 ( 
.A1(n_1053),
.A2(n_976),
.B(n_985),
.C(n_1023),
.Y(n_1115)
);

AO31x2_ASAP7_75t_L g1116 ( 
.A1(n_949),
.A2(n_993),
.A3(n_1064),
.B(n_1029),
.Y(n_1116)
);

AOI221xp5_ASAP7_75t_L g1117 ( 
.A1(n_985),
.A2(n_964),
.B1(n_991),
.B2(n_990),
.C(n_1012),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_1017),
.B(n_956),
.Y(n_1118)
);

CKINVDCx5p33_ASAP7_75t_R g1119 ( 
.A(n_1006),
.Y(n_1119)
);

A2O1A1Ixp33_ASAP7_75t_L g1120 ( 
.A1(n_1021),
.A2(n_1072),
.B(n_1031),
.C(n_948),
.Y(n_1120)
);

INVxp67_ASAP7_75t_SL g1121 ( 
.A(n_971),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_973),
.B(n_974),
.Y(n_1122)
);

AOI21xp33_ASAP7_75t_L g1123 ( 
.A1(n_970),
.A2(n_1076),
.B(n_1062),
.Y(n_1123)
);

AOI22xp5_ASAP7_75t_L g1124 ( 
.A1(n_1032),
.A2(n_1002),
.B1(n_1001),
.B2(n_1011),
.Y(n_1124)
);

OAI21x1_ASAP7_75t_L g1125 ( 
.A1(n_1038),
.A2(n_1027),
.B(n_1042),
.Y(n_1125)
);

BUFx6f_ASAP7_75t_L g1126 ( 
.A(n_954),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_1026),
.B(n_1008),
.Y(n_1127)
);

AOI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_1080),
.A2(n_947),
.B(n_1061),
.Y(n_1128)
);

AO21x2_ASAP7_75t_L g1129 ( 
.A1(n_1067),
.A2(n_1057),
.B(n_1077),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_1014),
.B(n_979),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_1000),
.B(n_1010),
.Y(n_1131)
);

OAI21xp5_ASAP7_75t_L g1132 ( 
.A1(n_1069),
.A2(n_1055),
.B(n_1056),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_1007),
.Y(n_1133)
);

AO32x2_ASAP7_75t_L g1134 ( 
.A1(n_1019),
.A2(n_1016),
.A3(n_1013),
.B1(n_982),
.B2(n_972),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_1022),
.B(n_1048),
.Y(n_1135)
);

INVx2_ASAP7_75t_L g1136 ( 
.A(n_1054),
.Y(n_1136)
);

OAI21x1_ASAP7_75t_L g1137 ( 
.A1(n_1052),
.A2(n_965),
.B(n_960),
.Y(n_1137)
);

A2O1A1Ixp33_ASAP7_75t_L g1138 ( 
.A1(n_1074),
.A2(n_1037),
.B(n_1019),
.C(n_1073),
.Y(n_1138)
);

A2O1A1Ixp33_ASAP7_75t_L g1139 ( 
.A1(n_1044),
.A2(n_980),
.B(n_978),
.C(n_1009),
.Y(n_1139)
);

O2A1O1Ixp33_ASAP7_75t_SL g1140 ( 
.A1(n_1068),
.A2(n_983),
.B(n_1050),
.C(n_1051),
.Y(n_1140)
);

CKINVDCx6p67_ASAP7_75t_R g1141 ( 
.A(n_987),
.Y(n_1141)
);

A2O1A1Ixp33_ASAP7_75t_L g1142 ( 
.A1(n_1066),
.A2(n_1004),
.B(n_1059),
.C(n_1063),
.Y(n_1142)
);

AOI21xp5_ASAP7_75t_L g1143 ( 
.A1(n_1013),
.A2(n_1020),
.B(n_1039),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_1028),
.B(n_1018),
.Y(n_1144)
);

INVxp67_ASAP7_75t_L g1145 ( 
.A(n_962),
.Y(n_1145)
);

INVx1_ASAP7_75t_SL g1146 ( 
.A(n_954),
.Y(n_1146)
);

OAI22xp5_ASAP7_75t_L g1147 ( 
.A1(n_972),
.A2(n_1041),
.B1(n_1035),
.B2(n_1046),
.Y(n_1147)
);

AND2x4_ASAP7_75t_L g1148 ( 
.A(n_1046),
.B(n_954),
.Y(n_1148)
);

OAI21x1_ASAP7_75t_L g1149 ( 
.A1(n_1041),
.A2(n_1035),
.B(n_1013),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_955),
.B(n_1025),
.Y(n_1150)
);

INVx3_ASAP7_75t_L g1151 ( 
.A(n_955),
.Y(n_1151)
);

AND2x2_ASAP7_75t_L g1152 ( 
.A(n_1025),
.B(n_1033),
.Y(n_1152)
);

OAI21x1_ASAP7_75t_L g1153 ( 
.A1(n_1025),
.A2(n_1033),
.B(n_1034),
.Y(n_1153)
);

AOI21xp5_ASAP7_75t_L g1154 ( 
.A1(n_1040),
.A2(n_773),
.B(n_1086),
.Y(n_1154)
);

O2A1O1Ixp33_ASAP7_75t_L g1155 ( 
.A1(n_1040),
.A2(n_1086),
.B(n_508),
.C(n_1078),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_1088),
.Y(n_1156)
);

NOR2xp67_ASAP7_75t_L g1157 ( 
.A(n_1088),
.B(n_914),
.Y(n_1157)
);

AOI21xp5_ASAP7_75t_L g1158 ( 
.A1(n_1086),
.A2(n_773),
.B(n_1089),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_975),
.B(n_387),
.Y(n_1159)
);

AOI21xp5_ASAP7_75t_L g1160 ( 
.A1(n_1086),
.A2(n_773),
.B(n_1089),
.Y(n_1160)
);

AOI21x1_ASAP7_75t_L g1161 ( 
.A1(n_986),
.A2(n_1089),
.B(n_993),
.Y(n_1161)
);

AO21x2_ASAP7_75t_L g1162 ( 
.A1(n_981),
.A2(n_1067),
.B(n_1080),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_952),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_SL g1164 ( 
.A(n_1078),
.B(n_977),
.Y(n_1164)
);

NOR2xp33_ASAP7_75t_L g1165 ( 
.A(n_968),
.B(n_724),
.Y(n_1165)
);

A2O1A1Ixp33_ASAP7_75t_L g1166 ( 
.A1(n_1078),
.A2(n_1086),
.B(n_508),
.C(n_450),
.Y(n_1166)
);

AND2x4_ASAP7_75t_L g1167 ( 
.A(n_988),
.B(n_953),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_975),
.B(n_387),
.Y(n_1168)
);

AOI22xp33_ASAP7_75t_L g1169 ( 
.A1(n_977),
.A2(n_742),
.B1(n_482),
.B2(n_665),
.Y(n_1169)
);

AND2x2_ASAP7_75t_L g1170 ( 
.A(n_957),
.B(n_665),
.Y(n_1170)
);

OAI21x1_ASAP7_75t_L g1171 ( 
.A1(n_1075),
.A2(n_986),
.B(n_993),
.Y(n_1171)
);

O2A1O1Ixp33_ASAP7_75t_L g1172 ( 
.A1(n_1086),
.A2(n_508),
.B(n_1078),
.C(n_1090),
.Y(n_1172)
);

O2A1O1Ixp33_ASAP7_75t_SL g1173 ( 
.A1(n_1086),
.A2(n_1053),
.B(n_982),
.C(n_1078),
.Y(n_1173)
);

A2O1A1Ixp33_ASAP7_75t_L g1174 ( 
.A1(n_1078),
.A2(n_1086),
.B(n_508),
.C(n_450),
.Y(n_1174)
);

NAND2x1_ASAP7_75t_L g1175 ( 
.A(n_1046),
.B(n_866),
.Y(n_1175)
);

AOI21xp5_ASAP7_75t_SL g1176 ( 
.A1(n_1086),
.A2(n_549),
.B(n_528),
.Y(n_1176)
);

CKINVDCx6p67_ASAP7_75t_R g1177 ( 
.A(n_1006),
.Y(n_1177)
);

BUFx6f_ASAP7_75t_L g1178 ( 
.A(n_1036),
.Y(n_1178)
);

AO31x2_ASAP7_75t_L g1179 ( 
.A1(n_981),
.A2(n_959),
.A3(n_1030),
.B(n_1058),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_952),
.Y(n_1180)
);

OAI21x1_ASAP7_75t_L g1181 ( 
.A1(n_1075),
.A2(n_986),
.B(n_993),
.Y(n_1181)
);

AOI21xp5_ASAP7_75t_L g1182 ( 
.A1(n_1086),
.A2(n_773),
.B(n_1089),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_952),
.Y(n_1183)
);

AOI21xp5_ASAP7_75t_L g1184 ( 
.A1(n_1086),
.A2(n_773),
.B(n_1089),
.Y(n_1184)
);

AOI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_1086),
.A2(n_773),
.B(n_1089),
.Y(n_1185)
);

CKINVDCx5p33_ASAP7_75t_R g1186 ( 
.A(n_1085),
.Y(n_1186)
);

BUFx2_ASAP7_75t_SL g1187 ( 
.A(n_967),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_975),
.B(n_387),
.Y(n_1188)
);

CKINVDCx5p33_ASAP7_75t_R g1189 ( 
.A(n_1085),
.Y(n_1189)
);

AND2x2_ASAP7_75t_L g1190 ( 
.A(n_957),
.B(n_665),
.Y(n_1190)
);

INVx2_ASAP7_75t_L g1191 ( 
.A(n_966),
.Y(n_1191)
);

OAI21xp5_ASAP7_75t_L g1192 ( 
.A1(n_1086),
.A2(n_1081),
.B(n_1045),
.Y(n_1192)
);

AOI22xp33_ASAP7_75t_L g1193 ( 
.A1(n_977),
.A2(n_742),
.B1(n_482),
.B2(n_665),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_975),
.B(n_387),
.Y(n_1194)
);

OA21x2_ASAP7_75t_L g1195 ( 
.A1(n_986),
.A2(n_1075),
.B(n_1080),
.Y(n_1195)
);

OAI21xp5_ASAP7_75t_L g1196 ( 
.A1(n_1086),
.A2(n_1081),
.B(n_1045),
.Y(n_1196)
);

NOR2xp33_ASAP7_75t_L g1197 ( 
.A(n_968),
.B(n_724),
.Y(n_1197)
);

NOR2xp33_ASAP7_75t_R g1198 ( 
.A(n_1085),
.B(n_765),
.Y(n_1198)
);

INVx2_ASAP7_75t_SL g1199 ( 
.A(n_953),
.Y(n_1199)
);

OAI21xp5_ASAP7_75t_SL g1200 ( 
.A1(n_977),
.A2(n_1003),
.B(n_1090),
.Y(n_1200)
);

NAND3xp33_ASAP7_75t_SL g1201 ( 
.A(n_977),
.B(n_434),
.C(n_317),
.Y(n_1201)
);

HB1xp67_ASAP7_75t_L g1202 ( 
.A(n_953),
.Y(n_1202)
);

OAI22xp5_ASAP7_75t_L g1203 ( 
.A1(n_1086),
.A2(n_508),
.B1(n_977),
.B2(n_598),
.Y(n_1203)
);

CKINVDCx20_ASAP7_75t_R g1204 ( 
.A(n_1085),
.Y(n_1204)
);

AO31x2_ASAP7_75t_L g1205 ( 
.A1(n_981),
.A2(n_959),
.A3(n_1030),
.B(n_1058),
.Y(n_1205)
);

NOR2xp33_ASAP7_75t_L g1206 ( 
.A(n_968),
.B(n_724),
.Y(n_1206)
);

O2A1O1Ixp33_ASAP7_75t_L g1207 ( 
.A1(n_1086),
.A2(n_508),
.B(n_1078),
.C(n_1090),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_952),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_952),
.Y(n_1209)
);

AOI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_1086),
.A2(n_773),
.B(n_1089),
.Y(n_1210)
);

AOI21xp5_ASAP7_75t_L g1211 ( 
.A1(n_1086),
.A2(n_773),
.B(n_1089),
.Y(n_1211)
);

CKINVDCx8_ASAP7_75t_R g1212 ( 
.A(n_1085),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_SL g1213 ( 
.A(n_1078),
.B(n_977),
.Y(n_1213)
);

BUFx10_ASAP7_75t_L g1214 ( 
.A(n_1085),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_952),
.Y(n_1215)
);

OAI21x1_ASAP7_75t_L g1216 ( 
.A1(n_1075),
.A2(n_986),
.B(n_993),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_952),
.Y(n_1217)
);

AOI21xp5_ASAP7_75t_L g1218 ( 
.A1(n_1086),
.A2(n_773),
.B(n_1089),
.Y(n_1218)
);

AO31x2_ASAP7_75t_L g1219 ( 
.A1(n_981),
.A2(n_959),
.A3(n_1030),
.B(n_1058),
.Y(n_1219)
);

OAI21xp5_ASAP7_75t_L g1220 ( 
.A1(n_1086),
.A2(n_1081),
.B(n_1045),
.Y(n_1220)
);

AO31x2_ASAP7_75t_L g1221 ( 
.A1(n_981),
.A2(n_959),
.A3(n_1030),
.B(n_1058),
.Y(n_1221)
);

OAI21x1_ASAP7_75t_L g1222 ( 
.A1(n_1075),
.A2(n_986),
.B(n_993),
.Y(n_1222)
);

AND2x2_ASAP7_75t_L g1223 ( 
.A(n_957),
.B(n_665),
.Y(n_1223)
);

AO31x2_ASAP7_75t_L g1224 ( 
.A1(n_981),
.A2(n_959),
.A3(n_1030),
.B(n_1058),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_952),
.Y(n_1225)
);

AOI22xp33_ASAP7_75t_L g1226 ( 
.A1(n_1169),
.A2(n_1193),
.B1(n_1117),
.B2(n_1201),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_1103),
.Y(n_1227)
);

OAI22xp5_ASAP7_75t_L g1228 ( 
.A1(n_1124),
.A2(n_1203),
.B1(n_1200),
.B2(n_1174),
.Y(n_1228)
);

NAND2x1p5_ASAP7_75t_L g1229 ( 
.A(n_1148),
.B(n_1175),
.Y(n_1229)
);

AOI22xp5_ASAP7_75t_L g1230 ( 
.A1(n_1200),
.A2(n_1099),
.B1(n_1124),
.B2(n_1164),
.Y(n_1230)
);

OAI22xp5_ASAP7_75t_L g1231 ( 
.A1(n_1166),
.A2(n_1093),
.B1(n_1213),
.B2(n_1097),
.Y(n_1231)
);

CKINVDCx11_ASAP7_75t_R g1232 ( 
.A(n_1212),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_L g1233 ( 
.A(n_1096),
.B(n_1159),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_1168),
.B(n_1188),
.Y(n_1234)
);

NAND2x1p5_ASAP7_75t_L g1235 ( 
.A(n_1148),
.B(n_1152),
.Y(n_1235)
);

NAND2xp33_ASAP7_75t_SL g1236 ( 
.A(n_1104),
.B(n_1178),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_L g1237 ( 
.A(n_1194),
.B(n_1107),
.Y(n_1237)
);

INVx6_ASAP7_75t_L g1238 ( 
.A(n_1106),
.Y(n_1238)
);

OAI22xp5_ASAP7_75t_L g1239 ( 
.A1(n_1192),
.A2(n_1196),
.B1(n_1220),
.B2(n_1110),
.Y(n_1239)
);

INVx6_ASAP7_75t_L g1240 ( 
.A(n_1106),
.Y(n_1240)
);

OAI22xp33_ASAP7_75t_L g1241 ( 
.A1(n_1192),
.A2(n_1220),
.B1(n_1196),
.B2(n_1113),
.Y(n_1241)
);

INVx3_ASAP7_75t_L g1242 ( 
.A(n_1126),
.Y(n_1242)
);

OAI22xp33_ASAP7_75t_L g1243 ( 
.A1(n_1113),
.A2(n_1110),
.B1(n_1094),
.B2(n_1118),
.Y(n_1243)
);

BUFx10_ASAP7_75t_L g1244 ( 
.A(n_1186),
.Y(n_1244)
);

INVx6_ASAP7_75t_L g1245 ( 
.A(n_1106),
.Y(n_1245)
);

INVx8_ASAP7_75t_L g1246 ( 
.A(n_1204),
.Y(n_1246)
);

OAI22xp33_ASAP7_75t_L g1247 ( 
.A1(n_1122),
.A2(n_1132),
.B1(n_1225),
.B2(n_1217),
.Y(n_1247)
);

BUFx4f_ASAP7_75t_SL g1248 ( 
.A(n_1177),
.Y(n_1248)
);

AOI22xp33_ASAP7_75t_SL g1249 ( 
.A1(n_1145),
.A2(n_1132),
.B1(n_1223),
.B2(n_1170),
.Y(n_1249)
);

AOI22xp33_ASAP7_75t_L g1250 ( 
.A1(n_1190),
.A2(n_1136),
.B1(n_1109),
.B2(n_1129),
.Y(n_1250)
);

INVx1_ASAP7_75t_SL g1251 ( 
.A(n_1091),
.Y(n_1251)
);

INVx4_ASAP7_75t_L g1252 ( 
.A(n_1104),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1163),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_L g1254 ( 
.A(n_1167),
.B(n_1202),
.Y(n_1254)
);

BUFx12f_ASAP7_75t_L g1255 ( 
.A(n_1112),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_L g1256 ( 
.A(n_1180),
.B(n_1183),
.Y(n_1256)
);

BUFx2_ASAP7_75t_SL g1257 ( 
.A(n_1108),
.Y(n_1257)
);

OAI21xp5_ASAP7_75t_SL g1258 ( 
.A1(n_1172),
.A2(n_1207),
.B(n_1115),
.Y(n_1258)
);

AOI22xp33_ASAP7_75t_L g1259 ( 
.A1(n_1129),
.A2(n_1121),
.B1(n_1208),
.B2(n_1215),
.Y(n_1259)
);

INVx4_ASAP7_75t_L g1260 ( 
.A(n_1104),
.Y(n_1260)
);

AOI22xp33_ASAP7_75t_SL g1261 ( 
.A1(n_1162),
.A2(n_1209),
.B1(n_1120),
.B2(n_1135),
.Y(n_1261)
);

CKINVDCx20_ASAP7_75t_R g1262 ( 
.A(n_1198),
.Y(n_1262)
);

INVx8_ASAP7_75t_L g1263 ( 
.A(n_1178),
.Y(n_1263)
);

CKINVDCx5p33_ASAP7_75t_R g1264 ( 
.A(n_1189),
.Y(n_1264)
);

AOI22xp33_ASAP7_75t_L g1265 ( 
.A1(n_1133),
.A2(n_1191),
.B1(n_1162),
.B2(n_1130),
.Y(n_1265)
);

AOI22xp33_ASAP7_75t_L g1266 ( 
.A1(n_1131),
.A2(n_1123),
.B1(n_1127),
.B2(n_1141),
.Y(n_1266)
);

BUFx6f_ASAP7_75t_L g1267 ( 
.A(n_1126),
.Y(n_1267)
);

BUFx12f_ASAP7_75t_L g1268 ( 
.A(n_1214),
.Y(n_1268)
);

CKINVDCx6p67_ASAP7_75t_R g1269 ( 
.A(n_1214),
.Y(n_1269)
);

CKINVDCx11_ASAP7_75t_R g1270 ( 
.A(n_1178),
.Y(n_1270)
);

CKINVDCx5p33_ASAP7_75t_R g1271 ( 
.A(n_1119),
.Y(n_1271)
);

OAI21xp5_ASAP7_75t_L g1272 ( 
.A1(n_1138),
.A2(n_1155),
.B(n_1105),
.Y(n_1272)
);

HB1xp67_ASAP7_75t_L g1273 ( 
.A(n_1095),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_1199),
.B(n_1165),
.Y(n_1274)
);

AOI22xp33_ASAP7_75t_SL g1275 ( 
.A1(n_1102),
.A2(n_1101),
.B1(n_1114),
.B2(n_1197),
.Y(n_1275)
);

CKINVDCx11_ASAP7_75t_R g1276 ( 
.A(n_1146),
.Y(n_1276)
);

CKINVDCx11_ASAP7_75t_R g1277 ( 
.A(n_1146),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1156),
.Y(n_1278)
);

BUFx2_ASAP7_75t_L g1279 ( 
.A(n_1144),
.Y(n_1279)
);

CKINVDCx11_ASAP7_75t_R g1280 ( 
.A(n_1187),
.Y(n_1280)
);

CKINVDCx11_ASAP7_75t_R g1281 ( 
.A(n_1147),
.Y(n_1281)
);

AOI22xp33_ASAP7_75t_SL g1282 ( 
.A1(n_1114),
.A2(n_1206),
.B1(n_1143),
.B2(n_1111),
.Y(n_1282)
);

CKINVDCx5p33_ASAP7_75t_R g1283 ( 
.A(n_1098),
.Y(n_1283)
);

INVxp67_ASAP7_75t_SL g1284 ( 
.A(n_1111),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_L g1285 ( 
.A(n_1157),
.B(n_1114),
.Y(n_1285)
);

CKINVDCx6p67_ASAP7_75t_R g1286 ( 
.A(n_1150),
.Y(n_1286)
);

BUFx12f_ASAP7_75t_L g1287 ( 
.A(n_1157),
.Y(n_1287)
);

AND2x2_ASAP7_75t_L g1288 ( 
.A(n_1151),
.B(n_1153),
.Y(n_1288)
);

CKINVDCx20_ASAP7_75t_R g1289 ( 
.A(n_1151),
.Y(n_1289)
);

OAI22xp5_ASAP7_75t_L g1290 ( 
.A1(n_1139),
.A2(n_1154),
.B1(n_1185),
.B2(n_1160),
.Y(n_1290)
);

CKINVDCx6p67_ASAP7_75t_R g1291 ( 
.A(n_1140),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1095),
.Y(n_1292)
);

AOI22xp33_ASAP7_75t_SL g1293 ( 
.A1(n_1158),
.A2(n_1218),
.B1(n_1182),
.B2(n_1211),
.Y(n_1293)
);

OAI22xp5_ASAP7_75t_L g1294 ( 
.A1(n_1184),
.A2(n_1210),
.B1(n_1128),
.B2(n_1176),
.Y(n_1294)
);

CKINVDCx20_ASAP7_75t_R g1295 ( 
.A(n_1195),
.Y(n_1295)
);

BUFx6f_ASAP7_75t_L g1296 ( 
.A(n_1149),
.Y(n_1296)
);

BUFx12f_ASAP7_75t_L g1297 ( 
.A(n_1142),
.Y(n_1297)
);

AOI22xp33_ASAP7_75t_L g1298 ( 
.A1(n_1137),
.A2(n_1134),
.B1(n_1100),
.B2(n_1125),
.Y(n_1298)
);

AOI22xp33_ASAP7_75t_L g1299 ( 
.A1(n_1134),
.A2(n_1092),
.B1(n_1224),
.B2(n_1221),
.Y(n_1299)
);

AND2x2_ASAP7_75t_L g1300 ( 
.A(n_1092),
.B(n_1224),
.Y(n_1300)
);

BUFx10_ASAP7_75t_L g1301 ( 
.A(n_1173),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1092),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1179),
.Y(n_1303)
);

CKINVDCx11_ASAP7_75t_R g1304 ( 
.A(n_1134),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1179),
.Y(n_1305)
);

OAI22xp33_ASAP7_75t_L g1306 ( 
.A1(n_1179),
.A2(n_1224),
.B1(n_1221),
.B2(n_1219),
.Y(n_1306)
);

INVx1_ASAP7_75t_SL g1307 ( 
.A(n_1171),
.Y(n_1307)
);

CKINVDCx11_ASAP7_75t_R g1308 ( 
.A(n_1116),
.Y(n_1308)
);

CKINVDCx11_ASAP7_75t_R g1309 ( 
.A(n_1116),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1205),
.Y(n_1310)
);

AOI22xp33_ASAP7_75t_L g1311 ( 
.A1(n_1205),
.A2(n_1219),
.B1(n_1221),
.B2(n_1222),
.Y(n_1311)
);

AOI22xp33_ASAP7_75t_L g1312 ( 
.A1(n_1205),
.A2(n_1219),
.B1(n_1181),
.B2(n_1216),
.Y(n_1312)
);

OAI22xp5_ASAP7_75t_L g1313 ( 
.A1(n_1161),
.A2(n_1124),
.B1(n_977),
.B2(n_1203),
.Y(n_1313)
);

AOI22xp33_ASAP7_75t_SL g1314 ( 
.A1(n_1203),
.A2(n_908),
.B1(n_902),
.B2(n_932),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1103),
.Y(n_1315)
);

INVx6_ASAP7_75t_L g1316 ( 
.A(n_1106),
.Y(n_1316)
);

OAI22xp5_ASAP7_75t_L g1317 ( 
.A1(n_1124),
.A2(n_977),
.B1(n_1203),
.B2(n_1086),
.Y(n_1317)
);

INVx1_ASAP7_75t_SL g1318 ( 
.A(n_1091),
.Y(n_1318)
);

CKINVDCx16_ASAP7_75t_R g1319 ( 
.A(n_1198),
.Y(n_1319)
);

CKINVDCx20_ASAP7_75t_R g1320 ( 
.A(n_1204),
.Y(n_1320)
);

OAI22xp33_ASAP7_75t_L g1321 ( 
.A1(n_1200),
.A2(n_1124),
.B1(n_977),
.B2(n_1203),
.Y(n_1321)
);

BUFx3_ASAP7_75t_L g1322 ( 
.A(n_1091),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1103),
.Y(n_1323)
);

OAI22xp5_ASAP7_75t_L g1324 ( 
.A1(n_1124),
.A2(n_977),
.B1(n_1203),
.B2(n_1086),
.Y(n_1324)
);

OAI21xp5_ASAP7_75t_L g1325 ( 
.A1(n_1166),
.A2(n_1174),
.B(n_1203),
.Y(n_1325)
);

AOI21xp33_ASAP7_75t_L g1326 ( 
.A1(n_1203),
.A2(n_1117),
.B(n_1097),
.Y(n_1326)
);

BUFx12f_ASAP7_75t_L g1327 ( 
.A(n_1112),
.Y(n_1327)
);

AOI22xp33_ASAP7_75t_L g1328 ( 
.A1(n_1169),
.A2(n_1193),
.B1(n_908),
.B2(n_902),
.Y(n_1328)
);

AOI22xp33_ASAP7_75t_L g1329 ( 
.A1(n_1169),
.A2(n_1193),
.B1(n_908),
.B2(n_902),
.Y(n_1329)
);

BUFx8_ASAP7_75t_SL g1330 ( 
.A(n_1204),
.Y(n_1330)
);

AOI22xp33_ASAP7_75t_L g1331 ( 
.A1(n_1169),
.A2(n_1193),
.B1(n_742),
.B2(n_1117),
.Y(n_1331)
);

CKINVDCx11_ASAP7_75t_R g1332 ( 
.A(n_1212),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1103),
.Y(n_1333)
);

BUFx12f_ASAP7_75t_L g1334 ( 
.A(n_1112),
.Y(n_1334)
);

OR2x2_ASAP7_75t_L g1335 ( 
.A(n_1107),
.B(n_1096),
.Y(n_1335)
);

INVxp67_ASAP7_75t_SL g1336 ( 
.A(n_1111),
.Y(n_1336)
);

BUFx4f_ASAP7_75t_SL g1337 ( 
.A(n_1204),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1103),
.Y(n_1338)
);

INVx1_ASAP7_75t_SL g1339 ( 
.A(n_1091),
.Y(n_1339)
);

AOI22xp33_ASAP7_75t_L g1340 ( 
.A1(n_1169),
.A2(n_1193),
.B1(n_908),
.B2(n_902),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1103),
.Y(n_1341)
);

OAI22xp5_ASAP7_75t_L g1342 ( 
.A1(n_1124),
.A2(n_977),
.B1(n_1203),
.B2(n_1086),
.Y(n_1342)
);

INVx8_ASAP7_75t_L g1343 ( 
.A(n_1106),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1273),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1273),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1292),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1302),
.Y(n_1347)
);

AND2x2_ASAP7_75t_L g1348 ( 
.A(n_1300),
.B(n_1299),
.Y(n_1348)
);

INVx3_ASAP7_75t_L g1349 ( 
.A(n_1296),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1303),
.Y(n_1350)
);

BUFx3_ASAP7_75t_L g1351 ( 
.A(n_1297),
.Y(n_1351)
);

INVx3_ASAP7_75t_SL g1352 ( 
.A(n_1291),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1305),
.Y(n_1353)
);

OAI21x1_ASAP7_75t_L g1354 ( 
.A1(n_1290),
.A2(n_1294),
.B(n_1298),
.Y(n_1354)
);

AOI21x1_ASAP7_75t_L g1355 ( 
.A1(n_1228),
.A2(n_1313),
.B(n_1231),
.Y(n_1355)
);

AND2x2_ASAP7_75t_L g1356 ( 
.A(n_1295),
.B(n_1282),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_L g1357 ( 
.A(n_1335),
.B(n_1233),
.Y(n_1357)
);

INVx2_ASAP7_75t_L g1358 ( 
.A(n_1227),
.Y(n_1358)
);

O2A1O1Ixp33_ASAP7_75t_SL g1359 ( 
.A1(n_1321),
.A2(n_1326),
.B(n_1241),
.C(n_1239),
.Y(n_1359)
);

OAI21x1_ASAP7_75t_L g1360 ( 
.A1(n_1312),
.A2(n_1325),
.B(n_1272),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1310),
.Y(n_1361)
);

INVx3_ASAP7_75t_L g1362 ( 
.A(n_1296),
.Y(n_1362)
);

AOI21xp5_ASAP7_75t_L g1363 ( 
.A1(n_1321),
.A2(n_1324),
.B(n_1342),
.Y(n_1363)
);

HB1xp67_ASAP7_75t_L g1364 ( 
.A(n_1256),
.Y(n_1364)
);

INVx3_ASAP7_75t_L g1365 ( 
.A(n_1296),
.Y(n_1365)
);

HB1xp67_ASAP7_75t_L g1366 ( 
.A(n_1278),
.Y(n_1366)
);

AOI21x1_ASAP7_75t_L g1367 ( 
.A1(n_1317),
.A2(n_1285),
.B(n_1288),
.Y(n_1367)
);

INVx2_ASAP7_75t_L g1368 ( 
.A(n_1253),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_L g1369 ( 
.A(n_1237),
.B(n_1234),
.Y(n_1369)
);

NAND2xp33_ASAP7_75t_L g1370 ( 
.A(n_1230),
.B(n_1343),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1315),
.Y(n_1371)
);

OR2x2_ASAP7_75t_L g1372 ( 
.A(n_1241),
.B(n_1306),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1323),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_L g1374 ( 
.A(n_1243),
.B(n_1251),
.Y(n_1374)
);

INVx2_ASAP7_75t_L g1375 ( 
.A(n_1333),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1338),
.Y(n_1376)
);

INVx2_ASAP7_75t_SL g1377 ( 
.A(n_1238),
.Y(n_1377)
);

HB1xp67_ASAP7_75t_L g1378 ( 
.A(n_1341),
.Y(n_1378)
);

INVx3_ASAP7_75t_L g1379 ( 
.A(n_1296),
.Y(n_1379)
);

OAI21x1_ASAP7_75t_L g1380 ( 
.A1(n_1311),
.A2(n_1336),
.B(n_1284),
.Y(n_1380)
);

OR2x2_ASAP7_75t_L g1381 ( 
.A(n_1306),
.B(n_1250),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1284),
.Y(n_1382)
);

OAI21x1_ASAP7_75t_L g1383 ( 
.A1(n_1336),
.A2(n_1265),
.B(n_1259),
.Y(n_1383)
);

NOR2x1_ASAP7_75t_L g1384 ( 
.A(n_1247),
.B(n_1243),
.Y(n_1384)
);

HB1xp67_ASAP7_75t_L g1385 ( 
.A(n_1254),
.Y(n_1385)
);

OR2x6_ASAP7_75t_L g1386 ( 
.A(n_1235),
.B(n_1229),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1247),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1259),
.Y(n_1388)
);

CKINVDCx5p33_ASAP7_75t_R g1389 ( 
.A(n_1232),
.Y(n_1389)
);

NOR2xp33_ASAP7_75t_L g1390 ( 
.A(n_1274),
.B(n_1337),
.Y(n_1390)
);

INVx1_ASAP7_75t_SL g1391 ( 
.A(n_1257),
.Y(n_1391)
);

AND2x2_ASAP7_75t_L g1392 ( 
.A(n_1282),
.B(n_1304),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1308),
.Y(n_1393)
);

AND2x2_ASAP7_75t_L g1394 ( 
.A(n_1309),
.B(n_1275),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1265),
.Y(n_1395)
);

HB1xp67_ASAP7_75t_L g1396 ( 
.A(n_1318),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1250),
.Y(n_1397)
);

CKINVDCx20_ASAP7_75t_R g1398 ( 
.A(n_1330),
.Y(n_1398)
);

INVx2_ASAP7_75t_L g1399 ( 
.A(n_1307),
.Y(n_1399)
);

INVx3_ASAP7_75t_L g1400 ( 
.A(n_1301),
.Y(n_1400)
);

AND2x2_ASAP7_75t_L g1401 ( 
.A(n_1275),
.B(n_1261),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1293),
.Y(n_1402)
);

AOI22xp33_ASAP7_75t_L g1403 ( 
.A1(n_1331),
.A2(n_1226),
.B1(n_1314),
.B2(n_1340),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1293),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1261),
.Y(n_1405)
);

A2O1A1Ixp33_ASAP7_75t_L g1406 ( 
.A1(n_1226),
.A2(n_1314),
.B(n_1328),
.C(n_1340),
.Y(n_1406)
);

BUFx2_ASAP7_75t_L g1407 ( 
.A(n_1322),
.Y(n_1407)
);

INVxp67_ASAP7_75t_L g1408 ( 
.A(n_1279),
.Y(n_1408)
);

OAI22xp33_ASAP7_75t_L g1409 ( 
.A1(n_1258),
.A2(n_1283),
.B1(n_1248),
.B2(n_1339),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1301),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1267),
.Y(n_1411)
);

AOI222xp33_ASAP7_75t_L g1412 ( 
.A1(n_1328),
.A2(n_1329),
.B1(n_1281),
.B2(n_1266),
.C1(n_1334),
.C2(n_1255),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1267),
.Y(n_1413)
);

NAND2xp5_ASAP7_75t_L g1414 ( 
.A(n_1249),
.B(n_1286),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1242),
.Y(n_1415)
);

AO31x2_ASAP7_75t_L g1416 ( 
.A1(n_1249),
.A2(n_1260),
.A3(n_1252),
.B(n_1329),
.Y(n_1416)
);

AOI22xp5_ASAP7_75t_L g1417 ( 
.A1(n_1289),
.A2(n_1236),
.B1(n_1270),
.B2(n_1276),
.Y(n_1417)
);

BUFx4f_ASAP7_75t_SL g1418 ( 
.A(n_1320),
.Y(n_1418)
);

OA21x2_ASAP7_75t_L g1419 ( 
.A1(n_1277),
.A2(n_1238),
.B(n_1240),
.Y(n_1419)
);

INVxp67_ASAP7_75t_SL g1420 ( 
.A(n_1287),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1245),
.Y(n_1421)
);

INVx1_ASAP7_75t_SL g1422 ( 
.A(n_1316),
.Y(n_1422)
);

OR2x6_ASAP7_75t_L g1423 ( 
.A(n_1343),
.B(n_1263),
.Y(n_1423)
);

AOI22xp33_ASAP7_75t_L g1424 ( 
.A1(n_1248),
.A2(n_1280),
.B1(n_1263),
.B2(n_1252),
.Y(n_1424)
);

AO32x1_ASAP7_75t_L g1425 ( 
.A1(n_1401),
.A2(n_1260),
.A3(n_1269),
.B1(n_1268),
.B2(n_1327),
.Y(n_1425)
);

AND2x2_ASAP7_75t_L g1426 ( 
.A(n_1356),
.B(n_1244),
.Y(n_1426)
);

AND2x2_ASAP7_75t_L g1427 ( 
.A(n_1356),
.B(n_1244),
.Y(n_1427)
);

AO21x2_ASAP7_75t_L g1428 ( 
.A1(n_1405),
.A2(n_1319),
.B(n_1246),
.Y(n_1428)
);

HB1xp67_ASAP7_75t_L g1429 ( 
.A(n_1378),
.Y(n_1429)
);

NOR2xp33_ASAP7_75t_L g1430 ( 
.A(n_1418),
.B(n_1337),
.Y(n_1430)
);

AND2x4_ASAP7_75t_L g1431 ( 
.A(n_1367),
.B(n_1262),
.Y(n_1431)
);

A2O1A1Ixp33_ASAP7_75t_L g1432 ( 
.A1(n_1384),
.A2(n_1246),
.B(n_1271),
.C(n_1264),
.Y(n_1432)
);

AND2x4_ASAP7_75t_L g1433 ( 
.A(n_1367),
.B(n_1332),
.Y(n_1433)
);

AND2x2_ASAP7_75t_L g1434 ( 
.A(n_1348),
.B(n_1246),
.Y(n_1434)
);

AOI221xp5_ASAP7_75t_L g1435 ( 
.A1(n_1403),
.A2(n_1406),
.B1(n_1359),
.B2(n_1405),
.C(n_1387),
.Y(n_1435)
);

A2O1A1Ixp33_ASAP7_75t_L g1436 ( 
.A1(n_1384),
.A2(n_1363),
.B(n_1401),
.C(n_1394),
.Y(n_1436)
);

BUFx3_ASAP7_75t_L g1437 ( 
.A(n_1419),
.Y(n_1437)
);

AOI22xp5_ASAP7_75t_L g1438 ( 
.A1(n_1412),
.A2(n_1372),
.B1(n_1374),
.B2(n_1394),
.Y(n_1438)
);

AND2x2_ASAP7_75t_L g1439 ( 
.A(n_1371),
.B(n_1373),
.Y(n_1439)
);

A2O1A1Ixp33_ASAP7_75t_SL g1440 ( 
.A1(n_1410),
.A2(n_1400),
.B(n_1390),
.C(n_1402),
.Y(n_1440)
);

AOI211xp5_ASAP7_75t_L g1441 ( 
.A1(n_1409),
.A2(n_1387),
.B(n_1392),
.C(n_1404),
.Y(n_1441)
);

AO32x2_ASAP7_75t_L g1442 ( 
.A1(n_1377),
.A2(n_1364),
.A3(n_1397),
.B1(n_1385),
.B2(n_1366),
.Y(n_1442)
);

AND2x2_ASAP7_75t_L g1443 ( 
.A(n_1373),
.B(n_1376),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_L g1444 ( 
.A(n_1408),
.B(n_1396),
.Y(n_1444)
);

AOI22xp5_ASAP7_75t_L g1445 ( 
.A1(n_1392),
.A2(n_1370),
.B1(n_1351),
.B2(n_1369),
.Y(n_1445)
);

OA21x2_ASAP7_75t_L g1446 ( 
.A1(n_1354),
.A2(n_1383),
.B(n_1380),
.Y(n_1446)
);

AND2x2_ASAP7_75t_L g1447 ( 
.A(n_1404),
.B(n_1358),
.Y(n_1447)
);

BUFx3_ASAP7_75t_L g1448 ( 
.A(n_1419),
.Y(n_1448)
);

OAI21xp5_ASAP7_75t_L g1449 ( 
.A1(n_1355),
.A2(n_1360),
.B(n_1410),
.Y(n_1449)
);

INVxp67_ASAP7_75t_L g1450 ( 
.A(n_1407),
.Y(n_1450)
);

AOI21xp5_ASAP7_75t_L g1451 ( 
.A1(n_1354),
.A2(n_1360),
.B(n_1400),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1346),
.Y(n_1452)
);

A2O1A1Ixp33_ASAP7_75t_L g1453 ( 
.A1(n_1381),
.A2(n_1414),
.B(n_1383),
.C(n_1417),
.Y(n_1453)
);

BUFx3_ASAP7_75t_L g1454 ( 
.A(n_1419),
.Y(n_1454)
);

HB1xp67_ASAP7_75t_L g1455 ( 
.A(n_1407),
.Y(n_1455)
);

NAND2xp5_ASAP7_75t_L g1456 ( 
.A(n_1357),
.B(n_1368),
.Y(n_1456)
);

AND2x2_ASAP7_75t_L g1457 ( 
.A(n_1375),
.B(n_1380),
.Y(n_1457)
);

OR2x2_ASAP7_75t_L g1458 ( 
.A(n_1381),
.B(n_1344),
.Y(n_1458)
);

OAI22xp5_ASAP7_75t_SL g1459 ( 
.A1(n_1352),
.A2(n_1417),
.B1(n_1398),
.B2(n_1424),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_L g1460 ( 
.A(n_1375),
.B(n_1391),
.Y(n_1460)
);

OR2x2_ASAP7_75t_L g1461 ( 
.A(n_1344),
.B(n_1345),
.Y(n_1461)
);

OAI21xp5_ASAP7_75t_L g1462 ( 
.A1(n_1355),
.A2(n_1400),
.B(n_1415),
.Y(n_1462)
);

OAI22xp5_ASAP7_75t_L g1463 ( 
.A1(n_1352),
.A2(n_1423),
.B1(n_1411),
.B2(n_1413),
.Y(n_1463)
);

OR2x2_ASAP7_75t_L g1464 ( 
.A(n_1345),
.B(n_1397),
.Y(n_1464)
);

NOR2xp33_ASAP7_75t_L g1465 ( 
.A(n_1352),
.B(n_1389),
.Y(n_1465)
);

BUFx3_ASAP7_75t_L g1466 ( 
.A(n_1419),
.Y(n_1466)
);

AND2x2_ASAP7_75t_L g1467 ( 
.A(n_1399),
.B(n_1382),
.Y(n_1467)
);

AOI22xp33_ASAP7_75t_SL g1468 ( 
.A1(n_1388),
.A2(n_1393),
.B1(n_1395),
.B2(n_1416),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1347),
.Y(n_1469)
);

NOR2xp33_ASAP7_75t_SL g1470 ( 
.A(n_1420),
.B(n_1422),
.Y(n_1470)
);

AND2x2_ASAP7_75t_L g1471 ( 
.A(n_1349),
.B(n_1365),
.Y(n_1471)
);

AND2x2_ASAP7_75t_L g1472 ( 
.A(n_1442),
.B(n_1379),
.Y(n_1472)
);

AND2x2_ASAP7_75t_L g1473 ( 
.A(n_1442),
.B(n_1457),
.Y(n_1473)
);

INVx2_ASAP7_75t_L g1474 ( 
.A(n_1457),
.Y(n_1474)
);

INVx2_ASAP7_75t_L g1475 ( 
.A(n_1452),
.Y(n_1475)
);

AND2x2_ASAP7_75t_L g1476 ( 
.A(n_1442),
.B(n_1365),
.Y(n_1476)
);

OAI22xp5_ASAP7_75t_L g1477 ( 
.A1(n_1436),
.A2(n_1393),
.B1(n_1386),
.B2(n_1421),
.Y(n_1477)
);

INVx2_ASAP7_75t_L g1478 ( 
.A(n_1452),
.Y(n_1478)
);

AOI22xp33_ASAP7_75t_L g1479 ( 
.A1(n_1435),
.A2(n_1350),
.B1(n_1353),
.B2(n_1361),
.Y(n_1479)
);

AND2x2_ASAP7_75t_L g1480 ( 
.A(n_1442),
.B(n_1362),
.Y(n_1480)
);

OR2x2_ASAP7_75t_L g1481 ( 
.A(n_1458),
.B(n_1416),
.Y(n_1481)
);

INVx2_ASAP7_75t_L g1482 ( 
.A(n_1469),
.Y(n_1482)
);

OR2x2_ASAP7_75t_L g1483 ( 
.A(n_1458),
.B(n_1416),
.Y(n_1483)
);

INVx2_ASAP7_75t_SL g1484 ( 
.A(n_1461),
.Y(n_1484)
);

INVx2_ASAP7_75t_L g1485 ( 
.A(n_1446),
.Y(n_1485)
);

INVx2_ASAP7_75t_L g1486 ( 
.A(n_1446),
.Y(n_1486)
);

OR2x2_ASAP7_75t_L g1487 ( 
.A(n_1461),
.B(n_1416),
.Y(n_1487)
);

BUFx3_ASAP7_75t_L g1488 ( 
.A(n_1433),
.Y(n_1488)
);

NAND2x1_ASAP7_75t_L g1489 ( 
.A(n_1433),
.B(n_1365),
.Y(n_1489)
);

AND2x2_ASAP7_75t_L g1490 ( 
.A(n_1439),
.B(n_1416),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_L g1491 ( 
.A(n_1429),
.B(n_1443),
.Y(n_1491)
);

INVx2_ASAP7_75t_SL g1492 ( 
.A(n_1433),
.Y(n_1492)
);

AND2x2_ASAP7_75t_L g1493 ( 
.A(n_1443),
.B(n_1416),
.Y(n_1493)
);

INVx2_ASAP7_75t_L g1494 ( 
.A(n_1446),
.Y(n_1494)
);

INVx2_ASAP7_75t_L g1495 ( 
.A(n_1446),
.Y(n_1495)
);

OR2x2_ASAP7_75t_L g1496 ( 
.A(n_1464),
.B(n_1361),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1490),
.B(n_1434),
.Y(n_1497)
);

INVx2_ASAP7_75t_L g1498 ( 
.A(n_1474),
.Y(n_1498)
);

AND2x2_ASAP7_75t_L g1499 ( 
.A(n_1490),
.B(n_1434),
.Y(n_1499)
);

AOI22xp5_ASAP7_75t_L g1500 ( 
.A1(n_1479),
.A2(n_1438),
.B1(n_1441),
.B2(n_1445),
.Y(n_1500)
);

AND2x2_ASAP7_75t_L g1501 ( 
.A(n_1490),
.B(n_1455),
.Y(n_1501)
);

INVx1_ASAP7_75t_SL g1502 ( 
.A(n_1496),
.Y(n_1502)
);

OR2x2_ASAP7_75t_L g1503 ( 
.A(n_1487),
.B(n_1464),
.Y(n_1503)
);

AOI33xp33_ASAP7_75t_L g1504 ( 
.A1(n_1473),
.A2(n_1468),
.A3(n_1426),
.B1(n_1427),
.B2(n_1438),
.B3(n_1431),
.Y(n_1504)
);

AND2x2_ASAP7_75t_L g1505 ( 
.A(n_1490),
.B(n_1493),
.Y(n_1505)
);

AND2x2_ASAP7_75t_L g1506 ( 
.A(n_1493),
.B(n_1473),
.Y(n_1506)
);

INVx3_ASAP7_75t_L g1507 ( 
.A(n_1488),
.Y(n_1507)
);

AND2x2_ASAP7_75t_L g1508 ( 
.A(n_1493),
.B(n_1471),
.Y(n_1508)
);

OR2x2_ASAP7_75t_L g1509 ( 
.A(n_1487),
.B(n_1460),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1475),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1475),
.Y(n_1511)
);

AND2x2_ASAP7_75t_L g1512 ( 
.A(n_1493),
.B(n_1471),
.Y(n_1512)
);

INVx5_ASAP7_75t_L g1513 ( 
.A(n_1472),
.Y(n_1513)
);

BUFx2_ASAP7_75t_L g1514 ( 
.A(n_1488),
.Y(n_1514)
);

BUFx2_ASAP7_75t_L g1515 ( 
.A(n_1488),
.Y(n_1515)
);

AND2x2_ASAP7_75t_L g1516 ( 
.A(n_1473),
.B(n_1472),
.Y(n_1516)
);

INVx2_ASAP7_75t_L g1517 ( 
.A(n_1474),
.Y(n_1517)
);

AOI221xp5_ASAP7_75t_L g1518 ( 
.A1(n_1473),
.A2(n_1453),
.B1(n_1449),
.B2(n_1432),
.C(n_1431),
.Y(n_1518)
);

AOI33xp33_ASAP7_75t_L g1519 ( 
.A1(n_1479),
.A2(n_1427),
.A3(n_1426),
.B1(n_1431),
.B2(n_1445),
.B3(n_1467),
.Y(n_1519)
);

NOR2xp33_ASAP7_75t_L g1520 ( 
.A(n_1491),
.B(n_1465),
.Y(n_1520)
);

NOR2xp67_ASAP7_75t_L g1521 ( 
.A(n_1492),
.B(n_1451),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1475),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_L g1523 ( 
.A(n_1484),
.B(n_1450),
.Y(n_1523)
);

AOI21xp5_ASAP7_75t_L g1524 ( 
.A1(n_1477),
.A2(n_1425),
.B(n_1440),
.Y(n_1524)
);

CKINVDCx5p33_ASAP7_75t_R g1525 ( 
.A(n_1491),
.Y(n_1525)
);

INVxp67_ASAP7_75t_SL g1526 ( 
.A(n_1485),
.Y(n_1526)
);

AOI221xp5_ASAP7_75t_L g1527 ( 
.A1(n_1487),
.A2(n_1459),
.B1(n_1444),
.B2(n_1447),
.C(n_1428),
.Y(n_1527)
);

INVxp67_ASAP7_75t_SL g1528 ( 
.A(n_1485),
.Y(n_1528)
);

OAI221xp5_ASAP7_75t_L g1529 ( 
.A1(n_1477),
.A2(n_1470),
.B1(n_1437),
.B2(n_1448),
.C(n_1454),
.Y(n_1529)
);

OAI31xp33_ASAP7_75t_L g1530 ( 
.A1(n_1477),
.A2(n_1466),
.A3(n_1454),
.B(n_1448),
.Y(n_1530)
);

INVx2_ASAP7_75t_L g1531 ( 
.A(n_1485),
.Y(n_1531)
);

OAI221xp5_ASAP7_75t_L g1532 ( 
.A1(n_1481),
.A2(n_1466),
.B1(n_1462),
.B2(n_1456),
.C(n_1463),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1510),
.Y(n_1533)
);

AND2x2_ASAP7_75t_L g1534 ( 
.A(n_1506),
.B(n_1472),
.Y(n_1534)
);

INVx2_ASAP7_75t_L g1535 ( 
.A(n_1498),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_L g1536 ( 
.A(n_1502),
.B(n_1484),
.Y(n_1536)
);

INVx2_ASAP7_75t_SL g1537 ( 
.A(n_1513),
.Y(n_1537)
);

AND2x2_ASAP7_75t_L g1538 ( 
.A(n_1506),
.B(n_1472),
.Y(n_1538)
);

INVx2_ASAP7_75t_L g1539 ( 
.A(n_1498),
.Y(n_1539)
);

AND2x2_ASAP7_75t_L g1540 ( 
.A(n_1506),
.B(n_1476),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1510),
.Y(n_1541)
);

NAND2x1_ASAP7_75t_L g1542 ( 
.A(n_1507),
.B(n_1492),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1511),
.Y(n_1543)
);

AND2x2_ASAP7_75t_L g1544 ( 
.A(n_1516),
.B(n_1476),
.Y(n_1544)
);

INVx2_ASAP7_75t_L g1545 ( 
.A(n_1498),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1511),
.Y(n_1546)
);

AND2x4_ASAP7_75t_L g1547 ( 
.A(n_1513),
.B(n_1488),
.Y(n_1547)
);

BUFx2_ASAP7_75t_L g1548 ( 
.A(n_1513),
.Y(n_1548)
);

NOR3xp33_ASAP7_75t_L g1549 ( 
.A(n_1518),
.B(n_1494),
.C(n_1485),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1516),
.B(n_1476),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_L g1551 ( 
.A(n_1502),
.B(n_1484),
.Y(n_1551)
);

AND2x2_ASAP7_75t_L g1552 ( 
.A(n_1516),
.B(n_1513),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1522),
.Y(n_1553)
);

AND2x4_ASAP7_75t_L g1554 ( 
.A(n_1513),
.B(n_1492),
.Y(n_1554)
);

OR2x2_ASAP7_75t_L g1555 ( 
.A(n_1505),
.B(n_1484),
.Y(n_1555)
);

AND2x2_ASAP7_75t_L g1556 ( 
.A(n_1513),
.B(n_1476),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_L g1557 ( 
.A(n_1505),
.B(n_1478),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1513),
.B(n_1480),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1513),
.B(n_1505),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1522),
.Y(n_1560)
);

AND2x2_ASAP7_75t_L g1561 ( 
.A(n_1508),
.B(n_1480),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1503),
.B(n_1478),
.Y(n_1562)
);

NOR2x1_ASAP7_75t_L g1563 ( 
.A(n_1507),
.B(n_1489),
.Y(n_1563)
);

AND2x2_ASAP7_75t_L g1564 ( 
.A(n_1508),
.B(n_1480),
.Y(n_1564)
);

NAND2xp5_ASAP7_75t_L g1565 ( 
.A(n_1503),
.B(n_1478),
.Y(n_1565)
);

INVx1_ASAP7_75t_SL g1566 ( 
.A(n_1514),
.Y(n_1566)
);

NAND2xp5_ASAP7_75t_L g1567 ( 
.A(n_1503),
.B(n_1482),
.Y(n_1567)
);

INVxp67_ASAP7_75t_SL g1568 ( 
.A(n_1526),
.Y(n_1568)
);

INVx2_ASAP7_75t_L g1569 ( 
.A(n_1517),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1508),
.B(n_1480),
.Y(n_1570)
);

AND2x2_ASAP7_75t_SL g1571 ( 
.A(n_1549),
.B(n_1518),
.Y(n_1571)
);

NAND2xp5_ASAP7_75t_L g1572 ( 
.A(n_1549),
.B(n_1519),
.Y(n_1572)
);

OR2x2_ASAP7_75t_L g1573 ( 
.A(n_1555),
.B(n_1509),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1533),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_L g1575 ( 
.A(n_1566),
.B(n_1501),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_L g1576 ( 
.A(n_1566),
.B(n_1501),
.Y(n_1576)
);

AND2x2_ASAP7_75t_L g1577 ( 
.A(n_1559),
.B(n_1514),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1559),
.B(n_1515),
.Y(n_1578)
);

OR2x2_ASAP7_75t_L g1579 ( 
.A(n_1555),
.B(n_1509),
.Y(n_1579)
);

INVxp67_ASAP7_75t_L g1580 ( 
.A(n_1536),
.Y(n_1580)
);

INVx2_ASAP7_75t_L g1581 ( 
.A(n_1555),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1533),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_L g1583 ( 
.A(n_1536),
.B(n_1501),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1546),
.Y(n_1584)
);

OR2x2_ASAP7_75t_L g1585 ( 
.A(n_1551),
.B(n_1509),
.Y(n_1585)
);

OR2x2_ASAP7_75t_L g1586 ( 
.A(n_1551),
.B(n_1523),
.Y(n_1586)
);

OR2x2_ASAP7_75t_L g1587 ( 
.A(n_1557),
.B(n_1523),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1546),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_L g1589 ( 
.A(n_1562),
.B(n_1525),
.Y(n_1589)
);

OR2x2_ASAP7_75t_L g1590 ( 
.A(n_1557),
.B(n_1517),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1562),
.B(n_1504),
.Y(n_1591)
);

AND2x2_ASAP7_75t_L g1592 ( 
.A(n_1559),
.B(n_1552),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_L g1593 ( 
.A(n_1565),
.B(n_1527),
.Y(n_1593)
);

NAND2xp67_ASAP7_75t_L g1594 ( 
.A(n_1552),
.B(n_1524),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1565),
.B(n_1527),
.Y(n_1595)
);

INVx2_ASAP7_75t_L g1596 ( 
.A(n_1535),
.Y(n_1596)
);

NOR2xp33_ASAP7_75t_L g1597 ( 
.A(n_1548),
.B(n_1520),
.Y(n_1597)
);

INVx2_ASAP7_75t_SL g1598 ( 
.A(n_1547),
.Y(n_1598)
);

OR2x2_ASAP7_75t_L g1599 ( 
.A(n_1567),
.B(n_1517),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1553),
.Y(n_1600)
);

AND2x2_ASAP7_75t_L g1601 ( 
.A(n_1552),
.B(n_1515),
.Y(n_1601)
);

BUFx2_ASAP7_75t_L g1602 ( 
.A(n_1548),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1553),
.Y(n_1603)
);

AOI22xp5_ASAP7_75t_L g1604 ( 
.A1(n_1534),
.A2(n_1500),
.B1(n_1428),
.B2(n_1529),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1560),
.Y(n_1605)
);

AND2x2_ASAP7_75t_L g1606 ( 
.A(n_1548),
.B(n_1507),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1567),
.B(n_1512),
.Y(n_1607)
);

INVx2_ASAP7_75t_SL g1608 ( 
.A(n_1547),
.Y(n_1608)
);

AND2x2_ASAP7_75t_L g1609 ( 
.A(n_1547),
.B(n_1534),
.Y(n_1609)
);

INVx2_ASAP7_75t_L g1610 ( 
.A(n_1535),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1560),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1541),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1574),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1582),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_SL g1615 ( 
.A(n_1571),
.B(n_1547),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1584),
.Y(n_1616)
);

AOI22xp33_ASAP7_75t_L g1617 ( 
.A1(n_1571),
.A2(n_1500),
.B1(n_1524),
.B2(n_1529),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1588),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_L g1619 ( 
.A(n_1572),
.B(n_1512),
.Y(n_1619)
);

OR2x2_ASAP7_75t_L g1620 ( 
.A(n_1591),
.B(n_1544),
.Y(n_1620)
);

INVxp67_ASAP7_75t_L g1621 ( 
.A(n_1602),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1600),
.Y(n_1622)
);

NOR2xp33_ASAP7_75t_L g1623 ( 
.A(n_1597),
.B(n_1430),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_L g1624 ( 
.A(n_1593),
.B(n_1512),
.Y(n_1624)
);

NOR2xp67_ASAP7_75t_L g1625 ( 
.A(n_1598),
.B(n_1537),
.Y(n_1625)
);

INVx2_ASAP7_75t_L g1626 ( 
.A(n_1609),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1603),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1605),
.Y(n_1628)
);

OR2x2_ASAP7_75t_L g1629 ( 
.A(n_1586),
.B(n_1544),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_L g1630 ( 
.A(n_1595),
.B(n_1497),
.Y(n_1630)
);

NOR2xp33_ASAP7_75t_L g1631 ( 
.A(n_1594),
.B(n_1542),
.Y(n_1631)
);

NAND4xp25_ASAP7_75t_L g1632 ( 
.A(n_1602),
.B(n_1556),
.C(n_1558),
.D(n_1563),
.Y(n_1632)
);

INVx2_ASAP7_75t_SL g1633 ( 
.A(n_1592),
.Y(n_1633)
);

OR2x2_ASAP7_75t_L g1634 ( 
.A(n_1586),
.B(n_1544),
.Y(n_1634)
);

INVx2_ASAP7_75t_L g1635 ( 
.A(n_1609),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1611),
.Y(n_1636)
);

NOR2xp33_ASAP7_75t_L g1637 ( 
.A(n_1589),
.B(n_1497),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1612),
.Y(n_1638)
);

AOI22xp5_ASAP7_75t_L g1639 ( 
.A1(n_1604),
.A2(n_1428),
.B1(n_1532),
.B2(n_1483),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_L g1640 ( 
.A(n_1580),
.B(n_1497),
.Y(n_1640)
);

AND2x4_ASAP7_75t_L g1641 ( 
.A(n_1598),
.B(n_1547),
.Y(n_1641)
);

NOR2xp33_ASAP7_75t_L g1642 ( 
.A(n_1594),
.B(n_1542),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_L g1643 ( 
.A(n_1581),
.B(n_1499),
.Y(n_1643)
);

INVxp67_ASAP7_75t_L g1644 ( 
.A(n_1596),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_L g1645 ( 
.A(n_1581),
.B(n_1573),
.Y(n_1645)
);

NOR2xp33_ASAP7_75t_SL g1646 ( 
.A(n_1577),
.B(n_1530),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_L g1647 ( 
.A(n_1573),
.B(n_1499),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1638),
.Y(n_1648)
);

AOI322xp5_ASAP7_75t_L g1649 ( 
.A1(n_1617),
.A2(n_1568),
.A3(n_1550),
.B1(n_1540),
.B2(n_1538),
.C1(n_1534),
.C2(n_1570),
.Y(n_1649)
);

AOI22xp5_ASAP7_75t_L g1650 ( 
.A1(n_1617),
.A2(n_1532),
.B1(n_1521),
.B2(n_1481),
.Y(n_1650)
);

NOR2xp33_ASAP7_75t_L g1651 ( 
.A(n_1623),
.B(n_1608),
.Y(n_1651)
);

AOI21xp5_ASAP7_75t_L g1652 ( 
.A1(n_1615),
.A2(n_1646),
.B(n_1642),
.Y(n_1652)
);

OR2x2_ASAP7_75t_L g1653 ( 
.A(n_1630),
.B(n_1585),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1613),
.Y(n_1654)
);

NAND2xp5_ASAP7_75t_L g1655 ( 
.A(n_1621),
.B(n_1575),
.Y(n_1655)
);

NOR2xp33_ASAP7_75t_L g1656 ( 
.A(n_1623),
.B(n_1608),
.Y(n_1656)
);

INVxp67_ASAP7_75t_L g1657 ( 
.A(n_1621),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_L g1658 ( 
.A(n_1619),
.B(n_1576),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_SL g1659 ( 
.A(n_1631),
.B(n_1554),
.Y(n_1659)
);

INVx2_ASAP7_75t_L g1660 ( 
.A(n_1641),
.Y(n_1660)
);

AND2x2_ASAP7_75t_L g1661 ( 
.A(n_1633),
.B(n_1626),
.Y(n_1661)
);

OAI22xp5_ASAP7_75t_L g1662 ( 
.A1(n_1624),
.A2(n_1554),
.B1(n_1579),
.B2(n_1537),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1614),
.Y(n_1663)
);

INVx2_ASAP7_75t_L g1664 ( 
.A(n_1641),
.Y(n_1664)
);

OR2x2_ASAP7_75t_L g1665 ( 
.A(n_1620),
.B(n_1585),
.Y(n_1665)
);

AOI32xp33_ASAP7_75t_L g1666 ( 
.A1(n_1631),
.A2(n_1568),
.A3(n_1540),
.B1(n_1538),
.B2(n_1550),
.Y(n_1666)
);

NOR2x1_ASAP7_75t_L g1667 ( 
.A(n_1632),
.B(n_1563),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1616),
.Y(n_1668)
);

OAI31xp33_ASAP7_75t_L g1669 ( 
.A1(n_1642),
.A2(n_1530),
.A3(n_1556),
.B(n_1558),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1618),
.Y(n_1670)
);

NOR2x1_ASAP7_75t_L g1671 ( 
.A(n_1625),
.B(n_1542),
.Y(n_1671)
);

INVx2_ASAP7_75t_L g1672 ( 
.A(n_1635),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_L g1673 ( 
.A(n_1651),
.B(n_1645),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1665),
.Y(n_1674)
);

AOI22xp5_ASAP7_75t_L g1675 ( 
.A1(n_1650),
.A2(n_1639),
.B1(n_1644),
.B2(n_1637),
.Y(n_1675)
);

AOI22xp5_ASAP7_75t_L g1676 ( 
.A1(n_1652),
.A2(n_1644),
.B1(n_1521),
.B2(n_1643),
.Y(n_1676)
);

OAI322xp33_ASAP7_75t_L g1677 ( 
.A1(n_1657),
.A2(n_1634),
.A3(n_1629),
.B1(n_1636),
.B2(n_1628),
.C1(n_1622),
.C2(n_1627),
.Y(n_1677)
);

AOI22xp5_ASAP7_75t_L g1678 ( 
.A1(n_1651),
.A2(n_1610),
.B1(n_1596),
.B2(n_1487),
.Y(n_1678)
);

AOI32xp33_ASAP7_75t_L g1679 ( 
.A1(n_1667),
.A2(n_1540),
.A3(n_1538),
.B1(n_1550),
.B2(n_1556),
.Y(n_1679)
);

OA21x2_ASAP7_75t_L g1680 ( 
.A1(n_1657),
.A2(n_1610),
.B(n_1606),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1672),
.Y(n_1681)
);

NAND2xp5_ASAP7_75t_L g1682 ( 
.A(n_1656),
.B(n_1647),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1656),
.B(n_1577),
.Y(n_1683)
);

NOR2xp67_ASAP7_75t_SL g1684 ( 
.A(n_1660),
.B(n_1492),
.Y(n_1684)
);

AND2x2_ASAP7_75t_L g1685 ( 
.A(n_1661),
.B(n_1664),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1672),
.Y(n_1686)
);

OAI22xp33_ASAP7_75t_L g1687 ( 
.A1(n_1653),
.A2(n_1658),
.B1(n_1537),
.B2(n_1481),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_L g1688 ( 
.A(n_1654),
.B(n_1640),
.Y(n_1688)
);

INVx2_ASAP7_75t_SL g1689 ( 
.A(n_1659),
.Y(n_1689)
);

INVxp67_ASAP7_75t_L g1690 ( 
.A(n_1655),
.Y(n_1690)
);

AOI221xp5_ASAP7_75t_SL g1691 ( 
.A1(n_1662),
.A2(n_1606),
.B1(n_1592),
.B2(n_1601),
.C(n_1578),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_L g1692 ( 
.A(n_1663),
.B(n_1579),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_L g1693 ( 
.A(n_1683),
.B(n_1668),
.Y(n_1693)
);

AOI211xp5_ASAP7_75t_L g1694 ( 
.A1(n_1677),
.A2(n_1669),
.B(n_1659),
.C(n_1670),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_L g1695 ( 
.A(n_1685),
.B(n_1648),
.Y(n_1695)
);

INVx2_ASAP7_75t_L g1696 ( 
.A(n_1680),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1674),
.Y(n_1697)
);

NAND2xp5_ASAP7_75t_L g1698 ( 
.A(n_1690),
.B(n_1673),
.Y(n_1698)
);

OAI21xp5_ASAP7_75t_L g1699 ( 
.A1(n_1680),
.A2(n_1649),
.B(n_1671),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1692),
.Y(n_1700)
);

HB1xp67_ASAP7_75t_L g1701 ( 
.A(n_1689),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1681),
.Y(n_1702)
);

A2O1A1Ixp33_ASAP7_75t_L g1703 ( 
.A1(n_1699),
.A2(n_1675),
.B(n_1678),
.C(n_1676),
.Y(n_1703)
);

AOI211xp5_ASAP7_75t_L g1704 ( 
.A1(n_1699),
.A2(n_1687),
.B(n_1688),
.C(n_1682),
.Y(n_1704)
);

HB1xp67_ASAP7_75t_SL g1705 ( 
.A(n_1701),
.Y(n_1705)
);

AOI221xp5_ASAP7_75t_L g1706 ( 
.A1(n_1696),
.A2(n_1686),
.B1(n_1678),
.B2(n_1691),
.C(n_1679),
.Y(n_1706)
);

OAI221xp5_ASAP7_75t_SL g1707 ( 
.A1(n_1694),
.A2(n_1666),
.B1(n_1684),
.B2(n_1590),
.C(n_1587),
.Y(n_1707)
);

NAND3xp33_ASAP7_75t_L g1708 ( 
.A(n_1697),
.B(n_1578),
.C(n_1601),
.Y(n_1708)
);

NAND3xp33_ASAP7_75t_SL g1709 ( 
.A(n_1698),
.B(n_1558),
.C(n_1587),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1695),
.Y(n_1710)
);

NOR3xp33_ASAP7_75t_L g1711 ( 
.A(n_1702),
.B(n_1599),
.C(n_1545),
.Y(n_1711)
);

OAI221xp5_ASAP7_75t_SL g1712 ( 
.A1(n_1703),
.A2(n_1700),
.B1(n_1693),
.B2(n_1599),
.C(n_1590),
.Y(n_1712)
);

AOI21xp5_ASAP7_75t_L g1713 ( 
.A1(n_1704),
.A2(n_1707),
.B(n_1706),
.Y(n_1713)
);

AOI21xp33_ASAP7_75t_L g1714 ( 
.A1(n_1710),
.A2(n_1535),
.B(n_1569),
.Y(n_1714)
);

NAND3xp33_ASAP7_75t_L g1715 ( 
.A(n_1711),
.B(n_1539),
.C(n_1535),
.Y(n_1715)
);

A2O1A1Ixp33_ASAP7_75t_L g1716 ( 
.A1(n_1708),
.A2(n_1528),
.B(n_1526),
.C(n_1531),
.Y(n_1716)
);

AOI211xp5_ASAP7_75t_L g1717 ( 
.A1(n_1713),
.A2(n_1712),
.B(n_1709),
.C(n_1714),
.Y(n_1717)
);

CKINVDCx16_ASAP7_75t_R g1718 ( 
.A(n_1716),
.Y(n_1718)
);

AOI222xp33_ASAP7_75t_L g1719 ( 
.A1(n_1715),
.A2(n_1705),
.B1(n_1528),
.B2(n_1495),
.C1(n_1494),
.C2(n_1485),
.Y(n_1719)
);

AOI31xp33_ASAP7_75t_L g1720 ( 
.A1(n_1713),
.A2(n_1554),
.A3(n_1583),
.B(n_1607),
.Y(n_1720)
);

OAI221xp5_ASAP7_75t_SL g1721 ( 
.A1(n_1713),
.A2(n_1561),
.B1(n_1564),
.B2(n_1570),
.C(n_1495),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1712),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1720),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1718),
.Y(n_1724)
);

CKINVDCx20_ASAP7_75t_R g1725 ( 
.A(n_1722),
.Y(n_1725)
);

NOR2x1_ASAP7_75t_L g1726 ( 
.A(n_1717),
.B(n_1554),
.Y(n_1726)
);

AND2x4_ASAP7_75t_L g1727 ( 
.A(n_1721),
.B(n_1554),
.Y(n_1727)
);

AND2x4_ASAP7_75t_L g1728 ( 
.A(n_1726),
.B(n_1507),
.Y(n_1728)
);

AND2x2_ASAP7_75t_L g1729 ( 
.A(n_1723),
.B(n_1719),
.Y(n_1729)
);

AOI221xp5_ASAP7_75t_L g1730 ( 
.A1(n_1724),
.A2(n_1531),
.B1(n_1486),
.B2(n_1495),
.C(n_1494),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1729),
.Y(n_1731)
);

OAI22xp5_ASAP7_75t_L g1732 ( 
.A1(n_1731),
.A2(n_1725),
.B1(n_1728),
.B2(n_1727),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1732),
.Y(n_1733)
);

INVx2_ASAP7_75t_L g1734 ( 
.A(n_1733),
.Y(n_1734)
);

OAI22xp33_ASAP7_75t_SL g1735 ( 
.A1(n_1734),
.A2(n_1730),
.B1(n_1569),
.B2(n_1545),
.Y(n_1735)
);

OAI21xp5_ASAP7_75t_L g1736 ( 
.A1(n_1735),
.A2(n_1539),
.B(n_1569),
.Y(n_1736)
);

AND2x2_ASAP7_75t_L g1737 ( 
.A(n_1736),
.B(n_1570),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1737),
.Y(n_1738)
);

OAI221xp5_ASAP7_75t_L g1739 ( 
.A1(n_1738),
.A2(n_1423),
.B1(n_1543),
.B2(n_1541),
.C(n_1545),
.Y(n_1739)
);

AOI211xp5_ASAP7_75t_L g1740 ( 
.A1(n_1739),
.A2(n_1543),
.B(n_1564),
.C(n_1561),
.Y(n_1740)
);


endmodule