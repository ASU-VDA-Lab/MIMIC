module fake_jpeg_21433_n_148 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_148);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_148;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_13),
.Y(n_48)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_5),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_4),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_29),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_20),
.Y(n_54)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_6),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_3),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_31),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

BUFx10_ASAP7_75t_L g59 ( 
.A(n_2),
.Y(n_59)
);

BUFx4f_ASAP7_75t_SL g60 ( 
.A(n_35),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_3),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_26),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_7),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_30),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_5),
.Y(n_65)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_19),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_37),
.Y(n_67)
);

BUFx24_ASAP7_75t_L g68 ( 
.A(n_0),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_1),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_1),
.Y(n_71)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_24),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_59),
.B(n_0),
.Y(n_74)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_74),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_68),
.Y(n_75)
);

INVx3_ASAP7_75t_SL g92 ( 
.A(n_75),
.Y(n_92)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_76),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_77),
.Y(n_86)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_68),
.Y(n_78)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_78),
.Y(n_90)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_71),
.Y(n_79)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_79),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_50),
.B(n_2),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_80),
.A2(n_61),
.B1(n_69),
.B2(n_63),
.Y(n_87)
);

BUFx24_ASAP7_75t_L g81 ( 
.A(n_60),
.Y(n_81)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_81),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_81),
.A2(n_49),
.B1(n_55),
.B2(n_72),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_83),
.A2(n_85),
.B1(n_59),
.B2(n_54),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_77),
.A2(n_52),
.B1(n_65),
.B2(n_66),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_87),
.B(n_71),
.Y(n_106)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_74),
.Y(n_89)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_89),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_88),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_93),
.B(n_97),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_82),
.B(n_62),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_95),
.B(n_99),
.Y(n_107)
);

BUFx2_ASAP7_75t_L g96 ( 
.A(n_86),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_90),
.B(n_56),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_83),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_98),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_85),
.B(n_58),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g116 ( 
.A1(n_100),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_91),
.A2(n_53),
.B1(n_57),
.B2(n_67),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_101),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_119)
);

INVx1_ASAP7_75t_SL g102 ( 
.A(n_86),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_102),
.B(n_106),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_92),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_103),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_92),
.A2(n_51),
.B1(n_48),
.B2(n_70),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_104),
.A2(n_105),
.B1(n_9),
.B2(n_11),
.Y(n_121)
);

OAI22xp33_ASAP7_75t_L g105 ( 
.A1(n_84),
.A2(n_70),
.B1(n_64),
.B2(n_73),
.Y(n_105)
);

AOI21xp33_ASAP7_75t_L g108 ( 
.A1(n_94),
.A2(n_60),
.B(n_59),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_108),
.A2(n_17),
.B(n_23),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_101),
.A2(n_73),
.B1(n_64),
.B2(n_22),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_110),
.A2(n_116),
.B1(n_121),
.B2(n_33),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_105),
.B(n_21),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_111),
.B(n_116),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_96),
.B(n_18),
.C(n_46),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_114),
.B(n_14),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_102),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_115),
.B(n_12),
.Y(n_122)
);

XNOR2x1_ASAP7_75t_SL g118 ( 
.A(n_94),
.B(n_8),
.Y(n_118)
);

AOI21xp33_ASAP7_75t_L g131 ( 
.A1(n_118),
.A2(n_34),
.B(n_36),
.Y(n_131)
);

AO21x2_ASAP7_75t_L g128 ( 
.A1(n_119),
.A2(n_25),
.B(n_27),
.Y(n_128)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_96),
.Y(n_120)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_120),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_122),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_123),
.A2(n_124),
.B(n_125),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_112),
.A2(n_15),
.B(n_16),
.Y(n_125)
);

OA21x2_ASAP7_75t_L g134 ( 
.A1(n_126),
.A2(n_128),
.B(n_131),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_117),
.B(n_28),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_129),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_130),
.A2(n_122),
.B1(n_107),
.B2(n_109),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_136),
.A2(n_112),
.B1(n_119),
.B2(n_113),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_133),
.Y(n_137)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_137),
.Y(n_139)
);

INVx2_ASAP7_75t_SL g140 ( 
.A(n_139),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_140),
.B(n_132),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_141),
.A2(n_132),
.B(n_135),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_142),
.B(n_138),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_143),
.B(n_128),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_144),
.B(n_128),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_145),
.B(n_134),
.Y(n_146)
);

AOI31xp33_ASAP7_75t_L g147 ( 
.A1(n_146),
.A2(n_127),
.A3(n_39),
.B(n_42),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_147),
.B(n_38),
.Y(n_148)
);


endmodule