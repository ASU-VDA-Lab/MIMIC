module fake_ibex_1153_n_1702 (n_151, n_85, n_84, n_64, n_171, n_103, n_204, n_274, n_130, n_177, n_76, n_273, n_309, n_330, n_9, n_328, n_293, n_124, n_37, n_256, n_193, n_108, n_165, n_86, n_70, n_255, n_175, n_59, n_28, n_125, n_304, n_191, n_5, n_62, n_71, n_153, n_194, n_249, n_334, n_312, n_239, n_94, n_134, n_88, n_142, n_226, n_258, n_40, n_90, n_17, n_74, n_176, n_58, n_43, n_216, n_33, n_166, n_163, n_114, n_236, n_34, n_15, n_24, n_189, n_280, n_317, n_105, n_187, n_1, n_154, n_182, n_196, n_326, n_327, n_89, n_50, n_144, n_170, n_270, n_113, n_117, n_265, n_158, n_259, n_276, n_210, n_220, n_91, n_287, n_54, n_243, n_19, n_228, n_147, n_251, n_244, n_73, n_310, n_323, n_143, n_106, n_8, n_224, n_183, n_67, n_333, n_110, n_306, n_47, n_169, n_10, n_21, n_242, n_278, n_316, n_16, n_60, n_7, n_109, n_127, n_121, n_48, n_325, n_57, n_301, n_296, n_120, n_168, n_155, n_315, n_13, n_122, n_116, n_0, n_289, n_12, n_150, n_286, n_321, n_133, n_51, n_215, n_279, n_49, n_235, n_22, n_136, n_261, n_30, n_221, n_102, n_52, n_99, n_269, n_156, n_126, n_25, n_104, n_45, n_141, n_222, n_186, n_295, n_331, n_230, n_96, n_185, n_290, n_174, n_157, n_219, n_246, n_31, n_146, n_207, n_167, n_128, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_205, n_139, n_275, n_98, n_129, n_267, n_245, n_229, n_209, n_82, n_263, n_27, n_299, n_87, n_262, n_75, n_137, n_173, n_180, n_201, n_14, n_257, n_77, n_44, n_66, n_305, n_307, n_192, n_140, n_4, n_6, n_100, n_179, n_206, n_329, n_26, n_188, n_200, n_199, n_308, n_135, n_283, n_111, n_36, n_18, n_322, n_53, n_227, n_115, n_11, n_248, n_92, n_101, n_190, n_138, n_214, n_238, n_332, n_211, n_218, n_314, n_132, n_277, n_225, n_272, n_23, n_223, n_95, n_285, n_288, n_247, n_320, n_55, n_291, n_318, n_63, n_161, n_237, n_29, n_203, n_268, n_148, n_2, n_233, n_118, n_164, n_38, n_198, n_264, n_217, n_324, n_78, n_20, n_69, n_39, n_178, n_303, n_93, n_162, n_240, n_282, n_61, n_266, n_42, n_294, n_112, n_46, n_284, n_80, n_172, n_250, n_313, n_119, n_72, n_319, n_195, n_212, n_311, n_97, n_197, n_181, n_131, n_123, n_260, n_302, n_297, n_41, n_252, n_83, n_32, n_107, n_149, n_254, n_213, n_271, n_241, n_68, n_292, n_79, n_81, n_35, n_159, n_202, n_231, n_298, n_160, n_184, n_56, n_232, n_281, n_1702);

input n_151;
input n_85;
input n_84;
input n_64;
input n_171;
input n_103;
input n_204;
input n_274;
input n_130;
input n_177;
input n_76;
input n_273;
input n_309;
input n_330;
input n_9;
input n_328;
input n_293;
input n_124;
input n_37;
input n_256;
input n_193;
input n_108;
input n_165;
input n_86;
input n_70;
input n_255;
input n_175;
input n_59;
input n_28;
input n_125;
input n_304;
input n_191;
input n_5;
input n_62;
input n_71;
input n_153;
input n_194;
input n_249;
input n_334;
input n_312;
input n_239;
input n_94;
input n_134;
input n_88;
input n_142;
input n_226;
input n_258;
input n_40;
input n_90;
input n_17;
input n_74;
input n_176;
input n_58;
input n_43;
input n_216;
input n_33;
input n_166;
input n_163;
input n_114;
input n_236;
input n_34;
input n_15;
input n_24;
input n_189;
input n_280;
input n_317;
input n_105;
input n_187;
input n_1;
input n_154;
input n_182;
input n_196;
input n_326;
input n_327;
input n_89;
input n_50;
input n_144;
input n_170;
input n_270;
input n_113;
input n_117;
input n_265;
input n_158;
input n_259;
input n_276;
input n_210;
input n_220;
input n_91;
input n_287;
input n_54;
input n_243;
input n_19;
input n_228;
input n_147;
input n_251;
input n_244;
input n_73;
input n_310;
input n_323;
input n_143;
input n_106;
input n_8;
input n_224;
input n_183;
input n_67;
input n_333;
input n_110;
input n_306;
input n_47;
input n_169;
input n_10;
input n_21;
input n_242;
input n_278;
input n_316;
input n_16;
input n_60;
input n_7;
input n_109;
input n_127;
input n_121;
input n_48;
input n_325;
input n_57;
input n_301;
input n_296;
input n_120;
input n_168;
input n_155;
input n_315;
input n_13;
input n_122;
input n_116;
input n_0;
input n_289;
input n_12;
input n_150;
input n_286;
input n_321;
input n_133;
input n_51;
input n_215;
input n_279;
input n_49;
input n_235;
input n_22;
input n_136;
input n_261;
input n_30;
input n_221;
input n_102;
input n_52;
input n_99;
input n_269;
input n_156;
input n_126;
input n_25;
input n_104;
input n_45;
input n_141;
input n_222;
input n_186;
input n_295;
input n_331;
input n_230;
input n_96;
input n_185;
input n_290;
input n_174;
input n_157;
input n_219;
input n_246;
input n_31;
input n_146;
input n_207;
input n_167;
input n_128;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_205;
input n_139;
input n_275;
input n_98;
input n_129;
input n_267;
input n_245;
input n_229;
input n_209;
input n_82;
input n_263;
input n_27;
input n_299;
input n_87;
input n_262;
input n_75;
input n_137;
input n_173;
input n_180;
input n_201;
input n_14;
input n_257;
input n_77;
input n_44;
input n_66;
input n_305;
input n_307;
input n_192;
input n_140;
input n_4;
input n_6;
input n_100;
input n_179;
input n_206;
input n_329;
input n_26;
input n_188;
input n_200;
input n_199;
input n_308;
input n_135;
input n_283;
input n_111;
input n_36;
input n_18;
input n_322;
input n_53;
input n_227;
input n_115;
input n_11;
input n_248;
input n_92;
input n_101;
input n_190;
input n_138;
input n_214;
input n_238;
input n_332;
input n_211;
input n_218;
input n_314;
input n_132;
input n_277;
input n_225;
input n_272;
input n_23;
input n_223;
input n_95;
input n_285;
input n_288;
input n_247;
input n_320;
input n_55;
input n_291;
input n_318;
input n_63;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_148;
input n_2;
input n_233;
input n_118;
input n_164;
input n_38;
input n_198;
input n_264;
input n_217;
input n_324;
input n_78;
input n_20;
input n_69;
input n_39;
input n_178;
input n_303;
input n_93;
input n_162;
input n_240;
input n_282;
input n_61;
input n_266;
input n_42;
input n_294;
input n_112;
input n_46;
input n_284;
input n_80;
input n_172;
input n_250;
input n_313;
input n_119;
input n_72;
input n_319;
input n_195;
input n_212;
input n_311;
input n_97;
input n_197;
input n_181;
input n_131;
input n_123;
input n_260;
input n_302;
input n_297;
input n_41;
input n_252;
input n_83;
input n_32;
input n_107;
input n_149;
input n_254;
input n_213;
input n_271;
input n_241;
input n_68;
input n_292;
input n_79;
input n_81;
input n_35;
input n_159;
input n_202;
input n_231;
input n_298;
input n_160;
input n_184;
input n_56;
input n_232;
input n_281;

output n_1702;

wire n_1084;
wire n_1474;
wire n_1295;
wire n_507;
wire n_992;
wire n_1582;
wire n_766;
wire n_1110;
wire n_1382;
wire n_1596;
wire n_926;
wire n_1079;
wire n_1100;
wire n_845;
wire n_446;
wire n_452;
wire n_1234;
wire n_1594;
wire n_773;
wire n_1469;
wire n_821;
wire n_873;
wire n_1227;
wire n_962;
wire n_1080;
wire n_862;
wire n_909;
wire n_957;
wire n_1652;
wire n_678;
wire n_969;
wire n_1125;
wire n_733;
wire n_622;
wire n_1226;
wire n_1034;
wire n_872;
wire n_1619;
wire n_457;
wire n_1666;
wire n_494;
wire n_930;
wire n_1044;
wire n_1492;
wire n_1134;
wire n_1478;
wire n_1684;
wire n_1614;
wire n_911;
wire n_652;
wire n_781;
wire n_475;
wire n_802;
wire n_1233;
wire n_1045;
wire n_500;
wire n_963;
wire n_376;
wire n_531;
wire n_1308;
wire n_556;
wire n_1138;
wire n_498;
wire n_708;
wire n_1096;
wire n_375;
wire n_1391;
wire n_667;
wire n_884;
wire n_850;
wire n_879;
wire n_723;
wire n_1144;
wire n_346;
wire n_1392;
wire n_1268;
wire n_739;
wire n_853;
wire n_504;
wire n_948;
wire n_1338;
wire n_875;
wire n_1307;
wire n_1327;
wire n_481;
wire n_876;
wire n_497;
wire n_711;
wire n_671;
wire n_989;
wire n_1668;
wire n_1641;
wire n_829;
wire n_825;
wire n_1480;
wire n_1463;
wire n_1681;
wire n_939;
wire n_1636;
wire n_1687;
wire n_655;
wire n_550;
wire n_557;
wire n_641;
wire n_527;
wire n_893;
wire n_1654;
wire n_496;
wire n_434;
wire n_1258;
wire n_1344;
wire n_1680;
wire n_835;
wire n_1195;
wire n_824;
wire n_441;
wire n_694;
wire n_523;
wire n_787;
wire n_614;
wire n_431;
wire n_1130;
wire n_1228;
wire n_1081;
wire n_374;
wire n_538;
wire n_1155;
wire n_1292;
wire n_459;
wire n_1576;
wire n_1664;
wire n_518;
wire n_852;
wire n_1427;
wire n_1133;
wire n_904;
wire n_355;
wire n_646;
wire n_448;
wire n_466;
wire n_1030;
wire n_1698;
wire n_1094;
wire n_1496;
wire n_715;
wire n_530;
wire n_1663;
wire n_1214;
wire n_1274;
wire n_420;
wire n_1606;
wire n_769;
wire n_1595;
wire n_1509;
wire n_1618;
wire n_1648;
wire n_857;
wire n_765;
wire n_1070;
wire n_777;
wire n_917;
wire n_968;
wire n_1253;
wire n_1306;
wire n_1484;
wire n_1493;
wire n_1313;
wire n_352;
wire n_558;
wire n_666;
wire n_1638;
wire n_1071;
wire n_1449;
wire n_793;
wire n_937;
wire n_1645;
wire n_973;
wire n_1038;
wire n_618;
wire n_1269;
wire n_662;
wire n_979;
wire n_1309;
wire n_1316;
wire n_1562;
wire n_1215;
wire n_629;
wire n_1445;
wire n_573;
wire n_359;
wire n_1466;
wire n_1412;
wire n_433;
wire n_439;
wire n_1672;
wire n_1007;
wire n_643;
wire n_1276;
wire n_1637;
wire n_841;
wire n_772;
wire n_810;
wire n_338;
wire n_1401;
wire n_369;
wire n_1588;
wire n_1301;
wire n_869;
wire n_1620;
wire n_1561;
wire n_718;
wire n_554;
wire n_553;
wire n_1078;
wire n_1219;
wire n_713;
wire n_1252;
wire n_1170;
wire n_605;
wire n_539;
wire n_630;
wire n_567;
wire n_745;
wire n_447;
wire n_564;
wire n_562;
wire n_1322;
wire n_1305;
wire n_795;
wire n_592;
wire n_1248;
wire n_762;
wire n_1388;
wire n_800;
wire n_706;
wire n_784;
wire n_684;
wire n_1653;
wire n_1375;
wire n_397;
wire n_1356;
wire n_894;
wire n_1118;
wire n_692;
wire n_709;
wire n_1296;
wire n_499;
wire n_702;
wire n_1326;
wire n_971;
wire n_451;
wire n_1350;
wire n_906;
wire n_1093;
wire n_978;
wire n_579;
wire n_899;
wire n_1019;
wire n_902;
wire n_1689;
wire n_1250;
wire n_1190;
wire n_1304;
wire n_744;
wire n_563;
wire n_1506;
wire n_881;
wire n_734;
wire n_1558;
wire n_1650;
wire n_1520;
wire n_1073;
wire n_1453;
wire n_1108;
wire n_382;
wire n_1423;
wire n_1239;
wire n_1370;
wire n_1209;
wire n_379;
wire n_551;
wire n_1616;
wire n_729;
wire n_1569;
wire n_1434;
wire n_603;
wire n_1649;
wire n_422;
wire n_1609;
wire n_391;
wire n_1613;
wire n_820;
wire n_805;
wire n_670;
wire n_1132;
wire n_892;
wire n_390;
wire n_1467;
wire n_544;
wire n_1281;
wire n_1447;
wire n_695;
wire n_1549;
wire n_639;
wire n_1531;
wire n_1332;
wire n_482;
wire n_1424;
wire n_870;
wire n_1610;
wire n_1298;
wire n_1387;
wire n_609;
wire n_1040;
wire n_476;
wire n_1159;
wire n_1368;
wire n_1154;
wire n_345;
wire n_455;
wire n_1701;
wire n_1243;
wire n_1121;
wire n_693;
wire n_406;
wire n_606;
wire n_737;
wire n_1571;
wire n_462;
wire n_1407;
wire n_1235;
wire n_1003;
wire n_889;
wire n_435;
wire n_396;
wire n_816;
wire n_1058;
wire n_399;
wire n_1543;
wire n_823;
wire n_1504;
wire n_1519;
wire n_1425;
wire n_1441;
wire n_657;
wire n_1156;
wire n_1293;
wire n_1360;
wire n_749;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_819;
wire n_822;
wire n_1042;
wire n_743;
wire n_754;
wire n_395;
wire n_1319;
wire n_389;
wire n_1553;
wire n_1041;
wire n_1090;
wire n_1196;
wire n_1182;
wire n_1271;
wire n_1031;
wire n_372;
wire n_981;
wire n_350;
wire n_398;
wire n_1591;
wire n_583;
wire n_1671;
wire n_1409;
wire n_1015;
wire n_663;
wire n_1377;
wire n_1583;
wire n_1521;
wire n_1152;
wire n_371;
wire n_1036;
wire n_974;
wire n_608;
wire n_864;
wire n_412;
wire n_959;
wire n_1106;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_449;
wire n_1634;
wire n_1552;
wire n_1452;
wire n_1318;
wire n_1508;
wire n_421;
wire n_738;
wire n_1217;
wire n_1189;
wire n_761;
wire n_748;
wire n_901;
wire n_1577;
wire n_340;
wire n_1255;
wire n_1700;
wire n_1218;
wire n_1181;
wire n_1140;
wire n_1056;
wire n_1283;
wire n_1446;
wire n_1487;
wire n_840;
wire n_1203;
wire n_1421;
wire n_561;
wire n_471;
wire n_846;
wire n_1237;
wire n_859;
wire n_965;
wire n_1109;
wire n_1633;
wire n_384;
wire n_1051;
wire n_1008;
wire n_458;
wire n_1498;
wire n_1053;
wire n_1656;
wire n_1207;
wire n_1076;
wire n_1032;
wire n_936;
wire n_469;
wire n_1589;
wire n_1210;
wire n_591;
wire n_1510;
wire n_1201;
wire n_1246;
wire n_1677;
wire n_732;
wire n_1236;
wire n_832;
wire n_590;
wire n_1568;
wire n_1184;
wire n_1477;
wire n_1364;
wire n_1540;
wire n_1676;
wire n_1013;
wire n_929;
wire n_637;
wire n_1136;
wire n_1075;
wire n_1249;
wire n_574;
wire n_515;
wire n_1229;
wire n_1440;
wire n_1490;
wire n_907;
wire n_1179;
wire n_1153;
wire n_669;
wire n_521;
wire n_1117;
wire n_1273;
wire n_1083;
wire n_1014;
wire n_724;
wire n_437;
wire n_938;
wire n_1178;
wire n_474;
wire n_878;
wire n_594;
wire n_1464;
wire n_1566;
wire n_944;
wire n_623;
wire n_585;
wire n_1334;
wire n_483;
wire n_1695;
wire n_1418;
wire n_1137;
wire n_660;
wire n_524;
wire n_1200;
wire n_1120;
wire n_576;
wire n_1602;
wire n_388;
wire n_1522;
wire n_1279;
wire n_931;
wire n_607;
wire n_827;
wire n_1064;
wire n_1408;
wire n_1028;
wire n_1264;
wire n_1146;
wire n_358;
wire n_488;
wire n_705;
wire n_1548;
wire n_429;
wire n_1682;
wire n_1608;
wire n_1009;
wire n_1260;
wire n_589;
wire n_472;
wire n_347;
wire n_847;
wire n_1436;
wire n_413;
wire n_1069;
wire n_1485;
wire n_1465;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_1232;
wire n_679;
wire n_1345;
wire n_696;
wire n_837;
wire n_1590;
wire n_640;
wire n_954;
wire n_363;
wire n_1628;
wire n_725;
wire n_596;
wire n_1545;
wire n_351;
wire n_456;
wire n_1471;
wire n_998;
wire n_1115;
wire n_1395;
wire n_801;
wire n_1479;
wire n_1046;
wire n_882;
wire n_942;
wire n_1627;
wire n_1431;
wire n_651;
wire n_721;
wire n_365;
wire n_814;
wire n_943;
wire n_1086;
wire n_1523;
wire n_1470;
wire n_444;
wire n_1593;
wire n_986;
wire n_495;
wire n_1420;
wire n_1699;
wire n_411;
wire n_927;
wire n_1563;
wire n_615;
wire n_803;
wire n_1615;
wire n_1087;
wire n_757;
wire n_1400;
wire n_712;
wire n_1539;
wire n_1599;
wire n_650;
wire n_409;
wire n_1575;
wire n_1448;
wire n_517;
wire n_817;
wire n_555;
wire n_337;
wire n_951;
wire n_468;
wire n_1580;
wire n_1574;
wire n_780;
wire n_502;
wire n_633;
wire n_726;
wire n_532;
wire n_1439;
wire n_863;
wire n_597;
wire n_1128;
wire n_1266;
wire n_1300;
wire n_807;
wire n_741;
wire n_430;
wire n_486;
wire n_1405;
wire n_997;
wire n_1428;
wire n_891;
wire n_1528;
wire n_1495;
wire n_717;
wire n_1357;
wire n_1512;
wire n_668;
wire n_871;
wire n_1339;
wire n_1544;
wire n_1426;
wire n_485;
wire n_1315;
wire n_1413;
wire n_811;
wire n_808;
wire n_945;
wire n_460;
wire n_1560;
wire n_1592;
wire n_1461;
wire n_461;
wire n_903;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_1378;
wire n_1048;
wire n_774;
wire n_588;
wire n_1430;
wire n_1251;
wire n_1247;
wire n_528;
wire n_836;
wire n_1475;
wire n_1263;
wire n_443;
wire n_1185;
wire n_1683;
wire n_344;
wire n_436;
wire n_1122;
wire n_628;
wire n_890;
wire n_874;
wire n_1505;
wire n_1163;
wire n_677;
wire n_1514;
wire n_964;
wire n_916;
wire n_503;
wire n_895;
wire n_687;
wire n_1035;
wire n_1535;
wire n_751;
wire n_1127;
wire n_932;
wire n_380;
wire n_947;
wire n_1004;
wire n_831;
wire n_778;
wire n_1254;
wire n_1148;
wire n_540;
wire n_1667;
wire n_1104;
wire n_1011;
wire n_1437;
wire n_529;
wire n_626;
wire n_1679;
wire n_1497;
wire n_1578;
wire n_1143;
wire n_418;
wire n_510;
wire n_972;
wire n_601;
wire n_610;
wire n_1444;
wire n_920;
wire n_664;
wire n_1067;
wire n_994;
wire n_545;
wire n_887;
wire n_1162;
wire n_634;
wire n_991;
wire n_961;
wire n_1223;
wire n_1349;
wire n_1331;
wire n_1323;
wire n_578;
wire n_432;
wire n_403;
wire n_1353;
wire n_423;
wire n_357;
wire n_1429;
wire n_1546;
wire n_1432;
wire n_1320;
wire n_996;
wire n_915;
wire n_1174;
wire n_1286;
wire n_1657;
wire n_542;
wire n_1294;
wire n_1601;
wire n_900;
wire n_1351;
wire n_377;
wire n_647;
wire n_1380;
wire n_1367;
wire n_1291;
wire n_1458;
wire n_1694;
wire n_1460;
wire n_1629;
wire n_1662;
wire n_1340;
wire n_339;
wire n_348;
wire n_1626;
wire n_674;
wire n_1660;
wire n_1643;
wire n_1670;
wire n_552;
wire n_1112;
wire n_1267;
wire n_1384;
wire n_1376;
wire n_1537;
wire n_1612;
wire n_703;
wire n_426;
wire n_1172;
wire n_1099;
wire n_598;
wire n_1422;
wire n_508;
wire n_453;
wire n_1527;
wire n_400;
wire n_1055;
wire n_1524;
wire n_673;
wire n_798;
wire n_404;
wire n_1177;
wire n_1025;
wire n_1517;
wire n_690;
wire n_1225;
wire n_982;
wire n_1624;
wire n_785;
wire n_604;
wire n_1598;
wire n_977;
wire n_719;
wire n_370;
wire n_1491;
wire n_716;
wire n_923;
wire n_642;
wire n_1607;
wire n_1625;
wire n_933;
wire n_1037;
wire n_464;
wire n_1348;
wire n_838;
wire n_1289;
wire n_1021;
wire n_746;
wire n_1557;
wire n_1188;
wire n_1567;
wire n_742;
wire n_1191;
wire n_1503;
wire n_1052;
wire n_789;
wire n_656;
wire n_602;
wire n_842;
wire n_767;
wire n_1617;
wire n_1587;
wire n_636;
wire n_1259;
wire n_490;
wire n_407;
wire n_595;
wire n_1001;
wire n_570;
wire n_1396;
wire n_1224;
wire n_356;
wire n_1538;
wire n_487;
wire n_349;
wire n_454;
wire n_1017;
wire n_730;
wire n_1456;
wire n_625;
wire n_619;
wire n_1124;
wire n_611;
wire n_1690;
wire n_1673;
wire n_922;
wire n_851;
wire n_993;
wire n_1135;
wire n_541;
wire n_613;
wire n_659;
wire n_1494;
wire n_1550;
wire n_1066;
wire n_1169;
wire n_648;
wire n_571;
wire n_830;
wire n_473;
wire n_1241;
wire n_445;
wire n_1072;
wire n_1231;
wire n_1173;
wire n_1208;
wire n_353;
wire n_1604;
wire n_1639;
wire n_826;
wire n_1337;
wire n_1647;
wire n_768;
wire n_839;
wire n_1278;
wire n_796;
wire n_797;
wire n_1006;
wire n_402;
wire n_1238;
wire n_1415;
wire n_976;
wire n_1063;
wire n_1270;
wire n_834;
wire n_1476;
wire n_935;
wire n_1603;
wire n_925;
wire n_1054;
wire n_722;
wire n_1644;
wire n_1406;
wire n_1489;
wire n_804;
wire n_484;
wire n_1455;
wire n_1642;
wire n_480;
wire n_354;
wire n_1057;
wire n_1473;
wire n_516;
wire n_1403;
wire n_1149;
wire n_1176;
wire n_1502;
wire n_1605;
wire n_506;
wire n_868;
wire n_1202;
wire n_1065;
wire n_1457;
wire n_905;
wire n_975;
wire n_675;
wire n_624;
wire n_463;
wire n_520;
wire n_934;
wire n_775;
wire n_512;
wire n_950;
wire n_685;
wire n_1222;
wire n_1630;
wire n_1198;
wire n_1311;
wire n_1261;
wire n_776;
wire n_1114;
wire n_818;
wire n_1167;
wire n_1282;
wire n_1321;
wire n_700;
wire n_360;
wire n_1107;
wire n_1573;
wire n_525;
wire n_815;
wire n_919;
wire n_535;
wire n_681;
wire n_415;
wire n_1411;
wire n_1139;
wire n_1018;
wire n_858;
wire n_385;
wire n_1324;
wire n_1669;
wire n_1501;
wire n_782;
wire n_616;
wire n_833;
wire n_1343;
wire n_1371;
wire n_1513;
wire n_728;
wire n_786;
wire n_362;
wire n_505;
wire n_1621;
wire n_1342;
wire n_501;
wire n_752;
wire n_958;
wire n_1175;
wire n_1416;
wire n_1659;
wire n_1221;
wire n_1047;
wire n_1515;
wire n_1374;
wire n_1435;
wire n_1688;
wire n_792;
wire n_1314;
wire n_1433;
wire n_575;
wire n_1242;
wire n_1119;
wire n_1085;
wire n_419;
wire n_885;
wire n_1530;
wire n_513;
wire n_877;
wire n_1088;
wire n_896;
wire n_1451;
wire n_1005;
wire n_1102;
wire n_631;
wire n_794;
wire n_1288;
wire n_1275;
wire n_985;
wire n_1165;
wire n_897;
wire n_1622;
wire n_393;
wire n_428;
wire n_697;
wire n_1105;
wire n_1459;
wire n_912;
wire n_1570;
wire n_424;
wire n_701;
wire n_995;
wire n_1000;
wire n_1256;
wire n_587;
wire n_1303;
wire n_1526;
wire n_764;
wire n_1507;
wire n_1206;
wire n_855;
wire n_812;
wire n_1050;
wire n_599;
wire n_1060;
wire n_1372;
wire n_756;
wire n_1565;
wire n_1257;
wire n_387;
wire n_1632;
wire n_688;
wire n_1542;
wire n_946;
wire n_1547;
wire n_707;
wire n_1362;
wire n_1586;
wire n_1097;
wire n_341;
wire n_621;
wire n_956;
wire n_790;
wire n_1541;
wire n_586;
wire n_1330;
wire n_638;
wire n_1697;
wire n_593;
wire n_1212;
wire n_1199;
wire n_1443;
wire n_478;
wire n_1585;
wire n_1564;
wire n_1631;
wire n_336;
wire n_1623;
wire n_861;
wire n_1389;
wire n_1131;
wire n_547;
wire n_727;
wire n_1077;
wire n_1554;
wire n_1481;
wire n_1584;
wire n_828;
wire n_1438;
wire n_753;
wire n_645;
wire n_747;
wire n_1147;
wire n_1363;
wire n_1691;
wire n_1098;
wire n_584;
wire n_1366;
wire n_1518;
wire n_1187;
wire n_1361;
wire n_1693;
wire n_698;
wire n_1061;
wire n_682;
wire n_1373;
wire n_1686;
wire n_1302;
wire n_383;
wire n_886;
wire n_1010;
wire n_883;
wire n_417;
wire n_755;
wire n_1029;
wire n_470;
wire n_770;
wire n_1572;
wire n_1635;
wire n_941;
wire n_1245;
wire n_1317;
wire n_632;
wire n_1329;
wire n_373;
wire n_854;
wire n_343;
wire n_714;
wire n_1297;
wire n_1369;
wire n_740;
wire n_386;
wire n_549;
wire n_533;
wire n_898;
wire n_928;
wire n_1285;
wire n_967;
wire n_736;
wire n_1529;
wire n_1381;
wire n_1597;
wire n_1103;
wire n_1161;
wire n_465;
wire n_1486;
wire n_1068;
wire n_617;
wire n_914;
wire n_526;
wire n_1024;
wire n_1141;
wire n_1197;
wire n_1168;
wire n_865;
wire n_569;
wire n_600;
wire n_1556;
wire n_1192;
wire n_1646;
wire n_1290;
wire n_987;
wire n_750;
wire n_1299;
wire n_665;
wire n_1101;
wire n_367;
wire n_880;
wire n_654;
wire n_731;
wire n_1336;
wire n_758;
wire n_1166;
wire n_720;
wire n_710;
wire n_1390;
wire n_1023;
wire n_568;
wire n_1358;
wire n_813;
wire n_1211;
wire n_1397;
wire n_1284;
wire n_1359;
wire n_1116;
wire n_791;
wire n_1532;
wire n_1419;
wire n_543;
wire n_580;
wire n_1685;
wire n_1082;
wire n_1213;
wire n_1193;
wire n_980;
wire n_849;
wire n_1488;
wire n_1074;
wire n_759;
wire n_1379;
wire n_953;
wire n_1180;
wire n_1462;
wire n_536;
wire n_1220;
wire n_467;
wire n_1398;
wire n_427;
wire n_1262;
wire n_442;
wire n_1692;
wire n_438;
wire n_1012;
wire n_689;
wire n_960;
wire n_1022;
wire n_676;
wire n_1240;
wire n_1183;
wire n_1204;
wire n_1151;
wire n_771;
wire n_999;
wire n_514;
wire n_1092;
wire n_560;
wire n_1658;
wire n_1386;
wire n_910;
wire n_635;
wire n_844;
wire n_1020;
wire n_783;
wire n_1142;
wire n_1385;
wire n_1062;
wire n_1230;
wire n_1027;
wire n_1516;
wire n_335;
wire n_1499;
wire n_1500;
wire n_966;
wire n_949;
wire n_704;
wire n_924;
wire n_1600;
wire n_477;
wire n_1661;
wire n_699;
wire n_368;
wire n_918;
wire n_672;
wire n_1039;
wire n_401;
wire n_1043;
wire n_1402;
wire n_735;
wire n_1450;
wire n_566;
wire n_416;
wire n_581;
wire n_1365;
wire n_1472;
wire n_1089;
wire n_392;
wire n_1536;
wire n_1049;
wire n_548;
wire n_1158;
wire n_763;
wire n_940;
wire n_1404;
wire n_546;
wire n_788;
wire n_410;
wire n_1160;
wire n_1442;
wire n_658;
wire n_1216;
wire n_1026;
wire n_366;
wire n_1454;
wire n_1033;
wire n_627;
wire n_990;
wire n_1383;
wire n_888;
wire n_1325;
wire n_582;
wire n_1483;
wire n_653;
wire n_1205;
wire n_843;
wire n_1059;
wire n_799;
wire n_691;
wire n_1581;
wire n_522;
wire n_479;
wire n_534;
wire n_511;
wire n_381;
wire n_1414;
wire n_1002;
wire n_1111;
wire n_1341;
wire n_405;
wire n_1310;
wire n_612;
wire n_1611;
wire n_955;
wire n_440;
wire n_1333;
wire n_342;
wire n_414;
wire n_378;
wire n_952;
wire n_1675;
wire n_1640;
wire n_1551;
wire n_1145;
wire n_1533;
wire n_1511;
wire n_537;
wire n_1113;
wire n_1651;
wire n_1468;
wire n_913;
wire n_509;
wire n_1164;
wire n_1354;
wire n_1277;
wire n_1696;
wire n_1016;
wire n_680;
wire n_1355;
wire n_809;
wire n_856;
wire n_779;
wire n_1559;
wire n_1579;
wire n_1280;
wire n_493;
wire n_1335;
wire n_519;
wire n_408;
wire n_361;
wire n_1665;
wire n_1091;
wire n_1678;
wire n_1287;
wire n_1482;
wire n_860;
wire n_1525;
wire n_661;
wire n_848;
wire n_683;
wire n_1150;
wire n_1194;
wire n_620;
wire n_1399;
wire n_450;
wire n_1674;
wire n_686;
wire n_572;
wire n_867;
wire n_983;
wire n_1417;
wire n_644;
wire n_577;
wire n_970;
wire n_491;
wire n_921;
wire n_489;
wire n_1534;
wire n_908;
wire n_1346;
wire n_565;
wire n_1123;
wire n_1272;
wire n_1393;
wire n_984;
wire n_1655;
wire n_394;
wire n_364;
wire n_1410;
wire n_988;
wire n_760;
wire n_1157;
wire n_806;
wire n_1186;
wire n_492;
wire n_649;
wire n_866;
wire n_559;
wire n_425;

INVx1_ASAP7_75t_L g335 ( 
.A(n_160),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_271),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_23),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_38),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_27),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_266),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_264),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_315),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_171),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_60),
.Y(n_344)
);

INVxp33_ASAP7_75t_L g345 ( 
.A(n_240),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_41),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_88),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_277),
.Y(n_348)
);

BUFx5_ASAP7_75t_L g349 ( 
.A(n_108),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_269),
.Y(n_350)
);

BUFx3_ASAP7_75t_L g351 ( 
.A(n_122),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_267),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_0),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_109),
.Y(n_354)
);

CKINVDCx14_ASAP7_75t_R g355 ( 
.A(n_255),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_163),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_234),
.Y(n_357)
);

BUFx3_ASAP7_75t_L g358 ( 
.A(n_60),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_310),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_161),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_130),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_254),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_290),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_166),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_176),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_21),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_208),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_211),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_295),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_101),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_307),
.Y(n_371)
);

BUFx6f_ASAP7_75t_L g372 ( 
.A(n_91),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_324),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_282),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_279),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_331),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_236),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_209),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_218),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_257),
.Y(n_380)
);

INVx2_ASAP7_75t_SL g381 ( 
.A(n_256),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_14),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_298),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_9),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_164),
.Y(n_385)
);

BUFx6f_ASAP7_75t_L g386 ( 
.A(n_15),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_233),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_205),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_241),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_247),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_73),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_232),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_273),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_242),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_5),
.Y(n_395)
);

INVx3_ASAP7_75t_L g396 ( 
.A(n_28),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_250),
.Y(n_397)
);

BUFx3_ASAP7_75t_L g398 ( 
.A(n_292),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_284),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_25),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_325),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_143),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_301),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_303),
.Y(n_404)
);

BUFx3_ASAP7_75t_L g405 ( 
.A(n_3),
.Y(n_405)
);

CKINVDCx16_ASAP7_75t_R g406 ( 
.A(n_170),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_308),
.Y(n_407)
);

BUFx6f_ASAP7_75t_L g408 ( 
.A(n_332),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_116),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_149),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_229),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_305),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_300),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_206),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_165),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_286),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_249),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_92),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_316),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_227),
.Y(n_420)
);

CKINVDCx16_ASAP7_75t_R g421 ( 
.A(n_145),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_13),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_132),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_244),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_34),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_8),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_304),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_302),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_181),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_291),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_93),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_322),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_86),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_180),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_294),
.Y(n_435)
);

INVxp67_ASAP7_75t_SL g436 ( 
.A(n_280),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_75),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_299),
.Y(n_438)
);

BUFx10_ASAP7_75t_L g439 ( 
.A(n_263),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_196),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_319),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_237),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_28),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_317),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_107),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_245),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_157),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_309),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_228),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_326),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_285),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_110),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_201),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_221),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_72),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_261),
.Y(n_456)
);

INVx1_ASAP7_75t_SL g457 ( 
.A(n_248),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_260),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_85),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_183),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_207),
.Y(n_461)
);

BUFx10_ASAP7_75t_L g462 ( 
.A(n_223),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_329),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_235),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_148),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g466 ( 
.A(n_7),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_142),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_84),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_117),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_313),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_199),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_281),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g473 ( 
.A(n_278),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_53),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_26),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_193),
.Y(n_476)
);

BUFx6f_ASAP7_75t_L g477 ( 
.A(n_76),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_274),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_39),
.Y(n_479)
);

BUFx8_ASAP7_75t_SL g480 ( 
.A(n_96),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_34),
.Y(n_481)
);

CKINVDCx20_ASAP7_75t_R g482 ( 
.A(n_314),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_184),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_321),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_231),
.Y(n_485)
);

CKINVDCx20_ASAP7_75t_R g486 ( 
.A(n_272),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_112),
.Y(n_487)
);

CKINVDCx14_ASAP7_75t_R g488 ( 
.A(n_51),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_262),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_75),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_220),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_126),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_150),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_212),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_252),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_57),
.Y(n_496)
);

BUFx5_ASAP7_75t_L g497 ( 
.A(n_198),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_251),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_118),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_330),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_253),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_318),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_98),
.Y(n_503)
);

CKINVDCx20_ASAP7_75t_R g504 ( 
.A(n_162),
.Y(n_504)
);

CKINVDCx20_ASAP7_75t_R g505 ( 
.A(n_224),
.Y(n_505)
);

BUFx10_ASAP7_75t_L g506 ( 
.A(n_238),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_225),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_293),
.Y(n_508)
);

INVx2_ASAP7_75t_SL g509 ( 
.A(n_296),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_195),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_258),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_57),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_134),
.Y(n_513)
);

BUFx3_ASAP7_75t_L g514 ( 
.A(n_312),
.Y(n_514)
);

CKINVDCx20_ASAP7_75t_R g515 ( 
.A(n_20),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_66),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_289),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_239),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_48),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_287),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_140),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_89),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_10),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_74),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_230),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_327),
.Y(n_526)
);

BUFx10_ASAP7_75t_L g527 ( 
.A(n_276),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_297),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_169),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_23),
.Y(n_530)
);

CKINVDCx20_ASAP7_75t_R g531 ( 
.A(n_270),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_288),
.Y(n_532)
);

BUFx3_ASAP7_75t_L g533 ( 
.A(n_10),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_101),
.Y(n_534)
);

BUFx10_ASAP7_75t_L g535 ( 
.A(n_203),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_78),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_323),
.Y(n_537)
);

BUFx3_ASAP7_75t_L g538 ( 
.A(n_333),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_89),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_306),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_190),
.Y(n_541)
);

HB1xp67_ASAP7_75t_L g542 ( 
.A(n_177),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_216),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_80),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_202),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_49),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_22),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_226),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_265),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_129),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_328),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_33),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_66),
.Y(n_553)
);

CKINVDCx20_ASAP7_75t_R g554 ( 
.A(n_311),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_147),
.Y(n_555)
);

BUFx3_ASAP7_75t_L g556 ( 
.A(n_144),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_8),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_204),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_275),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_36),
.Y(n_560)
);

BUFx10_ASAP7_75t_L g561 ( 
.A(n_13),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_243),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_86),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_77),
.Y(n_564)
);

INVx1_ASAP7_75t_SL g565 ( 
.A(n_2),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_268),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_259),
.Y(n_567)
);

INVx1_ASAP7_75t_SL g568 ( 
.A(n_85),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_81),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_246),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_79),
.Y(n_571)
);

CKINVDCx20_ASAP7_75t_R g572 ( 
.A(n_320),
.Y(n_572)
);

CKINVDCx20_ASAP7_75t_R g573 ( 
.A(n_194),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_215),
.Y(n_574)
);

HB1xp67_ASAP7_75t_L g575 ( 
.A(n_64),
.Y(n_575)
);

INVx2_ASAP7_75t_SL g576 ( 
.A(n_17),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_283),
.Y(n_577)
);

INVx1_ASAP7_75t_SL g578 ( 
.A(n_334),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_3),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_15),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_192),
.Y(n_581)
);

INVx3_ASAP7_75t_L g582 ( 
.A(n_79),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_61),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_189),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_178),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_36),
.Y(n_586)
);

CKINVDCx14_ASAP7_75t_R g587 ( 
.A(n_52),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_38),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_396),
.Y(n_589)
);

CKINVDCx20_ASAP7_75t_R g590 ( 
.A(n_587),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_336),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_396),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_575),
.B(n_0),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_401),
.Y(n_594)
);

NOR2xp67_ASAP7_75t_L g595 ( 
.A(n_582),
.B(n_1),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_410),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_413),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_582),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_542),
.Y(n_599)
);

CKINVDCx20_ASAP7_75t_R g600 ( 
.A(n_587),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_358),
.Y(n_601)
);

CKINVDCx20_ASAP7_75t_R g602 ( 
.A(n_488),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_453),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_358),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_405),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_405),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_533),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_533),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_473),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_479),
.Y(n_610)
);

CKINVDCx20_ASAP7_75t_R g611 ( 
.A(n_338),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_479),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_482),
.Y(n_613)
);

NOR2xp67_ASAP7_75t_L g614 ( 
.A(n_576),
.B(n_1),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_536),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_486),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_536),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_579),
.Y(n_618)
);

AND2x2_ASAP7_75t_L g619 ( 
.A(n_345),
.B(n_2),
.Y(n_619)
);

CKINVDCx20_ASAP7_75t_R g620 ( 
.A(n_344),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_L g621 ( 
.A(n_381),
.B(n_4),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_504),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_579),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_339),
.Y(n_624)
);

CKINVDCx20_ASAP7_75t_R g625 ( 
.A(n_347),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_505),
.Y(n_626)
);

CKINVDCx20_ASAP7_75t_R g627 ( 
.A(n_370),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_431),
.Y(n_628)
);

BUFx3_ASAP7_75t_L g629 ( 
.A(n_351),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_455),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_L g631 ( 
.A(n_509),
.B(n_4),
.Y(n_631)
);

BUFx6f_ASAP7_75t_L g632 ( 
.A(n_408),
.Y(n_632)
);

INVxp67_ASAP7_75t_L g633 ( 
.A(n_474),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_481),
.Y(n_634)
);

HB1xp67_ASAP7_75t_L g635 ( 
.A(n_337),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_531),
.Y(n_636)
);

NOR2xp33_ASAP7_75t_L g637 ( 
.A(n_335),
.B(n_5),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_554),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_490),
.Y(n_639)
);

CKINVDCx20_ASAP7_75t_R g640 ( 
.A(n_400),
.Y(n_640)
);

CKINVDCx20_ASAP7_75t_R g641 ( 
.A(n_466),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_496),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_516),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_572),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_519),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_523),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_534),
.Y(n_647)
);

CKINVDCx20_ASAP7_75t_R g648 ( 
.A(n_515),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_573),
.Y(n_649)
);

INVxp67_ASAP7_75t_L g650 ( 
.A(n_544),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_349),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_547),
.Y(n_652)
);

CKINVDCx16_ASAP7_75t_R g653 ( 
.A(n_406),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_557),
.Y(n_654)
);

CKINVDCx20_ASAP7_75t_R g655 ( 
.A(n_480),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_421),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_355),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_355),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_588),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_346),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_353),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_366),
.Y(n_662)
);

CKINVDCx20_ASAP7_75t_R g663 ( 
.A(n_561),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_580),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_382),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_583),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_586),
.Y(n_667)
);

CKINVDCx20_ASAP7_75t_R g668 ( 
.A(n_384),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_601),
.B(n_359),
.Y(n_669)
);

CKINVDCx20_ASAP7_75t_R g670 ( 
.A(n_620),
.Y(n_670)
);

AND2x2_ASAP7_75t_L g671 ( 
.A(n_653),
.B(n_561),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_591),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_589),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_594),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_592),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_596),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_629),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_598),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_599),
.B(n_391),
.Y(n_679)
);

CKINVDCx20_ASAP7_75t_R g680 ( 
.A(n_620),
.Y(n_680)
);

HB1xp67_ASAP7_75t_L g681 ( 
.A(n_635),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_597),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_604),
.Y(n_683)
);

CKINVDCx16_ASAP7_75t_R g684 ( 
.A(n_600),
.Y(n_684)
);

HB1xp67_ASAP7_75t_L g685 ( 
.A(n_659),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_605),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_629),
.B(n_395),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_603),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_606),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_607),
.Y(n_690)
);

INVx3_ASAP7_75t_L g691 ( 
.A(n_651),
.Y(n_691)
);

INVxp67_ASAP7_75t_L g692 ( 
.A(n_660),
.Y(n_692)
);

NOR2xp33_ASAP7_75t_R g693 ( 
.A(n_590),
.B(n_340),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_608),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_609),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_651),
.Y(n_696)
);

NOR2xp67_ASAP7_75t_L g697 ( 
.A(n_633),
.B(n_341),
.Y(n_697)
);

BUFx2_ASAP7_75t_L g698 ( 
.A(n_661),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_624),
.B(n_628),
.Y(n_699)
);

BUFx6f_ASAP7_75t_L g700 ( 
.A(n_632),
.Y(n_700)
);

OAI22xp5_ASAP7_75t_SL g701 ( 
.A1(n_625),
.A2(n_422),
.B1(n_425),
.B2(n_418),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_595),
.Y(n_702)
);

BUFx2_ASAP7_75t_L g703 ( 
.A(n_662),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_630),
.Y(n_704)
);

AOI22xp5_ASAP7_75t_L g705 ( 
.A1(n_650),
.A2(n_593),
.B1(n_619),
.B2(n_590),
.Y(n_705)
);

INVx1_ASAP7_75t_SL g706 ( 
.A(n_668),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_634),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_610),
.Y(n_708)
);

AND2x6_ASAP7_75t_L g709 ( 
.A(n_621),
.B(n_351),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_613),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_639),
.Y(n_711)
);

BUFx2_ASAP7_75t_L g712 ( 
.A(n_665),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_642),
.Y(n_713)
);

BUFx3_ASAP7_75t_L g714 ( 
.A(n_612),
.Y(n_714)
);

AND2x2_ASAP7_75t_L g715 ( 
.A(n_656),
.B(n_439),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_616),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_622),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_643),
.Y(n_718)
);

AND2x2_ASAP7_75t_L g719 ( 
.A(n_657),
.B(n_439),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_645),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_646),
.Y(n_721)
);

BUFx6f_ASAP7_75t_L g722 ( 
.A(n_632),
.Y(n_722)
);

BUFx6f_ASAP7_75t_L g723 ( 
.A(n_632),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_647),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_615),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_617),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_626),
.Y(n_727)
);

CKINVDCx16_ASAP7_75t_R g728 ( 
.A(n_602),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_658),
.B(n_426),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_618),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_636),
.Y(n_731)
);

INVx3_ASAP7_75t_L g732 ( 
.A(n_623),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_652),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_654),
.Y(n_734)
);

CKINVDCx5p33_ASAP7_75t_R g735 ( 
.A(n_638),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_SL g736 ( 
.A(n_664),
.B(n_462),
.Y(n_736)
);

INVxp67_ASAP7_75t_L g737 ( 
.A(n_644),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_666),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_SL g739 ( 
.A(n_667),
.B(n_462),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_614),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_649),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_611),
.Y(n_742)
);

AND2x2_ASAP7_75t_L g743 ( 
.A(n_663),
.B(n_506),
.Y(n_743)
);

CKINVDCx20_ASAP7_75t_R g744 ( 
.A(n_625),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_632),
.Y(n_745)
);

CKINVDCx20_ASAP7_75t_R g746 ( 
.A(n_627),
.Y(n_746)
);

INVxp67_ASAP7_75t_SL g747 ( 
.A(n_631),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_637),
.Y(n_748)
);

NAND2x1_ASAP7_75t_L g749 ( 
.A(n_663),
.B(n_342),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_655),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_648),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_627),
.Y(n_752)
);

INVxp67_ASAP7_75t_L g753 ( 
.A(n_640),
.Y(n_753)
);

INVx1_ASAP7_75t_SL g754 ( 
.A(n_640),
.Y(n_754)
);

BUFx8_ASAP7_75t_L g755 ( 
.A(n_641),
.Y(n_755)
);

HB1xp67_ASAP7_75t_L g756 ( 
.A(n_641),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_589),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_591),
.Y(n_758)
);

HB1xp67_ASAP7_75t_L g759 ( 
.A(n_635),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_599),
.B(n_433),
.Y(n_760)
);

CKINVDCx8_ASAP7_75t_R g761 ( 
.A(n_653),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_589),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_629),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_589),
.Y(n_764)
);

BUFx6f_ASAP7_75t_L g765 ( 
.A(n_632),
.Y(n_765)
);

INVx3_ASAP7_75t_L g766 ( 
.A(n_629),
.Y(n_766)
);

BUFx6f_ASAP7_75t_L g767 ( 
.A(n_632),
.Y(n_767)
);

AND2x4_ASAP7_75t_L g768 ( 
.A(n_599),
.B(n_372),
.Y(n_768)
);

BUFx6f_ASAP7_75t_L g769 ( 
.A(n_632),
.Y(n_769)
);

HB1xp67_ASAP7_75t_L g770 ( 
.A(n_635),
.Y(n_770)
);

AND2x6_ASAP7_75t_L g771 ( 
.A(n_619),
.B(n_398),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_591),
.Y(n_772)
);

INVx4_ASAP7_75t_L g773 ( 
.A(n_629),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_589),
.Y(n_774)
);

BUFx6f_ASAP7_75t_L g775 ( 
.A(n_632),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_589),
.Y(n_776)
);

BUFx6f_ASAP7_75t_L g777 ( 
.A(n_632),
.Y(n_777)
);

INVx4_ASAP7_75t_L g778 ( 
.A(n_629),
.Y(n_778)
);

CKINVDCx5p33_ASAP7_75t_R g779 ( 
.A(n_591),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_591),
.Y(n_780)
);

XNOR2x2_ASAP7_75t_L g781 ( 
.A(n_593),
.B(n_565),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_589),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_629),
.Y(n_783)
);

BUFx2_ASAP7_75t_L g784 ( 
.A(n_659),
.Y(n_784)
);

INVx3_ASAP7_75t_L g785 ( 
.A(n_629),
.Y(n_785)
);

CKINVDCx20_ASAP7_75t_R g786 ( 
.A(n_620),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_589),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_589),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_629),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_591),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_589),
.Y(n_791)
);

CKINVDCx5p33_ASAP7_75t_R g792 ( 
.A(n_591),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_589),
.Y(n_793)
);

CKINVDCx5p33_ASAP7_75t_R g794 ( 
.A(n_591),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_601),
.B(n_359),
.Y(n_795)
);

CKINVDCx5p33_ASAP7_75t_R g796 ( 
.A(n_591),
.Y(n_796)
);

INVx3_ASAP7_75t_L g797 ( 
.A(n_629),
.Y(n_797)
);

CKINVDCx5p33_ASAP7_75t_R g798 ( 
.A(n_591),
.Y(n_798)
);

NOR2xp33_ASAP7_75t_L g799 ( 
.A(n_599),
.B(n_348),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_591),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_589),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_589),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_589),
.Y(n_803)
);

AND2x6_ASAP7_75t_L g804 ( 
.A(n_619),
.B(n_398),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_591),
.Y(n_805)
);

CKINVDCx16_ASAP7_75t_R g806 ( 
.A(n_653),
.Y(n_806)
);

NOR2xp33_ASAP7_75t_R g807 ( 
.A(n_590),
.B(n_343),
.Y(n_807)
);

CKINVDCx5p33_ASAP7_75t_R g808 ( 
.A(n_591),
.Y(n_808)
);

CKINVDCx5p33_ASAP7_75t_R g809 ( 
.A(n_591),
.Y(n_809)
);

CKINVDCx20_ASAP7_75t_R g810 ( 
.A(n_620),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_589),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_589),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_629),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_766),
.Y(n_814)
);

AND2x4_ASAP7_75t_L g815 ( 
.A(n_736),
.B(n_568),
.Y(n_815)
);

INVx3_ASAP7_75t_L g816 ( 
.A(n_766),
.Y(n_816)
);

CKINVDCx5p33_ASAP7_75t_R g817 ( 
.A(n_742),
.Y(n_817)
);

BUFx6f_ASAP7_75t_L g818 ( 
.A(n_785),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_768),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_768),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_748),
.B(n_704),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_714),
.Y(n_822)
);

NOR2xp33_ASAP7_75t_L g823 ( 
.A(n_729),
.B(n_747),
.Y(n_823)
);

NOR2xp33_ASAP7_75t_L g824 ( 
.A(n_679),
.B(n_506),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_707),
.B(n_350),
.Y(n_825)
);

AOI22xp33_ASAP7_75t_L g826 ( 
.A1(n_771),
.A2(n_386),
.B1(n_477),
.B2(n_372),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_711),
.B(n_354),
.Y(n_827)
);

AND2x4_ASAP7_75t_L g828 ( 
.A(n_739),
.B(n_437),
.Y(n_828)
);

NOR2xp33_ASAP7_75t_L g829 ( 
.A(n_760),
.B(n_527),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_732),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_SL g831 ( 
.A(n_713),
.B(n_356),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_732),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_683),
.Y(n_833)
);

CKINVDCx5p33_ASAP7_75t_R g834 ( 
.A(n_751),
.Y(n_834)
);

OR2x6_ASAP7_75t_L g835 ( 
.A(n_737),
.B(n_372),
.Y(n_835)
);

NAND3xp33_ASAP7_75t_SL g836 ( 
.A(n_706),
.B(n_445),
.C(n_443),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_686),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_718),
.B(n_362),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_689),
.Y(n_839)
);

NOR2xp33_ASAP7_75t_L g840 ( 
.A(n_719),
.B(n_527),
.Y(n_840)
);

AND3x1_ASAP7_75t_L g841 ( 
.A(n_705),
.B(n_357),
.C(n_352),
.Y(n_841)
);

CKINVDCx5p33_ASAP7_75t_R g842 ( 
.A(n_755),
.Y(n_842)
);

AND2x4_ASAP7_75t_L g843 ( 
.A(n_740),
.B(n_459),
.Y(n_843)
);

INVx3_ASAP7_75t_L g844 ( 
.A(n_785),
.Y(n_844)
);

NOR2x1p5_ASAP7_75t_L g845 ( 
.A(n_749),
.B(n_468),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_690),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_694),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_708),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_725),
.Y(n_849)
);

BUFx6f_ASAP7_75t_L g850 ( 
.A(n_797),
.Y(n_850)
);

AND2x4_ASAP7_75t_L g851 ( 
.A(n_697),
.B(n_475),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_726),
.Y(n_852)
);

BUFx6f_ASAP7_75t_L g853 ( 
.A(n_797),
.Y(n_853)
);

INVx2_ASAP7_75t_L g854 ( 
.A(n_677),
.Y(n_854)
);

BUFx10_ASAP7_75t_L g855 ( 
.A(n_685),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_730),
.Y(n_856)
);

BUFx3_ASAP7_75t_L g857 ( 
.A(n_698),
.Y(n_857)
);

AOI22xp33_ASAP7_75t_L g858 ( 
.A1(n_771),
.A2(n_386),
.B1(n_477),
.B2(n_372),
.Y(n_858)
);

AOI22xp33_ASAP7_75t_L g859 ( 
.A1(n_771),
.A2(n_477),
.B1(n_386),
.B2(n_360),
.Y(n_859)
);

AND2x4_ASAP7_75t_L g860 ( 
.A(n_702),
.B(n_503),
.Y(n_860)
);

AND2x6_ASAP7_75t_L g861 ( 
.A(n_671),
.B(n_514),
.Y(n_861)
);

AND2x2_ASAP7_75t_SL g862 ( 
.A(n_806),
.B(n_386),
.Y(n_862)
);

AND2x2_ASAP7_75t_L g863 ( 
.A(n_681),
.B(n_512),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_763),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_673),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_783),
.Y(n_866)
);

INVx2_ASAP7_75t_L g867 ( 
.A(n_789),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_813),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_675),
.Y(n_869)
);

NOR2xp33_ASAP7_75t_L g870 ( 
.A(n_715),
.B(n_535),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_720),
.B(n_364),
.Y(n_871)
);

NOR2xp33_ASAP7_75t_L g872 ( 
.A(n_759),
.B(n_535),
.Y(n_872)
);

INVx3_ASAP7_75t_L g873 ( 
.A(n_773),
.Y(n_873)
);

NOR2xp33_ASAP7_75t_L g874 ( 
.A(n_770),
.B(n_457),
.Y(n_874)
);

NOR2xp33_ASAP7_75t_L g875 ( 
.A(n_721),
.B(n_578),
.Y(n_875)
);

AND2x6_ASAP7_75t_L g876 ( 
.A(n_743),
.B(n_514),
.Y(n_876)
);

NOR2xp33_ASAP7_75t_L g877 ( 
.A(n_724),
.B(n_733),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_678),
.Y(n_878)
);

AND2x2_ASAP7_75t_L g879 ( 
.A(n_703),
.B(n_522),
.Y(n_879)
);

BUFx3_ASAP7_75t_L g880 ( 
.A(n_712),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_773),
.Y(n_881)
);

OR2x2_ASAP7_75t_L g882 ( 
.A(n_706),
.B(n_524),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_778),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_757),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_762),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_778),
.Y(n_886)
);

NOR2xp33_ASAP7_75t_L g887 ( 
.A(n_734),
.B(n_367),
.Y(n_887)
);

CKINVDCx5p33_ASAP7_75t_R g888 ( 
.A(n_755),
.Y(n_888)
);

INVxp67_ASAP7_75t_L g889 ( 
.A(n_784),
.Y(n_889)
);

BUFx2_ASAP7_75t_L g890 ( 
.A(n_693),
.Y(n_890)
);

AND2x4_ASAP7_75t_L g891 ( 
.A(n_692),
.B(n_530),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_764),
.Y(n_892)
);

CKINVDCx5p33_ASAP7_75t_R g893 ( 
.A(n_670),
.Y(n_893)
);

INVx4_ASAP7_75t_L g894 ( 
.A(n_771),
.Y(n_894)
);

INVx2_ASAP7_75t_L g895 ( 
.A(n_691),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_738),
.B(n_368),
.Y(n_896)
);

INVx5_ASAP7_75t_L g897 ( 
.A(n_804),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_774),
.Y(n_898)
);

INVx4_ASAP7_75t_SL g899 ( 
.A(n_804),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_776),
.Y(n_900)
);

BUFx2_ASAP7_75t_L g901 ( 
.A(n_807),
.Y(n_901)
);

NOR2x1p5_ASAP7_75t_L g902 ( 
.A(n_672),
.B(n_539),
.Y(n_902)
);

HB1xp67_ASAP7_75t_L g903 ( 
.A(n_754),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_782),
.Y(n_904)
);

INVx3_ASAP7_75t_L g905 ( 
.A(n_787),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_SL g906 ( 
.A(n_699),
.B(n_369),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_SL g907 ( 
.A(n_699),
.B(n_371),
.Y(n_907)
);

INVx3_ASAP7_75t_L g908 ( 
.A(n_788),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_691),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_696),
.Y(n_910)
);

CKINVDCx5p33_ASAP7_75t_R g911 ( 
.A(n_680),
.Y(n_911)
);

INVx2_ASAP7_75t_L g912 ( 
.A(n_791),
.Y(n_912)
);

BUFx6f_ASAP7_75t_L g913 ( 
.A(n_804),
.Y(n_913)
);

AND2x2_ASAP7_75t_L g914 ( 
.A(n_705),
.B(n_546),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_SL g915 ( 
.A(n_687),
.B(n_374),
.Y(n_915)
);

CKINVDCx20_ASAP7_75t_R g916 ( 
.A(n_744),
.Y(n_916)
);

INVx2_ASAP7_75t_SL g917 ( 
.A(n_804),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_793),
.Y(n_918)
);

INVx3_ASAP7_75t_L g919 ( 
.A(n_801),
.Y(n_919)
);

INVx3_ASAP7_75t_L g920 ( 
.A(n_802),
.Y(n_920)
);

AND2x4_ASAP7_75t_SL g921 ( 
.A(n_756),
.B(n_477),
.Y(n_921)
);

AOI22xp5_ASAP7_75t_L g922 ( 
.A1(n_799),
.A2(n_552),
.B1(n_560),
.B2(n_553),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_803),
.B(n_375),
.Y(n_923)
);

AOI22xp5_ASAP7_75t_L g924 ( 
.A1(n_709),
.A2(n_563),
.B1(n_569),
.B2(n_564),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_812),
.Y(n_925)
);

INVx2_ASAP7_75t_L g926 ( 
.A(n_811),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_669),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_SL g928 ( 
.A(n_669),
.B(n_376),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_795),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_709),
.B(n_378),
.Y(n_930)
);

NOR2xp33_ASAP7_75t_L g931 ( 
.A(n_761),
.B(n_379),
.Y(n_931)
);

BUFx2_ASAP7_75t_L g932 ( 
.A(n_674),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_795),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_709),
.B(n_380),
.Y(n_934)
);

AND2x2_ASAP7_75t_L g935 ( 
.A(n_676),
.B(n_571),
.Y(n_935)
);

BUFx10_ASAP7_75t_L g936 ( 
.A(n_682),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_781),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_709),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_SL g939 ( 
.A(n_688),
.B(n_385),
.Y(n_939)
);

CKINVDCx5p33_ASAP7_75t_R g940 ( 
.A(n_746),
.Y(n_940)
);

AND2x2_ASAP7_75t_L g941 ( 
.A(n_695),
.B(n_710),
.Y(n_941)
);

AND2x2_ASAP7_75t_L g942 ( 
.A(n_716),
.B(n_436),
.Y(n_942)
);

AND2x4_ASAP7_75t_L g943 ( 
.A(n_717),
.B(n_727),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_745),
.Y(n_944)
);

BUFx6f_ASAP7_75t_L g945 ( 
.A(n_700),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_701),
.Y(n_946)
);

NOR2xp33_ASAP7_75t_L g947 ( 
.A(n_753),
.B(n_387),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_731),
.B(n_388),
.Y(n_948)
);

BUFx3_ASAP7_75t_L g949 ( 
.A(n_735),
.Y(n_949)
);

AND2x4_ASAP7_75t_L g950 ( 
.A(n_741),
.B(n_538),
.Y(n_950)
);

AND2x4_ASAP7_75t_L g951 ( 
.A(n_758),
.B(n_538),
.Y(n_951)
);

BUFx3_ASAP7_75t_L g952 ( 
.A(n_772),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_779),
.B(n_392),
.Y(n_953)
);

OR2x2_ASAP7_75t_L g954 ( 
.A(n_754),
.B(n_6),
.Y(n_954)
);

AO21x2_ASAP7_75t_L g955 ( 
.A1(n_752),
.A2(n_365),
.B(n_363),
.Y(n_955)
);

AND2x6_ASAP7_75t_L g956 ( 
.A(n_750),
.B(n_556),
.Y(n_956)
);

BUFx3_ASAP7_75t_L g957 ( 
.A(n_780),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_SL g958 ( 
.A(n_790),
.B(n_393),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_792),
.B(n_394),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_700),
.Y(n_960)
);

INVx3_ASAP7_75t_L g961 ( 
.A(n_700),
.Y(n_961)
);

AND2x6_ASAP7_75t_L g962 ( 
.A(n_722),
.B(n_556),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_722),
.Y(n_963)
);

BUFx6f_ASAP7_75t_L g964 ( 
.A(n_722),
.Y(n_964)
);

AND2x4_ASAP7_75t_L g965 ( 
.A(n_794),
.B(n_373),
.Y(n_965)
);

INVx3_ASAP7_75t_L g966 ( 
.A(n_723),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_796),
.B(n_397),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_798),
.B(n_399),
.Y(n_968)
);

INVx6_ASAP7_75t_L g969 ( 
.A(n_728),
.Y(n_969)
);

BUFx3_ASAP7_75t_L g970 ( 
.A(n_800),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_805),
.B(n_403),
.Y(n_971)
);

INVx1_ASAP7_75t_SL g972 ( 
.A(n_808),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_701),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_809),
.B(n_404),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_723),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_723),
.Y(n_976)
);

NAND2x1p5_ASAP7_75t_L g977 ( 
.A(n_684),
.B(n_377),
.Y(n_977)
);

INVx8_ASAP7_75t_L g978 ( 
.A(n_810),
.Y(n_978)
);

AND2x2_ASAP7_75t_SL g979 ( 
.A(n_786),
.B(n_383),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_765),
.B(n_407),
.Y(n_980)
);

NAND2xp33_ASAP7_75t_L g981 ( 
.A(n_765),
.B(n_349),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_765),
.Y(n_982)
);

NOR2xp33_ASAP7_75t_L g983 ( 
.A(n_767),
.B(n_411),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_767),
.Y(n_984)
);

AO22x2_ASAP7_75t_L g985 ( 
.A1(n_767),
.A2(n_389),
.B1(n_402),
.B2(n_390),
.Y(n_985)
);

INVx2_ASAP7_75t_L g986 ( 
.A(n_777),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_769),
.B(n_412),
.Y(n_987)
);

INVx2_ASAP7_75t_L g988 ( 
.A(n_777),
.Y(n_988)
);

AND2x4_ASAP7_75t_L g989 ( 
.A(n_769),
.B(n_409),
.Y(n_989)
);

BUFx3_ASAP7_75t_L g990 ( 
.A(n_769),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_SL g991 ( 
.A(n_775),
.B(n_414),
.Y(n_991)
);

AND2x4_ASAP7_75t_L g992 ( 
.A(n_775),
.B(n_415),
.Y(n_992)
);

INVx2_ASAP7_75t_L g993 ( 
.A(n_775),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_777),
.B(n_416),
.Y(n_994)
);

OR2x6_ASAP7_75t_L g995 ( 
.A(n_737),
.B(n_417),
.Y(n_995)
);

BUFx10_ASAP7_75t_L g996 ( 
.A(n_685),
.Y(n_996)
);

BUFx2_ASAP7_75t_L g997 ( 
.A(n_681),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_768),
.Y(n_998)
);

INVx2_ASAP7_75t_L g999 ( 
.A(n_766),
.Y(n_999)
);

NOR2xp33_ASAP7_75t_L g1000 ( 
.A(n_729),
.B(n_419),
.Y(n_1000)
);

OR2x2_ASAP7_75t_SL g1001 ( 
.A(n_728),
.B(n_430),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_768),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_768),
.Y(n_1003)
);

NOR2x1p5_ASAP7_75t_L g1004 ( 
.A(n_749),
.B(n_420),
.Y(n_1004)
);

INVx1_ASAP7_75t_SL g1005 ( 
.A(n_706),
.Y(n_1005)
);

INVx2_ASAP7_75t_L g1006 ( 
.A(n_766),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_768),
.Y(n_1007)
);

NAND2x1p5_ASAP7_75t_L g1008 ( 
.A(n_698),
.B(n_440),
.Y(n_1008)
);

OR2x2_ASAP7_75t_L g1009 ( 
.A(n_706),
.B(n_6),
.Y(n_1009)
);

OR2x6_ASAP7_75t_L g1010 ( 
.A(n_737),
.B(n_449),
.Y(n_1010)
);

OAI21xp33_ASAP7_75t_L g1011 ( 
.A1(n_799),
.A2(n_424),
.B(n_423),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_768),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_768),
.Y(n_1013)
);

INVx3_ASAP7_75t_L g1014 ( 
.A(n_766),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_748),
.B(n_429),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_SL g1016 ( 
.A(n_748),
.B(n_432),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_SL g1017 ( 
.A(n_748),
.B(n_434),
.Y(n_1017)
);

INVx3_ASAP7_75t_L g1018 ( 
.A(n_766),
.Y(n_1018)
);

INVx2_ASAP7_75t_L g1019 ( 
.A(n_766),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_768),
.Y(n_1020)
);

AND2x2_ASAP7_75t_L g1021 ( 
.A(n_681),
.B(n_435),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_748),
.B(n_441),
.Y(n_1022)
);

AND2x6_ASAP7_75t_L g1023 ( 
.A(n_671),
.B(n_451),
.Y(n_1023)
);

BUFx2_ASAP7_75t_L g1024 ( 
.A(n_681),
.Y(n_1024)
);

AND2x4_ASAP7_75t_L g1025 ( 
.A(n_736),
.B(n_454),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_768),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_748),
.B(n_442),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_732),
.Y(n_1028)
);

INVx2_ASAP7_75t_SL g1029 ( 
.A(n_681),
.Y(n_1029)
);

INVx4_ASAP7_75t_L g1030 ( 
.A(n_773),
.Y(n_1030)
);

INVx4_ASAP7_75t_L g1031 ( 
.A(n_773),
.Y(n_1031)
);

INVx3_ASAP7_75t_L g1032 ( 
.A(n_766),
.Y(n_1032)
);

HB1xp67_ASAP7_75t_L g1033 ( 
.A(n_681),
.Y(n_1033)
);

INVx2_ASAP7_75t_L g1034 ( 
.A(n_766),
.Y(n_1034)
);

INVx2_ASAP7_75t_L g1035 ( 
.A(n_766),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_927),
.B(n_458),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_929),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_933),
.B(n_444),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_925),
.B(n_460),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_925),
.B(n_461),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_865),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_869),
.Y(n_1042)
);

AND2x2_ASAP7_75t_SL g1043 ( 
.A(n_979),
.B(n_585),
.Y(n_1043)
);

INVx2_ASAP7_75t_SL g1044 ( 
.A(n_857),
.Y(n_1044)
);

NOR2xp33_ASAP7_75t_L g1045 ( 
.A(n_1029),
.B(n_446),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_SL g1046 ( 
.A(n_891),
.B(n_447),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_905),
.B(n_463),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_878),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_905),
.B(n_464),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_SL g1050 ( 
.A(n_891),
.B(n_913),
.Y(n_1050)
);

BUFx6f_ASAP7_75t_L g1051 ( 
.A(n_913),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_823),
.B(n_448),
.Y(n_1052)
);

NOR2xp33_ASAP7_75t_L g1053 ( 
.A(n_1033),
.B(n_450),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_884),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_885),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_821),
.B(n_452),
.Y(n_1056)
);

OR2x6_ASAP7_75t_L g1057 ( 
.A(n_880),
.B(n_465),
.Y(n_1057)
);

AOI22xp33_ASAP7_75t_L g1058 ( 
.A1(n_937),
.A2(n_476),
.B1(n_478),
.B2(n_470),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_877),
.B(n_456),
.Y(n_1059)
);

NOR2xp33_ASAP7_75t_L g1060 ( 
.A(n_997),
.B(n_467),
.Y(n_1060)
);

INVx2_ASAP7_75t_L g1061 ( 
.A(n_908),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_892),
.Y(n_1062)
);

AOI22xp5_ASAP7_75t_L g1063 ( 
.A1(n_841),
.A2(n_507),
.B1(n_513),
.B2(n_499),
.Y(n_1063)
);

NOR2xp33_ASAP7_75t_L g1064 ( 
.A(n_1024),
.B(n_469),
.Y(n_1064)
);

NOR2xp33_ASAP7_75t_L g1065 ( 
.A(n_828),
.B(n_471),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_SL g1066 ( 
.A(n_913),
.B(n_472),
.Y(n_1066)
);

CKINVDCx11_ASAP7_75t_R g1067 ( 
.A(n_936),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_908),
.B(n_483),
.Y(n_1068)
);

INVx2_ASAP7_75t_SL g1069 ( 
.A(n_855),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_919),
.B(n_484),
.Y(n_1070)
);

INVx2_ASAP7_75t_SL g1071 ( 
.A(n_855),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_919),
.B(n_485),
.Y(n_1072)
);

NOR2xp33_ASAP7_75t_L g1073 ( 
.A(n_828),
.B(n_487),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_898),
.Y(n_1074)
);

INVx2_ASAP7_75t_L g1075 ( 
.A(n_920),
.Y(n_1075)
);

BUFx2_ASAP7_75t_L g1076 ( 
.A(n_1005),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_SL g1077 ( 
.A(n_897),
.B(n_489),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_900),
.Y(n_1078)
);

AOI22xp5_ASAP7_75t_L g1079 ( 
.A1(n_1023),
.A2(n_528),
.B1(n_537),
.B2(n_526),
.Y(n_1079)
);

AOI22xp5_ASAP7_75t_L g1080 ( 
.A1(n_1023),
.A2(n_551),
.B1(n_559),
.B2(n_549),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_SL g1081 ( 
.A(n_897),
.B(n_491),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_920),
.B(n_492),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_912),
.B(n_493),
.Y(n_1083)
);

OAI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_1028),
.A2(n_570),
.B(n_562),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_904),
.Y(n_1085)
);

NOR2xp33_ASAP7_75t_L g1086 ( 
.A(n_889),
.B(n_495),
.Y(n_1086)
);

INVx1_ASAP7_75t_SL g1087 ( 
.A(n_903),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_918),
.Y(n_1088)
);

NOR3xp33_ASAP7_75t_L g1089 ( 
.A(n_946),
.B(n_973),
.C(n_836),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_926),
.B(n_833),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_SL g1091 ( 
.A(n_897),
.B(n_894),
.Y(n_1091)
);

NAND2x1_ASAP7_75t_L g1092 ( 
.A(n_894),
.B(n_361),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_837),
.B(n_498),
.Y(n_1093)
);

NOR2xp67_ASAP7_75t_L g1094 ( 
.A(n_842),
.B(n_7),
.Y(n_1094)
);

NOR2xp33_ASAP7_75t_L g1095 ( 
.A(n_863),
.B(n_500),
.Y(n_1095)
);

INVx2_ASAP7_75t_L g1096 ( 
.A(n_989),
.Y(n_1096)
);

AND2x6_ASAP7_75t_SL g1097 ( 
.A(n_943),
.B(n_574),
.Y(n_1097)
);

BUFx12f_ASAP7_75t_L g1098 ( 
.A(n_888),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_SL g1099 ( 
.A(n_996),
.B(n_917),
.Y(n_1099)
);

AOI22xp33_ASAP7_75t_L g1100 ( 
.A1(n_914),
.A2(n_584),
.B1(n_361),
.B2(n_428),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_839),
.B(n_427),
.Y(n_1101)
);

AOI22xp33_ASAP7_75t_L g1102 ( 
.A1(n_876),
.A2(n_427),
.B1(n_438),
.B2(n_428),
.Y(n_1102)
);

INVx2_ASAP7_75t_L g1103 ( 
.A(n_989),
.Y(n_1103)
);

OAI21xp5_ASAP7_75t_L g1104 ( 
.A1(n_1028),
.A2(n_494),
.B(n_438),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_846),
.B(n_501),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_819),
.Y(n_1106)
);

NOR2xp33_ASAP7_75t_L g1107 ( 
.A(n_1021),
.B(n_502),
.Y(n_1107)
);

AOI22xp33_ASAP7_75t_L g1108 ( 
.A1(n_876),
.A2(n_494),
.B1(n_548),
.B2(n_497),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_847),
.B(n_508),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_875),
.B(n_510),
.Y(n_1110)
);

NOR2xp33_ASAP7_75t_L g1111 ( 
.A(n_870),
.B(n_511),
.Y(n_1111)
);

AND2x2_ASAP7_75t_L g1112 ( 
.A(n_996),
.B(n_9),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_SL g1113 ( 
.A(n_1008),
.B(n_517),
.Y(n_1113)
);

CKINVDCx20_ASAP7_75t_R g1114 ( 
.A(n_916),
.Y(n_1114)
);

NOR2xp33_ASAP7_75t_L g1115 ( 
.A(n_879),
.B(n_518),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_820),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_SL g1117 ( 
.A(n_1025),
.B(n_520),
.Y(n_1117)
);

INVx2_ASAP7_75t_L g1118 ( 
.A(n_992),
.Y(n_1118)
);

NOR2xp33_ASAP7_75t_L g1119 ( 
.A(n_840),
.B(n_521),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_861),
.B(n_525),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_861),
.B(n_529),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_998),
.Y(n_1122)
);

AND2x4_ASAP7_75t_L g1123 ( 
.A(n_845),
.B(n_11),
.Y(n_1123)
);

INVx2_ASAP7_75t_SL g1124 ( 
.A(n_835),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_SL g1125 ( 
.A(n_1025),
.B(n_899),
.Y(n_1125)
);

INVx3_ASAP7_75t_L g1126 ( 
.A(n_1030),
.Y(n_1126)
);

AOI21xp5_ASAP7_75t_L g1127 ( 
.A1(n_1015),
.A2(n_548),
.B(n_540),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_861),
.B(n_532),
.Y(n_1128)
);

INVx4_ASAP7_75t_L g1129 ( 
.A(n_835),
.Y(n_1129)
);

INVx3_ASAP7_75t_L g1130 ( 
.A(n_1030),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_1002),
.Y(n_1131)
);

INVx2_ASAP7_75t_SL g1132 ( 
.A(n_921),
.Y(n_1132)
);

NOR2xp33_ASAP7_75t_L g1133 ( 
.A(n_965),
.B(n_541),
.Y(n_1133)
);

INVx3_ASAP7_75t_L g1134 ( 
.A(n_1031),
.Y(n_1134)
);

INVxp67_ASAP7_75t_L g1135 ( 
.A(n_932),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_861),
.B(n_543),
.Y(n_1136)
);

AOI22xp33_ASAP7_75t_L g1137 ( 
.A1(n_876),
.A2(n_497),
.B1(n_349),
.B2(n_545),
.Y(n_1137)
);

INVx2_ASAP7_75t_L g1138 ( 
.A(n_992),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_955),
.B(n_550),
.Y(n_1139)
);

INVx2_ASAP7_75t_L g1140 ( 
.A(n_818),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_SL g1141 ( 
.A(n_899),
.B(n_581),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_SL g1142 ( 
.A(n_965),
.B(n_555),
.Y(n_1142)
);

INVx2_ASAP7_75t_L g1143 ( 
.A(n_818),
.Y(n_1143)
);

AND2x2_ASAP7_75t_L g1144 ( 
.A(n_972),
.B(n_11),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_848),
.B(n_558),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_SL g1146 ( 
.A(n_930),
.B(n_577),
.Y(n_1146)
);

INVx2_ASAP7_75t_SL g1147 ( 
.A(n_995),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_SL g1148 ( 
.A(n_934),
.B(n_566),
.Y(n_1148)
);

OR2x6_ASAP7_75t_L g1149 ( 
.A(n_977),
.B(n_408),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_849),
.B(n_852),
.Y(n_1150)
);

NOR2xp33_ASAP7_75t_L g1151 ( 
.A(n_843),
.B(n_567),
.Y(n_1151)
);

AOI21xp5_ASAP7_75t_L g1152 ( 
.A1(n_1022),
.A2(n_408),
.B(n_349),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_856),
.B(n_349),
.Y(n_1153)
);

NAND3xp33_ASAP7_75t_SL g1154 ( 
.A(n_817),
.B(n_12),
.C(n_14),
.Y(n_1154)
);

BUFx3_ASAP7_75t_L g1155 ( 
.A(n_969),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_874),
.B(n_349),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_851),
.B(n_887),
.Y(n_1157)
);

INVx2_ASAP7_75t_L g1158 ( 
.A(n_818),
.Y(n_1158)
);

NOR2xp33_ASAP7_75t_L g1159 ( 
.A(n_843),
.B(n_12),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_1003),
.Y(n_1160)
);

O2A1O1Ixp33_ASAP7_75t_L g1161 ( 
.A1(n_954),
.A2(n_18),
.B(n_16),
.C(n_17),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_1007),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_851),
.B(n_497),
.Y(n_1163)
);

CKINVDCx5p33_ASAP7_75t_R g1164 ( 
.A(n_893),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_1012),
.Y(n_1165)
);

INVx2_ASAP7_75t_SL g1166 ( 
.A(n_995),
.Y(n_1166)
);

BUFx6f_ASAP7_75t_L g1167 ( 
.A(n_850),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_1027),
.B(n_497),
.Y(n_1168)
);

AOI21xp5_ASAP7_75t_L g1169 ( 
.A1(n_825),
.A2(n_408),
.B(n_497),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_876),
.B(n_497),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_SL g1171 ( 
.A(n_950),
.B(n_16),
.Y(n_1171)
);

AOI22xp5_ASAP7_75t_L g1172 ( 
.A1(n_1023),
.A2(n_20),
.B1(n_18),
.B2(n_19),
.Y(n_1172)
);

INVx2_ASAP7_75t_L g1173 ( 
.A(n_850),
.Y(n_1173)
);

AOI22xp33_ASAP7_75t_L g1174 ( 
.A1(n_1023),
.A2(n_22),
.B1(n_19),
.B2(n_21),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_815),
.B(n_24),
.Y(n_1175)
);

INVx2_ASAP7_75t_SL g1176 ( 
.A(n_1010),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_SL g1177 ( 
.A(n_950),
.B(n_24),
.Y(n_1177)
);

O2A1O1Ixp5_ASAP7_75t_L g1178 ( 
.A1(n_915),
.A2(n_113),
.B(n_114),
.C(n_111),
.Y(n_1178)
);

NOR2xp33_ASAP7_75t_L g1179 ( 
.A(n_860),
.B(n_25),
.Y(n_1179)
);

BUFx12f_ASAP7_75t_L g1180 ( 
.A(n_936),
.Y(n_1180)
);

AND2x6_ASAP7_75t_SL g1181 ( 
.A(n_943),
.B(n_26),
.Y(n_1181)
);

AND2x4_ASAP7_75t_L g1182 ( 
.A(n_1004),
.B(n_822),
.Y(n_1182)
);

BUFx3_ASAP7_75t_L g1183 ( 
.A(n_969),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_SL g1184 ( 
.A(n_951),
.B(n_850),
.Y(n_1184)
);

INVxp67_ASAP7_75t_L g1185 ( 
.A(n_882),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_1013),
.Y(n_1186)
);

O2A1O1Ixp33_ASAP7_75t_L g1187 ( 
.A1(n_1009),
.A2(n_30),
.B(n_27),
.C(n_29),
.Y(n_1187)
);

AND2x4_ASAP7_75t_SL g1188 ( 
.A(n_941),
.B(n_29),
.Y(n_1188)
);

AND2x2_ASAP7_75t_L g1189 ( 
.A(n_862),
.B(n_30),
.Y(n_1189)
);

AOI22xp33_ASAP7_75t_L g1190 ( 
.A1(n_985),
.A2(n_33),
.B1(n_31),
.B2(n_32),
.Y(n_1190)
);

INVx2_ASAP7_75t_L g1191 ( 
.A(n_853),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_815),
.B(n_31),
.Y(n_1192)
);

INVx2_ASAP7_75t_L g1193 ( 
.A(n_853),
.Y(n_1193)
);

INVx2_ASAP7_75t_L g1194 ( 
.A(n_853),
.Y(n_1194)
);

AOI22x1_ASAP7_75t_L g1195 ( 
.A1(n_938),
.A2(n_119),
.B1(n_120),
.B2(n_115),
.Y(n_1195)
);

AOI22xp5_ASAP7_75t_L g1196 ( 
.A1(n_860),
.A2(n_37),
.B1(n_32),
.B2(n_35),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_1000),
.B(n_35),
.Y(n_1197)
);

INVx2_ASAP7_75t_L g1198 ( 
.A(n_854),
.Y(n_1198)
);

OAI221xp5_ASAP7_75t_L g1199 ( 
.A1(n_922),
.A2(n_37),
.B1(n_39),
.B2(n_40),
.C(n_41),
.Y(n_1199)
);

NOR2xp33_ASAP7_75t_L g1200 ( 
.A(n_872),
.B(n_40),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_830),
.B(n_42),
.Y(n_1201)
);

AOI22xp5_ASAP7_75t_L g1202 ( 
.A1(n_942),
.A2(n_44),
.B1(n_42),
.B2(n_43),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_1020),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_1026),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_832),
.B(n_43),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_814),
.Y(n_1206)
);

INVx3_ASAP7_75t_L g1207 ( 
.A(n_1031),
.Y(n_1207)
);

CKINVDCx5p33_ASAP7_75t_R g1208 ( 
.A(n_911),
.Y(n_1208)
);

AOI22xp33_ASAP7_75t_L g1209 ( 
.A1(n_985),
.A2(n_46),
.B1(n_44),
.B2(n_45),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_924),
.B(n_45),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_999),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1006),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_824),
.B(n_46),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_829),
.B(n_47),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_827),
.B(n_47),
.Y(n_1215)
);

INVx2_ASAP7_75t_L g1216 ( 
.A(n_864),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_SL g1217 ( 
.A(n_951),
.B(n_48),
.Y(n_1217)
);

NOR2xp33_ASAP7_75t_L g1218 ( 
.A(n_935),
.B(n_49),
.Y(n_1218)
);

INVx2_ASAP7_75t_SL g1219 ( 
.A(n_1010),
.Y(n_1219)
);

CKINVDCx5p33_ASAP7_75t_R g1220 ( 
.A(n_940),
.Y(n_1220)
);

NOR2xp33_ASAP7_75t_L g1221 ( 
.A(n_947),
.B(n_50),
.Y(n_1221)
);

BUFx2_ASAP7_75t_L g1222 ( 
.A(n_1076),
.Y(n_1222)
);

AND2x2_ASAP7_75t_L g1223 ( 
.A(n_1087),
.B(n_949),
.Y(n_1223)
);

BUFx2_ASAP7_75t_L g1224 ( 
.A(n_1087),
.Y(n_1224)
);

INVx3_ASAP7_75t_SL g1225 ( 
.A(n_1164),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1037),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_1090),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_L g1228 ( 
.A(n_1089),
.B(n_838),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_L g1229 ( 
.A(n_1041),
.B(n_871),
.Y(n_1229)
);

NOR2xp33_ASAP7_75t_R g1230 ( 
.A(n_1067),
.B(n_834),
.Y(n_1230)
);

INVx2_ASAP7_75t_L g1231 ( 
.A(n_1042),
.Y(n_1231)
);

INVx2_ASAP7_75t_L g1232 ( 
.A(n_1048),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1054),
.Y(n_1233)
);

HB1xp67_ASAP7_75t_L g1234 ( 
.A(n_1044),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_1055),
.B(n_896),
.Y(n_1235)
);

NOR2xp33_ASAP7_75t_R g1236 ( 
.A(n_1114),
.B(n_978),
.Y(n_1236)
);

NOR2xp33_ASAP7_75t_L g1237 ( 
.A(n_1185),
.B(n_1001),
.Y(n_1237)
);

AOI22xp33_ASAP7_75t_L g1238 ( 
.A1(n_1043),
.A2(n_952),
.B1(n_970),
.B2(n_957),
.Y(n_1238)
);

AND2x4_ASAP7_75t_L g1239 ( 
.A(n_1069),
.B(n_1071),
.Y(n_1239)
);

NOR3xp33_ASAP7_75t_SL g1240 ( 
.A(n_1208),
.B(n_931),
.C(n_939),
.Y(n_1240)
);

BUFx3_ASAP7_75t_L g1241 ( 
.A(n_1180),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_L g1242 ( 
.A(n_1062),
.B(n_906),
.Y(n_1242)
);

AND2x2_ASAP7_75t_L g1243 ( 
.A(n_1057),
.B(n_890),
.Y(n_1243)
);

INVx2_ASAP7_75t_L g1244 ( 
.A(n_1074),
.Y(n_1244)
);

INVx3_ASAP7_75t_L g1245 ( 
.A(n_1126),
.Y(n_1245)
);

INVx3_ASAP7_75t_L g1246 ( 
.A(n_1126),
.Y(n_1246)
);

NOR3xp33_ASAP7_75t_SL g1247 ( 
.A(n_1220),
.B(n_958),
.C(n_953),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1078),
.Y(n_1248)
);

OR2x6_ASAP7_75t_L g1249 ( 
.A(n_1149),
.B(n_978),
.Y(n_1249)
);

CKINVDCx20_ASAP7_75t_R g1250 ( 
.A(n_1135),
.Y(n_1250)
);

INVx2_ASAP7_75t_L g1251 ( 
.A(n_1085),
.Y(n_1251)
);

INVx2_ASAP7_75t_L g1252 ( 
.A(n_1088),
.Y(n_1252)
);

NOR2xp33_ASAP7_75t_L g1253 ( 
.A(n_1147),
.B(n_901),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_L g1254 ( 
.A(n_1100),
.B(n_1036),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1150),
.Y(n_1255)
);

INVx4_ASAP7_75t_L g1256 ( 
.A(n_1149),
.Y(n_1256)
);

INVx2_ASAP7_75t_L g1257 ( 
.A(n_1106),
.Y(n_1257)
);

AND2x4_ASAP7_75t_SL g1258 ( 
.A(n_1149),
.B(n_816),
.Y(n_1258)
);

AOI22xp5_ASAP7_75t_L g1259 ( 
.A1(n_1166),
.A2(n_902),
.B1(n_956),
.B2(n_948),
.Y(n_1259)
);

INVx2_ASAP7_75t_L g1260 ( 
.A(n_1116),
.Y(n_1260)
);

INVx2_ASAP7_75t_L g1261 ( 
.A(n_1122),
.Y(n_1261)
);

NOR3xp33_ASAP7_75t_SL g1262 ( 
.A(n_1154),
.B(n_967),
.C(n_959),
.Y(n_1262)
);

INVx3_ASAP7_75t_SL g1263 ( 
.A(n_1057),
.Y(n_1263)
);

HB1xp67_ASAP7_75t_L g1264 ( 
.A(n_1057),
.Y(n_1264)
);

BUFx6f_ASAP7_75t_L g1265 ( 
.A(n_1051),
.Y(n_1265)
);

O2A1O1Ixp5_ASAP7_75t_L g1266 ( 
.A1(n_1197),
.A2(n_991),
.B(n_928),
.C(n_907),
.Y(n_1266)
);

NOR3xp33_ASAP7_75t_SL g1267 ( 
.A(n_1113),
.B(n_971),
.C(n_968),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1131),
.Y(n_1268)
);

AND2x2_ASAP7_75t_L g1269 ( 
.A(n_1176),
.B(n_974),
.Y(n_1269)
);

BUFx3_ASAP7_75t_L g1270 ( 
.A(n_1098),
.Y(n_1270)
);

INVx2_ASAP7_75t_L g1271 ( 
.A(n_1160),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_L g1272 ( 
.A(n_1036),
.B(n_923),
.Y(n_1272)
);

NOR3xp33_ASAP7_75t_SL g1273 ( 
.A(n_1046),
.B(n_1017),
.C(n_1016),
.Y(n_1273)
);

INVx2_ASAP7_75t_L g1274 ( 
.A(n_1162),
.Y(n_1274)
);

INVxp67_ASAP7_75t_L g1275 ( 
.A(n_1219),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1165),
.Y(n_1276)
);

CKINVDCx5p33_ASAP7_75t_R g1277 ( 
.A(n_1097),
.Y(n_1277)
);

BUFx4f_ASAP7_75t_L g1278 ( 
.A(n_1123),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_SL g1279 ( 
.A(n_1129),
.B(n_1011),
.Y(n_1279)
);

INVx5_ASAP7_75t_L g1280 ( 
.A(n_1129),
.Y(n_1280)
);

CKINVDCx5p33_ASAP7_75t_R g1281 ( 
.A(n_1155),
.Y(n_1281)
);

INVx1_ASAP7_75t_SL g1282 ( 
.A(n_1112),
.Y(n_1282)
);

INVx2_ASAP7_75t_L g1283 ( 
.A(n_1186),
.Y(n_1283)
);

OR2x6_ASAP7_75t_L g1284 ( 
.A(n_1183),
.B(n_831),
.Y(n_1284)
);

CKINVDCx20_ASAP7_75t_R g1285 ( 
.A(n_1188),
.Y(n_1285)
);

INVx1_ASAP7_75t_SL g1286 ( 
.A(n_1144),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_L g1287 ( 
.A(n_1175),
.B(n_956),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1203),
.Y(n_1288)
);

INVx1_ASAP7_75t_SL g1289 ( 
.A(n_1189),
.Y(n_1289)
);

NAND2xp33_ASAP7_75t_SL g1290 ( 
.A(n_1124),
.B(n_859),
.Y(n_1290)
);

BUFx6f_ASAP7_75t_L g1291 ( 
.A(n_1051),
.Y(n_1291)
);

BUFx6f_ASAP7_75t_L g1292 ( 
.A(n_1051),
.Y(n_1292)
);

AOI22xp5_ASAP7_75t_L g1293 ( 
.A1(n_1060),
.A2(n_956),
.B1(n_844),
.B2(n_816),
.Y(n_1293)
);

BUFx2_ASAP7_75t_L g1294 ( 
.A(n_1132),
.Y(n_1294)
);

BUFx3_ASAP7_75t_L g1295 ( 
.A(n_1182),
.Y(n_1295)
);

CKINVDCx5p33_ASAP7_75t_R g1296 ( 
.A(n_1181),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1204),
.Y(n_1297)
);

CKINVDCx5p33_ASAP7_75t_R g1298 ( 
.A(n_1123),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1201),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1201),
.Y(n_1300)
);

BUFx6f_ASAP7_75t_L g1301 ( 
.A(n_1167),
.Y(n_1301)
);

INVx2_ASAP7_75t_SL g1302 ( 
.A(n_1182),
.Y(n_1302)
);

AND2x4_ASAP7_75t_L g1303 ( 
.A(n_1050),
.B(n_844),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_L g1304 ( 
.A(n_1192),
.B(n_956),
.Y(n_1304)
);

CKINVDCx5p33_ASAP7_75t_R g1305 ( 
.A(n_1063),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_L g1306 ( 
.A(n_1157),
.B(n_1014),
.Y(n_1306)
);

HB1xp67_ASAP7_75t_L g1307 ( 
.A(n_1064),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1061),
.Y(n_1308)
);

INVx3_ASAP7_75t_SL g1309 ( 
.A(n_1184),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1075),
.Y(n_1310)
);

NOR3xp33_ASAP7_75t_SL g1311 ( 
.A(n_1199),
.B(n_1142),
.C(n_1073),
.Y(n_1311)
);

INVx2_ASAP7_75t_SL g1312 ( 
.A(n_1125),
.Y(n_1312)
);

OR2x2_ASAP7_75t_L g1313 ( 
.A(n_1053),
.B(n_1014),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_SL g1314 ( 
.A(n_1045),
.B(n_873),
.Y(n_1314)
);

BUFx6f_ASAP7_75t_L g1315 ( 
.A(n_1167),
.Y(n_1315)
);

OR2x2_ASAP7_75t_L g1316 ( 
.A(n_1086),
.B(n_1018),
.Y(n_1316)
);

INVx3_ASAP7_75t_L g1317 ( 
.A(n_1130),
.Y(n_1317)
);

INVx2_ASAP7_75t_SL g1318 ( 
.A(n_1099),
.Y(n_1318)
);

BUFx2_ASAP7_75t_L g1319 ( 
.A(n_1130),
.Y(n_1319)
);

NAND2xp5_ASAP7_75t_L g1320 ( 
.A(n_1218),
.B(n_1018),
.Y(n_1320)
);

AOI22xp5_ASAP7_75t_L g1321 ( 
.A1(n_1159),
.A2(n_1032),
.B1(n_1034),
.B2(n_1019),
.Y(n_1321)
);

BUFx6f_ASAP7_75t_L g1322 ( 
.A(n_1167),
.Y(n_1322)
);

INVx3_ASAP7_75t_L g1323 ( 
.A(n_1134),
.Y(n_1323)
);

NAND2x1p5_ASAP7_75t_L g1324 ( 
.A(n_1134),
.B(n_1207),
.Y(n_1324)
);

CKINVDCx5p33_ASAP7_75t_R g1325 ( 
.A(n_1179),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1205),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_L g1327 ( 
.A(n_1056),
.B(n_1032),
.Y(n_1327)
);

AND2x4_ASAP7_75t_L g1328 ( 
.A(n_1117),
.B(n_1035),
.Y(n_1328)
);

AND2x4_ASAP7_75t_L g1329 ( 
.A(n_1207),
.B(n_873),
.Y(n_1329)
);

BUFx2_ASAP7_75t_L g1330 ( 
.A(n_1068),
.Y(n_1330)
);

AND2x4_ASAP7_75t_SL g1331 ( 
.A(n_1079),
.B(n_895),
.Y(n_1331)
);

AND2x4_ASAP7_75t_L g1332 ( 
.A(n_1171),
.B(n_881),
.Y(n_1332)
);

NAND2x1p5_ASAP7_75t_L g1333 ( 
.A(n_1094),
.B(n_909),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1205),
.Y(n_1334)
);

AOI22xp33_ASAP7_75t_L g1335 ( 
.A1(n_1210),
.A2(n_1065),
.B1(n_1217),
.B2(n_1177),
.Y(n_1335)
);

NOR2x1p5_ASAP7_75t_L g1336 ( 
.A(n_1210),
.B(n_866),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1047),
.Y(n_1337)
);

INVx1_ASAP7_75t_SL g1338 ( 
.A(n_1047),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1049),
.Y(n_1339)
);

INVx1_ASAP7_75t_SL g1340 ( 
.A(n_1049),
.Y(n_1340)
);

AND2x2_ASAP7_75t_L g1341 ( 
.A(n_1095),
.B(n_867),
.Y(n_1341)
);

INVx2_ASAP7_75t_L g1342 ( 
.A(n_1096),
.Y(n_1342)
);

AND2x4_ASAP7_75t_L g1343 ( 
.A(n_1141),
.B(n_1206),
.Y(n_1343)
);

CKINVDCx16_ASAP7_75t_R g1344 ( 
.A(n_1080),
.Y(n_1344)
);

INVx4_ASAP7_75t_L g1345 ( 
.A(n_1198),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1101),
.Y(n_1346)
);

AND2x4_ASAP7_75t_L g1347 ( 
.A(n_1211),
.B(n_883),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_L g1348 ( 
.A(n_1058),
.B(n_910),
.Y(n_1348)
);

HB1xp67_ASAP7_75t_L g1349 ( 
.A(n_1103),
.Y(n_1349)
);

INVx2_ASAP7_75t_SL g1350 ( 
.A(n_1212),
.Y(n_1350)
);

NOR2xp33_ASAP7_75t_L g1351 ( 
.A(n_1115),
.B(n_886),
.Y(n_1351)
);

CKINVDCx5p33_ASAP7_75t_R g1352 ( 
.A(n_1196),
.Y(n_1352)
);

INVx2_ASAP7_75t_L g1353 ( 
.A(n_1118),
.Y(n_1353)
);

BUFx10_ASAP7_75t_L g1354 ( 
.A(n_1133),
.Y(n_1354)
);

INVx2_ASAP7_75t_L g1355 ( 
.A(n_1138),
.Y(n_1355)
);

BUFx3_ASAP7_75t_L g1356 ( 
.A(n_1216),
.Y(n_1356)
);

AOI22xp33_ASAP7_75t_L g1357 ( 
.A1(n_1107),
.A2(n_868),
.B1(n_858),
.B2(n_826),
.Y(n_1357)
);

HB1xp67_ASAP7_75t_L g1358 ( 
.A(n_1038),
.Y(n_1358)
);

AND2x6_ASAP7_75t_SL g1359 ( 
.A(n_1151),
.B(n_1200),
.Y(n_1359)
);

CKINVDCx5p33_ASAP7_75t_R g1360 ( 
.A(n_1202),
.Y(n_1360)
);

NAND2xp5_ASAP7_75t_L g1361 ( 
.A(n_1039),
.B(n_983),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1101),
.Y(n_1362)
);

AND2x2_ASAP7_75t_SL g1363 ( 
.A(n_1190),
.B(n_962),
.Y(n_1363)
);

OR2x2_ASAP7_75t_SL g1364 ( 
.A(n_1213),
.B(n_50),
.Y(n_1364)
);

BUFx6f_ASAP7_75t_L g1365 ( 
.A(n_1140),
.Y(n_1365)
);

BUFx6f_ASAP7_75t_L g1366 ( 
.A(n_1241),
.Y(n_1366)
);

AOI21xp5_ASAP7_75t_L g1367 ( 
.A1(n_1272),
.A2(n_1152),
.B(n_1169),
.Y(n_1367)
);

OAI21x1_ASAP7_75t_SL g1368 ( 
.A1(n_1256),
.A2(n_1209),
.B(n_1172),
.Y(n_1368)
);

AO31x2_ASAP7_75t_L g1369 ( 
.A1(n_1299),
.A2(n_1040),
.A3(n_1039),
.B(n_1168),
.Y(n_1369)
);

AO31x2_ASAP7_75t_L g1370 ( 
.A1(n_1300),
.A2(n_1040),
.A3(n_1221),
.B(n_1170),
.Y(n_1370)
);

AOI21xp5_ASAP7_75t_L g1371 ( 
.A1(n_1228),
.A2(n_1156),
.B(n_1163),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_L g1372 ( 
.A(n_1227),
.B(n_1213),
.Y(n_1372)
);

OAI21xp5_ASAP7_75t_L g1373 ( 
.A1(n_1254),
.A2(n_1340),
.B(n_1338),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_SL g1374 ( 
.A(n_1263),
.B(n_1102),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_L g1375 ( 
.A(n_1227),
.B(n_1214),
.Y(n_1375)
);

INVx2_ASAP7_75t_SL g1376 ( 
.A(n_1280),
.Y(n_1376)
);

AOI21xp5_ASAP7_75t_L g1377 ( 
.A1(n_1361),
.A2(n_1215),
.B(n_1214),
.Y(n_1377)
);

NAND2x1p5_ASAP7_75t_L g1378 ( 
.A(n_1256),
.B(n_1143),
.Y(n_1378)
);

OAI22xp5_ASAP7_75t_L g1379 ( 
.A1(n_1337),
.A2(n_1174),
.B1(n_1108),
.B2(n_1084),
.Y(n_1379)
);

HB1xp67_ASAP7_75t_L g1380 ( 
.A(n_1224),
.Y(n_1380)
);

AOI21xp5_ASAP7_75t_L g1381 ( 
.A1(n_1362),
.A2(n_1153),
.B(n_1092),
.Y(n_1381)
);

OR2x2_ASAP7_75t_L g1382 ( 
.A(n_1344),
.B(n_1093),
.Y(n_1382)
);

AO31x2_ASAP7_75t_L g1383 ( 
.A1(n_1326),
.A2(n_1139),
.A3(n_1173),
.B(n_1158),
.Y(n_1383)
);

AOI21x1_ASAP7_75t_L g1384 ( 
.A1(n_1287),
.A2(n_1104),
.B(n_1084),
.Y(n_1384)
);

OAI21x1_ASAP7_75t_L g1385 ( 
.A1(n_1304),
.A2(n_1195),
.B(n_1178),
.Y(n_1385)
);

OAI21xp5_ASAP7_75t_L g1386 ( 
.A1(n_1339),
.A2(n_1127),
.B(n_1052),
.Y(n_1386)
);

CKINVDCx6p67_ASAP7_75t_R g1387 ( 
.A(n_1225),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_L g1388 ( 
.A(n_1255),
.B(n_1111),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_L g1389 ( 
.A(n_1226),
.B(n_1119),
.Y(n_1389)
);

NAND2x1p5_ASAP7_75t_L g1390 ( 
.A(n_1280),
.B(n_1270),
.Y(n_1390)
);

OAI21x1_ASAP7_75t_L g1391 ( 
.A1(n_1362),
.A2(n_1104),
.B(n_1191),
.Y(n_1391)
);

OR2x2_ASAP7_75t_L g1392 ( 
.A(n_1222),
.B(n_1105),
.Y(n_1392)
);

NOR2x1_ASAP7_75t_L g1393 ( 
.A(n_1249),
.B(n_1187),
.Y(n_1393)
);

OAI21x1_ASAP7_75t_SL g1394 ( 
.A1(n_1346),
.A2(n_1161),
.B(n_1137),
.Y(n_1394)
);

OAI21xp5_ASAP7_75t_L g1395 ( 
.A1(n_1229),
.A2(n_1109),
.B(n_1059),
.Y(n_1395)
);

OAI21x1_ASAP7_75t_L g1396 ( 
.A1(n_1266),
.A2(n_1194),
.B(n_1193),
.Y(n_1396)
);

INVx3_ASAP7_75t_L g1397 ( 
.A(n_1249),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_L g1398 ( 
.A(n_1226),
.B(n_1110),
.Y(n_1398)
);

AOI21xp5_ASAP7_75t_L g1399 ( 
.A1(n_1334),
.A2(n_1327),
.B(n_1320),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1248),
.Y(n_1400)
);

AOI21xp5_ASAP7_75t_L g1401 ( 
.A1(n_1235),
.A2(n_1072),
.B(n_1070),
.Y(n_1401)
);

OAI21x1_ASAP7_75t_L g1402 ( 
.A1(n_1245),
.A2(n_1091),
.B(n_966),
.Y(n_1402)
);

OAI21xp5_ASAP7_75t_L g1403 ( 
.A1(n_1351),
.A2(n_1083),
.B(n_1082),
.Y(n_1403)
);

NAND3xp33_ASAP7_75t_L g1404 ( 
.A(n_1262),
.B(n_1121),
.C(n_1120),
.Y(n_1404)
);

OA22x2_ASAP7_75t_L g1405 ( 
.A1(n_1352),
.A2(n_1128),
.B1(n_1136),
.B2(n_1066),
.Y(n_1405)
);

BUFx10_ASAP7_75t_L g1406 ( 
.A(n_1239),
.Y(n_1406)
);

OA22x2_ASAP7_75t_L g1407 ( 
.A1(n_1264),
.A2(n_1148),
.B1(n_1146),
.B2(n_1081),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_L g1408 ( 
.A(n_1248),
.B(n_1145),
.Y(n_1408)
);

INVx1_ASAP7_75t_SL g1409 ( 
.A(n_1250),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1231),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_L g1411 ( 
.A(n_1360),
.B(n_1077),
.Y(n_1411)
);

AO31x2_ASAP7_75t_L g1412 ( 
.A1(n_1268),
.A2(n_960),
.A3(n_963),
.B(n_975),
.Y(n_1412)
);

AND2x2_ASAP7_75t_SL g1413 ( 
.A(n_1278),
.B(n_962),
.Y(n_1413)
);

NAND2xp5_ASAP7_75t_L g1414 ( 
.A(n_1233),
.B(n_980),
.Y(n_1414)
);

AO31x2_ASAP7_75t_L g1415 ( 
.A1(n_1268),
.A2(n_960),
.A3(n_963),
.B(n_976),
.Y(n_1415)
);

OAI21xp5_ASAP7_75t_L g1416 ( 
.A1(n_1348),
.A2(n_994),
.B(n_987),
.Y(n_1416)
);

A2O1A1Ixp33_ASAP7_75t_L g1417 ( 
.A1(n_1311),
.A2(n_981),
.B(n_944),
.C(n_990),
.Y(n_1417)
);

OAI21x1_ASAP7_75t_L g1418 ( 
.A1(n_1245),
.A2(n_966),
.B(n_961),
.Y(n_1418)
);

NAND2xp5_ASAP7_75t_L g1419 ( 
.A(n_1289),
.B(n_962),
.Y(n_1419)
);

AOI21xp5_ASAP7_75t_L g1420 ( 
.A1(n_1314),
.A2(n_984),
.B(n_982),
.Y(n_1420)
);

A2O1A1Ixp33_ASAP7_75t_L g1421 ( 
.A1(n_1336),
.A2(n_961),
.B(n_988),
.C(n_986),
.Y(n_1421)
);

BUFx6f_ASAP7_75t_L g1422 ( 
.A(n_1301),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1232),
.Y(n_1423)
);

INVx3_ASAP7_75t_L g1424 ( 
.A(n_1280),
.Y(n_1424)
);

AOI211x1_ASAP7_75t_L g1425 ( 
.A1(n_1279),
.A2(n_53),
.B(n_51),
.C(n_52),
.Y(n_1425)
);

AOI21xp33_ASAP7_75t_L g1426 ( 
.A1(n_1335),
.A2(n_993),
.B(n_964),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1244),
.Y(n_1427)
);

AOI21xp5_ASAP7_75t_L g1428 ( 
.A1(n_1290),
.A2(n_964),
.B(n_945),
.Y(n_1428)
);

NAND2xp5_ASAP7_75t_L g1429 ( 
.A(n_1358),
.B(n_962),
.Y(n_1429)
);

OAI21x1_ASAP7_75t_L g1430 ( 
.A1(n_1246),
.A2(n_964),
.B(n_945),
.Y(n_1430)
);

AOI21xp5_ASAP7_75t_L g1431 ( 
.A1(n_1306),
.A2(n_945),
.B(n_123),
.Y(n_1431)
);

OAI21x1_ASAP7_75t_L g1432 ( 
.A1(n_1246),
.A2(n_124),
.B(n_121),
.Y(n_1432)
);

OAI21xp5_ASAP7_75t_L g1433 ( 
.A1(n_1242),
.A2(n_54),
.B(n_55),
.Y(n_1433)
);

AOI21x1_ASAP7_75t_L g1434 ( 
.A1(n_1303),
.A2(n_127),
.B(n_125),
.Y(n_1434)
);

AOI21x1_ASAP7_75t_SL g1435 ( 
.A1(n_1332),
.A2(n_54),
.B(n_55),
.Y(n_1435)
);

OAI22xp5_ASAP7_75t_L g1436 ( 
.A1(n_1278),
.A2(n_59),
.B1(n_56),
.B2(n_58),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_L g1437 ( 
.A(n_1251),
.B(n_56),
.Y(n_1437)
);

AOI21xp5_ASAP7_75t_L g1438 ( 
.A1(n_1357),
.A2(n_1310),
.B(n_1308),
.Y(n_1438)
);

NOR2xp33_ASAP7_75t_SL g1439 ( 
.A(n_1285),
.B(n_58),
.Y(n_1439)
);

AND2x4_ASAP7_75t_L g1440 ( 
.A(n_1239),
.B(n_1223),
.Y(n_1440)
);

AOI21xp5_ASAP7_75t_L g1441 ( 
.A1(n_1308),
.A2(n_131),
.B(n_128),
.Y(n_1441)
);

OAI21x1_ASAP7_75t_L g1442 ( 
.A1(n_1317),
.A2(n_135),
.B(n_133),
.Y(n_1442)
);

OAI21x1_ASAP7_75t_L g1443 ( 
.A1(n_1317),
.A2(n_137),
.B(n_136),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_L g1444 ( 
.A(n_1252),
.B(n_59),
.Y(n_1444)
);

NAND3xp33_ASAP7_75t_L g1445 ( 
.A(n_1267),
.B(n_61),
.C(n_62),
.Y(n_1445)
);

OAI22xp5_ASAP7_75t_L g1446 ( 
.A1(n_1298),
.A2(n_64),
.B1(n_62),
.B2(n_63),
.Y(n_1446)
);

OAI21x1_ASAP7_75t_L g1447 ( 
.A1(n_1323),
.A2(n_139),
.B(n_138),
.Y(n_1447)
);

NOR4xp25_ASAP7_75t_L g1448 ( 
.A(n_1286),
.B(n_67),
.C(n_63),
.D(n_65),
.Y(n_1448)
);

AOI211x1_ASAP7_75t_L g1449 ( 
.A1(n_1341),
.A2(n_68),
.B(n_65),
.C(n_67),
.Y(n_1449)
);

BUFx12f_ASAP7_75t_L g1450 ( 
.A(n_1281),
.Y(n_1450)
);

AO21x1_ASAP7_75t_L g1451 ( 
.A1(n_1345),
.A2(n_68),
.B(n_69),
.Y(n_1451)
);

AOI21xp5_ASAP7_75t_L g1452 ( 
.A1(n_1310),
.A2(n_146),
.B(n_141),
.Y(n_1452)
);

OAI21x1_ASAP7_75t_L g1453 ( 
.A1(n_1323),
.A2(n_152),
.B(n_151),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_L g1454 ( 
.A(n_1276),
.B(n_69),
.Y(n_1454)
);

INVx2_ASAP7_75t_L g1455 ( 
.A(n_1400),
.Y(n_1455)
);

NAND2xp5_ASAP7_75t_L g1456 ( 
.A(n_1388),
.B(n_1305),
.Y(n_1456)
);

AOI21xp33_ASAP7_75t_SL g1457 ( 
.A1(n_1390),
.A2(n_1296),
.B(n_1277),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1410),
.Y(n_1458)
);

AOI21xp33_ASAP7_75t_L g1459 ( 
.A1(n_1405),
.A2(n_1282),
.B(n_1363),
.Y(n_1459)
);

AND2x4_ASAP7_75t_L g1460 ( 
.A(n_1422),
.B(n_1345),
.Y(n_1460)
);

NOR2xp33_ASAP7_75t_L g1461 ( 
.A(n_1382),
.B(n_1237),
.Y(n_1461)
);

OAI22xp5_ASAP7_75t_L g1462 ( 
.A1(n_1372),
.A2(n_1364),
.B1(n_1307),
.B2(n_1238),
.Y(n_1462)
);

AOI21xp5_ASAP7_75t_L g1463 ( 
.A1(n_1377),
.A2(n_1315),
.B(n_1301),
.Y(n_1463)
);

OAI21x1_ASAP7_75t_L g1464 ( 
.A1(n_1430),
.A2(n_1324),
.B(n_1333),
.Y(n_1464)
);

O2A1O1Ixp33_ASAP7_75t_SL g1465 ( 
.A1(n_1375),
.A2(n_1293),
.B(n_1316),
.C(n_1313),
.Y(n_1465)
);

OAI21x1_ASAP7_75t_L g1466 ( 
.A1(n_1385),
.A2(n_1297),
.B(n_1288),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1423),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1427),
.Y(n_1468)
);

BUFx2_ASAP7_75t_SL g1469 ( 
.A(n_1366),
.Y(n_1469)
);

INVx5_ASAP7_75t_L g1470 ( 
.A(n_1422),
.Y(n_1470)
);

AOI22xp33_ASAP7_75t_L g1471 ( 
.A1(n_1393),
.A2(n_1332),
.B1(n_1260),
.B2(n_1261),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1454),
.Y(n_1472)
);

OAI21x1_ASAP7_75t_L g1473 ( 
.A1(n_1428),
.A2(n_1271),
.B(n_1257),
.Y(n_1473)
);

OAI21x1_ASAP7_75t_L g1474 ( 
.A1(n_1391),
.A2(n_1283),
.B(n_1274),
.Y(n_1474)
);

OAI21x1_ASAP7_75t_L g1475 ( 
.A1(n_1396),
.A2(n_1353),
.B(n_1342),
.Y(n_1475)
);

NAND3xp33_ASAP7_75t_SL g1476 ( 
.A(n_1439),
.B(n_1230),
.C(n_1236),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1437),
.Y(n_1477)
);

AND2x2_ASAP7_75t_L g1478 ( 
.A(n_1440),
.B(n_1243),
.Y(n_1478)
);

OAI22xp33_ASAP7_75t_L g1479 ( 
.A1(n_1436),
.A2(n_1433),
.B1(n_1373),
.B2(n_1445),
.Y(n_1479)
);

AOI21x1_ASAP7_75t_L g1480 ( 
.A1(n_1384),
.A2(n_1303),
.B(n_1319),
.Y(n_1480)
);

AOI21xp5_ASAP7_75t_L g1481 ( 
.A1(n_1367),
.A2(n_1315),
.B(n_1301),
.Y(n_1481)
);

AO21x2_ASAP7_75t_L g1482 ( 
.A1(n_1438),
.A2(n_1321),
.B(n_1259),
.Y(n_1482)
);

AND2x4_ASAP7_75t_L g1483 ( 
.A(n_1422),
.B(n_1315),
.Y(n_1483)
);

AOI21xp5_ASAP7_75t_L g1484 ( 
.A1(n_1371),
.A2(n_1322),
.B(n_1291),
.Y(n_1484)
);

OAI21xp5_ASAP7_75t_L g1485 ( 
.A1(n_1401),
.A2(n_1273),
.B(n_1330),
.Y(n_1485)
);

OAI21x1_ASAP7_75t_L g1486 ( 
.A1(n_1402),
.A2(n_1355),
.B(n_1322),
.Y(n_1486)
);

INVx2_ASAP7_75t_L g1487 ( 
.A(n_1369),
.Y(n_1487)
);

BUFx2_ASAP7_75t_L g1488 ( 
.A(n_1440),
.Y(n_1488)
);

OAI21x1_ASAP7_75t_L g1489 ( 
.A1(n_1432),
.A2(n_1322),
.B(n_1291),
.Y(n_1489)
);

INVx2_ASAP7_75t_L g1490 ( 
.A(n_1369),
.Y(n_1490)
);

NAND2x1p5_ASAP7_75t_L g1491 ( 
.A(n_1413),
.B(n_1295),
.Y(n_1491)
);

NOR2xp33_ASAP7_75t_L g1492 ( 
.A(n_1389),
.B(n_1359),
.Y(n_1492)
);

AO21x2_ASAP7_75t_L g1493 ( 
.A1(n_1368),
.A2(n_1394),
.B(n_1451),
.Y(n_1493)
);

INVx1_ASAP7_75t_SL g1494 ( 
.A(n_1409),
.Y(n_1494)
);

AO31x2_ASAP7_75t_L g1495 ( 
.A1(n_1399),
.A2(n_1294),
.A3(n_1253),
.B(n_1291),
.Y(n_1495)
);

INVx2_ASAP7_75t_L g1496 ( 
.A(n_1369),
.Y(n_1496)
);

AOI22xp33_ASAP7_75t_L g1497 ( 
.A1(n_1379),
.A2(n_1343),
.B1(n_1349),
.B2(n_1328),
.Y(n_1497)
);

AND2x4_ASAP7_75t_L g1498 ( 
.A(n_1383),
.B(n_1265),
.Y(n_1498)
);

AO31x2_ASAP7_75t_L g1499 ( 
.A1(n_1381),
.A2(n_1292),
.A3(n_1265),
.B(n_1365),
.Y(n_1499)
);

AOI22xp33_ASAP7_75t_L g1500 ( 
.A1(n_1462),
.A2(n_1446),
.B1(n_1380),
.B2(n_1397),
.Y(n_1500)
);

OAI22xp5_ASAP7_75t_L g1501 ( 
.A1(n_1497),
.A2(n_1425),
.B1(n_1449),
.B2(n_1376),
.Y(n_1501)
);

AOI22xp33_ASAP7_75t_L g1502 ( 
.A1(n_1492),
.A2(n_1395),
.B1(n_1386),
.B2(n_1403),
.Y(n_1502)
);

AOI221xp5_ASAP7_75t_L g1503 ( 
.A1(n_1492),
.A2(n_1448),
.B1(n_1398),
.B2(n_1325),
.C(n_1408),
.Y(n_1503)
);

NAND2xp5_ASAP7_75t_SL g1504 ( 
.A(n_1479),
.B(n_1424),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1458),
.Y(n_1505)
);

NAND2xp5_ASAP7_75t_L g1506 ( 
.A(n_1467),
.B(n_1392),
.Y(n_1506)
);

OAI21x1_ASAP7_75t_L g1507 ( 
.A1(n_1489),
.A2(n_1435),
.B(n_1442),
.Y(n_1507)
);

BUFx4f_ASAP7_75t_L g1508 ( 
.A(n_1491),
.Y(n_1508)
);

BUFx6f_ASAP7_75t_L g1509 ( 
.A(n_1470),
.Y(n_1509)
);

BUFx12f_ASAP7_75t_L g1510 ( 
.A(n_1491),
.Y(n_1510)
);

INVx4_ASAP7_75t_L g1511 ( 
.A(n_1470),
.Y(n_1511)
);

NAND2xp33_ASAP7_75t_SL g1512 ( 
.A(n_1471),
.B(n_1247),
.Y(n_1512)
);

AOI22xp33_ASAP7_75t_L g1513 ( 
.A1(n_1497),
.A2(n_1374),
.B1(n_1407),
.B2(n_1444),
.Y(n_1513)
);

CKINVDCx20_ASAP7_75t_R g1514 ( 
.A(n_1469),
.Y(n_1514)
);

INVx2_ASAP7_75t_L g1515 ( 
.A(n_1487),
.Y(n_1515)
);

AND2x2_ASAP7_75t_L g1516 ( 
.A(n_1478),
.B(n_1406),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1468),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1455),
.Y(n_1518)
);

HB1xp67_ASAP7_75t_L g1519 ( 
.A(n_1455),
.Y(n_1519)
);

AOI22xp33_ASAP7_75t_SL g1520 ( 
.A1(n_1488),
.A2(n_1258),
.B1(n_1378),
.B2(n_1429),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1472),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1466),
.Y(n_1522)
);

AOI22xp33_ASAP7_75t_L g1523 ( 
.A1(n_1461),
.A2(n_1404),
.B1(n_1343),
.B2(n_1416),
.Y(n_1523)
);

CKINVDCx20_ASAP7_75t_R g1524 ( 
.A(n_1476),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_L g1525 ( 
.A(n_1461),
.B(n_1411),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1466),
.Y(n_1526)
);

AND2x2_ASAP7_75t_L g1527 ( 
.A(n_1456),
.B(n_70),
.Y(n_1527)
);

INVx4_ASAP7_75t_L g1528 ( 
.A(n_1470),
.Y(n_1528)
);

A2O1A1Ixp33_ASAP7_75t_L g1529 ( 
.A1(n_1485),
.A2(n_1447),
.B(n_1453),
.C(n_1443),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1477),
.Y(n_1530)
);

AOI22xp33_ASAP7_75t_SL g1531 ( 
.A1(n_1510),
.A2(n_1493),
.B1(n_1498),
.B2(n_1490),
.Y(n_1531)
);

AOI22xp33_ASAP7_75t_SL g1532 ( 
.A1(n_1510),
.A2(n_1508),
.B1(n_1524),
.B2(n_1511),
.Y(n_1532)
);

AOI221xp5_ASAP7_75t_L g1533 ( 
.A1(n_1502),
.A2(n_1459),
.B1(n_1479),
.B2(n_1494),
.C(n_1471),
.Y(n_1533)
);

AOI22xp33_ASAP7_75t_L g1534 ( 
.A1(n_1512),
.A2(n_1493),
.B1(n_1482),
.B2(n_1490),
.Y(n_1534)
);

AOI22xp5_ASAP7_75t_L g1535 ( 
.A1(n_1512),
.A2(n_1482),
.B1(n_1328),
.B2(n_1269),
.Y(n_1535)
);

OAI33xp33_ASAP7_75t_L g1536 ( 
.A1(n_1525),
.A2(n_1414),
.A3(n_1419),
.B1(n_1275),
.B2(n_1487),
.B3(n_1496),
.Y(n_1536)
);

AOI22xp33_ASAP7_75t_L g1537 ( 
.A1(n_1500),
.A2(n_1496),
.B1(n_1498),
.B2(n_1312),
.Y(n_1537)
);

AND2x2_ASAP7_75t_L g1538 ( 
.A(n_1521),
.B(n_1495),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1505),
.Y(n_1539)
);

AOI22xp33_ASAP7_75t_L g1540 ( 
.A1(n_1500),
.A2(n_1498),
.B1(n_1460),
.B2(n_1331),
.Y(n_1540)
);

AOI22xp33_ASAP7_75t_SL g1541 ( 
.A1(n_1508),
.A2(n_1460),
.B1(n_1470),
.B2(n_1464),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1517),
.Y(n_1542)
);

AOI22xp33_ASAP7_75t_L g1543 ( 
.A1(n_1502),
.A2(n_1460),
.B1(n_1354),
.B2(n_1309),
.Y(n_1543)
);

AOI22xp33_ASAP7_75t_L g1544 ( 
.A1(n_1513),
.A2(n_1503),
.B1(n_1504),
.B2(n_1527),
.Y(n_1544)
);

AOI22xp33_ASAP7_75t_SL g1545 ( 
.A1(n_1511),
.A2(n_1483),
.B1(n_1366),
.B2(n_1450),
.Y(n_1545)
);

INVxp67_ASAP7_75t_L g1546 ( 
.A(n_1519),
.Y(n_1546)
);

AOI211xp5_ASAP7_75t_SL g1547 ( 
.A1(n_1514),
.A2(n_1501),
.B(n_1465),
.C(n_1529),
.Y(n_1547)
);

AOI22xp33_ASAP7_75t_L g1548 ( 
.A1(n_1513),
.A2(n_1354),
.B1(n_1473),
.B2(n_1463),
.Y(n_1548)
);

CKINVDCx20_ASAP7_75t_R g1549 ( 
.A(n_1516),
.Y(n_1549)
);

AOI22xp33_ASAP7_75t_SL g1550 ( 
.A1(n_1528),
.A2(n_1483),
.B1(n_1234),
.B2(n_1474),
.Y(n_1550)
);

BUFx4f_ASAP7_75t_SL g1551 ( 
.A(n_1528),
.Y(n_1551)
);

INVxp67_ASAP7_75t_L g1552 ( 
.A(n_1530),
.Y(n_1552)
);

AOI22xp33_ASAP7_75t_L g1553 ( 
.A1(n_1504),
.A2(n_1523),
.B1(n_1506),
.B2(n_1520),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1518),
.Y(n_1554)
);

OR2x2_ASAP7_75t_L g1555 ( 
.A(n_1515),
.B(n_1495),
.Y(n_1555)
);

CKINVDCx5p33_ASAP7_75t_R g1556 ( 
.A(n_1509),
.Y(n_1556)
);

NOR2xp33_ASAP7_75t_L g1557 ( 
.A(n_1523),
.B(n_1465),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1538),
.B(n_1515),
.Y(n_1558)
);

INVxp33_ASAP7_75t_SL g1559 ( 
.A(n_1532),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_L g1560 ( 
.A(n_1554),
.B(n_1495),
.Y(n_1560)
);

AND2x2_ASAP7_75t_L g1561 ( 
.A(n_1555),
.B(n_1539),
.Y(n_1561)
);

INVx2_ASAP7_75t_L g1562 ( 
.A(n_1542),
.Y(n_1562)
);

INVxp67_ASAP7_75t_SL g1563 ( 
.A(n_1546),
.Y(n_1563)
);

INVx2_ASAP7_75t_L g1564 ( 
.A(n_1552),
.Y(n_1564)
);

INVx3_ASAP7_75t_L g1565 ( 
.A(n_1551),
.Y(n_1565)
);

OAI221xp5_ASAP7_75t_L g1566 ( 
.A1(n_1544),
.A2(n_1529),
.B1(n_1240),
.B2(n_1302),
.C(n_1318),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1531),
.Y(n_1567)
);

HB1xp67_ASAP7_75t_L g1568 ( 
.A(n_1556),
.Y(n_1568)
);

AND2x2_ASAP7_75t_L g1569 ( 
.A(n_1534),
.B(n_1522),
.Y(n_1569)
);

AOI22xp33_ASAP7_75t_L g1570 ( 
.A1(n_1557),
.A2(n_1509),
.B1(n_1526),
.B2(n_1426),
.Y(n_1570)
);

INVx4_ASAP7_75t_R g1571 ( 
.A(n_1541),
.Y(n_1571)
);

AND2x2_ASAP7_75t_L g1572 ( 
.A(n_1557),
.B(n_1495),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1550),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1535),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1537),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1548),
.Y(n_1576)
);

INVxp67_ASAP7_75t_L g1577 ( 
.A(n_1536),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1533),
.B(n_1480),
.Y(n_1578)
);

INVxp67_ASAP7_75t_L g1579 ( 
.A(n_1568),
.Y(n_1579)
);

AOI221xp5_ASAP7_75t_L g1580 ( 
.A1(n_1577),
.A2(n_1553),
.B1(n_1543),
.B2(n_1540),
.C(n_1457),
.Y(n_1580)
);

AOI22xp33_ASAP7_75t_L g1581 ( 
.A1(n_1559),
.A2(n_1549),
.B1(n_1545),
.B2(n_1509),
.Y(n_1581)
);

AOI33xp33_ASAP7_75t_L g1582 ( 
.A1(n_1567),
.A2(n_1547),
.A3(n_1350),
.B1(n_1347),
.B2(n_1549),
.B3(n_73),
.Y(n_1582)
);

AO21x2_ASAP7_75t_L g1583 ( 
.A1(n_1567),
.A2(n_1507),
.B(n_1481),
.Y(n_1583)
);

OAI22xp5_ASAP7_75t_L g1584 ( 
.A1(n_1566),
.A2(n_1509),
.B1(n_1387),
.B2(n_1483),
.Y(n_1584)
);

NOR3xp33_ASAP7_75t_SL g1585 ( 
.A(n_1566),
.B(n_1417),
.C(n_1441),
.Y(n_1585)
);

NOR2xp33_ASAP7_75t_R g1586 ( 
.A(n_1565),
.B(n_70),
.Y(n_1586)
);

INVx2_ASAP7_75t_SL g1587 ( 
.A(n_1565),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1562),
.Y(n_1588)
);

NAND3xp33_ASAP7_75t_L g1589 ( 
.A(n_1573),
.B(n_1484),
.C(n_1452),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1562),
.Y(n_1590)
);

OR2x2_ASAP7_75t_L g1591 ( 
.A(n_1561),
.B(n_1499),
.Y(n_1591)
);

OAI22xp5_ASAP7_75t_L g1592 ( 
.A1(n_1565),
.A2(n_1434),
.B1(n_1284),
.B2(n_1356),
.Y(n_1592)
);

INVx4_ASAP7_75t_L g1593 ( 
.A(n_1587),
.Y(n_1593)
);

AND2x2_ASAP7_75t_L g1594 ( 
.A(n_1591),
.B(n_1572),
.Y(n_1594)
);

INVx2_ASAP7_75t_L g1595 ( 
.A(n_1588),
.Y(n_1595)
);

OR2x2_ASAP7_75t_L g1596 ( 
.A(n_1590),
.B(n_1561),
.Y(n_1596)
);

NOR2x1_ASAP7_75t_L g1597 ( 
.A(n_1584),
.B(n_1565),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1579),
.B(n_1572),
.Y(n_1598)
);

OR2x2_ASAP7_75t_L g1599 ( 
.A(n_1583),
.B(n_1564),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1583),
.Y(n_1600)
);

AND2x2_ASAP7_75t_L g1601 ( 
.A(n_1581),
.B(n_1563),
.Y(n_1601)
);

AND2x2_ASAP7_75t_L g1602 ( 
.A(n_1580),
.B(n_1573),
.Y(n_1602)
);

AND2x2_ASAP7_75t_L g1603 ( 
.A(n_1586),
.B(n_1558),
.Y(n_1603)
);

INVxp67_ASAP7_75t_L g1604 ( 
.A(n_1589),
.Y(n_1604)
);

AND2x2_ASAP7_75t_L g1605 ( 
.A(n_1582),
.B(n_1558),
.Y(n_1605)
);

BUFx2_ASAP7_75t_L g1606 ( 
.A(n_1592),
.Y(n_1606)
);

OR2x2_ASAP7_75t_L g1607 ( 
.A(n_1592),
.B(n_1564),
.Y(n_1607)
);

AND2x2_ASAP7_75t_L g1608 ( 
.A(n_1585),
.B(n_1564),
.Y(n_1608)
);

OR2x2_ASAP7_75t_L g1609 ( 
.A(n_1596),
.B(n_1576),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1598),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_L g1611 ( 
.A(n_1605),
.B(n_1578),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1594),
.B(n_1576),
.Y(n_1612)
);

INVx2_ASAP7_75t_L g1613 ( 
.A(n_1595),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1598),
.Y(n_1614)
);

OR2x2_ASAP7_75t_L g1615 ( 
.A(n_1611),
.B(n_1609),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_L g1616 ( 
.A(n_1612),
.B(n_1602),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1610),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_1612),
.B(n_1602),
.Y(n_1618)
);

AOI31xp33_ASAP7_75t_L g1619 ( 
.A1(n_1616),
.A2(n_1597),
.A3(n_1604),
.B(n_1601),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1617),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1620),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1619),
.Y(n_1622)
);

NAND4xp25_ASAP7_75t_L g1623 ( 
.A(n_1620),
.B(n_1618),
.C(n_1606),
.D(n_1605),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1622),
.B(n_1615),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1621),
.Y(n_1625)
);

O2A1O1Ixp33_ASAP7_75t_L g1626 ( 
.A1(n_1623),
.A2(n_1608),
.B(n_1603),
.C(n_1600),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_L g1627 ( 
.A(n_1622),
.B(n_1614),
.Y(n_1627)
);

AND2x2_ASAP7_75t_SL g1628 ( 
.A(n_1622),
.B(n_1593),
.Y(n_1628)
);

INVx1_ASAP7_75t_SL g1629 ( 
.A(n_1621),
.Y(n_1629)
);

NAND4xp25_ASAP7_75t_L g1630 ( 
.A(n_1627),
.B(n_1593),
.C(n_1570),
.D(n_1575),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_L g1631 ( 
.A(n_1629),
.B(n_1626),
.Y(n_1631)
);

INVx5_ASAP7_75t_L g1632 ( 
.A(n_1628),
.Y(n_1632)
);

NAND3xp33_ASAP7_75t_L g1633 ( 
.A(n_1625),
.B(n_1593),
.C(n_1284),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1629),
.Y(n_1634)
);

NAND2x1_ASAP7_75t_SL g1635 ( 
.A(n_1624),
.B(n_1613),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_L g1636 ( 
.A(n_1624),
.B(n_1613),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_L g1637 ( 
.A(n_1624),
.B(n_1599),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1627),
.Y(n_1638)
);

NOR2x1_ASAP7_75t_L g1639 ( 
.A(n_1629),
.B(n_1607),
.Y(n_1639)
);

CKINVDCx6p67_ASAP7_75t_R g1640 ( 
.A(n_1632),
.Y(n_1640)
);

NAND3xp33_ASAP7_75t_SL g1641 ( 
.A(n_1634),
.B(n_1578),
.C(n_1575),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1636),
.Y(n_1642)
);

AOI21xp5_ASAP7_75t_L g1643 ( 
.A1(n_1631),
.A2(n_1595),
.B(n_1574),
.Y(n_1643)
);

AOI221xp5_ASAP7_75t_L g1644 ( 
.A1(n_1638),
.A2(n_1574),
.B1(n_1562),
.B2(n_1569),
.C(n_1560),
.Y(n_1644)
);

OR3x1_ASAP7_75t_L g1645 ( 
.A(n_1630),
.B(n_1571),
.C(n_71),
.Y(n_1645)
);

AOI221xp5_ASAP7_75t_L g1646 ( 
.A1(n_1633),
.A2(n_1569),
.B1(n_1560),
.B2(n_1329),
.C(n_1431),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1637),
.Y(n_1647)
);

AOI221x1_ASAP7_75t_L g1648 ( 
.A1(n_1632),
.A2(n_1421),
.B1(n_1329),
.B2(n_1347),
.C(n_1420),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_L g1649 ( 
.A(n_1635),
.B(n_80),
.Y(n_1649)
);

A2O1A1Ixp33_ASAP7_75t_L g1650 ( 
.A1(n_1639),
.A2(n_1486),
.B(n_1475),
.C(n_83),
.Y(n_1650)
);

NAND4xp25_ASAP7_75t_L g1651 ( 
.A(n_1631),
.B(n_81),
.C(n_82),
.D(n_83),
.Y(n_1651)
);

AND2x4_ASAP7_75t_L g1652 ( 
.A(n_1632),
.B(n_82),
.Y(n_1652)
);

AOI22xp5_ASAP7_75t_L g1653 ( 
.A1(n_1645),
.A2(n_1265),
.B1(n_1292),
.B2(n_1365),
.Y(n_1653)
);

OAI221xp5_ASAP7_75t_L g1654 ( 
.A1(n_1651),
.A2(n_87),
.B1(n_88),
.B2(n_90),
.C(n_91),
.Y(n_1654)
);

INVx2_ASAP7_75t_L g1655 ( 
.A(n_1652),
.Y(n_1655)
);

AOI32xp33_ASAP7_75t_L g1656 ( 
.A1(n_1642),
.A2(n_87),
.A3(n_90),
.B1(n_92),
.B2(n_93),
.Y(n_1656)
);

NOR2x1_ASAP7_75t_L g1657 ( 
.A(n_1647),
.B(n_94),
.Y(n_1657)
);

AND2x4_ASAP7_75t_L g1658 ( 
.A(n_1643),
.B(n_95),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_L g1659 ( 
.A(n_1648),
.B(n_96),
.Y(n_1659)
);

AND2x2_ASAP7_75t_L g1660 ( 
.A(n_1644),
.B(n_97),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_L g1661 ( 
.A(n_1650),
.B(n_97),
.Y(n_1661)
);

NOR2x1_ASAP7_75t_L g1662 ( 
.A(n_1641),
.B(n_98),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1646),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1649),
.Y(n_1664)
);

AOI22xp33_ASAP7_75t_L g1665 ( 
.A1(n_1640),
.A2(n_1365),
.B1(n_1292),
.B2(n_1418),
.Y(n_1665)
);

OR2x2_ASAP7_75t_L g1666 ( 
.A(n_1655),
.B(n_99),
.Y(n_1666)
);

OAI221xp5_ASAP7_75t_L g1667 ( 
.A1(n_1654),
.A2(n_100),
.B1(n_102),
.B2(n_103),
.C(n_104),
.Y(n_1667)
);

NOR2x1_ASAP7_75t_L g1668 ( 
.A(n_1657),
.B(n_100),
.Y(n_1668)
);

AO21x1_ASAP7_75t_L g1669 ( 
.A1(n_1664),
.A2(n_1658),
.B(n_1663),
.Y(n_1669)
);

NOR2x1p5_ASAP7_75t_L g1670 ( 
.A(n_1659),
.B(n_102),
.Y(n_1670)
);

NAND4xp75_ASAP7_75t_L g1671 ( 
.A(n_1662),
.B(n_103),
.C(n_104),
.D(n_105),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1661),
.Y(n_1672)
);

NAND3xp33_ASAP7_75t_SL g1673 ( 
.A(n_1656),
.B(n_106),
.C(n_153),
.Y(n_1673)
);

AOI211xp5_ASAP7_75t_L g1674 ( 
.A1(n_1660),
.A2(n_154),
.B(n_155),
.C(n_156),
.Y(n_1674)
);

AND3x4_ASAP7_75t_L g1675 ( 
.A(n_1665),
.B(n_1370),
.C(n_158),
.Y(n_1675)
);

NAND2x1p5_ASAP7_75t_L g1676 ( 
.A(n_1653),
.B(n_159),
.Y(n_1676)
);

AND4x1_ASAP7_75t_L g1677 ( 
.A(n_1674),
.B(n_167),
.C(n_168),
.D(n_172),
.Y(n_1677)
);

INVx3_ASAP7_75t_L g1678 ( 
.A(n_1666),
.Y(n_1678)
);

INVx2_ASAP7_75t_L g1679 ( 
.A(n_1676),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1671),
.Y(n_1680)
);

NOR3xp33_ASAP7_75t_L g1681 ( 
.A(n_1667),
.B(n_173),
.C(n_174),
.Y(n_1681)
);

XNOR2x1_ASAP7_75t_L g1682 ( 
.A(n_1670),
.B(n_175),
.Y(n_1682)
);

CKINVDCx16_ASAP7_75t_R g1683 ( 
.A(n_1673),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1682),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_L g1685 ( 
.A(n_1683),
.B(n_1668),
.Y(n_1685)
);

AO22x1_ASAP7_75t_L g1686 ( 
.A1(n_1681),
.A2(n_1672),
.B1(n_1675),
.B2(n_1669),
.Y(n_1686)
);

INVx1_ASAP7_75t_SL g1687 ( 
.A(n_1679),
.Y(n_1687)
);

AND2x2_ASAP7_75t_L g1688 ( 
.A(n_1678),
.B(n_1383),
.Y(n_1688)
);

XNOR2xp5_ASAP7_75t_L g1689 ( 
.A(n_1677),
.B(n_179),
.Y(n_1689)
);

XNOR2x1_ASAP7_75t_L g1690 ( 
.A(n_1689),
.B(n_1680),
.Y(n_1690)
);

BUFx24_ASAP7_75t_SL g1691 ( 
.A(n_1687),
.Y(n_1691)
);

NOR2x1_ASAP7_75t_L g1692 ( 
.A(n_1685),
.B(n_1684),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1688),
.Y(n_1693)
);

CKINVDCx20_ASAP7_75t_R g1694 ( 
.A(n_1691),
.Y(n_1694)
);

XNOR2xp5_ASAP7_75t_L g1695 ( 
.A(n_1690),
.B(n_1686),
.Y(n_1695)
);

CKINVDCx20_ASAP7_75t_R g1696 ( 
.A(n_1694),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1696),
.Y(n_1697)
);

AOI22xp33_ASAP7_75t_L g1698 ( 
.A1(n_1697),
.A2(n_1692),
.B1(n_1693),
.B2(n_1695),
.Y(n_1698)
);

AOI322xp5_ASAP7_75t_L g1699 ( 
.A1(n_1698),
.A2(n_1415),
.A3(n_1412),
.B1(n_1499),
.B2(n_186),
.C1(n_187),
.C2(n_188),
.Y(n_1699)
);

AOI322xp5_ASAP7_75t_L g1700 ( 
.A1(n_1698),
.A2(n_1412),
.A3(n_182),
.B1(n_185),
.B2(n_191),
.C1(n_197),
.C2(n_200),
.Y(n_1700)
);

AOI221xp5_ASAP7_75t_L g1701 ( 
.A1(n_1700),
.A2(n_210),
.B1(n_213),
.B2(n_214),
.C(n_217),
.Y(n_1701)
);

AOI211xp5_ASAP7_75t_L g1702 ( 
.A1(n_1701),
.A2(n_1699),
.B(n_219),
.C(n_222),
.Y(n_1702)
);


endmodule