module real_aes_4585_n_77 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_77);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_77;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_522;
wire n_485;
wire n_222;
wire n_287;
wire n_357;
wire n_503;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_580;
wire n_577;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_560;
wire n_260;
wire n_594;
wire n_97;
wire n_186;
wire n_138;
wire n_379;
wire n_374;
wire n_453;
wire n_235;
wire n_399;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_92;
wire n_519;
wire n_564;
wire n_573;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_570;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_231;
wire n_102;
wire n_547;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_582;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_93;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_323;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_368;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_250;
wire n_85;
wire n_605;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_87;
wire n_171;
wire n_78;
wire n_531;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_557;
wire n_488;
wire n_501;
wire n_251;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_589;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_526;
wire n_155;
wire n_243;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_446;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_266;
wire n_183;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_440;
wire n_525;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_566;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_597;
wire n_340;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_206;
wire n_307;
wire n_500;
wire n_601;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_91;
NAND2xp5_ASAP7_75t_L g291 ( .A(n_0), .B(n_271), .Y(n_291) );
CKINVDCx5p33_ASAP7_75t_R g307 ( .A(n_1), .Y(n_307) );
HB1xp67_ASAP7_75t_L g88 ( .A(n_2), .Y(n_88) );
HB1xp67_ASAP7_75t_L g87 ( .A(n_3), .Y(n_87) );
O2A1O1Ixp33_ASAP7_75t_SL g343 ( .A1(n_4), .A2(n_215), .B(n_344), .C(n_345), .Y(n_343) );
OAI22xp33_ASAP7_75t_L g296 ( .A1(n_5), .A2(n_62), .B1(n_214), .B2(n_243), .Y(n_296) );
AOI22xp33_ASAP7_75t_L g133 ( .A1(n_6), .A2(n_74), .B1(n_134), .B2(n_138), .Y(n_133) );
CKINVDCx5p33_ASAP7_75t_R g322 ( .A(n_7), .Y(n_322) );
OAI22xp5_ASAP7_75t_L g240 ( .A1(n_8), .A2(n_53), .B1(n_241), .B2(n_243), .Y(n_240) );
CKINVDCx5p33_ASAP7_75t_R g262 ( .A(n_9), .Y(n_262) );
INVx1_ASAP7_75t_L g121 ( .A(n_10), .Y(n_121) );
INVxp67_ASAP7_75t_L g162 ( .A(n_10), .Y(n_162) );
NOR2xp33_ASAP7_75t_L g173 ( .A(n_10), .B(n_55), .Y(n_173) );
AOI22xp5_ASAP7_75t_L g238 ( .A1(n_11), .A2(n_44), .B1(n_214), .B2(n_239), .Y(n_238) );
AOI22xp33_ASAP7_75t_L g177 ( .A1(n_12), .A2(n_34), .B1(n_178), .B2(n_179), .Y(n_177) );
OA21x2_ASAP7_75t_L g228 ( .A1(n_13), .A2(n_52), .B(n_229), .Y(n_228) );
OA21x2_ASAP7_75t_L g233 ( .A1(n_13), .A2(n_52), .B(n_229), .Y(n_233) );
NAND2xp5_ASAP7_75t_SL g117 ( .A(n_14), .B(n_105), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g317 ( .A(n_15), .Y(n_317) );
BUFx3_ASAP7_75t_L g186 ( .A(n_16), .Y(n_186) );
O2A1O1Ixp33_ASAP7_75t_L g349 ( .A1(n_17), .A2(n_297), .B(n_350), .C(n_351), .Y(n_349) );
OAI22xp33_ASAP7_75t_SL g294 ( .A1(n_18), .A2(n_32), .B1(n_214), .B2(n_261), .Y(n_294) );
AOI22xp33_ASAP7_75t_L g281 ( .A1(n_19), .A2(n_25), .B1(n_261), .B2(n_266), .Y(n_281) );
AOI22xp33_ASAP7_75t_L g153 ( .A1(n_20), .A2(n_26), .B1(n_154), .B2(n_155), .Y(n_153) );
BUFx6f_ASAP7_75t_L g105 ( .A(n_21), .Y(n_105) );
O2A1O1Ixp5_ASAP7_75t_L g209 ( .A1(n_22), .A2(n_210), .B(n_213), .C(n_215), .Y(n_209) );
AOI22xp33_ASAP7_75t_L g139 ( .A1(n_23), .A2(n_31), .B1(n_140), .B2(n_141), .Y(n_139) );
INVx1_ASAP7_75t_L g106 ( .A(n_24), .Y(n_106) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_24), .B(n_54), .Y(n_159) );
CKINVDCx5p33_ASAP7_75t_R g95 ( .A(n_27), .Y(n_95) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_28), .B(n_287), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_29), .B(n_151), .Y(n_150) );
CKINVDCx5p33_ASAP7_75t_R g347 ( .A(n_30), .Y(n_347) );
INVx1_ASAP7_75t_L g229 ( .A(n_33), .Y(n_229) );
HB1xp67_ASAP7_75t_L g197 ( .A(n_35), .Y(n_197) );
AND2x4_ASAP7_75t_L g225 ( .A(n_35), .B(n_195), .Y(n_225) );
AND2x4_ASAP7_75t_L g246 ( .A(n_35), .B(n_195), .Y(n_246) );
BUFx6f_ASAP7_75t_L g216 ( .A(n_36), .Y(n_216) );
CKINVDCx5p33_ASAP7_75t_R g305 ( .A(n_37), .Y(n_305) );
CKINVDCx5p33_ASAP7_75t_R g222 ( .A(n_38), .Y(n_222) );
INVx2_ASAP7_75t_L g267 ( .A(n_39), .Y(n_267) );
O2A1O1Ixp33_ASAP7_75t_L g319 ( .A1(n_40), .A2(n_215), .B(n_320), .C(n_321), .Y(n_319) );
CKINVDCx5p33_ASAP7_75t_R g304 ( .A(n_41), .Y(n_304) );
XNOR2xp5_ASAP7_75t_L g607 ( .A(n_42), .B(n_96), .Y(n_607) );
AOI22xp33_ASAP7_75t_L g99 ( .A1(n_43), .A2(n_67), .B1(n_100), .B2(n_124), .Y(n_99) );
AOI22xp5_ASAP7_75t_L g282 ( .A1(n_45), .A2(n_58), .B1(n_283), .B2(n_284), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_46), .B(n_247), .Y(n_309) );
OA22x2_ASAP7_75t_L g111 ( .A1(n_47), .A2(n_55), .B1(n_105), .B2(n_109), .Y(n_111) );
INVx1_ASAP7_75t_L g129 ( .A(n_47), .Y(n_129) );
CKINVDCx5p33_ASAP7_75t_R g80 ( .A(n_48), .Y(n_80) );
INVx1_ASAP7_75t_L g167 ( .A(n_49), .Y(n_167) );
CKINVDCx5p33_ASAP7_75t_R g308 ( .A(n_50), .Y(n_308) );
NAND2xp33_ASAP7_75t_R g248 ( .A(n_51), .B(n_233), .Y(n_248) );
AOI22xp33_ASAP7_75t_L g509 ( .A1(n_51), .A2(n_76), .B1(n_287), .B2(n_510), .Y(n_509) );
INVx1_ASAP7_75t_L g123 ( .A(n_54), .Y(n_123) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_54), .B(n_127), .Y(n_176) );
HB1xp67_ASAP7_75t_L g189 ( .A(n_54), .Y(n_189) );
OAI21xp33_ASAP7_75t_L g130 ( .A1(n_55), .A2(n_60), .B(n_131), .Y(n_130) );
CKINVDCx5p33_ASAP7_75t_R g265 ( .A(n_56), .Y(n_265) );
CKINVDCx5p33_ASAP7_75t_R g263 ( .A(n_57), .Y(n_263) );
HB1xp67_ASAP7_75t_L g84 ( .A(n_59), .Y(n_84) );
INVx1_ASAP7_75t_L g108 ( .A(n_60), .Y(n_108) );
NOR2xp33_ASAP7_75t_L g174 ( .A(n_60), .B(n_71), .Y(n_174) );
AOI22xp33_ASAP7_75t_L g142 ( .A1(n_61), .A2(n_69), .B1(n_143), .B2(n_146), .Y(n_142) );
BUFx6f_ASAP7_75t_L g212 ( .A(n_63), .Y(n_212) );
BUFx5_ASAP7_75t_L g214 ( .A(n_63), .Y(n_214) );
INVx1_ASAP7_75t_L g242 ( .A(n_63), .Y(n_242) );
INVx2_ASAP7_75t_L g355 ( .A(n_64), .Y(n_355) );
INVx2_ASAP7_75t_L g324 ( .A(n_65), .Y(n_324) );
CKINVDCx5p33_ASAP7_75t_R g352 ( .A(n_66), .Y(n_352) );
INVx2_ASAP7_75t_SL g195 ( .A(n_68), .Y(n_195) );
INVx1_ASAP7_75t_L g220 ( .A(n_70), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g115 ( .A(n_71), .B(n_116), .Y(n_115) );
AOI21xp33_ASAP7_75t_L g163 ( .A1(n_72), .A2(n_164), .B(n_166), .Y(n_163) );
INVx2_ASAP7_75t_L g231 ( .A(n_73), .Y(n_231) );
OAI21xp33_ASAP7_75t_SL g315 ( .A1(n_75), .A2(n_214), .B(n_316), .Y(n_315) );
INVxp67_ASAP7_75t_SL g269 ( .A(n_76), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_76), .B(n_287), .Y(n_378) );
AOI221xp5_ASAP7_75t_L g77 ( .A1(n_78), .A2(n_181), .B1(n_198), .B2(n_594), .C(n_600), .Y(n_77) );
XNOR2xp5_ASAP7_75t_L g78 ( .A(n_79), .B(n_92), .Y(n_78) );
OAI22xp5_ASAP7_75t_L g79 ( .A1(n_80), .A2(n_81), .B1(n_82), .B2(n_91), .Y(n_79) );
CKINVDCx5p33_ASAP7_75t_R g91 ( .A(n_80), .Y(n_91) );
CKINVDCx20_ASAP7_75t_R g81 ( .A(n_82), .Y(n_81) );
AOI22xp5_ASAP7_75t_L g82 ( .A1(n_83), .A2(n_84), .B1(n_85), .B2(n_86), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_84), .Y(n_83) );
INVx1_ASAP7_75t_L g85 ( .A(n_86), .Y(n_85) );
OAI22xp5_ASAP7_75t_L g86 ( .A1(n_87), .A2(n_88), .B1(n_89), .B2(n_90), .Y(n_86) );
INVx1_ASAP7_75t_L g90 ( .A(n_87), .Y(n_90) );
INVx1_ASAP7_75t_L g89 ( .A(n_88), .Y(n_89) );
AOI22xp5_ASAP7_75t_L g92 ( .A1(n_93), .A2(n_94), .B1(n_96), .B2(n_180), .Y(n_92) );
CKINVDCx5p33_ASAP7_75t_R g93 ( .A(n_94), .Y(n_93) );
HB1xp67_ASAP7_75t_L g94 ( .A(n_95), .Y(n_94) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_95), .B(n_214), .Y(n_213) );
INVx1_ASAP7_75t_L g180 ( .A(n_96), .Y(n_180) );
AOI22xp5_ASAP7_75t_SL g601 ( .A1(n_96), .A2(n_180), .B1(n_602), .B2(n_603), .Y(n_601) );
HB1xp67_ASAP7_75t_L g96 ( .A(n_97), .Y(n_96) );
NOR2xp67_ASAP7_75t_L g97 ( .A(n_98), .B(n_149), .Y(n_97) );
NAND4xp25_ASAP7_75t_L g98 ( .A(n_99), .B(n_133), .C(n_139), .D(n_142), .Y(n_98) );
AND2x4_ASAP7_75t_L g100 ( .A(n_101), .B(n_112), .Y(n_100) );
AND2x4_ASAP7_75t_L g140 ( .A(n_101), .B(n_136), .Y(n_140) );
AND2x4_ASAP7_75t_L g143 ( .A(n_101), .B(n_144), .Y(n_143) );
AND2x4_ASAP7_75t_L g146 ( .A(n_101), .B(n_147), .Y(n_146) );
AND2x4_ASAP7_75t_L g101 ( .A(n_102), .B(n_110), .Y(n_101) );
AND2x2_ASAP7_75t_L g165 ( .A(n_102), .B(n_111), .Y(n_165) );
INVx1_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
AND2x2_ASAP7_75t_L g135 ( .A(n_103), .B(n_111), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g103 ( .A(n_104), .B(n_107), .Y(n_103) );
NAND2xp33_ASAP7_75t_L g104 ( .A(n_105), .B(n_106), .Y(n_104) );
INVx2_ASAP7_75t_L g109 ( .A(n_105), .Y(n_109) );
INVx3_ASAP7_75t_L g116 ( .A(n_105), .Y(n_116) );
NAND2xp33_ASAP7_75t_L g122 ( .A(n_105), .B(n_123), .Y(n_122) );
INVx1_ASAP7_75t_L g131 ( .A(n_105), .Y(n_131) );
HB1xp67_ASAP7_75t_L g158 ( .A(n_105), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g128 ( .A(n_106), .B(n_129), .Y(n_128) );
INVxp67_ASAP7_75t_L g190 ( .A(n_106), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g107 ( .A(n_108), .B(n_109), .Y(n_107) );
OAI21xp5_ASAP7_75t_L g161 ( .A1(n_108), .A2(n_131), .B(n_162), .Y(n_161) );
INVx1_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
AND2x2_ASAP7_75t_L g160 ( .A(n_111), .B(n_161), .Y(n_160) );
INVx2_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
INVx2_ASAP7_75t_L g132 ( .A(n_113), .Y(n_132) );
OR2x2_ASAP7_75t_L g113 ( .A(n_114), .B(n_118), .Y(n_113) );
AND2x4_ASAP7_75t_L g136 ( .A(n_114), .B(n_137), .Y(n_136) );
AND2x4_ASAP7_75t_L g144 ( .A(n_114), .B(n_145), .Y(n_144) );
INVx2_ASAP7_75t_L g148 ( .A(n_114), .Y(n_148) );
AND2x2_ASAP7_75t_L g156 ( .A(n_114), .B(n_157), .Y(n_156) );
AND2x4_ASAP7_75t_L g114 ( .A(n_115), .B(n_117), .Y(n_114) );
NAND2xp5_ASAP7_75t_L g120 ( .A(n_116), .B(n_121), .Y(n_120) );
INVxp67_ASAP7_75t_L g127 ( .A(n_116), .Y(n_127) );
NAND3xp33_ASAP7_75t_L g175 ( .A(n_117), .B(n_126), .C(n_176), .Y(n_175) );
INVx1_ASAP7_75t_L g137 ( .A(n_118), .Y(n_137) );
INVx1_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVx1_ASAP7_75t_L g145 ( .A(n_119), .Y(n_145) );
AND2x2_ASAP7_75t_L g119 ( .A(n_120), .B(n_122), .Y(n_119) );
AND2x4_ASAP7_75t_L g124 ( .A(n_125), .B(n_132), .Y(n_124) );
AND2x4_ASAP7_75t_L g141 ( .A(n_125), .B(n_136), .Y(n_141) );
AND2x4_ASAP7_75t_L g179 ( .A(n_125), .B(n_147), .Y(n_179) );
AND2x2_ASAP7_75t_L g125 ( .A(n_126), .B(n_130), .Y(n_125) );
NAND2xp5_ASAP7_75t_L g126 ( .A(n_127), .B(n_128), .Y(n_126) );
HB1xp67_ASAP7_75t_L g191 ( .A(n_129), .Y(n_191) );
AND2x4_ASAP7_75t_L g138 ( .A(n_132), .B(n_135), .Y(n_138) );
AND2x4_ASAP7_75t_L g134 ( .A(n_135), .B(n_136), .Y(n_134) );
AND2x2_ASAP7_75t_L g152 ( .A(n_135), .B(n_147), .Y(n_152) );
AND2x4_ASAP7_75t_L g154 ( .A(n_135), .B(n_144), .Y(n_154) );
AND2x4_ASAP7_75t_L g164 ( .A(n_144), .B(n_165), .Y(n_164) );
AND2x4_ASAP7_75t_L g147 ( .A(n_145), .B(n_148), .Y(n_147) );
AND2x2_ASAP7_75t_L g178 ( .A(n_147), .B(n_165), .Y(n_178) );
NAND4xp25_ASAP7_75t_L g149 ( .A(n_150), .B(n_153), .C(n_163), .D(n_177), .Y(n_149) );
BUFx3_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
AND2x2_ASAP7_75t_L g155 ( .A(n_156), .B(n_160), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_158), .B(n_159), .Y(n_157) );
INVx1_ASAP7_75t_L g171 ( .A(n_158), .Y(n_171) );
HB1xp67_ASAP7_75t_L g187 ( .A(n_159), .Y(n_187) );
NOR2xp33_ASAP7_75t_L g166 ( .A(n_167), .B(n_168), .Y(n_166) );
INVx3_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
INVx3_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
AO21x2_ASAP7_75t_L g170 ( .A1(n_171), .A2(n_172), .B(n_175), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_173), .B(n_174), .Y(n_172) );
BUFx2_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
CKINVDCx5p33_ASAP7_75t_R g182 ( .A(n_183), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_184), .B(n_192), .Y(n_183) );
INVxp67_ASAP7_75t_SL g184 ( .A(n_185), .Y(n_184) );
AND2x2_ASAP7_75t_L g605 ( .A(n_185), .B(n_192), .Y(n_605) );
AOI211xp5_ASAP7_75t_L g185 ( .A1(n_186), .A2(n_187), .B(n_188), .C(n_191), .Y(n_185) );
NOR2xp33_ASAP7_75t_L g188 ( .A(n_189), .B(n_190), .Y(n_188) );
NOR2xp33_ASAP7_75t_L g192 ( .A(n_193), .B(n_196), .Y(n_192) );
OR2x2_ASAP7_75t_L g609 ( .A(n_193), .B(n_197), .Y(n_609) );
INVx1_ASAP7_75t_L g612 ( .A(n_193), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_193), .B(n_196), .Y(n_613) );
HB1xp67_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
HB1xp67_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
INVx1_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
INVx1_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
AND4x2_ASAP7_75t_L g201 ( .A(n_202), .B(n_452), .C(n_492), .D(n_561), .Y(n_201) );
NOR2x1_ASAP7_75t_L g202 ( .A(n_203), .B(n_390), .Y(n_202) );
NAND2xp5_ASAP7_75t_SL g203 ( .A(n_204), .B(n_370), .Y(n_203) );
O2A1O1Ixp33_ASAP7_75t_L g204 ( .A1(n_205), .A2(n_249), .B(n_273), .C(n_325), .Y(n_204) );
AND2x2_ASAP7_75t_L g384 ( .A(n_205), .B(n_385), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_205), .B(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g438 ( .A(n_205), .Y(n_438) );
AND2x2_ASAP7_75t_L g458 ( .A(n_205), .B(n_327), .Y(n_458) );
AND2x2_ASAP7_75t_L g560 ( .A(n_205), .B(n_541), .Y(n_560) );
AND2x4_ASAP7_75t_L g205 ( .A(n_206), .B(n_234), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_206), .B(n_377), .Y(n_376) );
OR2x2_ASAP7_75t_L g586 ( .A(n_206), .B(n_525), .Y(n_586) );
INVx2_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
AND2x2_ASAP7_75t_L g357 ( .A(n_207), .B(n_358), .Y(n_357) );
INVx2_ASAP7_75t_L g364 ( .A(n_207), .Y(n_364) );
BUFx2_ASAP7_75t_R g424 ( .A(n_207), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_207), .B(n_341), .Y(n_533) );
AND2x2_ASAP7_75t_L g537 ( .A(n_207), .B(n_340), .Y(n_537) );
AO21x2_ASAP7_75t_L g207 ( .A1(n_208), .A2(n_226), .B(n_230), .Y(n_207) );
NOR3xp33_ASAP7_75t_L g208 ( .A(n_209), .B(n_217), .C(n_224), .Y(n_208) );
INVx1_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
INVx1_ASAP7_75t_L g218 ( .A(n_211), .Y(n_218) );
INVx1_ASAP7_75t_L g320 ( .A(n_211), .Y(n_320) );
INVx3_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
INVx2_ASAP7_75t_L g239 ( .A(n_212), .Y(n_239) );
INVx2_ASAP7_75t_L g243 ( .A(n_212), .Y(n_243) );
INVx6_ASAP7_75t_L g261 ( .A(n_212), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_214), .B(n_222), .Y(n_221) );
AOI22xp5_ASAP7_75t_L g260 ( .A1(n_214), .A2(n_261), .B1(n_262), .B2(n_263), .Y(n_260) );
AOI22xp33_ASAP7_75t_SL g303 ( .A1(n_214), .A2(n_261), .B1(n_304), .B2(n_305), .Y(n_303) );
AOI22xp33_ASAP7_75t_L g306 ( .A1(n_214), .A2(n_239), .B1(n_307), .B2(n_308), .Y(n_306) );
NAND2xp5_ASAP7_75t_SL g316 ( .A(n_214), .B(n_317), .Y(n_316) );
AOI22xp5_ASAP7_75t_L g237 ( .A1(n_215), .A2(n_223), .B1(n_238), .B2(n_240), .Y(n_237) );
OAI22xp33_ASAP7_75t_L g259 ( .A1(n_215), .A2(n_223), .B1(n_260), .B2(n_264), .Y(n_259) );
OAI221xp5_ASAP7_75t_L g302 ( .A1(n_215), .A2(n_246), .B1(n_297), .B2(n_303), .C(n_306), .Y(n_302) );
INVx1_ASAP7_75t_L g383 ( .A(n_215), .Y(n_383) );
BUFx6f_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_216), .B(n_220), .Y(n_219) );
INVx4_ASAP7_75t_L g223 ( .A(n_216), .Y(n_223) );
BUFx6f_ASAP7_75t_L g280 ( .A(n_216), .Y(n_280) );
INVx1_ASAP7_75t_L g285 ( .A(n_216), .Y(n_285) );
NAND2xp5_ASAP7_75t_SL g293 ( .A(n_216), .B(n_294), .Y(n_293) );
INVx3_ASAP7_75t_L g297 ( .A(n_216), .Y(n_297) );
OAI22xp5_ASAP7_75t_L g217 ( .A1(n_218), .A2(n_219), .B1(n_221), .B2(n_223), .Y(n_217) );
INVx2_ASAP7_75t_L g318 ( .A(n_223), .Y(n_318) );
NOR2xp33_ASAP7_75t_SL g353 ( .A(n_224), .B(n_271), .Y(n_353) );
AOI221xp5_ASAP7_75t_L g380 ( .A1(n_224), .A2(n_318), .B1(n_381), .B2(n_382), .C(n_383), .Y(n_380) );
INVx4_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_225), .B(n_257), .Y(n_278) );
AND2x2_ASAP7_75t_L g312 ( .A(n_225), .B(n_313), .Y(n_312) );
NAND2xp5_ASAP7_75t_SL g379 ( .A(n_226), .B(n_380), .Y(n_379) );
BUFx3_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
INVx3_ASAP7_75t_L g247 ( .A(n_227), .Y(n_247) );
NOR2xp33_ASAP7_75t_L g323 ( .A(n_227), .B(n_324), .Y(n_323) );
INVx2_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
INVx4_ASAP7_75t_L g272 ( .A(n_228), .Y(n_272) );
BUFx3_ASAP7_75t_L g334 ( .A(n_228), .Y(n_334) );
NOR2xp33_ASAP7_75t_L g230 ( .A(n_231), .B(n_232), .Y(n_230) );
INVx1_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
BUFx3_ASAP7_75t_L g258 ( .A(n_233), .Y(n_258) );
INVx1_ASAP7_75t_L g313 ( .A(n_233), .Y(n_313) );
INVx2_ASAP7_75t_L g511 ( .A(n_233), .Y(n_511) );
INVx1_ASAP7_75t_SL g251 ( .A(n_234), .Y(n_251) );
INVx1_ASAP7_75t_L g365 ( .A(n_234), .Y(n_365) );
AND2x2_ASAP7_75t_L g447 ( .A(n_234), .B(n_340), .Y(n_447) );
INVx2_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
INVx1_ASAP7_75t_L g358 ( .A(n_235), .Y(n_358) );
HB1xp67_ASAP7_75t_L g374 ( .A(n_235), .Y(n_374) );
AND2x2_ASAP7_75t_L g462 ( .A(n_235), .B(n_364), .Y(n_462) );
AND2x2_ASAP7_75t_L g534 ( .A(n_235), .B(n_254), .Y(n_534) );
AND2x2_ASAP7_75t_L g235 ( .A(n_236), .B(n_248), .Y(n_235) );
AND2x2_ASAP7_75t_L g508 ( .A(n_236), .B(n_509), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_237), .B(n_244), .Y(n_236) );
AOI22xp5_ASAP7_75t_L g264 ( .A1(n_239), .A2(n_265), .B1(n_266), .B2(n_267), .Y(n_264) );
INVx1_ASAP7_75t_L g350 ( .A(n_239), .Y(n_350) );
INVx2_ASAP7_75t_L g283 ( .A(n_241), .Y(n_283) );
INVx2_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
INVx2_ASAP7_75t_L g266 ( .A(n_242), .Y(n_266) );
NOR2xp67_ASAP7_75t_L g244 ( .A(n_245), .B(n_247), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
BUFx6f_ASAP7_75t_L g256 ( .A(n_246), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_246), .B(n_272), .Y(n_298) );
INVxp67_ASAP7_75t_SL g249 ( .A(n_250), .Y(n_249) );
OR2x2_ASAP7_75t_L g250 ( .A(n_251), .B(n_252), .Y(n_250) );
NOR2xp33_ASAP7_75t_L g583 ( .A(n_252), .B(n_356), .Y(n_583) );
INVx2_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
AND2x4_ASAP7_75t_L g449 ( .A(n_254), .B(n_341), .Y(n_449) );
OAI21x1_ASAP7_75t_L g254 ( .A1(n_255), .A2(n_259), .B(n_268), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_256), .B(n_257), .Y(n_255) );
AND2x2_ASAP7_75t_L g595 ( .A(n_256), .B(n_596), .Y(n_595) );
INVx1_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
INVx1_ASAP7_75t_L g381 ( .A(n_260), .Y(n_381) );
INVx2_ASAP7_75t_SL g284 ( .A(n_261), .Y(n_284) );
INVx2_ASAP7_75t_L g346 ( .A(n_261), .Y(n_346) );
INVx1_ASAP7_75t_L g615 ( .A(n_262), .Y(n_615) );
INVx1_ASAP7_75t_L g382 ( .A(n_264), .Y(n_382) );
NAND2xp5_ASAP7_75t_SL g321 ( .A(n_266), .B(n_322), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_266), .B(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g602 ( .A(n_267), .Y(n_602) );
OR2x2_ASAP7_75t_L g268 ( .A(n_269), .B(n_270), .Y(n_268) );
INVx2_ASAP7_75t_L g301 ( .A(n_270), .Y(n_301) );
INVx2_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
INVx2_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
INVx2_ASAP7_75t_L g287 ( .A(n_272), .Y(n_287) );
NOR2xp33_ASAP7_75t_SL g354 ( .A(n_272), .B(n_355), .Y(n_354) );
INVxp67_ASAP7_75t_SL g273 ( .A(n_274), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_275), .B(n_288), .Y(n_274) );
AND2x4_ASAP7_75t_L g367 ( .A(n_275), .B(n_368), .Y(n_367) );
INVx2_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
AND2x2_ASAP7_75t_L g451 ( .A(n_276), .B(n_420), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_276), .B(n_445), .Y(n_464) );
OR2x2_ASAP7_75t_L g568 ( .A(n_276), .B(n_524), .Y(n_568) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
INVx2_ASAP7_75t_L g404 ( .A(n_277), .Y(n_404) );
OAI21x1_ASAP7_75t_L g277 ( .A1(n_278), .A2(n_279), .B(n_286), .Y(n_277) );
INVx1_ASAP7_75t_L g332 ( .A(n_279), .Y(n_332) );
OA22x2_ASAP7_75t_L g279 ( .A1(n_280), .A2(n_281), .B1(n_282), .B2(n_285), .Y(n_279) );
INVx4_ASAP7_75t_L g598 ( .A(n_280), .Y(n_598) );
INVx1_ASAP7_75t_L g344 ( .A(n_283), .Y(n_344) );
INVx1_ASAP7_75t_L g335 ( .A(n_286), .Y(n_335) );
BUFx2_ASAP7_75t_SL g432 ( .A(n_288), .Y(n_432) );
NOR2xp67_ASAP7_75t_L g288 ( .A(n_289), .B(n_299), .Y(n_288) );
INVx1_ASAP7_75t_L g387 ( .A(n_289), .Y(n_387) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
INVx2_ASAP7_75t_L g369 ( .A(n_290), .Y(n_369) );
INVx3_ASAP7_75t_L g406 ( .A(n_290), .Y(n_406) );
AND2x2_ASAP7_75t_L g441 ( .A(n_290), .B(n_407), .Y(n_441) );
AND2x2_ASAP7_75t_L g471 ( .A(n_290), .B(n_310), .Y(n_471) );
AND2x4_ASAP7_75t_L g290 ( .A(n_291), .B(n_292), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_293), .B(n_295), .Y(n_292) );
AOI21xp5_ASAP7_75t_L g295 ( .A1(n_296), .A2(n_297), .B(n_298), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_300), .B(n_310), .Y(n_299) );
INVx2_ASAP7_75t_L g336 ( .A(n_300), .Y(n_336) );
INVx2_ASAP7_75t_L g389 ( .A(n_300), .Y(n_389) );
OA21x2_ASAP7_75t_L g300 ( .A1(n_301), .A2(n_302), .B(n_309), .Y(n_300) );
OA21x2_ASAP7_75t_L g407 ( .A1(n_301), .A2(n_302), .B(n_309), .Y(n_407) );
INVx1_ASAP7_75t_L g328 ( .A(n_310), .Y(n_328) );
AND2x2_ASAP7_75t_L g388 ( .A(n_310), .B(n_389), .Y(n_388) );
OR2x2_ASAP7_75t_L g414 ( .A(n_310), .B(n_369), .Y(n_414) );
INVx2_ASAP7_75t_L g420 ( .A(n_310), .Y(n_420) );
AND2x2_ASAP7_75t_L g445 ( .A(n_310), .B(n_406), .Y(n_445) );
BUFx2_ASAP7_75t_L g514 ( .A(n_310), .Y(n_514) );
INVx2_ASAP7_75t_L g525 ( .A(n_310), .Y(n_525) );
INVx3_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
AOI21x1_ASAP7_75t_L g311 ( .A1(n_312), .A2(n_314), .B(n_323), .Y(n_311) );
AOI21xp5_ASAP7_75t_L g314 ( .A1(n_315), .A2(n_318), .B(n_319), .Y(n_314) );
OAI22xp5_ASAP7_75t_L g325 ( .A1(n_326), .A2(n_337), .B1(n_359), .B2(n_366), .Y(n_325) );
OR2x2_ASAP7_75t_L g326 ( .A(n_327), .B(n_329), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
INVx2_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
AND2x2_ASAP7_75t_L g426 ( .A(n_330), .B(n_419), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_330), .B(n_471), .Y(n_470) );
INVx2_ASAP7_75t_SL g520 ( .A(n_330), .Y(n_520) );
AND2x4_ASAP7_75t_L g330 ( .A(n_331), .B(n_336), .Y(n_330) );
OR2x2_ASAP7_75t_L g412 ( .A(n_331), .B(n_407), .Y(n_412) );
AOI21xp5_ASAP7_75t_L g331 ( .A1(n_332), .A2(n_333), .B(n_335), .Y(n_331) );
INVx3_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
AND2x4_ASAP7_75t_L g368 ( .A(n_336), .B(n_369), .Y(n_368) );
NAND3xp33_ASAP7_75t_L g392 ( .A(n_337), .B(n_393), .C(n_397), .Y(n_392) );
OR2x2_ASAP7_75t_L g337 ( .A(n_338), .B(n_356), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
OR2x2_ASAP7_75t_L g375 ( .A(n_339), .B(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
INVx2_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
AND2x2_ASAP7_75t_L g385 ( .A(n_341), .B(n_377), .Y(n_385) );
INVx1_ASAP7_75t_L g396 ( .A(n_341), .Y(n_396) );
HB1xp67_ASAP7_75t_L g400 ( .A(n_341), .Y(n_400) );
OR2x2_ASAP7_75t_L g429 ( .A(n_341), .B(n_377), .Y(n_429) );
INVx1_ASAP7_75t_L g466 ( .A(n_341), .Y(n_466) );
HB1xp67_ASAP7_75t_L g588 ( .A(n_341), .Y(n_588) );
AO31x2_ASAP7_75t_L g341 ( .A1(n_342), .A2(n_348), .A3(n_353), .B(n_354), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_346), .B(n_347), .Y(n_345) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
HB1xp67_ASAP7_75t_L g599 ( .A(n_350), .Y(n_599) );
OR2x2_ASAP7_75t_L g415 ( .A(n_356), .B(n_416), .Y(n_415) );
INVx2_ASAP7_75t_SL g356 ( .A(n_357), .Y(n_356) );
AND2x4_ASAP7_75t_L g427 ( .A(n_357), .B(n_428), .Y(n_427) );
AND2x2_ASAP7_75t_L g436 ( .A(n_357), .B(n_385), .Y(n_436) );
AND2x4_ASAP7_75t_L g472 ( .A(n_357), .B(n_449), .Y(n_472) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
BUFx2_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
OR2x2_ASAP7_75t_L g517 ( .A(n_362), .B(n_400), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_363), .B(n_365), .Y(n_362) );
NOR2xp33_ASAP7_75t_L g557 ( .A(n_363), .B(n_377), .Y(n_557) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
HB1xp67_ASAP7_75t_L g491 ( .A(n_364), .Y(n_491) );
AND2x2_ASAP7_75t_L g542 ( .A(n_364), .B(n_507), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_366), .B(n_470), .Y(n_469) );
INVx2_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
AND2x2_ASAP7_75t_L g549 ( .A(n_367), .B(n_502), .Y(n_549) );
NAND2x1p5_ASAP7_75t_L g513 ( .A(n_368), .B(n_514), .Y(n_513) );
NAND2x1p5_ASAP7_75t_L g559 ( .A(n_368), .B(n_554), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_368), .B(n_451), .Y(n_572) );
AND2x2_ASAP7_75t_L g434 ( .A(n_369), .B(n_404), .Y(n_434) );
OAI21xp5_ASAP7_75t_L g370 ( .A1(n_371), .A2(n_384), .B(n_386), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
OR2x2_ASAP7_75t_L g372 ( .A(n_373), .B(n_375), .Y(n_372) );
AND2x2_ASAP7_75t_L g394 ( .A(n_373), .B(n_395), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_373), .B(n_449), .Y(n_448) );
OR2x2_ASAP7_75t_L g475 ( .A(n_373), .B(n_476), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_373), .B(n_528), .Y(n_527) );
INVx2_ASAP7_75t_SL g373 ( .A(n_374), .Y(n_373) );
INVx2_ASAP7_75t_L g521 ( .A(n_375), .Y(n_521) );
INVx1_ASAP7_75t_L g592 ( .A(n_376), .Y(n_592) );
AND2x2_ASAP7_75t_L g395 ( .A(n_377), .B(n_396), .Y(n_395) );
HB1xp67_ASAP7_75t_L g481 ( .A(n_377), .Y(n_481) );
AND2x2_ASAP7_75t_L g377 ( .A(n_378), .B(n_379), .Y(n_377) );
AND2x2_ASAP7_75t_L g507 ( .A(n_379), .B(n_508), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_385), .B(n_424), .Y(n_423) );
BUFx6f_ASAP7_75t_L g528 ( .A(n_385), .Y(n_528) );
AOI22xp5_ASAP7_75t_SL g467 ( .A1(n_386), .A2(n_468), .B1(n_469), .B2(n_472), .Y(n_467) );
AND2x4_ASAP7_75t_L g386 ( .A(n_387), .B(n_388), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_391), .B(n_425), .Y(n_390) );
AOI21xp5_ASAP7_75t_L g391 ( .A1(n_392), .A2(n_401), .B(n_408), .Y(n_391) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g439 ( .A(n_395), .Y(n_439) );
OR2x2_ASAP7_75t_L g505 ( .A(n_396), .B(n_506), .Y(n_505) );
AND2x2_ASAP7_75t_L g577 ( .A(n_396), .B(n_534), .Y(n_577) );
INVxp67_ASAP7_75t_SL g468 ( .A(n_397), .Y(n_468) );
BUFx3_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVxp67_ASAP7_75t_L g416 ( .A(n_399), .Y(n_416) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
AND2x2_ASAP7_75t_L g401 ( .A(n_402), .B(n_405), .Y(n_401) );
A2O1A1Ixp33_ASAP7_75t_L g473 ( .A1(n_402), .A2(n_471), .B(n_474), .C(n_477), .Y(n_473) );
OR2x2_ASAP7_75t_L g546 ( .A(n_402), .B(n_414), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_402), .B(n_405), .Y(n_580) );
AND2x2_ASAP7_75t_L g593 ( .A(n_402), .B(n_441), .Y(n_593) );
INVx3_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
AND2x4_ASAP7_75t_L g501 ( .A(n_403), .B(n_405), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_403), .B(n_441), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_403), .B(n_445), .Y(n_564) );
AND2x2_ASAP7_75t_L g569 ( .A(n_403), .B(n_471), .Y(n_569) );
INVx3_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g457 ( .A(n_404), .Y(n_457) );
AND2x2_ASAP7_75t_L g575 ( .A(n_404), .B(n_407), .Y(n_575) );
AND2x2_ASAP7_75t_L g482 ( .A(n_405), .B(n_451), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_405), .B(n_514), .Y(n_545) );
AND2x4_ASAP7_75t_L g405 ( .A(n_406), .B(n_407), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_406), .B(n_525), .Y(n_524) );
AND2x2_ASAP7_75t_L g456 ( .A(n_407), .B(n_457), .Y(n_456) );
OAI22xp5_ASAP7_75t_SL g408 ( .A1(n_409), .A2(n_415), .B1(n_417), .B2(n_421), .Y(n_408) );
INVx2_ASAP7_75t_SL g409 ( .A(n_410), .Y(n_409) );
AND2x2_ASAP7_75t_L g410 ( .A(n_411), .B(n_413), .Y(n_410) );
AND2x2_ASAP7_75t_L g418 ( .A(n_411), .B(n_419), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_411), .B(n_554), .Y(n_553) );
INVx2_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g443 ( .A(n_412), .Y(n_443) );
INVx2_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_SL g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g502 ( .A(n_419), .Y(n_502) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
AND2x2_ASAP7_75t_L g485 ( .A(n_420), .B(n_434), .Y(n_485) );
AND2x2_ASAP7_75t_L g487 ( .A(n_420), .B(n_441), .Y(n_487) );
INVx1_ASAP7_75t_L g555 ( .A(n_420), .Y(n_555) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
AOI22xp5_ASAP7_75t_L g566 ( .A1(n_422), .A2(n_560), .B1(n_567), .B2(n_569), .Y(n_566) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g497 ( .A(n_424), .Y(n_497) );
AOI211xp5_ASAP7_75t_SL g425 ( .A1(n_426), .A2(n_427), .B(n_430), .C(n_437), .Y(n_425) );
NOR2x1_ASAP7_75t_L g565 ( .A(n_427), .B(n_531), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_428), .B(n_497), .Y(n_496) );
INVx2_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
AOI21xp33_ASAP7_75t_L g430 ( .A1(n_431), .A2(n_433), .B(n_435), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
OAI332xp33_ASAP7_75t_L g437 ( .A1(n_438), .A2(n_439), .A3(n_440), .B1(n_442), .B2(n_444), .B3(n_446), .C1(n_448), .C2(n_450), .Y(n_437) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
AOI22xp5_ASAP7_75t_L g530 ( .A1(n_441), .A2(n_531), .B1(n_535), .B2(n_536), .Y(n_530) );
INVxp67_ASAP7_75t_SL g535 ( .A(n_442), .Y(n_535) );
INVx2_ASAP7_75t_SL g442 ( .A(n_443), .Y(n_442) );
INVx2_ASAP7_75t_SL g590 ( .A(n_444), .Y(n_590) );
INVx2_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
AND2x2_ASAP7_75t_L g556 ( .A(n_447), .B(n_557), .Y(n_556) );
AND2x2_ASAP7_75t_L g591 ( .A(n_447), .B(n_592), .Y(n_591) );
INVx2_ASAP7_75t_SL g476 ( .A(n_449), .Y(n_476) );
AND2x2_ASAP7_75t_L g477 ( .A(n_449), .B(n_462), .Y(n_477) );
INVx2_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
AND4x1_ASAP7_75t_L g452 ( .A(n_453), .B(n_467), .C(n_473), .D(n_478), .Y(n_452) );
A2O1A1Ixp33_ASAP7_75t_L g453 ( .A1(n_454), .A2(n_458), .B(n_459), .C(n_465), .Y(n_453) );
INVxp67_ASAP7_75t_SL g454 ( .A(n_455), .Y(n_454) );
OAI321xp33_ASAP7_75t_L g581 ( .A1(n_455), .A2(n_522), .A3(n_535), .B1(n_582), .B2(n_584), .C(n_589), .Y(n_581) );
INVx3_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVxp67_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_461), .B(n_463), .Y(n_460) );
BUFx2_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx1_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVx1_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx2_ASAP7_75t_SL g541 ( .A(n_466), .Y(n_541) );
INVx2_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
AOI21xp5_ASAP7_75t_L g483 ( .A1(n_476), .A2(n_484), .B(n_486), .Y(n_483) );
A2O1A1Ixp33_ASAP7_75t_L g478 ( .A1(n_479), .A2(n_482), .B(n_483), .C(n_488), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
INVxp67_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
INVx1_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
AOI22xp33_ASAP7_75t_L g503 ( .A1(n_487), .A2(n_504), .B1(n_512), .B2(n_515), .Y(n_503) );
INVxp67_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
HB1xp67_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
HB1xp67_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
NOR2x1_ASAP7_75t_L g492 ( .A(n_493), .B(n_529), .Y(n_492) );
OAI211xp5_ASAP7_75t_SL g493 ( .A1(n_494), .A2(n_498), .B(n_503), .C(n_518), .Y(n_493) );
INVxp67_ASAP7_75t_SL g494 ( .A(n_495), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
INVx1_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_501), .B(n_502), .Y(n_500) );
OR2x2_ASAP7_75t_L g573 ( .A(n_502), .B(n_574), .Y(n_573) );
INVx2_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
NOR2xp33_ASAP7_75t_L g579 ( .A(n_505), .B(n_580), .Y(n_579) );
OR2x2_ASAP7_75t_L g587 ( .A(n_506), .B(n_588), .Y(n_587) );
INVx1_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
INVx2_ASAP7_75t_L g548 ( .A(n_507), .Y(n_548) );
INVx1_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
INVx1_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
INVx1_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
HB1xp67_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
AOI32xp33_ASAP7_75t_L g518 ( .A1(n_519), .A2(n_521), .A3(n_522), .B1(n_523), .B2(n_526), .Y(n_518) );
INVx2_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
INVx1_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
INVx2_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
NAND3xp33_ASAP7_75t_SL g529 ( .A(n_530), .B(n_538), .C(n_550), .Y(n_529) );
AND2x4_ASAP7_75t_L g531 ( .A(n_532), .B(n_534), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
AND2x2_ASAP7_75t_L g536 ( .A(n_534), .B(n_537), .Y(n_536) );
AOI22xp33_ASAP7_75t_L g589 ( .A1(n_534), .A2(n_590), .B1(n_591), .B2(n_593), .Y(n_589) );
AOI22xp33_ASAP7_75t_L g538 ( .A1(n_539), .A2(n_543), .B1(n_547), .B2(n_549), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
NAND2x1p5_ASAP7_75t_SL g540 ( .A(n_541), .B(n_542), .Y(n_540) );
NAND3xp33_ASAP7_75t_L g543 ( .A(n_544), .B(n_545), .C(n_546), .Y(n_543) );
A2O1A1Ixp33_ASAP7_75t_L g562 ( .A1(n_546), .A2(n_563), .B(n_565), .C(n_566), .Y(n_562) );
INVx1_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
AOI22xp5_ASAP7_75t_L g550 ( .A1(n_551), .A2(n_556), .B1(n_558), .B2(n_560), .Y(n_550) );
BUFx2_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
INVx2_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
INVx1_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
NOR3xp33_ASAP7_75t_L g561 ( .A(n_562), .B(n_570), .C(n_581), .Y(n_561) );
BUFx2_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
INVx1_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
A2O1A1Ixp33_ASAP7_75t_L g570 ( .A1(n_571), .A2(n_573), .B(n_576), .C(n_578), .Y(n_570) );
HB1xp67_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
INVx1_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
INVx1_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
INVxp67_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
NOR2x1_ASAP7_75t_L g585 ( .A(n_586), .B(n_587), .Y(n_585) );
BUFx2_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
OA21x2_ASAP7_75t_L g611 ( .A1(n_596), .A2(n_612), .B(n_613), .Y(n_611) );
NOR2xp33_ASAP7_75t_L g596 ( .A(n_597), .B(n_599), .Y(n_596) );
HB1xp67_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
OAI222xp33_ASAP7_75t_L g600 ( .A1(n_601), .A2(n_604), .B1(n_606), .B2(n_608), .C1(n_610), .C2(n_614), .Y(n_600) );
CKINVDCx20_ASAP7_75t_R g603 ( .A(n_602), .Y(n_603) );
INVx1_ASAP7_75t_SL g604 ( .A(n_605), .Y(n_604) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
BUFx2_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
BUFx2_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
INVx1_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
endmodule