module fake_jpeg_1425_n_80 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_80);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_80;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_24),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_20),
.B(n_0),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_28),
.B(n_30),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_26),
.Y(n_29)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_21),
.B(n_0),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_31),
.B(n_23),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_L g32 ( 
.A1(n_29),
.A2(n_26),
.B1(n_24),
.B2(n_25),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_27),
.B(n_22),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_37),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_31),
.B(n_23),
.Y(n_36)
);

NOR2x1_ASAP7_75t_L g41 ( 
.A(n_36),
.B(n_31),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g39 ( 
.A(n_37),
.Y(n_39)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

BUFx12f_ASAP7_75t_SL g49 ( 
.A(n_41),
.Y(n_49)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_38),
.Y(n_42)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

INVx13_ASAP7_75t_L g51 ( 
.A(n_45),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_41),
.B(n_33),
.Y(n_47)
);

NOR3xp33_ASAP7_75t_L g57 ( 
.A(n_47),
.B(n_43),
.C(n_12),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_43),
.A2(n_38),
.B1(n_31),
.B2(n_3),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_52),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_47),
.B(n_44),
.C(n_13),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_54),
.B(n_1),
.C(n_2),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_46),
.B(n_44),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_55),
.B(n_56),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_52),
.Y(n_56)
);

NAND3xp33_ASAP7_75t_L g66 ( 
.A(n_57),
.B(n_58),
.C(n_59),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_48),
.B(n_1),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_50),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_53),
.A2(n_49),
.B1(n_51),
.B2(n_3),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_61),
.B(n_4),
.Y(n_69)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_57),
.Y(n_62)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_62),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_63),
.B(n_65),
.C(n_2),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_56),
.A2(n_49),
.B1(n_51),
.B2(n_5),
.Y(n_64)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_64),
.Y(n_71)
);

XOR2xp5_ASAP7_75t_L g65 ( 
.A(n_55),
.B(n_15),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_67),
.B(n_4),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_69),
.B(n_70),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_60),
.B(n_17),
.C(n_19),
.Y(n_70)
);

XOR2xp5_ASAP7_75t_L g72 ( 
.A(n_68),
.B(n_65),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_L g75 ( 
.A(n_72),
.B(n_73),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_L g76 ( 
.A(n_72),
.B(n_71),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_76),
.B(n_75),
.Y(n_77)
);

OAI21x1_ASAP7_75t_L g78 ( 
.A1(n_77),
.A2(n_74),
.B(n_66),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_78),
.A2(n_66),
.B(n_10),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g80 ( 
.A1(n_79),
.A2(n_14),
.B(n_18),
.Y(n_80)
);


endmodule