module fake_jpeg_28442_n_35 (n_3, n_2, n_1, n_0, n_4, n_5, n_35);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_35;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_20;
wire n_18;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

BUFx6f_ASAP7_75t_L g6 ( 
.A(n_2),
.Y(n_6)
);

OR2x2_ASAP7_75t_L g7 ( 
.A(n_4),
.B(n_5),
.Y(n_7)
);

INVx3_ASAP7_75t_SL g8 ( 
.A(n_5),
.Y(n_8)
);

INVx3_ASAP7_75t_L g9 ( 
.A(n_0),
.Y(n_9)
);

BUFx12f_ASAP7_75t_L g10 ( 
.A(n_2),
.Y(n_10)
);

BUFx12f_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_9),
.Y(n_12)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g13 ( 
.A(n_7),
.B(n_3),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_13),
.B(n_15),
.Y(n_18)
);

AOI22xp33_ASAP7_75t_L g14 ( 
.A1(n_6),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_14)
);

OAI22xp5_ASAP7_75t_L g19 ( 
.A1(n_14),
.A2(n_8),
.B1(n_6),
.B2(n_1),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_7),
.B(n_4),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_16),
.B(n_10),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_11),
.B(n_1),
.Y(n_17)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_17),
.B(n_11),
.C(n_8),
.Y(n_21)
);

AOI21xp5_ASAP7_75t_L g23 ( 
.A1(n_19),
.A2(n_21),
.B(n_17),
.Y(n_23)
);

NAND3xp33_ASAP7_75t_SL g26 ( 
.A(n_22),
.B(n_10),
.C(n_11),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g28 ( 
.A(n_23),
.B(n_24),
.C(n_25),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_20),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_L g25 ( 
.A1(n_18),
.A2(n_15),
.B(n_12),
.Y(n_25)
);

XOR2xp5_ASAP7_75t_L g27 ( 
.A(n_26),
.B(n_21),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_27),
.B(n_10),
.Y(n_30)
);

FAx1_ASAP7_75t_SL g29 ( 
.A(n_28),
.B(n_11),
.CI(n_10),
.CON(n_29),
.SN(n_29)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_29),
.B(n_30),
.Y(n_32)
);

XNOR2xp5_ASAP7_75t_L g31 ( 
.A(n_30),
.B(n_27),
.Y(n_31)
);

AOI21xp5_ASAP7_75t_L g33 ( 
.A1(n_31),
.A2(n_32),
.B(n_29),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g34 ( 
.A(n_33),
.B(n_29),
.C(n_31),
.Y(n_34)
);

XOR2xp5_ASAP7_75t_L g35 ( 
.A(n_34),
.B(n_29),
.Y(n_35)
);


endmodule