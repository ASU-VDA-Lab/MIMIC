module fake_jpeg_19904_n_407 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_407);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_407;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVxp33_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_11),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_5),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_11),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_13),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

BUFx4f_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_10),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_44),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_45),
.Y(n_94)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_46),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_34),
.B(n_14),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_47),
.B(n_50),
.Y(n_89)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_21),
.Y(n_48)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_48),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_20),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_49),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_34),
.B(n_14),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_18),
.B(n_13),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_51),
.B(n_54),
.Y(n_93)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_19),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g112 ( 
.A(n_52),
.Y(n_112)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_17),
.Y(n_53)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_53),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_17),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_20),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_55),
.Y(n_119)
);

OR2x2_ASAP7_75t_L g56 ( 
.A(n_18),
.B(n_0),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_56),
.B(n_61),
.Y(n_96)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_57),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_58),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

INVx6_ASAP7_75t_L g131 ( 
.A(n_59),
.Y(n_131)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_26),
.Y(n_60)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_60),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_17),
.Y(n_61)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_26),
.Y(n_62)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_62),
.Y(n_91)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_17),
.Y(n_63)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_63),
.Y(n_109)
);

INVx13_ASAP7_75t_L g64 ( 
.A(n_15),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_64),
.B(n_65),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_22),
.B(n_0),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

INVx6_ASAP7_75t_L g138 ( 
.A(n_66),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

BUFx2_ASAP7_75t_L g92 ( 
.A(n_67),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_19),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_68),
.B(n_71),
.Y(n_124)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_38),
.Y(n_69)
);

BUFx2_ASAP7_75t_SL g139 ( 
.A(n_69),
.Y(n_139)
);

BUFx4f_ASAP7_75t_SL g70 ( 
.A(n_19),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_70),
.B(n_82),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_22),
.B(n_0),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_19),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g136 ( 
.A(n_72),
.Y(n_136)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_26),
.Y(n_73)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_73),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_19),
.Y(n_74)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_74),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_40),
.B(n_2),
.C(n_3),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_75),
.B(n_24),
.C(n_37),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_25),
.B(n_2),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_76),
.B(n_78),
.Y(n_127)
);

BUFx10_ASAP7_75t_L g77 ( 
.A(n_29),
.Y(n_77)
);

INVx13_ASAP7_75t_L g106 ( 
.A(n_77),
.Y(n_106)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_40),
.Y(n_78)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_40),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_79),
.B(n_80),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_25),
.B(n_3),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_40),
.Y(n_81)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_81),
.Y(n_101)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_40),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_36),
.Y(n_83)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_83),
.Y(n_116)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_33),
.Y(n_84)
);

HB1xp67_ASAP7_75t_L g111 ( 
.A(n_84),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_27),
.B(n_3),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_85),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_21),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_86),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_36),
.Y(n_87)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_87),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_56),
.A2(n_23),
.B1(n_39),
.B2(n_27),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_97),
.A2(n_104),
.B1(n_114),
.B2(n_120),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_46),
.A2(n_23),
.B1(n_33),
.B2(n_29),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_100),
.A2(n_107),
.B1(n_108),
.B2(n_77),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_57),
.A2(n_23),
.B1(n_33),
.B2(n_32),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_60),
.A2(n_29),
.B1(n_32),
.B2(n_39),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_62),
.A2(n_73),
.B1(n_63),
.B2(n_53),
.Y(n_108)
);

NAND2x1_ASAP7_75t_L g110 ( 
.A(n_75),
.B(n_64),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_110),
.B(n_115),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_66),
.A2(n_24),
.B1(n_37),
.B2(n_35),
.Y(n_114)
);

OA22x2_ASAP7_75t_L g117 ( 
.A1(n_82),
.A2(n_35),
.B1(n_31),
.B2(n_30),
.Y(n_117)
);

OA22x2_ASAP7_75t_L g140 ( 
.A1(n_117),
.A2(n_59),
.B1(n_58),
.B2(n_67),
.Y(n_140)
);

AND2x2_ASAP7_75t_SL g118 ( 
.A(n_45),
.B(n_16),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_118),
.B(n_121),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_L g120 ( 
.A1(n_48),
.A2(n_31),
.B1(n_30),
.B2(n_28),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_44),
.B(n_28),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g122 ( 
.A1(n_69),
.A2(n_43),
.B1(n_36),
.B2(n_42),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_122),
.A2(n_132),
.B1(n_8),
.B2(n_9),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_49),
.B(n_43),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_126),
.B(n_134),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_84),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_130),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_79),
.A2(n_43),
.B1(n_42),
.B2(n_16),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_55),
.B(n_4),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_140),
.A2(n_162),
.B(n_169),
.Y(n_197)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_135),
.Y(n_142)
);

BUFx2_ASAP7_75t_L g195 ( 
.A(n_142),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_89),
.B(n_87),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_143),
.B(n_171),
.Y(n_190)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_123),
.Y(n_144)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_144),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_125),
.B(n_113),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_146),
.B(n_150),
.Y(n_194)
);

OAI22xp33_ASAP7_75t_L g147 ( 
.A1(n_126),
.A2(n_70),
.B1(n_81),
.B2(n_74),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_147),
.A2(n_164),
.B1(n_170),
.B2(n_177),
.Y(n_218)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_88),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g205 ( 
.A(n_148),
.Y(n_205)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_123),
.Y(n_149)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_149),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_129),
.B(n_70),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_93),
.B(n_83),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_151),
.B(n_152),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_124),
.B(n_52),
.Y(n_152)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_139),
.Y(n_154)
);

INVx5_ASAP7_75t_L g210 ( 
.A(n_154),
.Y(n_210)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_135),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_155),
.B(n_156),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_105),
.B(n_52),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_95),
.Y(n_157)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_157),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_127),
.B(n_78),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_158),
.B(n_159),
.Y(n_219)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_88),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_98),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_160),
.B(n_161),
.Y(n_222)
);

INVx13_ASAP7_75t_L g161 ( 
.A(n_121),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_110),
.B(n_78),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_96),
.B(n_115),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_163),
.B(n_165),
.Y(n_223)
);

BUFx16f_ASAP7_75t_L g165 ( 
.A(n_112),
.Y(n_165)
);

INVx5_ASAP7_75t_L g166 ( 
.A(n_102),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_166),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_95),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_167),
.Y(n_208)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_117),
.B(n_72),
.Y(n_169)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_112),
.Y(n_171)
);

BUFx2_ASAP7_75t_L g172 ( 
.A(n_112),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_172),
.B(n_176),
.Y(n_224)
);

AOI21xp33_ASAP7_75t_L g173 ( 
.A1(n_137),
.A2(n_4),
.B(n_8),
.Y(n_173)
);

OR2x2_ASAP7_75t_SL g215 ( 
.A(n_173),
.B(n_179),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_L g221 ( 
.A1(n_174),
.A2(n_92),
.B1(n_106),
.B2(n_136),
.Y(n_221)
);

OA22x2_ASAP7_75t_L g175 ( 
.A1(n_128),
.A2(n_77),
.B1(n_9),
.B2(n_10),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_175),
.A2(n_130),
.B1(n_174),
.B2(n_153),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_134),
.B(n_77),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_L g177 ( 
.A1(n_128),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_177)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_94),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_178),
.B(n_182),
.Y(n_200)
);

AOI21xp33_ASAP7_75t_L g179 ( 
.A1(n_117),
.A2(n_11),
.B(n_116),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_98),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_180),
.B(n_181),
.Y(n_226)
);

BUFx2_ASAP7_75t_L g181 ( 
.A(n_99),
.Y(n_181)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_94),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_116),
.Y(n_183)
);

AND2x2_ASAP7_75t_SL g212 ( 
.A(n_183),
.B(n_119),
.Y(n_212)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_136),
.Y(n_184)
);

AND2x2_ASAP7_75t_L g204 ( 
.A(n_184),
.B(n_103),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_117),
.B(n_114),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_185),
.B(n_186),
.Y(n_189)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_101),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_187),
.A2(n_188),
.B1(n_216),
.B2(n_217),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_153),
.A2(n_131),
.B1(n_138),
.B2(n_101),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_168),
.B(n_118),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_191),
.B(n_192),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_145),
.B(n_118),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_169),
.A2(n_111),
.B(n_133),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_198),
.A2(n_175),
.B(n_92),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_SL g201 ( 
.A(n_141),
.B(n_162),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_SL g261 ( 
.A(n_201),
.B(n_225),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_141),
.B(n_133),
.C(n_109),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_203),
.B(n_165),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_204),
.A2(n_211),
.B(n_212),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_141),
.B(n_138),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_206),
.B(n_214),
.Y(n_243)
);

AND2x6_ASAP7_75t_L g209 ( 
.A(n_162),
.B(n_109),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_209),
.B(n_147),
.Y(n_227)
);

AND2x2_ASAP7_75t_L g211 ( 
.A(n_140),
.B(n_131),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_169),
.B(n_119),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_140),
.A2(n_90),
.B1(n_91),
.B2(n_102),
.Y(n_216)
);

OAI22xp33_ASAP7_75t_L g217 ( 
.A1(n_161),
.A2(n_90),
.B1(n_91),
.B2(n_103),
.Y(n_217)
);

AND2x2_ASAP7_75t_SL g220 ( 
.A(n_140),
.B(n_99),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_220),
.B(n_197),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_221),
.A2(n_220),
.B1(n_216),
.B2(n_211),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_164),
.B(n_106),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_227),
.B(n_231),
.Y(n_279)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_226),
.Y(n_228)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_228),
.Y(n_269)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_226),
.Y(n_230)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_230),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_223),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_219),
.B(n_166),
.Y(n_232)
);

CKINVDCx14_ASAP7_75t_R g283 ( 
.A(n_232),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_218),
.A2(n_175),
.B1(n_142),
.B2(n_155),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_233),
.A2(n_245),
.B1(n_246),
.B2(n_254),
.Y(n_273)
);

HB1xp67_ASAP7_75t_L g234 ( 
.A(n_193),
.Y(n_234)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_234),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_207),
.B(n_154),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_235),
.B(n_238),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_236),
.A2(n_198),
.B1(n_201),
.B2(n_203),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_199),
.Y(n_238)
);

AOI32xp33_ASAP7_75t_L g239 ( 
.A1(n_209),
.A2(n_175),
.A3(n_149),
.B1(n_144),
.B2(n_171),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_239),
.B(n_242),
.Y(n_280)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_195),
.Y(n_240)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_240),
.Y(n_272)
);

BUFx2_ASAP7_75t_L g241 ( 
.A(n_195),
.Y(n_241)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_241),
.Y(n_281)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_195),
.Y(n_242)
);

INVx13_ASAP7_75t_L g244 ( 
.A(n_206),
.Y(n_244)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_244),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_218),
.A2(n_184),
.B1(n_178),
.B2(n_182),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_189),
.A2(n_181),
.B1(n_167),
.B2(n_157),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_199),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_247),
.B(n_252),
.Y(n_262)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_200),
.Y(n_249)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_249),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_202),
.Y(n_250)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_250),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_251),
.B(n_261),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_194),
.Y(n_252)
);

AND2x2_ASAP7_75t_L g264 ( 
.A(n_253),
.B(n_188),
.Y(n_264)
);

OAI22xp33_ASAP7_75t_SL g254 ( 
.A1(n_220),
.A2(n_165),
.B1(n_172),
.B2(n_211),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_196),
.B(n_205),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_255),
.Y(n_265)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_200),
.Y(n_256)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_256),
.Y(n_290)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_200),
.Y(n_257)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_257),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_258),
.B(n_260),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_205),
.B(n_190),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_259),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_213),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_264),
.A2(n_246),
.B1(n_256),
.B2(n_237),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_270),
.A2(n_271),
.B(n_243),
.Y(n_296)
);

A2O1A1O1Ixp25_ASAP7_75t_L g271 ( 
.A1(n_236),
.A2(n_215),
.B(n_225),
.C(n_197),
.D(n_189),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_274),
.B(n_192),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_240),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_277),
.B(n_286),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_229),
.B(n_191),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_282),
.B(n_289),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_233),
.A2(n_187),
.B1(n_214),
.B2(n_215),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_284),
.A2(n_285),
.B1(n_237),
.B2(n_253),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_245),
.A2(n_224),
.B1(n_217),
.B2(n_190),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_238),
.Y(n_286)
);

AND2x2_ASAP7_75t_L g287 ( 
.A(n_249),
.B(n_224),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_287),
.A2(n_248),
.B(n_257),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_229),
.B(n_222),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_L g292 ( 
.A1(n_280),
.A2(n_258),
.B(n_243),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_L g339 ( 
.A1(n_292),
.A2(n_299),
.B(n_312),
.Y(n_339)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_262),
.Y(n_293)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_293),
.Y(n_320)
);

OR2x2_ASAP7_75t_L g294 ( 
.A(n_268),
.B(n_284),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_294),
.B(n_301),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_SL g328 ( 
.A(n_296),
.B(n_305),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_297),
.A2(n_311),
.B1(n_264),
.B2(n_287),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_267),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_298),
.B(n_309),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_289),
.B(n_230),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_282),
.B(n_228),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_302),
.B(n_306),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_274),
.B(n_251),
.C(n_261),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_303),
.B(n_269),
.C(n_290),
.Y(n_332)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_262),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_304),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_263),
.B(n_231),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_266),
.Y(n_307)
);

CKINVDCx16_ASAP7_75t_R g318 ( 
.A(n_307),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_276),
.B(n_265),
.Y(n_308)
);

CKINVDCx16_ASAP7_75t_R g333 ( 
.A(n_308),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_266),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_310),
.B(n_313),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_264),
.A2(n_239),
.B1(n_252),
.B2(n_244),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_L g312 ( 
.A1(n_270),
.A2(n_248),
.B(n_247),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_283),
.B(n_260),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_272),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_314),
.Y(n_324)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_272),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_315),
.A2(n_317),
.B1(n_281),
.B2(n_242),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g316 ( 
.A(n_279),
.Y(n_316)
);

INVx2_ASAP7_75t_SL g325 ( 
.A(n_316),
.Y(n_325)
);

INVx2_ASAP7_75t_SL g317 ( 
.A(n_281),
.Y(n_317)
);

FAx1_ASAP7_75t_SL g319 ( 
.A(n_296),
.B(n_287),
.CI(n_271),
.CON(n_319),
.SN(n_319)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_319),
.B(n_295),
.Y(n_353)
);

CKINVDCx14_ASAP7_75t_R g352 ( 
.A(n_322),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_323),
.B(n_330),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_297),
.A2(n_273),
.B1(n_275),
.B2(n_268),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_293),
.A2(n_273),
.B1(n_275),
.B2(n_263),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_331),
.B(n_336),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_332),
.B(n_334),
.Y(n_342)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_303),
.B(n_285),
.Y(n_334)
);

NOR2xp67_ASAP7_75t_R g335 ( 
.A(n_312),
.B(n_291),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_SL g356 ( 
.A(n_335),
.B(n_212),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_304),
.A2(n_291),
.B1(n_290),
.B2(n_278),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_SL g337 ( 
.A(n_303),
.B(n_278),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_337),
.A2(n_312),
.B1(n_292),
.B2(n_305),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_326),
.A2(n_309),
.B1(n_294),
.B2(n_311),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_340),
.A2(n_347),
.B1(n_348),
.B2(n_331),
.Y(n_363)
);

XOR2xp5_ASAP7_75t_L g361 ( 
.A(n_341),
.B(n_350),
.Y(n_361)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_338),
.Y(n_343)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_343),
.Y(n_358)
);

OAI21xp5_ASAP7_75t_SL g345 ( 
.A1(n_335),
.A2(n_299),
.B(n_300),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_345),
.B(n_346),
.Y(n_364)
);

OAI21xp5_ASAP7_75t_SL g346 ( 
.A1(n_323),
.A2(n_300),
.B(n_310),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_321),
.A2(n_294),
.B1(n_301),
.B2(n_314),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_321),
.A2(n_306),
.B1(n_302),
.B2(n_295),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_332),
.B(n_305),
.C(n_292),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_349),
.B(n_355),
.C(n_339),
.Y(n_369)
);

OAI21xp5_ASAP7_75t_SL g350 ( 
.A1(n_324),
.A2(n_313),
.B(n_307),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_327),
.Y(n_351)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_351),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_SL g362 ( 
.A(n_353),
.B(n_329),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_334),
.B(n_315),
.C(n_308),
.Y(n_355)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_356),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_327),
.B(n_212),
.Y(n_357)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_357),
.Y(n_365)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_362),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_363),
.A2(n_366),
.B1(n_367),
.B2(n_371),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_352),
.A2(n_320),
.B1(n_330),
.B2(n_328),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_344),
.A2(n_320),
.B1(n_339),
.B2(n_336),
.Y(n_367)
);

INVxp33_ASAP7_75t_L g368 ( 
.A(n_347),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_368),
.B(n_348),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_369),
.B(n_355),
.C(n_342),
.Y(n_372)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_350),
.Y(n_370)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_370),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_344),
.A2(n_322),
.B1(n_333),
.B2(n_319),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_372),
.B(n_349),
.C(n_342),
.Y(n_383)
);

BUFx3_ASAP7_75t_L g375 ( 
.A(n_358),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_375),
.B(n_377),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_369),
.A2(n_360),
.B1(n_361),
.B2(n_359),
.Y(n_376)
);

OAI21xp5_ASAP7_75t_L g384 ( 
.A1(n_376),
.A2(n_361),
.B(n_345),
.Y(n_384)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_365),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_371),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_378),
.B(n_380),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_SL g380 ( 
.A(n_364),
.B(n_346),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_363),
.A2(n_354),
.B1(n_340),
.B2(n_357),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_381),
.B(n_367),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_SL g391 ( 
.A(n_382),
.B(n_354),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_SL g394 ( 
.A(n_383),
.B(n_389),
.Y(n_394)
);

AOI21xp5_ASAP7_75t_L g393 ( 
.A1(n_384),
.A2(n_385),
.B(n_386),
.Y(n_393)
);

AND2x2_ASAP7_75t_L g385 ( 
.A(n_373),
.B(n_364),
.Y(n_385)
);

OAI21xp5_ASAP7_75t_SL g386 ( 
.A1(n_374),
.A2(n_318),
.B(n_366),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_SL g388 ( 
.A(n_376),
.B(n_325),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_L g395 ( 
.A1(n_388),
.A2(n_379),
.B1(n_381),
.B2(n_368),
.Y(n_395)
);

AO21x1_ASAP7_75t_L g397 ( 
.A1(n_391),
.A2(n_325),
.B(n_375),
.Y(n_397)
);

OAI21xp5_ASAP7_75t_L g392 ( 
.A1(n_388),
.A2(n_372),
.B(n_341),
.Y(n_392)
);

AOI322xp5_ASAP7_75t_L g401 ( 
.A1(n_392),
.A2(n_395),
.A3(n_397),
.B1(n_288),
.B2(n_317),
.C1(n_213),
.C2(n_250),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_390),
.B(n_379),
.C(n_337),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_SL g398 ( 
.A(n_396),
.B(n_387),
.Y(n_398)
);

AOI322xp5_ASAP7_75t_L g403 ( 
.A1(n_398),
.A2(n_399),
.A3(n_401),
.B1(n_317),
.B2(n_204),
.C1(n_210),
.C2(n_241),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_L g399 ( 
.A1(n_393),
.A2(n_325),
.B1(n_319),
.B2(n_328),
.Y(n_399)
);

A2O1A1O1Ixp25_ASAP7_75t_L g400 ( 
.A1(n_394),
.A2(n_317),
.B(n_193),
.C(n_288),
.D(n_250),
.Y(n_400)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_400),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_403),
.B(n_208),
.C(n_204),
.Y(n_404)
);

AOI21xp5_ASAP7_75t_L g406 ( 
.A1(n_404),
.A2(n_405),
.B(n_202),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_402),
.B(n_208),
.C(n_210),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_L g407 ( 
.A(n_406),
.B(n_241),
.Y(n_407)
);


endmodule