module fake_jpeg_28482_n_167 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_167);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_167;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g51 ( 
.A(n_23),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_40),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_34),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_43),
.B(n_14),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_49),
.Y(n_57)
);

CKINVDCx5p33_ASAP7_75t_R g58 ( 
.A(n_8),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_31),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_8),
.Y(n_60)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_29),
.Y(n_62)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_7),
.Y(n_63)
);

INVx1_ASAP7_75t_SL g64 ( 
.A(n_24),
.Y(n_64)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_27),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_12),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_4),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_25),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_37),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_22),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_10),
.Y(n_71)
);

OR2x2_ASAP7_75t_L g72 ( 
.A(n_64),
.B(n_0),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_72),
.B(n_74),
.Y(n_93)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_63),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_73),
.B(n_75),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_56),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_67),
.Y(n_76)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_76),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_60),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_77),
.A2(n_64),
.B1(n_59),
.B2(n_71),
.Y(n_82)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_60),
.Y(n_78)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_78),
.Y(n_94)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_51),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_79),
.B(n_80),
.Y(n_81)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_53),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_82),
.A2(n_59),
.B1(n_62),
.B2(n_57),
.Y(n_103)
);

OAI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_76),
.A2(n_65),
.B1(n_55),
.B2(n_71),
.Y(n_83)
);

OAI21xp33_ASAP7_75t_SL g98 ( 
.A1(n_83),
.A2(n_65),
.B(n_84),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_79),
.B(n_66),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_86),
.B(n_89),
.Y(n_96)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_78),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_87),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_73),
.Y(n_88)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_88),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_80),
.B(n_52),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_72),
.B(n_59),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_90),
.B(n_3),
.Y(n_111)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_75),
.Y(n_91)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_91),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_78),
.Y(n_92)
);

HB1xp67_ASAP7_75t_L g95 ( 
.A(n_92),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_98),
.A2(n_92),
.B1(n_6),
.B2(n_7),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_81),
.B(n_70),
.C(n_68),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_99),
.B(n_100),
.C(n_4),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_81),
.B(n_70),
.C(n_69),
.Y(n_100)
);

INVx1_ASAP7_75t_SL g101 ( 
.A(n_88),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_101),
.B(n_108),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_103),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_93),
.B(n_58),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_104),
.B(n_105),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_90),
.B(n_54),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_91),
.Y(n_106)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_106),
.Y(n_134)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_84),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_107),
.B(n_16),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_85),
.B(n_1),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_94),
.B(n_61),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_109),
.B(n_61),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_94),
.B(n_2),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_110),
.B(n_111),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_87),
.B(n_3),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_113),
.B(n_15),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_117),
.B(n_118),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_119),
.A2(n_121),
.B1(n_122),
.B2(n_123),
.Y(n_147)
);

BUFx2_ASAP7_75t_L g120 ( 
.A(n_97),
.Y(n_120)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_120),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_103),
.A2(n_5),
.B1(n_6),
.B2(n_9),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_98),
.A2(n_5),
.B1(n_9),
.B2(n_10),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_102),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_123)
);

AND2x2_ASAP7_75t_SL g124 ( 
.A(n_108),
.B(n_32),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_124),
.B(n_38),
.Y(n_143)
);

OR2x2_ASAP7_75t_L g125 ( 
.A(n_96),
.B(n_11),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_125),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_126),
.A2(n_129),
.B(n_132),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_127),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_95),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_128),
.Y(n_135)
);

BUFx5_ASAP7_75t_L g130 ( 
.A(n_97),
.Y(n_130)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_130),
.Y(n_145)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_95),
.Y(n_131)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_131),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_112),
.A2(n_20),
.B1(n_21),
.B2(n_26),
.Y(n_132)
);

OAI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_98),
.A2(n_28),
.B1(n_30),
.B2(n_33),
.Y(n_133)
);

AND2x2_ASAP7_75t_SL g148 ( 
.A(n_133),
.B(n_47),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_120),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_137),
.B(n_148),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_114),
.B(n_35),
.C(n_36),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_139),
.B(n_143),
.C(n_146),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_114),
.A2(n_41),
.B(n_42),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_144),
.A2(n_125),
.B(n_124),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_115),
.B(n_46),
.Y(n_146)
);

NOR2x1_ASAP7_75t_L g150 ( 
.A(n_116),
.B(n_48),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_150),
.B(n_50),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_151),
.B(n_157),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_136),
.A2(n_133),
.B(n_134),
.Y(n_152)
);

AO21x1_ASAP7_75t_L g160 ( 
.A1(n_152),
.A2(n_140),
.B(n_138),
.Y(n_160)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_149),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_154),
.B(n_155),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_145),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_160),
.A2(n_153),
.B1(n_148),
.B2(n_147),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_161),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_162),
.B(n_159),
.Y(n_163)
);

AOI322xp5_ASAP7_75t_L g164 ( 
.A1(n_163),
.A2(n_135),
.A3(n_157),
.B1(n_158),
.B2(n_141),
.C1(n_146),
.C2(n_142),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_164),
.B(n_139),
.C(n_143),
.Y(n_165)
);

HB1xp67_ASAP7_75t_L g166 ( 
.A(n_165),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_166),
.B(n_156),
.C(n_150),
.Y(n_167)
);


endmodule