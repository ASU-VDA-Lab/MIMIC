module fake_jpeg_5904_n_228 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_228);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_228;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_9),
.Y(n_15)
);

INVxp67_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx5_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

HB1xp67_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

CKINVDCx16_ASAP7_75t_R g31 ( 
.A(n_4),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_32),
.B(n_36),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_15),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_33),
.B(n_30),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

HB1xp67_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

BUFx2_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_38),
.A2(n_20),
.B1(n_18),
.B2(n_17),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_40),
.B(n_41),
.Y(n_62)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_43),
.B(n_56),
.Y(n_81)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_44),
.B(n_50),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_48),
.A2(n_54),
.B1(n_58),
.B2(n_0),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_36),
.A2(n_18),
.B1(n_24),
.B2(n_15),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_49),
.A2(n_51),
.B1(n_29),
.B2(n_22),
.Y(n_78)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_32),
.A2(n_18),
.B1(n_24),
.B2(n_21),
.Y(n_51)
);

OAI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_36),
.A2(n_19),
.B1(n_21),
.B2(n_26),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_53),
.A2(n_38),
.B1(n_29),
.B2(n_22),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_32),
.A2(n_31),
.B1(n_26),
.B2(n_19),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_55),
.B(n_59),
.Y(n_82)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_40),
.A2(n_31),
.B1(n_30),
.B2(n_25),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_60),
.B(n_61),
.Y(n_83)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_40),
.B(n_16),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_63),
.B(n_25),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_65),
.B(n_28),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_66),
.A2(n_74),
.B1(n_47),
.B2(n_44),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_57),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_68),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_62),
.B(n_39),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_69),
.B(n_75),
.Y(n_92)
);

OR2x4_ASAP7_75t_L g70 ( 
.A(n_63),
.B(n_34),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_70),
.A2(n_79),
.B(n_45),
.Y(n_105)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_57),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_71),
.B(n_73),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_62),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_72),
.B(n_75),
.Y(n_91)
);

BUFx2_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

OAI22xp33_ASAP7_75t_L g74 ( 
.A1(n_49),
.A2(n_34),
.B1(n_35),
.B2(n_42),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_50),
.B(n_38),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_63),
.A2(n_38),
.B1(n_35),
.B2(n_42),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_76),
.A2(n_47),
.B1(n_56),
.B2(n_43),
.Y(n_86)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_52),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_77),
.B(n_84),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_78),
.A2(n_80),
.B1(n_1),
.B2(n_3),
.Y(n_107)
);

O2A1O1Ixp33_ASAP7_75t_L g79 ( 
.A1(n_46),
.A2(n_35),
.B(n_39),
.C(n_29),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_55),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_59),
.B(n_1),
.Y(n_85)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_85),
.Y(n_89)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_86),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_78),
.A2(n_70),
.B1(n_72),
.B2(n_69),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_88),
.B(n_28),
.Y(n_125)
);

HB1xp67_ASAP7_75t_L g90 ( 
.A(n_68),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_90),
.B(n_94),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_92),
.B(n_100),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_93),
.B(n_95),
.Y(n_126)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_83),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_67),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_96),
.B(n_98),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g97 ( 
.A(n_80),
.B(n_39),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_97),
.B(n_67),
.C(n_77),
.Y(n_112)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_81),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_76),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_99),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_82),
.B(n_60),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_65),
.Y(n_102)
);

INVx13_ASAP7_75t_L g111 ( 
.A(n_102),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_82),
.B(n_39),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_103),
.B(n_73),
.Y(n_130)
);

AO22x1_ASAP7_75t_SL g104 ( 
.A1(n_66),
.A2(n_45),
.B1(n_61),
.B2(n_22),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_104),
.A2(n_105),
.B(n_85),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_107),
.B(n_108),
.Y(n_127)
);

OR2x2_ASAP7_75t_L g108 ( 
.A(n_84),
.B(n_39),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_109),
.A2(n_115),
.B(n_117),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_112),
.B(n_125),
.C(n_130),
.Y(n_137)
);

OR2x2_ASAP7_75t_L g113 ( 
.A(n_96),
.B(n_79),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_113),
.B(n_104),
.Y(n_141)
);

INVx13_ASAP7_75t_L g114 ( 
.A(n_98),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_114),
.B(n_116),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_105),
.A2(n_79),
.B(n_64),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_106),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_92),
.A2(n_64),
.B(n_28),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_91),
.A2(n_103),
.B(n_97),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_119),
.A2(n_123),
.B(n_129),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_91),
.A2(n_64),
.B(n_28),
.Y(n_123)
);

AND2x6_ASAP7_75t_L g124 ( 
.A(n_88),
.B(n_64),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g133 ( 
.A(n_124),
.Y(n_133)
);

INVx13_ASAP7_75t_L g128 ( 
.A(n_94),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_128),
.B(n_100),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_99),
.A2(n_73),
.B(n_71),
.Y(n_129)
);

A2O1A1O1Ixp25_ASAP7_75t_L g134 ( 
.A1(n_124),
.A2(n_125),
.B(n_127),
.C(n_119),
.D(n_109),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_134),
.A2(n_141),
.B(n_142),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_135),
.B(n_144),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_SL g136 ( 
.A(n_124),
.B(n_95),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_136),
.B(n_123),
.C(n_116),
.Y(n_163)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_113),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_139),
.B(n_140),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_120),
.A2(n_104),
.B1(n_86),
.B2(n_101),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_115),
.A2(n_101),
.B(n_108),
.Y(n_142)
);

XNOR2x2_ASAP7_75t_SL g143 ( 
.A(n_113),
.B(n_95),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_143),
.B(n_111),
.Y(n_166)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_118),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_121),
.B(n_89),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_145),
.B(n_146),
.Y(n_155)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_121),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_120),
.A2(n_102),
.B1(n_89),
.B2(n_71),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_147),
.A2(n_149),
.B1(n_127),
.B2(n_117),
.Y(n_156)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_118),
.Y(n_148)
);

INVxp33_ASAP7_75t_L g162 ( 
.A(n_148),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_122),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_128),
.B(n_68),
.Y(n_150)
);

CKINVDCx14_ASAP7_75t_R g164 ( 
.A(n_150),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_128),
.B(n_114),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_151),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_143),
.B(n_130),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_153),
.A2(n_131),
.B(n_138),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_156),
.B(n_168),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_146),
.B(n_130),
.Y(n_157)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_157),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_139),
.A2(n_126),
.B1(n_112),
.B2(n_125),
.Y(n_159)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_159),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_132),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_160),
.B(n_165),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_133),
.A2(n_126),
.B1(n_112),
.B2(n_129),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_161),
.A2(n_134),
.B1(n_141),
.B2(n_142),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_163),
.B(n_137),
.C(n_138),
.Y(n_171)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_145),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_166),
.B(n_110),
.Y(n_182)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_147),
.Y(n_167)
);

INVx13_ASAP7_75t_L g179 ( 
.A(n_167),
.Y(n_179)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_140),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_171),
.B(n_172),
.C(n_178),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_157),
.B(n_137),
.C(n_136),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_154),
.A2(n_131),
.B(n_133),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_174),
.A2(n_176),
.B(n_180),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_177),
.B(n_182),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_158),
.B(n_110),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_168),
.A2(n_149),
.B(n_111),
.Y(n_180)
);

MAJx2_ASAP7_75t_L g181 ( 
.A(n_158),
.B(n_111),
.C(n_114),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_181),
.B(n_166),
.C(n_159),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_155),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_183),
.B(n_155),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_173),
.A2(n_167),
.B1(n_152),
.B2(n_160),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_186),
.A2(n_184),
.B1(n_164),
.B2(n_170),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_175),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_188),
.B(n_189),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_183),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_173),
.A2(n_163),
.B1(n_161),
.B2(n_165),
.Y(n_190)
);

O2A1O1Ixp33_ASAP7_75t_L g198 ( 
.A1(n_190),
.A2(n_194),
.B(n_177),
.C(n_184),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_170),
.B(n_152),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_192),
.B(n_169),
.C(n_180),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_193),
.A2(n_174),
.B(n_181),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_171),
.B(n_153),
.C(n_156),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_195),
.B(n_179),
.C(n_87),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_178),
.B(n_162),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_196),
.B(n_182),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_197),
.A2(n_200),
.B(n_203),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_198),
.B(n_201),
.Y(n_206)
);

MAJx2_ASAP7_75t_L g199 ( 
.A(n_187),
.B(n_176),
.C(n_153),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_199),
.A2(n_204),
.B(n_3),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_186),
.B(n_172),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_205),
.B(n_87),
.C(n_5),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_198),
.A2(n_193),
.B1(n_195),
.B2(n_190),
.Y(n_207)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_207),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_202),
.A2(n_185),
.B(n_191),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_209),
.B(n_211),
.Y(n_215)
);

OAI221xp5_ASAP7_75t_L g210 ( 
.A1(n_199),
.A2(n_205),
.B1(n_185),
.B2(n_179),
.C(n_191),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_210),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_212),
.B(n_6),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_206),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_213),
.B(n_217),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_216),
.B(n_208),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_211),
.B(n_7),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_218),
.A2(n_7),
.B(n_8),
.Y(n_220)
);

O2A1O1Ixp33_ASAP7_75t_L g223 ( 
.A1(n_219),
.A2(n_222),
.B(n_215),
.C(n_213),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_220),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_L g222 ( 
.A1(n_214),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_222)
);

AOI322xp5_ASAP7_75t_L g227 ( 
.A1(n_223),
.A2(n_224),
.A3(n_12),
.B1(n_14),
.B2(n_220),
.C1(n_124),
.C2(n_169),
.Y(n_227)
);

OAI21x1_ASAP7_75t_L g224 ( 
.A1(n_221),
.A2(n_9),
.B(n_11),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_225),
.B(n_12),
.C(n_13),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_226),
.B(n_227),
.Y(n_228)
);


endmodule