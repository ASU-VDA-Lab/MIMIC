module fake_jpeg_12079_n_22 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_22);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_22;

wire n_13;
wire n_21;
wire n_10;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_16;
wire n_9;
wire n_11;
wire n_17;
wire n_12;
wire n_8;
wire n_15;
wire n_7;

INVx4_ASAP7_75t_L g7 ( 
.A(n_3),
.Y(n_7)
);

NOR2xp33_ASAP7_75t_SL g8 ( 
.A(n_3),
.B(n_0),
.Y(n_8)
);

NOR2xp33_ASAP7_75t_L g9 ( 
.A(n_5),
.B(n_4),
.Y(n_9)
);

NAND2xp5_ASAP7_75t_L g10 ( 
.A(n_5),
.B(n_2),
.Y(n_10)
);

AOI21xp33_ASAP7_75t_L g11 ( 
.A1(n_4),
.A2(n_6),
.B(n_1),
.Y(n_11)
);

INVx4_ASAP7_75t_SL g12 ( 
.A(n_2),
.Y(n_12)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

OAI21xp5_ASAP7_75t_L g15 ( 
.A1(n_10),
.A2(n_13),
.B(n_9),
.Y(n_15)
);

AOI322xp5_ASAP7_75t_SL g20 ( 
.A1(n_15),
.A2(n_16),
.A3(n_17),
.B1(n_18),
.B2(n_12),
.C1(n_10),
.C2(n_8),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_10),
.B(n_13),
.Y(n_16)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_11),
.B(n_14),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_14),
.B(n_7),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_SL g19 ( 
.A1(n_17),
.A2(n_7),
.B1(n_12),
.B2(n_8),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_19),
.B(n_20),
.Y(n_21)
);

INVxp33_ASAP7_75t_SL g22 ( 
.A(n_21),
.Y(n_22)
);


endmodule