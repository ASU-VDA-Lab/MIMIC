module fake_jpeg_12315_n_616 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_616);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_616;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_596;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_442;
wire n_299;
wire n_300;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_384;
wire n_296;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_11),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_0),
.B(n_4),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx16f_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

CKINVDCx14_ASAP7_75t_R g38 ( 
.A(n_13),
.Y(n_38)
);

INVx1_ASAP7_75t_SL g39 ( 
.A(n_18),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_9),
.B(n_8),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_12),
.Y(n_43)
);

BUFx4f_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_3),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_11),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_12),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_16),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_11),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_6),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_9),
.Y(n_53)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_2),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_0),
.Y(n_55)
);

CKINVDCx14_ASAP7_75t_R g56 ( 
.A(n_3),
.Y(n_56)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_4),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g58 ( 
.A(n_2),
.Y(n_58)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_13),
.Y(n_59)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_7),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_3),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_62),
.Y(n_138)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_19),
.Y(n_63)
);

BUFx10_ASAP7_75t_L g198 ( 
.A(n_63),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_25),
.B(n_9),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_64),
.B(n_93),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_40),
.B(n_7),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_65),
.B(n_82),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_20),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_66),
.Y(n_136)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_67),
.Y(n_140)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_68),
.Y(n_141)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_19),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_69),
.Y(n_184)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_33),
.Y(n_70)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_70),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_20),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_71),
.Y(n_145)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_60),
.Y(n_72)
);

BUFx2_ASAP7_75t_L g160 ( 
.A(n_72),
.Y(n_160)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_30),
.Y(n_73)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_73),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_20),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_74),
.Y(n_147)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_30),
.Y(n_75)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_75),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_26),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_76),
.Y(n_164)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_26),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_77),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_26),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_78),
.Y(n_187)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_28),
.Y(n_79)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_79),
.Y(n_146)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_30),
.Y(n_80)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_80),
.Y(n_135)
);

BUFx12f_ASAP7_75t_L g81 ( 
.A(n_60),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g197 ( 
.A(n_81),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_40),
.B(n_7),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_32),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_83),
.Y(n_203)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_32),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_84),
.Y(n_211)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_33),
.Y(n_85)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_85),
.Y(n_149)
);

INVx11_ASAP7_75t_L g86 ( 
.A(n_56),
.Y(n_86)
);

INVx8_ASAP7_75t_L g167 ( 
.A(n_86),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_32),
.Y(n_87)
);

INVx6_ASAP7_75t_L g139 ( 
.A(n_87),
.Y(n_139)
);

BUFx24_ASAP7_75t_L g88 ( 
.A(n_38),
.Y(n_88)
);

INVx3_ASAP7_75t_SL g152 ( 
.A(n_88),
.Y(n_152)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_36),
.Y(n_89)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_89),
.Y(n_158)
);

NAND2xp33_ASAP7_75t_SL g90 ( 
.A(n_39),
.B(n_18),
.Y(n_90)
);

NAND2xp33_ASAP7_75t_SL g154 ( 
.A(n_90),
.B(n_121),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_48),
.Y(n_91)
);

INVx6_ASAP7_75t_L g189 ( 
.A(n_91),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_48),
.Y(n_92)
);

INVx3_ASAP7_75t_SL g162 ( 
.A(n_92),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_21),
.B(n_18),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_39),
.B(n_7),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_94),
.B(n_126),
.Y(n_192)
);

BUFx2_ASAP7_75t_L g95 ( 
.A(n_31),
.Y(n_95)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_95),
.Y(n_150)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_24),
.Y(n_96)
);

INVx5_ASAP7_75t_L g132 ( 
.A(n_96),
.Y(n_132)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_28),
.Y(n_97)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_97),
.Y(n_151)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_48),
.Y(n_98)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_98),
.Y(n_173)
);

INVx13_ASAP7_75t_L g99 ( 
.A(n_58),
.Y(n_99)
);

INVx2_ASAP7_75t_SL g133 ( 
.A(n_99),
.Y(n_133)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_34),
.Y(n_100)
);

INVx5_ASAP7_75t_L g161 ( 
.A(n_100),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_51),
.Y(n_101)
);

INVx5_ASAP7_75t_L g166 ( 
.A(n_101),
.Y(n_166)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_42),
.Y(n_102)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_102),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_51),
.Y(n_103)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_103),
.Y(n_159)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_42),
.Y(n_104)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_104),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_51),
.Y(n_105)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_105),
.Y(n_176)
);

BUFx2_ASAP7_75t_L g106 ( 
.A(n_31),
.Y(n_106)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_106),
.Y(n_181)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_34),
.Y(n_107)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_107),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_54),
.Y(n_108)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_108),
.Y(n_178)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_47),
.Y(n_109)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_109),
.Y(n_186)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_24),
.Y(n_110)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_110),
.Y(n_142)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_27),
.Y(n_111)
);

INVx4_ASAP7_75t_L g206 ( 
.A(n_111),
.Y(n_206)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_43),
.Y(n_112)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_112),
.Y(n_188)
);

INVx11_ASAP7_75t_L g113 ( 
.A(n_58),
.Y(n_113)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_113),
.Y(n_195)
);

INVx8_ASAP7_75t_L g114 ( 
.A(n_43),
.Y(n_114)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_114),
.Y(n_148)
);

INVx8_ASAP7_75t_L g115 ( 
.A(n_59),
.Y(n_115)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_115),
.Y(n_157)
);

BUFx12f_ASAP7_75t_L g116 ( 
.A(n_22),
.Y(n_116)
);

INVx4_ASAP7_75t_L g199 ( 
.A(n_116),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_54),
.Y(n_117)
);

INVx4_ASAP7_75t_L g210 ( 
.A(n_117),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_59),
.Y(n_118)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_118),
.Y(n_190)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_27),
.Y(n_119)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_119),
.Y(n_193)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_36),
.Y(n_120)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_120),
.Y(n_174)
);

BUFx3_ASAP7_75t_L g121 ( 
.A(n_27),
.Y(n_121)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_27),
.Y(n_122)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_122),
.Y(n_194)
);

INVx8_ASAP7_75t_L g123 ( 
.A(n_57),
.Y(n_123)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_123),
.Y(n_202)
);

INVx5_ASAP7_75t_L g124 ( 
.A(n_57),
.Y(n_124)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_124),
.Y(n_204)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_37),
.Y(n_125)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_125),
.Y(n_182)
);

BUFx12f_ASAP7_75t_L g126 ( 
.A(n_22),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_47),
.Y(n_127)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_127),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_47),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_128),
.B(n_47),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_94),
.A2(n_23),
.B1(n_52),
.B2(n_49),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_129),
.A2(n_170),
.B1(n_41),
.B2(n_35),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_88),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_134),
.B(n_143),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_65),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_82),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_153),
.B(n_168),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_112),
.A2(n_23),
.B1(n_52),
.B2(n_49),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_155),
.A2(n_83),
.B1(n_76),
.B2(n_101),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_95),
.A2(n_29),
.B1(n_50),
.B2(n_46),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g268 ( 
.A(n_156),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_72),
.A2(n_106),
.B1(n_123),
.B2(n_81),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_163),
.A2(n_171),
.B1(n_185),
.B2(n_200),
.Y(n_243)
);

AND2x2_ASAP7_75t_L g239 ( 
.A(n_165),
.B(n_172),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_99),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_116),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_169),
.B(n_201),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_L g170 ( 
.A1(n_107),
.A2(n_61),
.B1(n_55),
.B2(n_35),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_81),
.A2(n_29),
.B1(n_50),
.B2(n_46),
.Y(n_171)
);

AND2x2_ASAP7_75t_SL g172 ( 
.A(n_116),
.B(n_29),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_126),
.B(n_21),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_175),
.B(n_205),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_100),
.A2(n_29),
.B1(n_46),
.B2(n_50),
.Y(n_185)
);

AO22x2_ASAP7_75t_L g191 ( 
.A1(n_77),
.A2(n_61),
.B1(n_55),
.B2(n_41),
.Y(n_191)
);

AO22x2_ASAP7_75t_L g270 ( 
.A1(n_191),
.A2(n_1),
.B1(n_17),
.B2(n_5),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_114),
.A2(n_50),
.B1(n_46),
.B2(n_53),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_126),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_98),
.B(n_53),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_115),
.B(n_45),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_208),
.B(n_209),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_127),
.Y(n_209)
);

BUFx12f_ASAP7_75t_L g212 ( 
.A(n_197),
.Y(n_212)
);

INVx1_ASAP7_75t_SL g302 ( 
.A(n_212),
.Y(n_302)
);

BUFx3_ASAP7_75t_L g213 ( 
.A(n_197),
.Y(n_213)
);

INVx3_ASAP7_75t_L g287 ( 
.A(n_213),
.Y(n_287)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_137),
.Y(n_214)
);

INVx1_ASAP7_75t_SL g330 ( 
.A(n_214),
.Y(n_330)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_167),
.Y(n_215)
);

HB1xp67_ASAP7_75t_L g308 ( 
.A(n_215),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_144),
.B(n_45),
.Y(n_216)
);

NAND3xp33_ASAP7_75t_L g339 ( 
.A(n_216),
.B(n_249),
.C(n_252),
.Y(n_339)
);

INVx6_ASAP7_75t_L g218 ( 
.A(n_164),
.Y(n_218)
);

INVx3_ASAP7_75t_L g301 ( 
.A(n_218),
.Y(n_301)
);

BUFx2_ASAP7_75t_L g219 ( 
.A(n_161),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g342 ( 
.A(n_219),
.Y(n_342)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_138),
.Y(n_222)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_222),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_149),
.B(n_128),
.C(n_118),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_223),
.B(n_271),
.C(n_162),
.Y(n_334)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_158),
.Y(n_224)
);

BUFx2_ASAP7_75t_SL g315 ( 
.A(n_224),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_225),
.A2(n_284),
.B1(n_162),
.B2(n_189),
.Y(n_291)
);

INVx5_ASAP7_75t_L g226 ( 
.A(n_178),
.Y(n_226)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_226),
.Y(n_304)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_140),
.Y(n_227)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_227),
.Y(n_306)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_141),
.Y(n_228)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_228),
.Y(n_331)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_164),
.Y(n_229)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_229),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_196),
.B(n_37),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g316 ( 
.A(n_230),
.B(n_234),
.Y(n_316)
);

INVx4_ASAP7_75t_L g231 ( 
.A(n_148),
.Y(n_231)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_231),
.Y(n_340)
);

INVx4_ASAP7_75t_L g232 ( 
.A(n_157),
.Y(n_232)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_232),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_192),
.A2(n_87),
.B1(n_105),
.B2(n_103),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_233),
.A2(n_256),
.B1(n_257),
.B2(n_273),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_196),
.B(n_17),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_173),
.Y(n_235)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_235),
.Y(n_290)
);

BUFx2_ASAP7_75t_L g236 ( 
.A(n_132),
.Y(n_236)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_236),
.Y(n_293)
);

INVx1_ASAP7_75t_SL g237 ( 
.A(n_172),
.Y(n_237)
);

AND2x2_ASAP7_75t_L g311 ( 
.A(n_237),
.B(n_244),
.Y(n_311)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_174),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_238),
.B(n_240),
.Y(n_288)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_182),
.Y(n_240)
);

INVx4_ASAP7_75t_L g241 ( 
.A(n_150),
.Y(n_241)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_241),
.Y(n_312)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_183),
.Y(n_242)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_242),
.Y(n_319)
);

INVx1_ASAP7_75t_SL g244 ( 
.A(n_160),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_186),
.Y(n_245)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_245),
.Y(n_323)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_146),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_246),
.B(n_260),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_247),
.A2(n_203),
.B1(n_147),
.B2(n_195),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_191),
.B(n_15),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_SL g250 ( 
.A1(n_160),
.A2(n_108),
.B1(n_117),
.B2(n_210),
.Y(n_250)
);

OAI22x1_ASAP7_75t_L g324 ( 
.A1(n_250),
.A2(n_254),
.B1(n_275),
.B2(n_279),
.Y(n_324)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_190),
.Y(n_251)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_251),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_191),
.B(n_14),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_187),
.Y(n_253)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_253),
.Y(n_337)
);

AOI22xp33_ASAP7_75t_SL g254 ( 
.A1(n_178),
.A2(n_74),
.B1(n_71),
.B2(n_66),
.Y(n_254)
);

AND2x2_ASAP7_75t_L g255 ( 
.A(n_152),
.B(n_91),
.Y(n_255)
);

CKINVDCx14_ASAP7_75t_R g327 ( 
.A(n_255),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_185),
.A2(n_92),
.B1(n_78),
.B2(n_2),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_170),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_257)
);

AND2x4_ASAP7_75t_SL g259 ( 
.A(n_154),
.B(n_0),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g296 ( 
.A(n_259),
.Y(n_296)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_151),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_198),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_261),
.B(n_265),
.Y(n_299)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_188),
.Y(n_262)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_262),
.Y(n_344)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_177),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_263),
.B(n_264),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_180),
.B(n_10),
.Y(n_264)
);

AND2x2_ASAP7_75t_L g265 ( 
.A(n_152),
.B(n_17),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_130),
.B(n_131),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_266),
.B(n_269),
.Y(n_314)
);

INVx4_ASAP7_75t_L g267 ( 
.A(n_181),
.Y(n_267)
);

INVx11_ASAP7_75t_L g321 ( 
.A(n_267),
.Y(n_321)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_207),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_270),
.B(n_17),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_142),
.B(n_10),
.C(n_4),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_199),
.B(n_12),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_272),
.B(n_274),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_200),
.A2(n_1),
.B1(n_5),
.B2(n_6),
.Y(n_273)
);

INVx1_ASAP7_75t_SL g274 ( 
.A(n_135),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_SL g275 ( 
.A1(n_210),
.A2(n_6),
.B1(n_10),
.B2(n_12),
.Y(n_275)
);

INVx6_ASAP7_75t_L g276 ( 
.A(n_187),
.Y(n_276)
);

INVxp33_ASAP7_75t_L g313 ( 
.A(n_276),
.Y(n_313)
);

INVx3_ASAP7_75t_L g277 ( 
.A(n_202),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_277),
.Y(n_295)
);

BUFx3_ASAP7_75t_L g278 ( 
.A(n_133),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_278),
.B(n_280),
.Y(n_328)
);

AOI22xp33_ASAP7_75t_SL g279 ( 
.A1(n_204),
.A2(n_6),
.B1(n_15),
.B2(n_16),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_194),
.Y(n_280)
);

INVx1_ASAP7_75t_SL g281 ( 
.A(n_193),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_281),
.B(n_282),
.Y(n_343)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_133),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_159),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_283),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_163),
.A2(n_1),
.B1(n_15),
.B2(n_16),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_159),
.Y(n_285)
);

AOI22xp33_ASAP7_75t_SL g338 ( 
.A1(n_285),
.A2(n_195),
.B1(n_147),
.B2(n_145),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_L g371 ( 
.A1(n_291),
.A2(n_292),
.B1(n_303),
.B2(n_244),
.Y(n_371)
);

AOI22xp33_ASAP7_75t_L g292 ( 
.A1(n_268),
.A2(n_176),
.B1(n_189),
.B2(n_139),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_220),
.B(n_199),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_298),
.B(n_310),
.Y(n_346)
);

AOI22xp33_ASAP7_75t_L g303 ( 
.A1(n_257),
.A2(n_176),
.B1(n_139),
.B2(n_211),
.Y(n_303)
);

AND2x2_ASAP7_75t_L g350 ( 
.A(n_305),
.B(n_334),
.Y(n_350)
);

OAI32xp33_ASAP7_75t_L g307 ( 
.A1(n_221),
.A2(n_167),
.A3(n_211),
.B1(n_179),
.B2(n_206),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_307),
.B(n_203),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_259),
.B(n_239),
.Y(n_310)
);

O2A1O1Ixp33_ASAP7_75t_L g317 ( 
.A1(n_259),
.A2(n_184),
.B(n_198),
.C(n_171),
.Y(n_317)
);

A2O1A1Ixp33_ASAP7_75t_SL g354 ( 
.A1(n_317),
.A2(n_256),
.B(n_284),
.C(n_254),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_239),
.B(n_179),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g353 ( 
.A(n_318),
.B(n_322),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_270),
.B(n_136),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_217),
.B(n_166),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_SL g375 ( 
.A(n_325),
.B(n_278),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_270),
.B(n_223),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_326),
.B(n_329),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_270),
.B(n_136),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_237),
.B(n_145),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g369 ( 
.A(n_332),
.B(n_215),
.Y(n_369)
);

AOI21xp5_ASAP7_75t_L g333 ( 
.A1(n_243),
.A2(n_184),
.B(n_198),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_L g345 ( 
.A1(n_333),
.A2(n_243),
.B(n_250),
.Y(n_345)
);

INVxp67_ASAP7_75t_L g352 ( 
.A(n_338),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_341),
.A2(n_255),
.B1(n_276),
.B2(n_218),
.Y(n_358)
);

OAI21xp5_ASAP7_75t_SL g409 ( 
.A1(n_345),
.A2(n_354),
.B(n_311),
.Y(n_409)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_290),
.Y(n_347)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_347),
.Y(n_393)
);

INVx5_ASAP7_75t_L g348 ( 
.A(n_301),
.Y(n_348)
);

INVx3_ASAP7_75t_L g404 ( 
.A(n_348),
.Y(n_404)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_290),
.Y(n_349)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_349),
.Y(n_403)
);

INVx4_ASAP7_75t_L g351 ( 
.A(n_301),
.Y(n_351)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_351),
.Y(n_421)
);

INVx3_ASAP7_75t_L g355 ( 
.A(n_335),
.Y(n_355)
);

INVx2_ASAP7_75t_SL g390 ( 
.A(n_355),
.Y(n_390)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_319),
.Y(n_356)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_356),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_L g357 ( 
.A1(n_294),
.A2(n_247),
.B1(n_275),
.B2(n_248),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_357),
.A2(n_368),
.B1(n_370),
.B2(n_379),
.Y(n_405)
);

AND2x2_ASAP7_75t_L g396 ( 
.A(n_358),
.B(n_363),
.Y(n_396)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_319),
.Y(n_359)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_359),
.Y(n_420)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_344),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_361),
.B(n_364),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_322),
.A2(n_273),
.B1(n_232),
.B2(n_231),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_L g399 ( 
.A1(n_362),
.A2(n_365),
.B1(n_381),
.B2(n_358),
.Y(n_399)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_344),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_329),
.A2(n_277),
.B1(n_262),
.B2(n_242),
.Y(n_365)
);

OAI21xp33_ASAP7_75t_L g366 ( 
.A1(n_310),
.A2(n_265),
.B(n_258),
.Y(n_366)
);

INVxp67_ASAP7_75t_L g397 ( 
.A(n_366),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_325),
.B(n_274),
.Y(n_367)
);

INVxp67_ASAP7_75t_L g425 ( 
.A(n_367),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_326),
.A2(n_279),
.B1(n_271),
.B2(n_235),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_SL g394 ( 
.A(n_369),
.B(n_318),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_294),
.A2(n_253),
.B1(n_229),
.B2(n_283),
.Y(n_370)
);

AOI22xp33_ASAP7_75t_L g398 ( 
.A1(n_371),
.A2(n_377),
.B1(n_330),
.B2(n_314),
.Y(n_398)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_315),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_372),
.B(n_373),
.Y(n_411)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_293),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_288),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_374),
.B(n_378),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_SL g400 ( 
.A(n_375),
.B(n_376),
.Y(n_400)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_323),
.Y(n_376)
);

INVxp33_ASAP7_75t_L g377 ( 
.A(n_343),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_323),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_SL g379 ( 
.A1(n_291),
.A2(n_267),
.B1(n_241),
.B2(n_219),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_293),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_380),
.B(n_382),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_341),
.A2(n_226),
.B1(n_281),
.B2(n_236),
.Y(n_381)
);

INVxp67_ASAP7_75t_L g382 ( 
.A(n_328),
.Y(n_382)
);

XOR2xp5_ASAP7_75t_L g383 ( 
.A(n_298),
.B(n_213),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_383),
.B(n_311),
.C(n_314),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_288),
.B(n_212),
.Y(n_384)
);

CKINVDCx16_ASAP7_75t_R g419 ( 
.A(n_384),
.Y(n_419)
);

OAI22xp33_ASAP7_75t_SL g385 ( 
.A1(n_307),
.A2(n_333),
.B1(n_339),
.B2(n_334),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_SL g412 ( 
.A1(n_385),
.A2(n_350),
.B1(n_368),
.B2(n_346),
.Y(n_412)
);

OAI21xp5_ASAP7_75t_SL g386 ( 
.A1(n_296),
.A2(n_212),
.B(n_327),
.Y(n_386)
);

OAI21xp5_ASAP7_75t_L g401 ( 
.A1(n_386),
.A2(n_317),
.B(n_311),
.Y(n_401)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_336),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_387),
.B(n_295),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_316),
.B(n_330),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_388),
.Y(n_395)
);

HB1xp67_ASAP7_75t_L g389 ( 
.A(n_286),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_389),
.Y(n_418)
);

XNOR2x1_ASAP7_75t_SL g392 ( 
.A(n_350),
.B(n_296),
.Y(n_392)
);

XOR2xp5_ASAP7_75t_L g433 ( 
.A(n_392),
.B(n_394),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_398),
.B(n_379),
.Y(n_446)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_399),
.Y(n_432)
);

OAI21xp5_ASAP7_75t_SL g444 ( 
.A1(n_401),
.A2(n_412),
.B(n_423),
.Y(n_444)
);

AOI22xp33_ASAP7_75t_SL g406 ( 
.A1(n_352),
.A2(n_324),
.B1(n_287),
.B2(n_286),
.Y(n_406)
);

OAI22x1_ASAP7_75t_L g451 ( 
.A1(n_406),
.A2(n_354),
.B1(n_287),
.B2(n_351),
.Y(n_451)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_357),
.A2(n_324),
.B1(n_305),
.B2(n_332),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_SL g448 ( 
.A1(n_408),
.A2(n_415),
.B1(n_424),
.B2(n_381),
.Y(n_448)
);

AOI21xp5_ASAP7_75t_L g430 ( 
.A1(n_409),
.A2(n_426),
.B(n_369),
.Y(n_430)
);

XOR2xp5_ASAP7_75t_L g410 ( 
.A(n_360),
.B(n_297),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_410),
.B(n_427),
.C(n_386),
.Y(n_429)
);

XOR2xp5_ASAP7_75t_L g436 ( 
.A(n_413),
.B(n_427),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_L g414 ( 
.A1(n_362),
.A2(n_320),
.B1(n_297),
.B2(n_299),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_414),
.A2(n_422),
.B1(n_382),
.B2(n_375),
.Y(n_440)
);

AOI22xp5_ASAP7_75t_L g415 ( 
.A1(n_370),
.A2(n_313),
.B1(n_337),
.B2(n_295),
.Y(n_415)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_417),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_L g422 ( 
.A1(n_353),
.A2(n_320),
.B1(n_337),
.B2(n_289),
.Y(n_422)
);

OAI21xp33_ASAP7_75t_SL g423 ( 
.A1(n_345),
.A2(n_352),
.B(n_346),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_350),
.A2(n_335),
.B1(n_340),
.B2(n_309),
.Y(n_424)
);

NAND2x1p5_ASAP7_75t_L g426 ( 
.A(n_360),
.B(n_289),
.Y(n_426)
);

XOR2xp5_ASAP7_75t_L g427 ( 
.A(n_383),
.B(n_308),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_SL g428 ( 
.A(n_395),
.B(n_374),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_SL g464 ( 
.A(n_428),
.B(n_442),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_L g475 ( 
.A(n_429),
.B(n_413),
.Y(n_475)
);

OAI21xp5_ASAP7_75t_SL g478 ( 
.A1(n_430),
.A2(n_451),
.B(n_405),
.Y(n_478)
);

CKINVDCx16_ASAP7_75t_R g431 ( 
.A(n_417),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_431),
.B(n_434),
.Y(n_477)
);

CKINVDCx14_ASAP7_75t_R g434 ( 
.A(n_400),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_436),
.B(n_445),
.C(n_452),
.Y(n_469)
);

CKINVDCx16_ASAP7_75t_R g437 ( 
.A(n_411),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_437),
.B(n_441),
.Y(n_484)
);

BUFx12f_ASAP7_75t_L g438 ( 
.A(n_418),
.Y(n_438)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_438),
.Y(n_489)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_402),
.Y(n_439)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_439),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_SL g482 ( 
.A(n_440),
.B(n_422),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_391),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_391),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_402),
.Y(n_443)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_443),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_394),
.B(n_354),
.C(n_387),
.Y(n_445)
);

INVxp67_ASAP7_75t_L g466 ( 
.A(n_446),
.Y(n_466)
);

AOI22xp5_ASAP7_75t_L g447 ( 
.A1(n_396),
.A2(n_354),
.B1(n_365),
.B2(n_349),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_SL g479 ( 
.A1(n_447),
.A2(n_424),
.B1(n_415),
.B2(n_416),
.Y(n_479)
);

AOI22xp5_ASAP7_75t_L g493 ( 
.A1(n_448),
.A2(n_456),
.B1(n_399),
.B2(n_419),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_SL g449 ( 
.A(n_395),
.B(n_372),
.Y(n_449)
);

INVxp67_ASAP7_75t_L g472 ( 
.A(n_449),
.Y(n_472)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_393),
.Y(n_450)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_450),
.Y(n_476)
);

XNOR2xp5_ASAP7_75t_L g452 ( 
.A(n_410),
.B(n_376),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_416),
.Y(n_453)
);

CKINVDCx20_ASAP7_75t_R g491 ( 
.A(n_453),
.Y(n_491)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_393),
.Y(n_454)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_454),
.Y(n_483)
);

OAI32xp33_ASAP7_75t_L g455 ( 
.A1(n_396),
.A2(n_378),
.A3(n_354),
.B1(n_347),
.B2(n_361),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_455),
.B(n_457),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_SL g456 ( 
.A1(n_408),
.A2(n_359),
.B1(n_364),
.B2(n_356),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_403),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_L g458 ( 
.A(n_392),
.B(n_336),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_458),
.B(n_459),
.C(n_426),
.Y(n_487)
);

XOR2xp5_ASAP7_75t_L g459 ( 
.A(n_394),
.B(n_312),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_403),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_460),
.B(n_461),
.Y(n_474)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_420),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_420),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_462),
.B(n_461),
.Y(n_486)
);

AOI21xp5_ASAP7_75t_L g463 ( 
.A1(n_444),
.A2(n_409),
.B(n_401),
.Y(n_463)
);

OAI21xp5_ASAP7_75t_SL g499 ( 
.A1(n_463),
.A2(n_492),
.B(n_460),
.Y(n_499)
);

BUFx24_ASAP7_75t_SL g465 ( 
.A(n_440),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_465),
.B(n_456),
.Y(n_500)
);

OAI22xp5_ASAP7_75t_L g471 ( 
.A1(n_432),
.A2(n_405),
.B1(n_412),
.B2(n_423),
.Y(n_471)
);

AOI22xp5_ASAP7_75t_L g517 ( 
.A1(n_471),
.A2(n_479),
.B1(n_480),
.B2(n_485),
.Y(n_517)
);

CKINVDCx16_ASAP7_75t_R g473 ( 
.A(n_447),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_473),
.B(n_455),
.Y(n_503)
);

XOR2xp5_ASAP7_75t_L g501 ( 
.A(n_475),
.B(n_487),
.Y(n_501)
);

AOI21xp5_ASAP7_75t_L g514 ( 
.A1(n_478),
.A2(n_481),
.B(n_463),
.Y(n_514)
);

OAI22xp5_ASAP7_75t_SL g480 ( 
.A1(n_432),
.A2(n_445),
.B1(n_435),
.B2(n_430),
.Y(n_480)
);

OAI21xp5_ASAP7_75t_L g481 ( 
.A1(n_444),
.A2(n_396),
.B(n_400),
.Y(n_481)
);

OAI22xp5_ASAP7_75t_L g494 ( 
.A1(n_482),
.A2(n_493),
.B1(n_446),
.B2(n_448),
.Y(n_494)
);

OAI22xp5_ASAP7_75t_L g485 ( 
.A1(n_435),
.A2(n_425),
.B1(n_419),
.B2(n_418),
.Y(n_485)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_486),
.Y(n_512)
);

XNOR2xp5_ASAP7_75t_L g488 ( 
.A(n_436),
.B(n_426),
.Y(n_488)
);

XOR2xp5_ASAP7_75t_L g520 ( 
.A(n_488),
.B(n_312),
.Y(n_520)
);

HB1xp67_ASAP7_75t_L g490 ( 
.A(n_439),
.Y(n_490)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_490),
.Y(n_498)
);

AND2x2_ASAP7_75t_L g492 ( 
.A(n_443),
.B(n_411),
.Y(n_492)
);

AOI22xp5_ASAP7_75t_L g527 ( 
.A1(n_494),
.A2(n_479),
.B1(n_466),
.B2(n_470),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_469),
.B(n_429),
.C(n_459),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_495),
.B(n_502),
.C(n_508),
.Y(n_523)
);

XNOR2xp5_ASAP7_75t_L g496 ( 
.A(n_469),
.B(n_452),
.Y(n_496)
);

XNOR2xp5_ASAP7_75t_L g538 ( 
.A(n_496),
.B(n_509),
.Y(n_538)
);

OAI22xp5_ASAP7_75t_L g497 ( 
.A1(n_472),
.A2(n_397),
.B1(n_462),
.B2(n_454),
.Y(n_497)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_497),
.Y(n_526)
);

XOR2xp5_ASAP7_75t_L g534 ( 
.A(n_499),
.B(n_507),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_SL g529 ( 
.A(n_500),
.B(n_505),
.Y(n_529)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_475),
.B(n_458),
.C(n_433),
.Y(n_502)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_503),
.Y(n_530)
);

OAI22xp5_ASAP7_75t_L g504 ( 
.A1(n_493),
.A2(n_464),
.B1(n_482),
.B2(n_477),
.Y(n_504)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_504),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_464),
.B(n_414),
.Y(n_505)
);

INVxp67_ASAP7_75t_SL g506 ( 
.A(n_484),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_506),
.B(n_518),
.Y(n_535)
);

XNOR2xp5_ASAP7_75t_SL g507 ( 
.A(n_488),
.B(n_433),
.Y(n_507)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_487),
.B(n_451),
.C(n_407),
.Y(n_508)
);

XNOR2xp5_ASAP7_75t_L g509 ( 
.A(n_480),
.B(n_457),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_491),
.B(n_438),
.Y(n_510)
);

CKINVDCx20_ASAP7_75t_R g528 ( 
.A(n_510),
.Y(n_528)
);

XNOR2xp5_ASAP7_75t_SL g511 ( 
.A(n_471),
.B(n_468),
.Y(n_511)
);

XOR2xp5_ASAP7_75t_L g536 ( 
.A(n_511),
.B(n_514),
.Y(n_536)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_485),
.B(n_407),
.C(n_450),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_513),
.B(n_515),
.C(n_519),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_492),
.B(n_421),
.C(n_404),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_474),
.Y(n_516)
);

INVx1_ASAP7_75t_SL g543 ( 
.A(n_516),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_SL g518 ( 
.A(n_491),
.B(n_316),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_492),
.B(n_421),
.C(n_404),
.Y(n_519)
);

XOR2xp5_ASAP7_75t_L g540 ( 
.A(n_520),
.B(n_483),
.Y(n_540)
);

AOI21xp5_ASAP7_75t_L g521 ( 
.A1(n_478),
.A2(n_438),
.B(n_390),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_521),
.B(n_489),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_510),
.B(n_467),
.Y(n_522)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_522),
.Y(n_547)
);

OAI22x1_ASAP7_75t_L g525 ( 
.A1(n_517),
.A2(n_473),
.B1(n_468),
.B2(n_467),
.Y(n_525)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_525),
.Y(n_552)
);

OAI22xp5_ASAP7_75t_SL g560 ( 
.A1(n_527),
.A2(n_539),
.B1(n_543),
.B2(n_522),
.Y(n_560)
);

OAI22xp5_ASAP7_75t_SL g531 ( 
.A1(n_517),
.A2(n_481),
.B1(n_470),
.B2(n_486),
.Y(n_531)
);

AOI22xp5_ASAP7_75t_L g545 ( 
.A1(n_531),
.A2(n_541),
.B1(n_542),
.B2(n_498),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_498),
.B(n_489),
.Y(n_533)
);

CKINVDCx20_ASAP7_75t_R g562 ( 
.A(n_533),
.Y(n_562)
);

AOI21x1_ASAP7_75t_SL g548 ( 
.A1(n_537),
.A2(n_499),
.B(n_533),
.Y(n_548)
);

AOI22xp5_ASAP7_75t_L g539 ( 
.A1(n_512),
.A2(n_474),
.B1(n_476),
.B2(n_483),
.Y(n_539)
);

XOR2xp5_ASAP7_75t_L g549 ( 
.A(n_540),
.B(n_520),
.Y(n_549)
);

OAI22xp5_ASAP7_75t_SL g541 ( 
.A1(n_503),
.A2(n_476),
.B1(n_438),
.B2(n_390),
.Y(n_541)
);

OAI22xp5_ASAP7_75t_SL g542 ( 
.A1(n_516),
.A2(n_390),
.B1(n_380),
.B2(n_373),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g544 ( 
.A(n_509),
.B(n_348),
.Y(n_544)
);

CKINVDCx14_ASAP7_75t_R g555 ( 
.A(n_544),
.Y(n_555)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_545),
.Y(n_565)
);

AOI22xp5_ASAP7_75t_L g546 ( 
.A1(n_532),
.A2(n_508),
.B1(n_513),
.B2(n_511),
.Y(n_546)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_546),
.Y(n_568)
);

INVx11_ASAP7_75t_L g577 ( 
.A(n_548),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_L g564 ( 
.A(n_549),
.B(n_560),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_524),
.B(n_529),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_SL g578 ( 
.A(n_550),
.B(n_557),
.Y(n_578)
);

MAJIxp5_ASAP7_75t_L g551 ( 
.A(n_524),
.B(n_501),
.C(n_496),
.Y(n_551)
);

MAJIxp5_ASAP7_75t_L g569 ( 
.A(n_551),
.B(n_554),
.C(n_556),
.Y(n_569)
);

XNOR2xp5_ASAP7_75t_L g553 ( 
.A(n_538),
.B(n_501),
.Y(n_553)
);

NOR2xp33_ASAP7_75t_L g579 ( 
.A(n_553),
.B(n_558),
.Y(n_579)
);

XOR2xp5_ASAP7_75t_L g554 ( 
.A(n_538),
.B(n_507),
.Y(n_554)
);

MAJIxp5_ASAP7_75t_L g556 ( 
.A(n_523),
.B(n_495),
.C(n_540),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_535),
.B(n_519),
.Y(n_557)
);

XNOR2xp5_ASAP7_75t_L g558 ( 
.A(n_523),
.B(n_502),
.Y(n_558)
);

XOR2xp5_ASAP7_75t_L g559 ( 
.A(n_534),
.B(n_514),
.Y(n_559)
);

MAJIxp5_ASAP7_75t_L g572 ( 
.A(n_559),
.B(n_534),
.C(n_525),
.Y(n_572)
);

OA22x2_ASAP7_75t_L g561 ( 
.A1(n_528),
.A2(n_521),
.B1(n_515),
.B2(n_355),
.Y(n_561)
);

NOR2xp33_ASAP7_75t_L g566 ( 
.A(n_561),
.B(n_563),
.Y(n_566)
);

AOI22xp5_ASAP7_75t_L g563 ( 
.A1(n_532),
.A2(n_340),
.B1(n_342),
.B2(n_309),
.Y(n_563)
);

AOI21xp5_ASAP7_75t_L g567 ( 
.A1(n_552),
.A2(n_526),
.B(n_530),
.Y(n_567)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_567),
.Y(n_582)
);

NOR2xp67_ASAP7_75t_R g570 ( 
.A(n_562),
.B(n_543),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_SL g585 ( 
.A(n_570),
.B(n_571),
.Y(n_585)
);

NOR2xp33_ASAP7_75t_L g571 ( 
.A(n_555),
.B(n_531),
.Y(n_571)
);

MAJx2_ASAP7_75t_L g583 ( 
.A(n_572),
.B(n_561),
.C(n_559),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_L g573 ( 
.A(n_556),
.B(n_551),
.Y(n_573)
);

NOR2xp33_ASAP7_75t_SL g588 ( 
.A(n_573),
.B(n_554),
.Y(n_588)
);

AOI21xp5_ASAP7_75t_L g574 ( 
.A1(n_547),
.A2(n_530),
.B(n_536),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_574),
.B(n_302),
.Y(n_589)
);

MAJIxp5_ASAP7_75t_L g575 ( 
.A(n_553),
.B(n_536),
.C(n_541),
.Y(n_575)
);

MAJIxp5_ASAP7_75t_L g587 ( 
.A(n_575),
.B(n_576),
.C(n_549),
.Y(n_587)
);

MAJIxp5_ASAP7_75t_L g576 ( 
.A(n_558),
.B(n_527),
.C(n_539),
.Y(n_576)
);

NOR2xp33_ASAP7_75t_L g580 ( 
.A(n_578),
.B(n_546),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_580),
.B(n_581),
.Y(n_593)
);

NOR2xp33_ASAP7_75t_L g581 ( 
.A(n_578),
.B(n_563),
.Y(n_581)
);

AO21x1_ASAP7_75t_L g595 ( 
.A1(n_583),
.A2(n_568),
.B(n_570),
.Y(n_595)
);

AOI22xp5_ASAP7_75t_SL g584 ( 
.A1(n_572),
.A2(n_561),
.B1(n_545),
.B2(n_548),
.Y(n_584)
);

OAI211xp5_ASAP7_75t_L g594 ( 
.A1(n_584),
.A2(n_589),
.B(n_590),
.C(n_574),
.Y(n_594)
);

NOR2xp33_ASAP7_75t_L g586 ( 
.A(n_576),
.B(n_542),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_586),
.B(n_587),
.Y(n_598)
);

NOR2xp33_ASAP7_75t_SL g596 ( 
.A(n_588),
.B(n_579),
.Y(n_596)
);

INVx11_ASAP7_75t_L g590 ( 
.A(n_577),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_565),
.B(n_342),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_SL g592 ( 
.A(n_591),
.B(n_566),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_592),
.B(n_594),
.Y(n_601)
);

AOI21xp5_ASAP7_75t_L g605 ( 
.A1(n_595),
.A2(n_597),
.B(n_599),
.Y(n_605)
);

INVxp33_ASAP7_75t_L g606 ( 
.A(n_596),
.Y(n_606)
);

AOI21xp5_ASAP7_75t_L g597 ( 
.A1(n_590),
.A2(n_568),
.B(n_569),
.Y(n_597)
);

OAI21xp5_ASAP7_75t_L g599 ( 
.A1(n_585),
.A2(n_577),
.B(n_569),
.Y(n_599)
);

NOR2xp33_ASAP7_75t_L g600 ( 
.A(n_582),
.B(n_565),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_L g603 ( 
.A(n_600),
.B(n_564),
.Y(n_603)
);

OAI21xp5_ASAP7_75t_SL g602 ( 
.A1(n_598),
.A2(n_587),
.B(n_584),
.Y(n_602)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_602),
.Y(n_609)
);

MAJIxp5_ASAP7_75t_L g607 ( 
.A(n_603),
.B(n_604),
.C(n_592),
.Y(n_607)
);

MAJIxp5_ASAP7_75t_L g604 ( 
.A(n_593),
.B(n_567),
.C(n_583),
.Y(n_604)
);

AOI21xp5_ASAP7_75t_L g612 ( 
.A1(n_607),
.A2(n_608),
.B(n_610),
.Y(n_612)
);

A2O1A1O1Ixp25_ASAP7_75t_L g608 ( 
.A1(n_601),
.A2(n_575),
.B(n_591),
.C(n_589),
.D(n_321),
.Y(n_608)
);

MAJIxp5_ASAP7_75t_L g610 ( 
.A(n_606),
.B(n_302),
.C(n_304),
.Y(n_610)
);

MAJIxp5_ASAP7_75t_L g611 ( 
.A(n_609),
.B(n_605),
.C(n_304),
.Y(n_611)
);

A2O1A1Ixp33_ASAP7_75t_L g613 ( 
.A1(n_611),
.A2(n_321),
.B(n_306),
.C(n_300),
.Y(n_613)
);

OAI21xp5_ASAP7_75t_L g614 ( 
.A1(n_613),
.A2(n_612),
.B(n_306),
.Y(n_614)
);

MAJIxp5_ASAP7_75t_L g615 ( 
.A(n_614),
.B(n_300),
.C(n_331),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_SL g616 ( 
.A(n_615),
.B(n_331),
.Y(n_616)
);


endmodule