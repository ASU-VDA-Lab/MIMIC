module fake_ariane_3215_n_2935 (n_295, n_356, n_556, n_170, n_190, n_160, n_64, n_180, n_119, n_124, n_386, n_307, n_516, n_589, n_332, n_581, n_294, n_197, n_463, n_176, n_34, n_404, n_172, n_347, n_423, n_183, n_469, n_479, n_373, n_299, n_541, n_499, n_12, n_564, n_133, n_66, n_205, n_341, n_71, n_109, n_245, n_421, n_96, n_549, n_522, n_319, n_49, n_20, n_416, n_283, n_50, n_187, n_525, n_367, n_345, n_374, n_318, n_103, n_244, n_226, n_220, n_261, n_36, n_370, n_189, n_72, n_286, n_443, n_586, n_57, n_424, n_528, n_584, n_387, n_406, n_117, n_139, n_524, n_85, n_130, n_349, n_391, n_466, n_346, n_214, n_348, n_552, n_2, n_462, n_32, n_410, n_379, n_445, n_515, n_138, n_162, n_264, n_137, n_122, n_198, n_232, n_52, n_441, n_568, n_385, n_73, n_327, n_77, n_372, n_377, n_15, n_396, n_23, n_399, n_554, n_520, n_87, n_279, n_207, n_363, n_354, n_41, n_140, n_419, n_151, n_28, n_146, n_230, n_270, n_194, n_154, n_338, n_142, n_285, n_473, n_186, n_202, n_145, n_193, n_500, n_59, n_336, n_315, n_311, n_239, n_402, n_35, n_272, n_54, n_8, n_339, n_487, n_167, n_90, n_38, n_422, n_47, n_153, n_18, n_269, n_75, n_158, n_69, n_259, n_95, n_446, n_553, n_143, n_566, n_578, n_152, n_405, n_557, n_120, n_169, n_106, n_173, n_242, n_309, n_320, n_115, n_331, n_559, n_401, n_485, n_267, n_495, n_504, n_483, n_335, n_435, n_350, n_291, n_344, n_381, n_426, n_433, n_481, n_398, n_62, n_210, n_200, n_529, n_502, n_166, n_253, n_561, n_218, n_79, n_3, n_271, n_465, n_486, n_507, n_247, n_569, n_567, n_91, n_240, n_369, n_128, n_224, n_44, n_82, n_31, n_547, n_420, n_562, n_518, n_439, n_222, n_478, n_510, n_256, n_326, n_227, n_48, n_188, n_323, n_550, n_330, n_400, n_11, n_129, n_126, n_282, n_328, n_368, n_277, n_248, n_301, n_467, n_432, n_545, n_536, n_293, n_228, n_325, n_276, n_93, n_427, n_108, n_587, n_497, n_303, n_442, n_168, n_81, n_1, n_206, n_352, n_538, n_576, n_511, n_238, n_365, n_429, n_455, n_588, n_136, n_334, n_192, n_488, n_300, n_533, n_505, n_14, n_163, n_88, n_141, n_390, n_498, n_104, n_501, n_438, n_314, n_16, n_440, n_273, n_305, n_539, n_312, n_233, n_56, n_60, n_388, n_333, n_449, n_413, n_392, n_376, n_512, n_579, n_459, n_221, n_321, n_86, n_361, n_458, n_89, n_149, n_383, n_237, n_175, n_453, n_74, n_491, n_19, n_40, n_181, n_570, n_53, n_260, n_362, n_543, n_310, n_236, n_565, n_281, n_24, n_7, n_461, n_209, n_262, n_490, n_17, n_225, n_235, n_464, n_575, n_546, n_297, n_503, n_290, n_527, n_46, n_84, n_371, n_199, n_107, n_217, n_452, n_178, n_42, n_551, n_308, n_417, n_201, n_70, n_572, n_343, n_10, n_414, n_571, n_287, n_302, n_380, n_6, n_582, n_94, n_284, n_4, n_448, n_249, n_534, n_37, n_58, n_65, n_123, n_212, n_355, n_444, n_278, n_255, n_560, n_450, n_257, n_148, n_451, n_475, n_135, n_409, n_171, n_519, n_384, n_468, n_61, n_526, n_102, n_182, n_482, n_316, n_196, n_125, n_43, n_577, n_407, n_13, n_27, n_254, n_476, n_460, n_219, n_55, n_535, n_231, n_366, n_555, n_234, n_492, n_574, n_280, n_215, n_252, n_161, n_454, n_298, n_532, n_68, n_415, n_78, n_63, n_99, n_540, n_216, n_544, n_5, n_514, n_418, n_537, n_223, n_403, n_25, n_83, n_389, n_513, n_288, n_179, n_395, n_195, n_213, n_110, n_304, n_67, n_509, n_583, n_306, n_313, n_92, n_430, n_493, n_203, n_378, n_436, n_150, n_98, n_375, n_113, n_114, n_33, n_324, n_585, n_337, n_437, n_111, n_21, n_274, n_472, n_296, n_265, n_208, n_456, n_156, n_292, n_174, n_275, n_100, n_132, n_147, n_204, n_521, n_51, n_496, n_76, n_342, n_26, n_246, n_517, n_530, n_0, n_428, n_159, n_358, n_105, n_580, n_30, n_494, n_131, n_263, n_434, n_360, n_563, n_229, n_394, n_250, n_165, n_144, n_317, n_101, n_243, n_134, n_329, n_185, n_340, n_289, n_9, n_112, n_45, n_542, n_548, n_523, n_268, n_266, n_470, n_457, n_164, n_157, n_184, n_177, n_477, n_364, n_258, n_425, n_431, n_508, n_118, n_121, n_411, n_484, n_353, n_22, n_241, n_29, n_357, n_412, n_447, n_191, n_382, n_489, n_80, n_480, n_211, n_97, n_408, n_322, n_251, n_506, n_558, n_116, n_397, n_471, n_351, n_39, n_393, n_474, n_359, n_155, n_573, n_127, n_531, n_2935);

input n_295;
input n_356;
input n_556;
input n_170;
input n_190;
input n_160;
input n_64;
input n_180;
input n_119;
input n_124;
input n_386;
input n_307;
input n_516;
input n_589;
input n_332;
input n_581;
input n_294;
input n_197;
input n_463;
input n_176;
input n_34;
input n_404;
input n_172;
input n_347;
input n_423;
input n_183;
input n_469;
input n_479;
input n_373;
input n_299;
input n_541;
input n_499;
input n_12;
input n_564;
input n_133;
input n_66;
input n_205;
input n_341;
input n_71;
input n_109;
input n_245;
input n_421;
input n_96;
input n_549;
input n_522;
input n_319;
input n_49;
input n_20;
input n_416;
input n_283;
input n_50;
input n_187;
input n_525;
input n_367;
input n_345;
input n_374;
input n_318;
input n_103;
input n_244;
input n_226;
input n_220;
input n_261;
input n_36;
input n_370;
input n_189;
input n_72;
input n_286;
input n_443;
input n_586;
input n_57;
input n_424;
input n_528;
input n_584;
input n_387;
input n_406;
input n_117;
input n_139;
input n_524;
input n_85;
input n_130;
input n_349;
input n_391;
input n_466;
input n_346;
input n_214;
input n_348;
input n_552;
input n_2;
input n_462;
input n_32;
input n_410;
input n_379;
input n_445;
input n_515;
input n_138;
input n_162;
input n_264;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_441;
input n_568;
input n_385;
input n_73;
input n_327;
input n_77;
input n_372;
input n_377;
input n_15;
input n_396;
input n_23;
input n_399;
input n_554;
input n_520;
input n_87;
input n_279;
input n_207;
input n_363;
input n_354;
input n_41;
input n_140;
input n_419;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_154;
input n_338;
input n_142;
input n_285;
input n_473;
input n_186;
input n_202;
input n_145;
input n_193;
input n_500;
input n_59;
input n_336;
input n_315;
input n_311;
input n_239;
input n_402;
input n_35;
input n_272;
input n_54;
input n_8;
input n_339;
input n_487;
input n_167;
input n_90;
input n_38;
input n_422;
input n_47;
input n_153;
input n_18;
input n_269;
input n_75;
input n_158;
input n_69;
input n_259;
input n_95;
input n_446;
input n_553;
input n_143;
input n_566;
input n_578;
input n_152;
input n_405;
input n_557;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_309;
input n_320;
input n_115;
input n_331;
input n_559;
input n_401;
input n_485;
input n_267;
input n_495;
input n_504;
input n_483;
input n_335;
input n_435;
input n_350;
input n_291;
input n_344;
input n_381;
input n_426;
input n_433;
input n_481;
input n_398;
input n_62;
input n_210;
input n_200;
input n_529;
input n_502;
input n_166;
input n_253;
input n_561;
input n_218;
input n_79;
input n_3;
input n_271;
input n_465;
input n_486;
input n_507;
input n_247;
input n_569;
input n_567;
input n_91;
input n_240;
input n_369;
input n_128;
input n_224;
input n_44;
input n_82;
input n_31;
input n_547;
input n_420;
input n_562;
input n_518;
input n_439;
input n_222;
input n_478;
input n_510;
input n_256;
input n_326;
input n_227;
input n_48;
input n_188;
input n_323;
input n_550;
input n_330;
input n_400;
input n_11;
input n_129;
input n_126;
input n_282;
input n_328;
input n_368;
input n_277;
input n_248;
input n_301;
input n_467;
input n_432;
input n_545;
input n_536;
input n_293;
input n_228;
input n_325;
input n_276;
input n_93;
input n_427;
input n_108;
input n_587;
input n_497;
input n_303;
input n_442;
input n_168;
input n_81;
input n_1;
input n_206;
input n_352;
input n_538;
input n_576;
input n_511;
input n_238;
input n_365;
input n_429;
input n_455;
input n_588;
input n_136;
input n_334;
input n_192;
input n_488;
input n_300;
input n_533;
input n_505;
input n_14;
input n_163;
input n_88;
input n_141;
input n_390;
input n_498;
input n_104;
input n_501;
input n_438;
input n_314;
input n_16;
input n_440;
input n_273;
input n_305;
input n_539;
input n_312;
input n_233;
input n_56;
input n_60;
input n_388;
input n_333;
input n_449;
input n_413;
input n_392;
input n_376;
input n_512;
input n_579;
input n_459;
input n_221;
input n_321;
input n_86;
input n_361;
input n_458;
input n_89;
input n_149;
input n_383;
input n_237;
input n_175;
input n_453;
input n_74;
input n_491;
input n_19;
input n_40;
input n_181;
input n_570;
input n_53;
input n_260;
input n_362;
input n_543;
input n_310;
input n_236;
input n_565;
input n_281;
input n_24;
input n_7;
input n_461;
input n_209;
input n_262;
input n_490;
input n_17;
input n_225;
input n_235;
input n_464;
input n_575;
input n_546;
input n_297;
input n_503;
input n_290;
input n_527;
input n_46;
input n_84;
input n_371;
input n_199;
input n_107;
input n_217;
input n_452;
input n_178;
input n_42;
input n_551;
input n_308;
input n_417;
input n_201;
input n_70;
input n_572;
input n_343;
input n_10;
input n_414;
input n_571;
input n_287;
input n_302;
input n_380;
input n_6;
input n_582;
input n_94;
input n_284;
input n_4;
input n_448;
input n_249;
input n_534;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_355;
input n_444;
input n_278;
input n_255;
input n_560;
input n_450;
input n_257;
input n_148;
input n_451;
input n_475;
input n_135;
input n_409;
input n_171;
input n_519;
input n_384;
input n_468;
input n_61;
input n_526;
input n_102;
input n_182;
input n_482;
input n_316;
input n_196;
input n_125;
input n_43;
input n_577;
input n_407;
input n_13;
input n_27;
input n_254;
input n_476;
input n_460;
input n_219;
input n_55;
input n_535;
input n_231;
input n_366;
input n_555;
input n_234;
input n_492;
input n_574;
input n_280;
input n_215;
input n_252;
input n_161;
input n_454;
input n_298;
input n_532;
input n_68;
input n_415;
input n_78;
input n_63;
input n_99;
input n_540;
input n_216;
input n_544;
input n_5;
input n_514;
input n_418;
input n_537;
input n_223;
input n_403;
input n_25;
input n_83;
input n_389;
input n_513;
input n_288;
input n_179;
input n_395;
input n_195;
input n_213;
input n_110;
input n_304;
input n_67;
input n_509;
input n_583;
input n_306;
input n_313;
input n_92;
input n_430;
input n_493;
input n_203;
input n_378;
input n_436;
input n_150;
input n_98;
input n_375;
input n_113;
input n_114;
input n_33;
input n_324;
input n_585;
input n_337;
input n_437;
input n_111;
input n_21;
input n_274;
input n_472;
input n_296;
input n_265;
input n_208;
input n_456;
input n_156;
input n_292;
input n_174;
input n_275;
input n_100;
input n_132;
input n_147;
input n_204;
input n_521;
input n_51;
input n_496;
input n_76;
input n_342;
input n_26;
input n_246;
input n_517;
input n_530;
input n_0;
input n_428;
input n_159;
input n_358;
input n_105;
input n_580;
input n_30;
input n_494;
input n_131;
input n_263;
input n_434;
input n_360;
input n_563;
input n_229;
input n_394;
input n_250;
input n_165;
input n_144;
input n_317;
input n_101;
input n_243;
input n_134;
input n_329;
input n_185;
input n_340;
input n_289;
input n_9;
input n_112;
input n_45;
input n_542;
input n_548;
input n_523;
input n_268;
input n_266;
input n_470;
input n_457;
input n_164;
input n_157;
input n_184;
input n_177;
input n_477;
input n_364;
input n_258;
input n_425;
input n_431;
input n_508;
input n_118;
input n_121;
input n_411;
input n_484;
input n_353;
input n_22;
input n_241;
input n_29;
input n_357;
input n_412;
input n_447;
input n_191;
input n_382;
input n_489;
input n_80;
input n_480;
input n_211;
input n_97;
input n_408;
input n_322;
input n_251;
input n_506;
input n_558;
input n_116;
input n_397;
input n_471;
input n_351;
input n_39;
input n_393;
input n_474;
input n_359;
input n_155;
input n_573;
input n_127;
input n_531;

output n_2935;

wire n_2752;
wire n_913;
wire n_1681;
wire n_2163;
wire n_1486;
wire n_1507;
wire n_1938;
wire n_2484;
wire n_2866;
wire n_1174;
wire n_2346;
wire n_1469;
wire n_691;
wire n_1353;
wire n_2679;
wire n_1355;
wire n_2131;
wire n_2559;
wire n_2500;
wire n_2509;
wire n_1383;
wire n_2182;
wire n_603;
wire n_2135;
wire n_2334;
wire n_2680;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_2879;
wire n_610;
wire n_1713;
wire n_1436;
wire n_2407;
wire n_690;
wire n_2818;
wire n_1109;
wire n_1430;
wire n_2537;
wire n_2002;
wire n_1463;
wire n_2243;
wire n_1238;
wire n_2694;
wire n_2011;
wire n_2729;
wire n_1515;
wire n_1837;
wire n_817;
wire n_924;
wire n_781;
wire n_2013;
wire n_2786;
wire n_1566;
wire n_2837;
wire n_717;
wire n_2006;
wire n_952;
wire n_864;
wire n_2446;
wire n_1096;
wire n_1379;
wire n_2436;
wire n_2376;
wire n_2367;
wire n_2671;
wire n_2790;
wire n_1706;
wire n_2207;
wire n_2461;
wire n_2702;
wire n_2731;
wire n_1214;
wire n_634;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_2042;
wire n_2123;
wire n_1853;
wire n_764;
wire n_1503;
wire n_2238;
wire n_2529;
wire n_2374;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_2380;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_2646;
wire n_737;
wire n_1298;
wire n_2653;
wire n_1745;
wire n_2873;
wire n_1366;
wire n_2084;
wire n_2278;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_2482;
wire n_1682;
wire n_2750;
wire n_1836;
wire n_870;
wire n_2547;
wire n_1453;
wire n_958;
wire n_945;
wire n_2554;
wire n_2248;
wire n_813;
wire n_1985;
wire n_2288;
wire n_2621;
wire n_2908;
wire n_995;
wire n_2579;
wire n_1909;
wire n_2156;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_2323;
wire n_1073;
wire n_2844;
wire n_1979;
wire n_1277;
wire n_2107;
wire n_1746;
wire n_1761;
wire n_829;
wire n_1062;
wire n_738;
wire n_1690;
wire n_2221;
wire n_2807;
wire n_672;
wire n_740;
wire n_1283;
wire n_2317;
wire n_2838;
wire n_1974;
wire n_2906;
wire n_1736;
wire n_1018;
wire n_2342;
wire n_2200;
wire n_2781;
wire n_2442;
wire n_2735;
wire n_953;
wire n_1364;
wire n_2390;
wire n_1888;
wire n_1224;
wire n_2109;
wire n_1425;
wire n_2634;
wire n_2709;
wire n_625;
wire n_2322;
wire n_2746;
wire n_1107;
wire n_2832;
wire n_1688;
wire n_989;
wire n_645;
wire n_1944;
wire n_2233;
wire n_2370;
wire n_2663;
wire n_2914;
wire n_1988;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_2149;
wire n_2277;
wire n_1428;
wire n_1284;
wire n_2878;
wire n_1241;
wire n_821;
wire n_770;
wire n_1514;
wire n_2539;
wire n_1528;
wire n_901;
wire n_2782;
wire n_2078;
wire n_1145;
wire n_971;
wire n_2359;
wire n_2201;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_1207;
wire n_786;
wire n_1404;
wire n_868;
wire n_2232;
wire n_1847;
wire n_2458;
wire n_2779;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_2227;
wire n_2301;
wire n_1539;
wire n_2859;
wire n_2847;
wire n_884;
wire n_1851;
wire n_2162;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_2192;
wire n_1676;
wire n_1085;
wire n_1636;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_1977;
wire n_693;
wire n_863;
wire n_2650;
wire n_1254;
wire n_929;
wire n_2433;
wire n_1703;
wire n_899;
wire n_2332;
wire n_2391;
wire n_611;
wire n_1295;
wire n_2060;
wire n_1850;
wire n_2004;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_2571;
wire n_2427;
wire n_2885;
wire n_661;
wire n_2098;
wire n_2616;
wire n_1751;
wire n_2874;
wire n_2867;
wire n_1917;
wire n_2456;
wire n_2769;
wire n_1924;
wire n_1560;
wire n_1654;
wire n_2341;
wire n_2899;
wire n_1548;
wire n_1811;
wire n_2045;
wire n_2575;
wire n_2722;
wire n_1396;
wire n_1230;
wire n_612;
wire n_1840;
wire n_2739;
wire n_1597;
wire n_1771;
wire n_2902;
wire n_1544;
wire n_844;
wire n_1012;
wire n_1267;
wire n_2061;
wire n_2685;
wire n_2094;
wire n_2512;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_2382;
wire n_2043;
wire n_780;
wire n_2349;
wire n_1918;
wire n_2788;
wire n_1443;
wire n_1021;
wire n_2595;
wire n_1465;
wire n_2686;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_2727;
wire n_942;
wire n_1437;
wire n_2077;
wire n_1378;
wire n_1121;
wire n_1416;
wire n_2909;
wire n_1461;
wire n_2717;
wire n_1391;
wire n_1947;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_2527;
wire n_1112;
wire n_1159;
wire n_700;
wire n_772;
wire n_1216;
wire n_2759;
wire n_1245;
wire n_2743;
wire n_1669;
wire n_1675;
wire n_2466;
wire n_676;
wire n_2038;
wire n_2263;
wire n_2800;
wire n_2568;
wire n_2116;
wire n_2271;
wire n_2145;
wire n_2326;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_2806;
wire n_1716;
wire n_1872;
wire n_1585;
wire n_2281;
wire n_1432;
wire n_2245;
wire n_1108;
wire n_1590;
wire n_851;
wire n_1351;
wire n_2216;
wire n_1274;
wire n_2426;
wire n_652;
wire n_1819;
wire n_947;
wire n_2134;
wire n_1260;
wire n_930;
wire n_1179;
wire n_2703;
wire n_696;
wire n_1442;
wire n_2926;
wire n_2620;
wire n_798;
wire n_1833;
wire n_1691;
wire n_916;
wire n_1386;
wire n_2810;
wire n_1884;
wire n_912;
wire n_1555;
wire n_1842;
wire n_2549;
wire n_2499;
wire n_1253;
wire n_1468;
wire n_762;
wire n_1661;
wire n_2791;
wire n_2683;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_2855;
wire n_2166;
wire n_2848;
wire n_1692;
wire n_2611;
wire n_1562;
wire n_2748;
wire n_2185;
wire n_2398;
wire n_1376;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_2015;
wire n_2925;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_2202;
wire n_2072;
wire n_2415;
wire n_2693;
wire n_2877;
wire n_2922;
wire n_2871;
wire n_2930;
wire n_2745;
wire n_2087;
wire n_669;
wire n_1491;
wire n_931;
wire n_2628;
wire n_619;
wire n_967;
wire n_1083;
wire n_2161;
wire n_1418;
wire n_746;
wire n_1357;
wire n_1079;
wire n_1787;
wire n_2462;
wire n_1389;
wire n_2155;
wire n_2659;
wire n_615;
wire n_1139;
wire n_2836;
wire n_2439;
wire n_2864;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_2172;
wire n_2601;
wire n_892;
wire n_1880;
wire n_959;
wire n_2365;
wire n_2257;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_2219;
wire n_1855;
wire n_2100;
wire n_2333;
wire n_1623;
wire n_990;
wire n_1903;
wire n_867;
wire n_2147;
wire n_2435;
wire n_1226;
wire n_2224;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_2825;
wire n_2888;
wire n_1970;
wire n_1920;
wire n_2083;
wire n_815;
wire n_2167;
wire n_2293;
wire n_2753;
wire n_1340;
wire n_2668;
wire n_1240;
wire n_2921;
wire n_1087;
wire n_2701;
wire n_2400;
wire n_632;
wire n_650;
wire n_2388;
wire n_2273;
wire n_2712;
wire n_1433;
wire n_1911;
wire n_2567;
wire n_2557;
wire n_2695;
wire n_2898;
wire n_1908;
wire n_1825;
wire n_1155;
wire n_2598;
wire n_1071;
wire n_2755;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_2795;
wire n_2682;
wire n_1841;
wire n_1680;
wire n_2066;
wire n_2302;
wire n_2762;
wire n_964;
wire n_1627;
wire n_2220;
wire n_2294;
wire n_2274;
wire n_2895;
wire n_2903;
wire n_974;
wire n_1731;
wire n_799;
wire n_1147;
wire n_2829;
wire n_2378;
wire n_2467;
wire n_2768;
wire n_1914;
wire n_965;
wire n_2253;
wire n_934;
wire n_2213;
wire n_1447;
wire n_2363;
wire n_1220;
wire n_2019;
wire n_698;
wire n_2728;
wire n_2130;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_2160;
wire n_1992;
wire n_2924;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_2507;
wire n_2142;
wire n_1633;
wire n_2625;
wire n_2896;
wire n_1913;
wire n_2069;
wire n_2495;
wire n_1058;
wire n_2328;
wire n_2434;
wire n_1042;
wire n_1234;
wire n_2311;
wire n_1578;
wire n_2261;
wire n_1455;
wire n_2287;
wire n_836;
wire n_2223;
wire n_1279;
wire n_2473;
wire n_2144;
wire n_2511;
wire n_1029;
wire n_2649;
wire n_1247;
wire n_760;
wire n_2438;
wire n_1568;
wire n_2919;
wire n_1483;
wire n_1363;
wire n_2681;
wire n_1111;
wire n_1689;
wire n_970;
wire n_2535;
wire n_713;
wire n_1255;
wire n_2632;
wire n_1646;
wire n_598;
wire n_2262;
wire n_2565;
wire n_1237;
wire n_927;
wire n_1095;
wire n_1728;
wire n_2335;
wire n_706;
wire n_2120;
wire n_2631;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_2860;
wire n_2041;
wire n_2113;
wire n_1933;
wire n_1651;
wire n_2697;
wire n_1387;
wire n_1263;
wire n_1817;
wire n_2404;
wire n_2168;
wire n_2757;
wire n_2312;
wire n_670;
wire n_2677;
wire n_1826;
wire n_2834;
wire n_2483;
wire n_1951;
wire n_2490;
wire n_1032;
wire n_1217;
wire n_2558;
wire n_1496;
wire n_637;
wire n_1592;
wire n_2812;
wire n_2662;
wire n_1259;
wire n_2801;
wire n_1177;
wire n_2655;
wire n_1231;
wire n_2132;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_2718;
wire n_720;
wire n_926;
wire n_1943;
wire n_2687;
wire n_2296;
wire n_1802;
wire n_2178;
wire n_2112;
wire n_2765;
wire n_1163;
wire n_2640;
wire n_2811;
wire n_1795;
wire n_1384;
wire n_2237;
wire n_2146;
wire n_1868;
wire n_1501;
wire n_2241;
wire n_2373;
wire n_1173;
wire n_2350;
wire n_1068;
wire n_1198;
wire n_2531;
wire n_1570;
wire n_2099;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_2187;
wire n_1413;
wire n_2617;
wire n_2481;
wire n_2129;
wire n_855;
wire n_2327;
wire n_808;
wire n_1365;
wire n_2476;
wire n_2814;
wire n_2059;
wire n_2437;
wire n_2636;
wire n_1439;
wire n_814;
wire n_2074;
wire n_1665;
wire n_1287;
wire n_2841;
wire n_1611;
wire n_2122;
wire n_2399;
wire n_1414;
wire n_1134;
wire n_2067;
wire n_1484;
wire n_1901;
wire n_647;
wire n_2055;
wire n_2027;
wire n_2932;
wire n_1423;
wire n_2117;
wire n_600;
wire n_1609;
wire n_1053;
wire n_2822;
wire n_1939;
wire n_2308;
wire n_2242;
wire n_1906;
wire n_1899;
wire n_2195;
wire n_2194;
wire n_1467;
wire n_1828;
wire n_2159;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_2267;
wire n_1105;
wire n_677;
wire n_604;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_2102;
wire n_681;
wire n_874;
wire n_2286;
wire n_2023;
wire n_1278;
wire n_707;
wire n_983;
wire n_2783;
wire n_2599;
wire n_699;
wire n_590;
wire n_2075;
wire n_727;
wire n_1726;
wire n_2523;
wire n_1945;
wire n_1015;
wire n_2418;
wire n_1377;
wire n_1162;
wire n_1614;
wire n_2031;
wire n_2496;
wire n_2118;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_2853;
wire n_1098;
wire n_1490;
wire n_2338;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_2225;
wire n_986;
wire n_1104;
wire n_1963;
wire n_2802;
wire n_729;
wire n_887;
wire n_2057;
wire n_2218;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_2593;
wire n_1693;
wire n_2125;
wire n_2716;
wire n_1132;
wire n_1156;
wire n_2741;
wire n_2184;
wire n_2714;
wire n_1823;
wire n_2861;
wire n_2780;
wire n_1120;
wire n_1202;
wire n_627;
wire n_2254;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_2033;
wire n_2618;
wire n_1402;
wire n_957;
wire n_1242;
wire n_2754;
wire n_2707;
wire n_2774;
wire n_2849;
wire n_1607;
wire n_1489;
wire n_2799;
wire n_1218;
wire n_2756;
wire n_2217;
wire n_2226;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_2214;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_2763;
wire n_2256;
wire n_1189;
wire n_1089;
wire n_1859;
wire n_2660;
wire n_1502;
wire n_1523;
wire n_2190;
wire n_1478;
wire n_2732;
wire n_1883;
wire n_2516;
wire n_2776;
wire n_2555;
wire n_1969;
wire n_2708;
wire n_735;
wire n_1005;
wire n_2379;
wire n_1294;
wire n_2661;
wire n_1667;
wire n_845;
wire n_888;
wire n_2894;
wire n_2300;
wire n_1649;
wire n_2452;
wire n_1677;
wire n_2470;
wire n_1927;
wire n_1297;
wire n_2827;
wire n_1708;
wire n_1222;
wire n_2284;
wire n_1844;
wire n_2283;
wire n_2526;
wire n_1957;
wire n_1953;
wire n_2643;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_1919;
wire n_710;
wire n_1791;
wire n_2508;
wire n_2124;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_2594;
wire n_2266;
wire n_2449;
wire n_890;
wire n_842;
wire n_1898;
wire n_1741;
wire n_745;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_1975;
wire n_1373;
wire n_1081;
wire n_742;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_2119;
wire n_2742;
wire n_769;
wire n_1797;
wire n_2366;
wire n_2493;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_832;
wire n_744;
wire n_1895;
wire n_2821;
wire n_2690;
wire n_2474;
wire n_2623;
wire n_982;
wire n_1800;
wire n_915;
wire n_1075;
wire n_2008;
wire n_1331;
wire n_1890;
wire n_2904;
wire n_1529;
wire n_1227;
wire n_2127;
wire n_655;
wire n_1734;
wire n_1860;
wire n_2785;
wire n_2460;
wire n_2840;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_2448;
wire n_2211;
wire n_2292;
wire n_2480;
wire n_606;
wire n_951;
wire n_2772;
wire n_1700;
wire n_862;
wire n_2637;
wire n_659;
wire n_1332;
wire n_2306;
wire n_1854;
wire n_666;
wire n_1747;
wire n_2071;
wire n_2424;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_2414;
wire n_2082;
wire n_2893;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_2389;
wire n_1309;
wire n_999;
wire n_2280;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_2737;
wire n_1867;
wire n_852;
wire n_1394;
wire n_2916;
wire n_2576;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_2696;
wire n_2140;
wire n_1748;
wire n_1301;
wire n_873;
wire n_2157;
wire n_1966;
wire n_1243;
wire n_2171;
wire n_2468;
wire n_1400;
wire n_2035;
wire n_2614;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_2581;
wire n_1783;
wire n_608;
wire n_2494;
wire n_1538;
wire n_2831;
wire n_2457;
wire n_2128;
wire n_1037;
wire n_1329;
wire n_1993;
wire n_1545;
wire n_2629;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_2540;
wire n_1605;
wire n_1078;
wire n_2486;
wire n_1897;
wire n_2520;
wire n_2137;
wire n_1161;
wire n_2489;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_1191;
wire n_618;
wire n_2492;
wire n_736;
wire n_1025;
wire n_1215;
wire n_1449;
wire n_2337;
wire n_2265;
wire n_687;
wire n_2900;
wire n_797;
wire n_2026;
wire n_2912;
wire n_1786;
wire n_2627;
wire n_1327;
wire n_1475;
wire n_642;
wire n_2106;
wire n_1804;
wire n_1406;
wire n_595;
wire n_1405;
wire n_2684;
wire n_2726;
wire n_602;
wire n_2622;
wire n_2272;
wire n_1757;
wire n_592;
wire n_1499;
wire n_1318;
wire n_854;
wire n_2091;
wire n_1632;
wire n_1769;
wire n_1929;
wire n_1950;
wire n_2264;
wire n_2691;
wire n_805;
wire n_2032;
wire n_2090;
wire n_2929;
wire n_1658;
wire n_2249;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_1596;
wire n_2348;
wire n_2656;
wire n_1281;
wire n_2364;
wire n_1997;
wire n_2574;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_1733;
wire n_1476;
wire n_1524;
wire n_1856;
wire n_2016;
wire n_2667;
wire n_2725;
wire n_2928;
wire n_1118;
wire n_943;
wire n_678;
wire n_2905;
wire n_2884;
wire n_651;
wire n_2850;
wire n_1874;
wire n_1293;
wire n_961;
wire n_1046;
wire n_1807;
wire n_1123;
wire n_726;
wire n_1657;
wire n_878;
wire n_2857;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_2307;
wire n_1488;
wire n_985;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_2295;
wire n_2730;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_2412;
wire n_2720;
wire n_1352;
wire n_2405;
wire n_2815;
wire n_1824;
wire n_643;
wire n_2606;
wire n_2700;
wire n_1492;
wire n_2383;
wire n_2764;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_2633;
wire n_2416;
wire n_819;
wire n_2386;
wire n_2907;
wire n_1971;
wire n_1324;
wire n_1429;
wire n_2064;
wire n_2353;
wire n_2528;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_2325;
wire n_1130;
wire n_1450;
wire n_756;
wire n_2022;
wire n_1016;
wire n_2298;
wire n_1149;
wire n_1505;
wire n_2408;
wire n_2698;
wire n_2320;
wire n_979;
wire n_2329;
wire n_2570;
wire n_1642;
wire n_2417;
wire n_2789;
wire n_2525;
wire n_1815;
wire n_2813;
wire n_897;
wire n_2546;
wire n_949;
wire n_2454;
wire n_1493;
wire n_2890;
wire n_2911;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_2354;
wire n_1864;
wire n_2760;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_2368;
wire n_802;
wire n_1151;
wire n_960;
wire n_2352;
wire n_2502;
wire n_1256;
wire n_714;
wire n_2170;
wire n_790;
wire n_2244;
wire n_2143;
wire n_2393;
wire n_725;
wire n_2377;
wire n_1577;
wire n_1448;
wire n_2198;
wire n_1009;
wire n_2652;
wire n_1133;
wire n_883;
wire n_1852;
wire n_801;
wire n_1286;
wire n_2612;
wire n_818;
wire n_1685;
wire n_779;
wire n_2410;
wire n_2314;
wire n_2477;
wire n_2279;
wire n_594;
wire n_2222;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_2076;
wire n_2133;
wire n_2203;
wire n_833;
wire n_1426;
wire n_2250;
wire n_2497;
wire n_2247;
wire n_2230;
wire n_879;
wire n_1117;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_2001;
wire n_1047;
wire n_2506;
wire n_1472;
wire n_2413;
wire n_1593;
wire n_2610;
wire n_1050;
wire n_2626;
wire n_2158;
wire n_2578;
wire n_2607;
wire n_2285;
wire n_2892;
wire n_1201;
wire n_1288;
wire n_2605;
wire n_858;
wire n_2804;
wire n_1185;
wire n_2475;
wire n_2796;
wire n_2173;
wire n_2715;
wire n_1035;
wire n_1143;
wire n_2665;
wire n_2070;
wire n_2136;
wire n_2771;
wire n_1090;
wire n_2403;
wire n_1367;
wire n_2044;
wire n_928;
wire n_1153;
wire n_1103;
wire n_825;
wire n_732;
wire n_2619;
wire n_1565;
wire n_1192;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_2854;
wire n_1291;
wire n_2020;
wire n_748;
wire n_2310;
wire n_1045;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_2711;
wire n_1881;
wire n_2635;
wire n_988;
wire n_914;
wire n_689;
wire n_1116;
wire n_1958;
wire n_2747;
wire n_1511;
wire n_2177;
wire n_2713;
wire n_1422;
wire n_2766;
wire n_1965;
wire n_644;
wire n_1197;
wire n_2820;
wire n_2613;
wire n_1165;
wire n_2934;
wire n_1641;
wire n_2845;
wire n_1517;
wire n_2036;
wire n_843;
wire n_2647;
wire n_638;
wire n_2003;
wire n_2533;
wire n_2210;
wire n_1307;
wire n_1128;
wire n_2053;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_2343;
wire n_775;
wire n_667;
wire n_2419;
wire n_1049;
wire n_2330;
wire n_2826;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_2777;
wire n_2450;
wire n_2411;
wire n_1356;
wire n_1341;
wire n_2234;
wire n_2309;
wire n_1504;
wire n_1955;
wire n_2110;
wire n_2431;
wire n_1773;
wire n_1440;
wire n_2666;
wire n_1370;
wire n_1603;
wire n_728;
wire n_2401;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_2588;
wire n_2863;
wire n_2331;
wire n_935;
wire n_2886;
wire n_2478;
wire n_685;
wire n_911;
wire n_2658;
wire n_623;
wire n_2608;
wire n_2920;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_1534;
wire n_1948;
wire n_2767;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_2396;
wire n_1362;
wire n_1559;
wire n_2121;
wire n_2692;
wire n_601;
wire n_683;
wire n_628;
wire n_1300;
wire n_1960;
wire n_2068;
wire n_743;
wire n_1194;
wire n_2862;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_2553;
wire n_2645;
wire n_907;
wire n_2749;
wire n_1454;
wire n_2592;
wire n_660;
wire n_2459;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_2566;
wire n_2751;
wire n_1968;
wire n_918;
wire n_1885;
wire n_639;
wire n_673;
wire n_2842;
wire n_2833;
wire n_2196;
wire n_1038;
wire n_2371;
wire n_1978;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_593;
wire n_1695;
wire n_2560;
wire n_1164;
wire n_2313;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_2609;
wire n_2561;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_1653;
wire n_872;
wire n_2882;
wire n_2303;
wire n_2669;
wire n_1157;
wire n_1584;
wire n_848;
wire n_1664;
wire n_629;
wire n_1739;
wire n_2642;
wire n_1814;
wire n_2154;
wire n_2441;
wire n_2236;
wire n_1789;
wire n_763;
wire n_1986;
wire n_2174;
wire n_2688;
wire n_692;
wire n_2624;
wire n_2054;
wire n_1857;
wire n_2315;
wire n_984;
wire n_1687;
wire n_2073;
wire n_2150;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_2498;
wire n_800;
wire n_2638;
wire n_2046;
wire n_1910;
wire n_1816;
wire n_2803;
wire n_1756;
wire n_2887;
wire n_1606;
wire n_2189;
wire n_621;
wire n_2648;
wire n_1587;
wire n_2093;
wire n_2340;
wire n_2018;
wire n_2672;
wire n_1772;
wire n_2444;
wire n_2602;
wire n_1014;
wire n_724;
wire n_2204;
wire n_2931;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_1311;
wire n_2199;
wire n_2881;
wire n_1956;
wire n_1589;
wire n_2151;
wire n_1100;
wire n_875;
wire n_1617;
wire n_2455;
wire n_827;
wire n_2600;
wire n_2231;
wire n_697;
wire n_2828;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_2305;
wire n_880;
wire n_793;
wire n_2114;
wire n_2927;
wire n_1175;
wire n_2289;
wire n_2530;
wire n_2299;
wire n_751;
wire n_1027;
wire n_1070;
wire n_2406;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_2883;
wire n_1221;
wire n_1785;
wire n_1262;
wire n_792;
wire n_1942;
wire n_2180;
wire n_1579;
wire n_2809;
wire n_2181;
wire n_2014;
wire n_975;
wire n_1645;
wire n_923;
wire n_1381;
wire n_1124;
wire n_2870;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_2889;
wire n_2276;
wire n_1805;
wire n_2282;
wire n_981;
wire n_2910;
wire n_2141;
wire n_1110;
wire n_1758;
wire n_2503;
wire n_2270;
wire n_2443;
wire n_1407;
wire n_2465;
wire n_1204;
wire n_2865;
wire n_1554;
wire n_994;
wire n_2428;
wire n_2586;
wire n_1360;
wire n_973;
wire n_2858;
wire n_972;
wire n_2251;
wire n_2923;
wire n_2843;
wire n_856;
wire n_2572;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_1679;
wire n_2872;
wire n_2126;
wire n_1952;
wire n_2425;
wire n_2394;
wire n_1858;
wire n_1678;
wire n_2589;
wire n_1482;
wire n_1361;
wire n_2356;
wire n_1601;
wire n_1057;
wire n_2487;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_2534;
wire n_2488;
wire n_1509;
wire n_828;
wire n_1411;
wire n_1359;
wire n_1721;
wire n_2564;
wire n_2591;
wire n_653;
wire n_1445;
wire n_1317;
wire n_2050;
wire n_2197;
wire n_783;
wire n_2550;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_2385;
wire n_2387;
wire n_1008;
wire n_1024;
wire n_830;
wire n_2291;
wire n_2816;
wire n_1980;
wire n_2518;
wire n_987;
wire n_936;
wire n_2510;
wire n_1620;
wire n_2501;
wire n_2542;
wire n_1385;
wire n_1525;
wire n_2793;
wire n_1998;
wire n_2165;
wire n_2675;
wire n_2604;
wire n_1775;
wire n_788;
wire n_908;
wire n_2639;
wire n_1036;
wire n_2169;
wire n_2603;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_2630;
wire n_591;
wire n_2794;
wire n_969;
wire n_2028;
wire n_919;
wire n_1663;
wire n_2901;
wire n_2092;
wire n_2175;
wire n_1625;
wire n_2086;
wire n_2773;
wire n_2817;
wire n_1926;
wire n_2402;
wire n_1458;
wire n_1630;
wire n_679;
wire n_663;
wire n_1720;
wire n_2409;
wire n_2176;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_1358;
wire n_1200;
wire n_826;
wire n_2808;
wire n_2453;
wire n_2344;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_940;
wire n_2392;
wire n_1537;
wire n_2138;
wire n_2065;
wire n_2543;
wire n_2321;
wire n_1077;
wire n_2597;
wire n_607;
wire n_956;
wire n_1930;
wire n_765;
wire n_1809;
wire n_2787;
wire n_1904;
wire n_1843;
wire n_2000;
wire n_2805;
wire n_1268;
wire n_2676;
wire n_2758;
wire n_2395;
wire n_917;
wire n_2868;
wire n_2723;
wire n_1271;
wire n_2096;
wire n_2440;
wire n_2556;
wire n_2186;
wire n_1530;
wire n_2215;
wire n_2770;
wire n_631;
wire n_1170;
wire n_2724;
wire n_2258;
wire n_1261;
wire n_2471;
wire n_702;
wire n_898;
wire n_857;
wire n_1067;
wire n_968;
wire n_1235;
wire n_1323;
wire n_2584;
wire n_2375;
wire n_1462;
wire n_1937;
wire n_2012;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_733;
wire n_761;
wire n_2212;
wire n_731;
wire n_1813;
wire n_2268;
wire n_1452;
wire n_2835;
wire n_1573;
wire n_2734;
wire n_668;
wire n_2569;
wire n_758;
wire n_2252;
wire n_2111;
wire n_2420;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_784;
wire n_648;
wire n_816;
wire n_2897;
wire n_1322;
wire n_2583;
wire n_2918;
wire n_1473;
wire n_835;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_2651;
wire n_753;
wire n_2445;
wire n_2733;
wire n_1770;
wire n_701;
wire n_1003;
wire n_2469;
wire n_1125;
wire n_2103;
wire n_2358;
wire n_1710;
wire n_1865;
wire n_2522;
wire n_2641;
wire n_2463;
wire n_1344;
wire n_2355;
wire n_1390;
wire n_2580;
wire n_2699;
wire n_1792;
wire n_2062;
wire n_1141;
wire n_1629;
wire n_1640;
wire n_822;
wire n_1094;
wire n_1459;
wire n_840;
wire n_2153;
wire n_2324;
wire n_1510;
wire n_2710;
wire n_2505;
wire n_2139;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_2397;
wire n_2521;
wire n_1727;
wire n_2740;
wire n_2235;
wire n_1991;
wire n_1575;
wire n_2721;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_2615;
wire n_614;
wire n_2775;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_2351;
wire n_2260;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_2206;
wire n_2784;
wire n_2541;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_2347;
wire n_1152;
wire n_2657;
wire n_2538;
wire n_2034;
wire n_1845;
wire n_2447;
wire n_1934;
wire n_2101;
wire n_2577;
wire n_921;
wire n_2362;
wire n_1615;
wire n_1236;
wire n_2104;
wire n_1265;
wire n_1576;
wire n_2105;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_2372;
wire n_2552;
wire n_1409;
wire n_1588;
wire n_1148;
wire n_1684;
wire n_1673;
wire n_2422;
wire n_2704;
wire n_1334;
wire n_654;
wire n_2290;
wire n_2933;
wire n_2856;
wire n_2088;
wire n_1275;
wire n_904;
wire n_2005;
wire n_2048;
wire n_1696;
wire n_1875;
wire n_1059;
wire n_684;
wire n_2429;
wire n_2108;
wire n_2736;
wire n_1039;
wire n_2246;
wire n_1150;
wire n_977;
wire n_2339;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_2532;
wire n_2191;
wire n_1497;
wire n_1866;
wire n_2472;
wire n_2664;
wire n_2705;
wire n_2056;
wire n_2852;
wire n_1136;
wire n_2515;
wire n_1782;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_838;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_2519;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_2360;
wire n_1393;
wire n_723;
wire n_2240;
wire n_658;
wire n_630;
wire n_1369;
wire n_2846;
wire n_1781;
wire n_709;
wire n_2917;
wire n_2544;
wire n_809;
wire n_2085;
wire n_2432;
wire n_1686;
wire n_1964;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_2188;
wire n_1982;
wire n_2097;
wire n_662;
wire n_641;
wire n_2430;
wire n_2504;
wire n_910;
wire n_741;
wire n_1410;
wire n_939;
wire n_2297;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_1223;
wire n_2545;
wire n_1768;
wire n_2513;
wire n_2193;
wire n_2369;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_2451;
wire n_2115;
wire n_2913;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_922;
wire n_1004;
wire n_1810;
wire n_2587;
wire n_1347;
wire n_2839;
wire n_860;
wire n_1043;
wire n_2869;
wire n_1923;
wire n_2670;
wire n_1764;
wire n_2674;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_2644;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_2148;
wire n_1946;
wire n_774;
wire n_933;
wire n_1779;
wire n_2562;
wire n_596;
wire n_954;
wire n_2051;
wire n_1168;
wire n_1821;
wire n_1310;
wire n_656;
wire n_2673;
wire n_664;
wire n_1591;
wire n_2585;
wire n_1229;
wire n_1683;
wire n_2582;
wire n_2548;
wire n_1896;
wire n_2164;
wire n_1732;
wire n_2381;
wire n_2744;
wire n_1967;
wire n_2384;
wire n_2678;
wire n_2179;
wire n_1280;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_2052;
wire n_2485;
wire n_1063;
wire n_2205;
wire n_2275;
wire n_991;
wire n_2183;
wire n_2563;
wire n_1724;
wire n_1670;
wire n_1799;
wire n_1707;
wire n_2080;
wire n_2058;
wire n_1126;
wire n_2761;
wire n_2357;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_2875;
wire n_1639;
wire n_2209;
wire n_2421;
wire n_1302;
wire n_1000;
wire n_626;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_2047;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_2792;
wire n_1634;
wire n_2596;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_2269;
wire n_1474;
wire n_2081;
wire n_937;
wire n_2536;
wire n_2524;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_1702;
wire n_1794;
wire n_1375;
wire n_1232;
wire n_1211;
wire n_1368;
wire n_996;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_2891;
wire n_2318;
wire n_1827;
wire n_866;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1722;
wire n_1001;
wire n_2361;
wire n_1115;
wire n_2229;
wire n_2819;
wire n_2880;
wire n_1339;
wire n_1644;
wire n_1002;
wire n_1051;
wire n_2551;
wire n_1102;
wire n_719;
wire n_2255;
wire n_1252;
wire n_1129;
wire n_2239;
wire n_1464;
wire n_1296;
wire n_773;
wire n_2798;
wire n_2316;
wire n_2464;
wire n_1010;
wire n_2830;
wire n_882;
wire n_2706;
wire n_2304;
wire n_1249;
wire n_1871;
wire n_803;
wire n_2514;
wire n_718;
wire n_1434;
wire n_1905;
wire n_1569;
wire n_2573;
wire n_2336;
wire n_1662;
wire n_1299;
wire n_1870;
wire n_2063;
wire n_1925;
wire n_782;
wire n_2915;
wire n_2654;
wire n_2491;
wire n_1861;
wire n_2079;
wire n_1228;
wire n_2319;
wire n_2152;
wire n_2517;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_2259;
wire n_849;
wire n_2095;
wire n_2719;
wire n_2738;
wire n_1820;
wire n_2590;
wire n_2876;
wire n_2797;
wire n_1251;
wire n_1989;
wire n_1421;
wire n_2208;
wire n_2423;
wire n_2689;
wire n_2778;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_2228;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_2479;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2824;
wire n_2037;
wire n_1308;
wire n_796;
wire n_2851;
wire n_2823;
wire n_2345;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_2089;
wire n_1487;
wire n_675;

INVx1_ASAP7_75t_L g590 ( 
.A(n_102),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_556),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_496),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_527),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_255),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_290),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_33),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_429),
.Y(n_597)
);

INVx1_ASAP7_75t_SL g598 ( 
.A(n_279),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_131),
.Y(n_599)
);

BUFx10_ASAP7_75t_L g600 ( 
.A(n_262),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_3),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_373),
.Y(n_602)
);

CKINVDCx20_ASAP7_75t_R g603 ( 
.A(n_263),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_493),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_243),
.Y(n_605)
);

CKINVDCx20_ASAP7_75t_R g606 ( 
.A(n_484),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_63),
.Y(n_607)
);

INVx2_ASAP7_75t_SL g608 ( 
.A(n_542),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_580),
.Y(n_609)
);

CKINVDCx16_ASAP7_75t_R g610 ( 
.A(n_286),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_449),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_248),
.Y(n_612)
);

HB1xp67_ASAP7_75t_L g613 ( 
.A(n_118),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_213),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_93),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_225),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_177),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_150),
.Y(n_618)
);

INVx2_ASAP7_75t_SL g619 ( 
.A(n_185),
.Y(n_619)
);

INVx1_ASAP7_75t_SL g620 ( 
.A(n_98),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_451),
.Y(n_621)
);

CKINVDCx20_ASAP7_75t_R g622 ( 
.A(n_139),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_285),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_7),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_420),
.Y(n_625)
);

BUFx10_ASAP7_75t_L g626 ( 
.A(n_407),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_449),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_1),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_116),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_575),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_203),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_346),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_37),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_398),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_176),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_81),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_161),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_557),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_339),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_573),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_563),
.Y(n_641)
);

HB1xp67_ASAP7_75t_L g642 ( 
.A(n_494),
.Y(n_642)
);

BUFx3_ASAP7_75t_L g643 ( 
.A(n_396),
.Y(n_643)
);

BUFx3_ASAP7_75t_L g644 ( 
.A(n_92),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_555),
.Y(n_645)
);

CKINVDCx5p33_ASAP7_75t_R g646 ( 
.A(n_89),
.Y(n_646)
);

INVxp67_ASAP7_75t_L g647 ( 
.A(n_76),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_32),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_231),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_349),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_413),
.Y(n_651)
);

CKINVDCx20_ASAP7_75t_R g652 ( 
.A(n_175),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_528),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_60),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_124),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_413),
.Y(n_656)
);

BUFx5_ASAP7_75t_L g657 ( 
.A(n_434),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_98),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_380),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_525),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_297),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_315),
.Y(n_662)
);

INVx1_ASAP7_75t_SL g663 ( 
.A(n_400),
.Y(n_663)
);

CKINVDCx20_ASAP7_75t_R g664 ( 
.A(n_583),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_360),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_43),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_560),
.Y(n_667)
);

INVx1_ASAP7_75t_SL g668 ( 
.A(n_273),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_215),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_351),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_88),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_484),
.Y(n_672)
);

CKINVDCx16_ASAP7_75t_R g673 ( 
.A(n_533),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_534),
.Y(n_674)
);

CKINVDCx20_ASAP7_75t_R g675 ( 
.A(n_473),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_284),
.Y(n_676)
);

CKINVDCx20_ASAP7_75t_R g677 ( 
.A(n_20),
.Y(n_677)
);

BUFx10_ASAP7_75t_L g678 ( 
.A(n_397),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_202),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_407),
.Y(n_680)
);

CKINVDCx16_ASAP7_75t_R g681 ( 
.A(n_549),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_115),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_539),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_295),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_544),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_128),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_25),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_52),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_587),
.Y(n_689)
);

CKINVDCx20_ASAP7_75t_R g690 ( 
.A(n_448),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_396),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_356),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_516),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_180),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_141),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_544),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_140),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_64),
.Y(n_698)
);

INVx2_ASAP7_75t_SL g699 ( 
.A(n_165),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_270),
.Y(n_700)
);

BUFx3_ASAP7_75t_L g701 ( 
.A(n_360),
.Y(n_701)
);

BUFx6f_ASAP7_75t_L g702 ( 
.A(n_356),
.Y(n_702)
);

INVx1_ASAP7_75t_SL g703 ( 
.A(n_40),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_430),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_186),
.Y(n_705)
);

INVx1_ASAP7_75t_SL g706 ( 
.A(n_94),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_208),
.Y(n_707)
);

INVx1_ASAP7_75t_SL g708 ( 
.A(n_345),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_561),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_180),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_7),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_461),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_461),
.Y(n_713)
);

INVx2_ASAP7_75t_SL g714 ( 
.A(n_93),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_254),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_113),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_511),
.Y(n_717)
);

CKINVDCx5p33_ASAP7_75t_R g718 ( 
.A(n_324),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_412),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_305),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_405),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_100),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_274),
.Y(n_723)
);

CKINVDCx20_ASAP7_75t_R g724 ( 
.A(n_565),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_51),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_552),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_173),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_284),
.Y(n_728)
);

BUFx10_ASAP7_75t_L g729 ( 
.A(n_509),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_394),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_65),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_429),
.Y(n_732)
);

BUFx3_ASAP7_75t_L g733 ( 
.A(n_540),
.Y(n_733)
);

BUFx5_ASAP7_75t_L g734 ( 
.A(n_572),
.Y(n_734)
);

CKINVDCx5p33_ASAP7_75t_R g735 ( 
.A(n_279),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_234),
.Y(n_736)
);

CKINVDCx20_ASAP7_75t_R g737 ( 
.A(n_378),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_522),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_134),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_40),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_90),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_432),
.Y(n_742)
);

INVx1_ASAP7_75t_SL g743 ( 
.A(n_64),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_526),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_249),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_306),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_246),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_450),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_440),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_398),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_167),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_11),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_376),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_147),
.Y(n_754)
);

CKINVDCx5p33_ASAP7_75t_R g755 ( 
.A(n_472),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_300),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_478),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_148),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_532),
.Y(n_759)
);

BUFx2_ASAP7_75t_L g760 ( 
.A(n_18),
.Y(n_760)
);

CKINVDCx16_ASAP7_75t_R g761 ( 
.A(n_335),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_388),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_233),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_547),
.Y(n_764)
);

INVx2_ASAP7_75t_L g765 ( 
.A(n_291),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_310),
.Y(n_766)
);

CKINVDCx20_ASAP7_75t_R g767 ( 
.A(n_307),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_177),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_26),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_480),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_182),
.Y(n_771)
);

BUFx2_ASAP7_75t_L g772 ( 
.A(n_497),
.Y(n_772)
);

CKINVDCx5p33_ASAP7_75t_R g773 ( 
.A(n_446),
.Y(n_773)
);

CKINVDCx5p33_ASAP7_75t_R g774 ( 
.A(n_543),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_47),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_503),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_564),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_554),
.Y(n_778)
);

BUFx3_ASAP7_75t_L g779 ( 
.A(n_20),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_370),
.Y(n_780)
);

BUFx2_ASAP7_75t_L g781 ( 
.A(n_430),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_371),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_303),
.Y(n_783)
);

CKINVDCx20_ASAP7_75t_R g784 ( 
.A(n_218),
.Y(n_784)
);

CKINVDCx5p33_ASAP7_75t_R g785 ( 
.A(n_384),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_204),
.Y(n_786)
);

CKINVDCx14_ASAP7_75t_R g787 ( 
.A(n_411),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_173),
.Y(n_788)
);

BUFx2_ASAP7_75t_L g789 ( 
.A(n_115),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_86),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_91),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_529),
.Y(n_792)
);

CKINVDCx5p33_ASAP7_75t_R g793 ( 
.A(n_280),
.Y(n_793)
);

INVx1_ASAP7_75t_SL g794 ( 
.A(n_277),
.Y(n_794)
);

CKINVDCx14_ASAP7_75t_R g795 ( 
.A(n_17),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_125),
.Y(n_796)
);

INVx1_ASAP7_75t_SL g797 ( 
.A(n_54),
.Y(n_797)
);

INVx2_ASAP7_75t_SL g798 ( 
.A(n_425),
.Y(n_798)
);

BUFx3_ASAP7_75t_L g799 ( 
.A(n_162),
.Y(n_799)
);

INVx3_ASAP7_75t_L g800 ( 
.A(n_567),
.Y(n_800)
);

CKINVDCx20_ASAP7_75t_R g801 ( 
.A(n_110),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_343),
.Y(n_802)
);

CKINVDCx5p33_ASAP7_75t_R g803 ( 
.A(n_353),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_26),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_432),
.Y(n_805)
);

BUFx6f_ASAP7_75t_L g806 ( 
.A(n_239),
.Y(n_806)
);

CKINVDCx20_ASAP7_75t_R g807 ( 
.A(n_258),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_251),
.Y(n_808)
);

CKINVDCx5p33_ASAP7_75t_R g809 ( 
.A(n_559),
.Y(n_809)
);

CKINVDCx5p33_ASAP7_75t_R g810 ( 
.A(n_72),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_447),
.Y(n_811)
);

CKINVDCx5p33_ASAP7_75t_R g812 ( 
.A(n_528),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_469),
.Y(n_813)
);

BUFx3_ASAP7_75t_L g814 ( 
.A(n_225),
.Y(n_814)
);

CKINVDCx5p33_ASAP7_75t_R g815 ( 
.A(n_34),
.Y(n_815)
);

INVx1_ASAP7_75t_SL g816 ( 
.A(n_282),
.Y(n_816)
);

CKINVDCx5p33_ASAP7_75t_R g817 ( 
.A(n_198),
.Y(n_817)
);

CKINVDCx5p33_ASAP7_75t_R g818 ( 
.A(n_378),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_459),
.Y(n_819)
);

INVx2_ASAP7_75t_SL g820 ( 
.A(n_495),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_91),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_585),
.Y(n_822)
);

CKINVDCx5p33_ASAP7_75t_R g823 ( 
.A(n_289),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_531),
.Y(n_824)
);

CKINVDCx5p33_ASAP7_75t_R g825 ( 
.A(n_285),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_331),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_176),
.Y(n_827)
);

CKINVDCx20_ASAP7_75t_R g828 ( 
.A(n_244),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_389),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_462),
.Y(n_830)
);

CKINVDCx5p33_ASAP7_75t_R g831 ( 
.A(n_441),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_6),
.Y(n_832)
);

CKINVDCx5p33_ASAP7_75t_R g833 ( 
.A(n_148),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_538),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_230),
.Y(n_835)
);

CKINVDCx5p33_ASAP7_75t_R g836 ( 
.A(n_527),
.Y(n_836)
);

CKINVDCx5p33_ASAP7_75t_R g837 ( 
.A(n_58),
.Y(n_837)
);

CKINVDCx5p33_ASAP7_75t_R g838 ( 
.A(n_324),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_16),
.Y(n_839)
);

BUFx10_ASAP7_75t_L g840 ( 
.A(n_531),
.Y(n_840)
);

CKINVDCx5p33_ASAP7_75t_R g841 ( 
.A(n_537),
.Y(n_841)
);

CKINVDCx5p33_ASAP7_75t_R g842 ( 
.A(n_410),
.Y(n_842)
);

CKINVDCx5p33_ASAP7_75t_R g843 ( 
.A(n_242),
.Y(n_843)
);

CKINVDCx5p33_ASAP7_75t_R g844 ( 
.A(n_349),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_259),
.Y(n_845)
);

CKINVDCx5p33_ASAP7_75t_R g846 ( 
.A(n_576),
.Y(n_846)
);

BUFx2_ASAP7_75t_L g847 ( 
.A(n_128),
.Y(n_847)
);

CKINVDCx5p33_ASAP7_75t_R g848 ( 
.A(n_106),
.Y(n_848)
);

CKINVDCx5p33_ASAP7_75t_R g849 ( 
.A(n_381),
.Y(n_849)
);

CKINVDCx5p33_ASAP7_75t_R g850 ( 
.A(n_127),
.Y(n_850)
);

CKINVDCx5p33_ASAP7_75t_R g851 ( 
.A(n_301),
.Y(n_851)
);

CKINVDCx5p33_ASAP7_75t_R g852 ( 
.A(n_466),
.Y(n_852)
);

CKINVDCx5p33_ASAP7_75t_R g853 ( 
.A(n_397),
.Y(n_853)
);

CKINVDCx5p33_ASAP7_75t_R g854 ( 
.A(n_582),
.Y(n_854)
);

CKINVDCx5p33_ASAP7_75t_R g855 ( 
.A(n_427),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_568),
.Y(n_856)
);

CKINVDCx5p33_ASAP7_75t_R g857 ( 
.A(n_145),
.Y(n_857)
);

BUFx6f_ASAP7_75t_L g858 ( 
.A(n_8),
.Y(n_858)
);

CKINVDCx5p33_ASAP7_75t_R g859 ( 
.A(n_491),
.Y(n_859)
);

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_24),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_532),
.Y(n_861)
);

CKINVDCx5p33_ASAP7_75t_R g862 ( 
.A(n_421),
.Y(n_862)
);

CKINVDCx5p33_ASAP7_75t_R g863 ( 
.A(n_305),
.Y(n_863)
);

BUFx3_ASAP7_75t_L g864 ( 
.A(n_286),
.Y(n_864)
);

BUFx6f_ASAP7_75t_L g865 ( 
.A(n_66),
.Y(n_865)
);

BUFx6f_ASAP7_75t_L g866 ( 
.A(n_139),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_221),
.Y(n_867)
);

BUFx10_ASAP7_75t_L g868 ( 
.A(n_332),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_363),
.Y(n_869)
);

CKINVDCx5p33_ASAP7_75t_R g870 ( 
.A(n_146),
.Y(n_870)
);

CKINVDCx20_ASAP7_75t_R g871 ( 
.A(n_418),
.Y(n_871)
);

CKINVDCx5p33_ASAP7_75t_R g872 ( 
.A(n_10),
.Y(n_872)
);

CKINVDCx5p33_ASAP7_75t_R g873 ( 
.A(n_256),
.Y(n_873)
);

CKINVDCx5p33_ASAP7_75t_R g874 ( 
.A(n_546),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_223),
.Y(n_875)
);

CKINVDCx5p33_ASAP7_75t_R g876 ( 
.A(n_551),
.Y(n_876)
);

CKINVDCx5p33_ASAP7_75t_R g877 ( 
.A(n_391),
.Y(n_877)
);

CKINVDCx5p33_ASAP7_75t_R g878 ( 
.A(n_445),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_118),
.Y(n_879)
);

CKINVDCx5p33_ASAP7_75t_R g880 ( 
.A(n_537),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_439),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_490),
.Y(n_882)
);

INVx1_ASAP7_75t_SL g883 ( 
.A(n_168),
.Y(n_883)
);

CKINVDCx20_ASAP7_75t_R g884 ( 
.A(n_224),
.Y(n_884)
);

BUFx5_ASAP7_75t_L g885 ( 
.A(n_482),
.Y(n_885)
);

CKINVDCx5p33_ASAP7_75t_R g886 ( 
.A(n_70),
.Y(n_886)
);

CKINVDCx5p33_ASAP7_75t_R g887 ( 
.A(n_485),
.Y(n_887)
);

CKINVDCx5p33_ASAP7_75t_R g888 ( 
.A(n_335),
.Y(n_888)
);

CKINVDCx5p33_ASAP7_75t_R g889 ( 
.A(n_581),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_278),
.Y(n_890)
);

CKINVDCx5p33_ASAP7_75t_R g891 ( 
.A(n_558),
.Y(n_891)
);

CKINVDCx20_ASAP7_75t_R g892 ( 
.A(n_5),
.Y(n_892)
);

CKINVDCx5p33_ASAP7_75t_R g893 ( 
.A(n_492),
.Y(n_893)
);

CKINVDCx5p33_ASAP7_75t_R g894 ( 
.A(n_35),
.Y(n_894)
);

CKINVDCx16_ASAP7_75t_R g895 ( 
.A(n_464),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_347),
.Y(n_896)
);

BUFx3_ASAP7_75t_L g897 ( 
.A(n_43),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_282),
.Y(n_898)
);

CKINVDCx5p33_ASAP7_75t_R g899 ( 
.A(n_492),
.Y(n_899)
);

CKINVDCx5p33_ASAP7_75t_R g900 ( 
.A(n_456),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_301),
.Y(n_901)
);

CKINVDCx5p33_ASAP7_75t_R g902 ( 
.A(n_316),
.Y(n_902)
);

CKINVDCx5p33_ASAP7_75t_R g903 ( 
.A(n_422),
.Y(n_903)
);

CKINVDCx5p33_ASAP7_75t_R g904 ( 
.A(n_553),
.Y(n_904)
);

CKINVDCx5p33_ASAP7_75t_R g905 ( 
.A(n_264),
.Y(n_905)
);

CKINVDCx20_ASAP7_75t_R g906 ( 
.A(n_210),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_283),
.Y(n_907)
);

CKINVDCx5p33_ASAP7_75t_R g908 ( 
.A(n_337),
.Y(n_908)
);

CKINVDCx5p33_ASAP7_75t_R g909 ( 
.A(n_386),
.Y(n_909)
);

CKINVDCx5p33_ASAP7_75t_R g910 ( 
.A(n_226),
.Y(n_910)
);

CKINVDCx5p33_ASAP7_75t_R g911 ( 
.A(n_21),
.Y(n_911)
);

CKINVDCx5p33_ASAP7_75t_R g912 ( 
.A(n_274),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_376),
.Y(n_913)
);

INVx2_ASAP7_75t_L g914 ( 
.A(n_491),
.Y(n_914)
);

CKINVDCx5p33_ASAP7_75t_R g915 ( 
.A(n_56),
.Y(n_915)
);

CKINVDCx20_ASAP7_75t_R g916 ( 
.A(n_411),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_21),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_441),
.Y(n_918)
);

CKINVDCx20_ASAP7_75t_R g919 ( 
.A(n_263),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_271),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_12),
.Y(n_921)
);

CKINVDCx5p33_ASAP7_75t_R g922 ( 
.A(n_498),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_550),
.Y(n_923)
);

CKINVDCx20_ASAP7_75t_R g924 ( 
.A(n_339),
.Y(n_924)
);

CKINVDCx5p33_ASAP7_75t_R g925 ( 
.A(n_50),
.Y(n_925)
);

INVx3_ASAP7_75t_L g926 ( 
.A(n_230),
.Y(n_926)
);

CKINVDCx5p33_ASAP7_75t_R g927 ( 
.A(n_566),
.Y(n_927)
);

CKINVDCx5p33_ASAP7_75t_R g928 ( 
.A(n_111),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_522),
.Y(n_929)
);

CKINVDCx5p33_ASAP7_75t_R g930 ( 
.A(n_250),
.Y(n_930)
);

CKINVDCx5p33_ASAP7_75t_R g931 ( 
.A(n_586),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_269),
.Y(n_932)
);

CKINVDCx5p33_ASAP7_75t_R g933 ( 
.A(n_95),
.Y(n_933)
);

CKINVDCx5p33_ASAP7_75t_R g934 ( 
.A(n_267),
.Y(n_934)
);

CKINVDCx5p33_ASAP7_75t_R g935 ( 
.A(n_387),
.Y(n_935)
);

CKINVDCx20_ASAP7_75t_R g936 ( 
.A(n_120),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_472),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_71),
.Y(n_938)
);

CKINVDCx5p33_ASAP7_75t_R g939 ( 
.A(n_63),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_370),
.Y(n_940)
);

CKINVDCx5p33_ASAP7_75t_R g941 ( 
.A(n_23),
.Y(n_941)
);

CKINVDCx5p33_ASAP7_75t_R g942 ( 
.A(n_584),
.Y(n_942)
);

BUFx3_ASAP7_75t_L g943 ( 
.A(n_291),
.Y(n_943)
);

CKINVDCx5p33_ASAP7_75t_R g944 ( 
.A(n_82),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_545),
.Y(n_945)
);

CKINVDCx5p33_ASAP7_75t_R g946 ( 
.A(n_466),
.Y(n_946)
);

CKINVDCx5p33_ASAP7_75t_R g947 ( 
.A(n_137),
.Y(n_947)
);

CKINVDCx5p33_ASAP7_75t_R g948 ( 
.A(n_60),
.Y(n_948)
);

CKINVDCx5p33_ASAP7_75t_R g949 ( 
.A(n_342),
.Y(n_949)
);

CKINVDCx5p33_ASAP7_75t_R g950 ( 
.A(n_379),
.Y(n_950)
);

HB1xp67_ASAP7_75t_L g951 ( 
.A(n_403),
.Y(n_951)
);

CKINVDCx5p33_ASAP7_75t_R g952 ( 
.A(n_577),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_278),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_464),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_330),
.Y(n_955)
);

INVx2_ASAP7_75t_L g956 ( 
.A(n_292),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_241),
.Y(n_957)
);

BUFx3_ASAP7_75t_L g958 ( 
.A(n_479),
.Y(n_958)
);

INVx2_ASAP7_75t_L g959 ( 
.A(n_244),
.Y(n_959)
);

CKINVDCx5p33_ASAP7_75t_R g960 ( 
.A(n_355),
.Y(n_960)
);

CKINVDCx5p33_ASAP7_75t_R g961 ( 
.A(n_123),
.Y(n_961)
);

CKINVDCx5p33_ASAP7_75t_R g962 ( 
.A(n_453),
.Y(n_962)
);

CKINVDCx5p33_ASAP7_75t_R g963 ( 
.A(n_493),
.Y(n_963)
);

CKINVDCx5p33_ASAP7_75t_R g964 ( 
.A(n_46),
.Y(n_964)
);

CKINVDCx5p33_ASAP7_75t_R g965 ( 
.A(n_507),
.Y(n_965)
);

CKINVDCx5p33_ASAP7_75t_R g966 ( 
.A(n_530),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_578),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_535),
.Y(n_968)
);

INVx2_ASAP7_75t_L g969 ( 
.A(n_463),
.Y(n_969)
);

CKINVDCx5p33_ASAP7_75t_R g970 ( 
.A(n_41),
.Y(n_970)
);

INVx1_ASAP7_75t_SL g971 ( 
.A(n_394),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_570),
.Y(n_972)
);

CKINVDCx5p33_ASAP7_75t_R g973 ( 
.A(n_47),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_120),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_571),
.Y(n_975)
);

CKINVDCx5p33_ASAP7_75t_R g976 ( 
.A(n_191),
.Y(n_976)
);

CKINVDCx5p33_ASAP7_75t_R g977 ( 
.A(n_100),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_206),
.Y(n_978)
);

CKINVDCx5p33_ASAP7_75t_R g979 ( 
.A(n_138),
.Y(n_979)
);

CKINVDCx5p33_ASAP7_75t_R g980 ( 
.A(n_337),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_211),
.Y(n_981)
);

INVx2_ASAP7_75t_L g982 ( 
.A(n_157),
.Y(n_982)
);

CKINVDCx16_ASAP7_75t_R g983 ( 
.A(n_402),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_548),
.Y(n_984)
);

CKINVDCx5p33_ASAP7_75t_R g985 ( 
.A(n_478),
.Y(n_985)
);

CKINVDCx5p33_ASAP7_75t_R g986 ( 
.A(n_500),
.Y(n_986)
);

CKINVDCx5p33_ASAP7_75t_R g987 ( 
.A(n_521),
.Y(n_987)
);

CKINVDCx5p33_ASAP7_75t_R g988 ( 
.A(n_552),
.Y(n_988)
);

CKINVDCx5p33_ASAP7_75t_R g989 ( 
.A(n_488),
.Y(n_989)
);

CKINVDCx5p33_ASAP7_75t_R g990 ( 
.A(n_494),
.Y(n_990)
);

CKINVDCx5p33_ASAP7_75t_R g991 ( 
.A(n_37),
.Y(n_991)
);

CKINVDCx5p33_ASAP7_75t_R g992 ( 
.A(n_309),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_588),
.Y(n_993)
);

INVx2_ASAP7_75t_L g994 ( 
.A(n_512),
.Y(n_994)
);

CKINVDCx5p33_ASAP7_75t_R g995 ( 
.A(n_579),
.Y(n_995)
);

CKINVDCx5p33_ASAP7_75t_R g996 ( 
.A(n_547),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_505),
.Y(n_997)
);

INVx2_ASAP7_75t_SL g998 ( 
.A(n_212),
.Y(n_998)
);

BUFx6f_ASAP7_75t_L g999 ( 
.A(n_256),
.Y(n_999)
);

BUFx6f_ASAP7_75t_L g1000 ( 
.A(n_92),
.Y(n_1000)
);

CKINVDCx5p33_ASAP7_75t_R g1001 ( 
.A(n_574),
.Y(n_1001)
);

CKINVDCx5p33_ASAP7_75t_R g1002 ( 
.A(n_425),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_419),
.Y(n_1003)
);

CKINVDCx5p33_ASAP7_75t_R g1004 ( 
.A(n_53),
.Y(n_1004)
);

CKINVDCx5p33_ASAP7_75t_R g1005 ( 
.A(n_198),
.Y(n_1005)
);

CKINVDCx5p33_ASAP7_75t_R g1006 ( 
.A(n_560),
.Y(n_1006)
);

CKINVDCx5p33_ASAP7_75t_R g1007 ( 
.A(n_536),
.Y(n_1007)
);

BUFx10_ASAP7_75t_L g1008 ( 
.A(n_440),
.Y(n_1008)
);

CKINVDCx5p33_ASAP7_75t_R g1009 ( 
.A(n_16),
.Y(n_1009)
);

CKINVDCx5p33_ASAP7_75t_R g1010 ( 
.A(n_541),
.Y(n_1010)
);

CKINVDCx5p33_ASAP7_75t_R g1011 ( 
.A(n_167),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_589),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_124),
.Y(n_1013)
);

INVx2_ASAP7_75t_SL g1014 ( 
.A(n_207),
.Y(n_1014)
);

CKINVDCx20_ASAP7_75t_R g1015 ( 
.A(n_161),
.Y(n_1015)
);

CKINVDCx5p33_ASAP7_75t_R g1016 ( 
.A(n_350),
.Y(n_1016)
);

CKINVDCx5p33_ASAP7_75t_R g1017 ( 
.A(n_482),
.Y(n_1017)
);

CKINVDCx5p33_ASAP7_75t_R g1018 ( 
.A(n_524),
.Y(n_1018)
);

BUFx2_ASAP7_75t_L g1019 ( 
.A(n_29),
.Y(n_1019)
);

INVxp67_ASAP7_75t_SL g1020 ( 
.A(n_569),
.Y(n_1020)
);

CKINVDCx5p33_ASAP7_75t_R g1021 ( 
.A(n_73),
.Y(n_1021)
);

CKINVDCx5p33_ASAP7_75t_R g1022 ( 
.A(n_469),
.Y(n_1022)
);

CKINVDCx5p33_ASAP7_75t_R g1023 ( 
.A(n_333),
.Y(n_1023)
);

CKINVDCx5p33_ASAP7_75t_R g1024 ( 
.A(n_302),
.Y(n_1024)
);

CKINVDCx5p33_ASAP7_75t_R g1025 ( 
.A(n_471),
.Y(n_1025)
);

CKINVDCx5p33_ASAP7_75t_R g1026 ( 
.A(n_73),
.Y(n_1026)
);

CKINVDCx5p33_ASAP7_75t_R g1027 ( 
.A(n_401),
.Y(n_1027)
);

INVx1_ASAP7_75t_SL g1028 ( 
.A(n_314),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_657),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_926),
.Y(n_1030)
);

INVx2_ASAP7_75t_L g1031 ( 
.A(n_657),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_926),
.Y(n_1032)
);

CKINVDCx5p33_ASAP7_75t_R g1033 ( 
.A(n_787),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_926),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_926),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_643),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_643),
.Y(n_1037)
);

CKINVDCx20_ASAP7_75t_R g1038 ( 
.A(n_795),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_657),
.Y(n_1039)
);

INVxp33_ASAP7_75t_L g1040 ( 
.A(n_613),
.Y(n_1040)
);

HB1xp67_ASAP7_75t_L g1041 ( 
.A(n_760),
.Y(n_1041)
);

CKINVDCx20_ASAP7_75t_R g1042 ( 
.A(n_664),
.Y(n_1042)
);

BUFx5_ASAP7_75t_L g1043 ( 
.A(n_640),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_657),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_657),
.Y(n_1045)
);

CKINVDCx5p33_ASAP7_75t_R g1046 ( 
.A(n_610),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_657),
.Y(n_1047)
);

INVxp67_ASAP7_75t_SL g1048 ( 
.A(n_643),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_657),
.Y(n_1049)
);

BUFx3_ASAP7_75t_L g1050 ( 
.A(n_640),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_657),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_657),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_885),
.Y(n_1053)
);

CKINVDCx20_ASAP7_75t_R g1054 ( 
.A(n_724),
.Y(n_1054)
);

CKINVDCx5p33_ASAP7_75t_R g1055 ( 
.A(n_610),
.Y(n_1055)
);

INVx2_ASAP7_75t_SL g1056 ( 
.A(n_644),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_885),
.Y(n_1057)
);

CKINVDCx20_ASAP7_75t_R g1058 ( 
.A(n_603),
.Y(n_1058)
);

HB1xp67_ASAP7_75t_L g1059 ( 
.A(n_760),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_644),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_644),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_885),
.Y(n_1062)
);

CKINVDCx16_ASAP7_75t_R g1063 ( 
.A(n_673),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_701),
.Y(n_1064)
);

CKINVDCx20_ASAP7_75t_R g1065 ( 
.A(n_606),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_885),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_701),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_701),
.Y(n_1068)
);

BUFx2_ASAP7_75t_L g1069 ( 
.A(n_772),
.Y(n_1069)
);

INVxp67_ASAP7_75t_SL g1070 ( 
.A(n_733),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_733),
.Y(n_1071)
);

INVx2_ASAP7_75t_L g1072 ( 
.A(n_885),
.Y(n_1072)
);

INVx2_ASAP7_75t_L g1073 ( 
.A(n_885),
.Y(n_1073)
);

CKINVDCx5p33_ASAP7_75t_R g1074 ( 
.A(n_673),
.Y(n_1074)
);

INVxp33_ASAP7_75t_SL g1075 ( 
.A(n_642),
.Y(n_1075)
);

INVx2_ASAP7_75t_L g1076 ( 
.A(n_885),
.Y(n_1076)
);

CKINVDCx5p33_ASAP7_75t_R g1077 ( 
.A(n_681),
.Y(n_1077)
);

INVxp67_ASAP7_75t_SL g1078 ( 
.A(n_733),
.Y(n_1078)
);

CKINVDCx5p33_ASAP7_75t_R g1079 ( 
.A(n_681),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_885),
.Y(n_1080)
);

INVxp67_ASAP7_75t_SL g1081 ( 
.A(n_779),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_779),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_885),
.Y(n_1083)
);

CKINVDCx5p33_ASAP7_75t_R g1084 ( 
.A(n_761),
.Y(n_1084)
);

CKINVDCx5p33_ASAP7_75t_R g1085 ( 
.A(n_761),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_779),
.Y(n_1086)
);

BUFx2_ASAP7_75t_L g1087 ( 
.A(n_772),
.Y(n_1087)
);

HB1xp67_ASAP7_75t_L g1088 ( 
.A(n_781),
.Y(n_1088)
);

CKINVDCx16_ASAP7_75t_R g1089 ( 
.A(n_895),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_799),
.Y(n_1090)
);

CKINVDCx20_ASAP7_75t_R g1091 ( 
.A(n_622),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_822),
.Y(n_1092)
);

CKINVDCx20_ASAP7_75t_R g1093 ( 
.A(n_652),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_822),
.Y(n_1094)
);

INVxp33_ASAP7_75t_L g1095 ( 
.A(n_951),
.Y(n_1095)
);

INVxp33_ASAP7_75t_SL g1096 ( 
.A(n_781),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_967),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_967),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_972),
.Y(n_1099)
);

CKINVDCx5p33_ASAP7_75t_R g1100 ( 
.A(n_895),
.Y(n_1100)
);

CKINVDCx20_ASAP7_75t_R g1101 ( 
.A(n_675),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_972),
.Y(n_1102)
);

INVxp67_ASAP7_75t_SL g1103 ( 
.A(n_799),
.Y(n_1103)
);

INVx4_ASAP7_75t_L g1104 ( 
.A(n_1050),
.Y(n_1104)
);

CKINVDCx5p33_ASAP7_75t_R g1105 ( 
.A(n_1042),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_1029),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_1030),
.B(n_975),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_1029),
.Y(n_1108)
);

NAND3xp33_ASAP7_75t_L g1109 ( 
.A(n_1092),
.B(n_595),
.C(n_594),
.Y(n_1109)
);

CKINVDCx16_ASAP7_75t_R g1110 ( 
.A(n_1063),
.Y(n_1110)
);

OAI21x1_ASAP7_75t_L g1111 ( 
.A1(n_1031),
.A2(n_1073),
.B(n_1072),
.Y(n_1111)
);

AND2x4_ASAP7_75t_L g1112 ( 
.A(n_1050),
.B(n_1092),
.Y(n_1112)
);

CKINVDCx6p67_ASAP7_75t_R g1113 ( 
.A(n_1089),
.Y(n_1113)
);

INVx4_ASAP7_75t_L g1114 ( 
.A(n_1043),
.Y(n_1114)
);

INVxp67_ASAP7_75t_L g1115 ( 
.A(n_1041),
.Y(n_1115)
);

BUFx2_ASAP7_75t_L g1116 ( 
.A(n_1046),
.Y(n_1116)
);

AND2x2_ASAP7_75t_L g1117 ( 
.A(n_1094),
.B(n_799),
.Y(n_1117)
);

INVx2_ASAP7_75t_L g1118 ( 
.A(n_1031),
.Y(n_1118)
);

BUFx6f_ASAP7_75t_L g1119 ( 
.A(n_1072),
.Y(n_1119)
);

BUFx8_ASAP7_75t_SL g1120 ( 
.A(n_1058),
.Y(n_1120)
);

OA21x2_ASAP7_75t_L g1121 ( 
.A1(n_1094),
.A2(n_993),
.B(n_975),
.Y(n_1121)
);

AND2x4_ASAP7_75t_L g1122 ( 
.A(n_1097),
.B(n_814),
.Y(n_1122)
);

BUFx2_ASAP7_75t_L g1123 ( 
.A(n_1046),
.Y(n_1123)
);

INVx2_ASAP7_75t_L g1124 ( 
.A(n_1073),
.Y(n_1124)
);

INVx2_ASAP7_75t_L g1125 ( 
.A(n_1076),
.Y(n_1125)
);

BUFx6f_ASAP7_75t_L g1126 ( 
.A(n_1076),
.Y(n_1126)
);

AND2x2_ASAP7_75t_L g1127 ( 
.A(n_1097),
.B(n_814),
.Y(n_1127)
);

OAI21x1_ASAP7_75t_L g1128 ( 
.A1(n_1039),
.A2(n_800),
.B(n_630),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_1039),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_1044),
.Y(n_1130)
);

AND2x4_ASAP7_75t_L g1131 ( 
.A(n_1098),
.B(n_814),
.Y(n_1131)
);

INVx3_ASAP7_75t_L g1132 ( 
.A(n_1044),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_1045),
.Y(n_1133)
);

INVx3_ASAP7_75t_L g1134 ( 
.A(n_1045),
.Y(n_1134)
);

AND2x2_ASAP7_75t_L g1135 ( 
.A(n_1098),
.B(n_1099),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_SL g1136 ( 
.A(n_1033),
.B(n_702),
.Y(n_1136)
);

BUFx8_ASAP7_75t_L g1137 ( 
.A(n_1069),
.Y(n_1137)
);

OAI22xp5_ASAP7_75t_L g1138 ( 
.A1(n_1096),
.A2(n_983),
.B1(n_690),
.B2(n_737),
.Y(n_1138)
);

BUFx6f_ASAP7_75t_L g1139 ( 
.A(n_1047),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_1047),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_1049),
.Y(n_1141)
);

INVx3_ASAP7_75t_L g1142 ( 
.A(n_1049),
.Y(n_1142)
);

INVx2_ASAP7_75t_L g1143 ( 
.A(n_1051),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_1032),
.B(n_993),
.Y(n_1144)
);

AOI22xp5_ASAP7_75t_SL g1145 ( 
.A1(n_1065),
.A2(n_767),
.B1(n_784),
.B2(n_677),
.Y(n_1145)
);

INVx2_ASAP7_75t_L g1146 ( 
.A(n_1051),
.Y(n_1146)
);

AND2x4_ASAP7_75t_L g1147 ( 
.A(n_1099),
.B(n_864),
.Y(n_1147)
);

INVx2_ASAP7_75t_L g1148 ( 
.A(n_1052),
.Y(n_1148)
);

OA21x2_ASAP7_75t_L g1149 ( 
.A1(n_1102),
.A2(n_1012),
.B(n_856),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_1053),
.Y(n_1150)
);

OAI21x1_ASAP7_75t_L g1151 ( 
.A1(n_1053),
.A2(n_800),
.B(n_630),
.Y(n_1151)
);

INVx2_ASAP7_75t_L g1152 ( 
.A(n_1057),
.Y(n_1152)
);

OAI21x1_ASAP7_75t_L g1153 ( 
.A1(n_1057),
.A2(n_1066),
.B(n_1062),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_1062),
.Y(n_1154)
);

INVx4_ASAP7_75t_L g1155 ( 
.A(n_1043),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_1066),
.Y(n_1156)
);

AND2x2_ASAP7_75t_SL g1157 ( 
.A(n_1102),
.B(n_630),
.Y(n_1157)
);

NOR2x1_ASAP7_75t_L g1158 ( 
.A(n_1036),
.B(n_1012),
.Y(n_1158)
);

INVx4_ASAP7_75t_L g1159 ( 
.A(n_1043),
.Y(n_1159)
);

OAI22x1_ASAP7_75t_R g1160 ( 
.A1(n_1091),
.A2(n_807),
.B1(n_828),
.B2(n_801),
.Y(n_1160)
);

INVx2_ASAP7_75t_L g1161 ( 
.A(n_1080),
.Y(n_1161)
);

INVx2_ASAP7_75t_L g1162 ( 
.A(n_1080),
.Y(n_1162)
);

INVx2_ASAP7_75t_L g1163 ( 
.A(n_1083),
.Y(n_1163)
);

CKINVDCx20_ASAP7_75t_R g1164 ( 
.A(n_1120),
.Y(n_1164)
);

CKINVDCx5p33_ASAP7_75t_R g1165 ( 
.A(n_1120),
.Y(n_1165)
);

CKINVDCx5p33_ASAP7_75t_R g1166 ( 
.A(n_1105),
.Y(n_1166)
);

OAI22xp5_ASAP7_75t_SL g1167 ( 
.A1(n_1138),
.A2(n_1101),
.B1(n_1093),
.B2(n_884),
.Y(n_1167)
);

BUFx6f_ASAP7_75t_L g1168 ( 
.A(n_1119),
.Y(n_1168)
);

CKINVDCx5p33_ASAP7_75t_R g1169 ( 
.A(n_1113),
.Y(n_1169)
);

CKINVDCx5p33_ASAP7_75t_R g1170 ( 
.A(n_1113),
.Y(n_1170)
);

CKINVDCx20_ASAP7_75t_R g1171 ( 
.A(n_1113),
.Y(n_1171)
);

HB1xp67_ASAP7_75t_L g1172 ( 
.A(n_1110),
.Y(n_1172)
);

NOR2xp33_ASAP7_75t_R g1173 ( 
.A(n_1110),
.B(n_1054),
.Y(n_1173)
);

CKINVDCx5p33_ASAP7_75t_R g1174 ( 
.A(n_1137),
.Y(n_1174)
);

INVx3_ASAP7_75t_L g1175 ( 
.A(n_1132),
.Y(n_1175)
);

NOR2xp67_ASAP7_75t_L g1176 ( 
.A(n_1115),
.B(n_1055),
.Y(n_1176)
);

INVx2_ASAP7_75t_L g1177 ( 
.A(n_1111),
.Y(n_1177)
);

CKINVDCx5p33_ASAP7_75t_R g1178 ( 
.A(n_1137),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_1135),
.Y(n_1179)
);

CKINVDCx5p33_ASAP7_75t_R g1180 ( 
.A(n_1137),
.Y(n_1180)
);

NOR2xp67_ASAP7_75t_L g1181 ( 
.A(n_1115),
.B(n_1055),
.Y(n_1181)
);

CKINVDCx5p33_ASAP7_75t_R g1182 ( 
.A(n_1137),
.Y(n_1182)
);

CKINVDCx5p33_ASAP7_75t_R g1183 ( 
.A(n_1137),
.Y(n_1183)
);

NOR2xp33_ASAP7_75t_R g1184 ( 
.A(n_1116),
.B(n_1033),
.Y(n_1184)
);

CKINVDCx16_ASAP7_75t_R g1185 ( 
.A(n_1160),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_1135),
.Y(n_1186)
);

CKINVDCx5p33_ASAP7_75t_R g1187 ( 
.A(n_1116),
.Y(n_1187)
);

CKINVDCx5p33_ASAP7_75t_R g1188 ( 
.A(n_1116),
.Y(n_1188)
);

CKINVDCx20_ASAP7_75t_R g1189 ( 
.A(n_1123),
.Y(n_1189)
);

NOR2xp33_ASAP7_75t_R g1190 ( 
.A(n_1123),
.B(n_1074),
.Y(n_1190)
);

NOR2xp33_ASAP7_75t_L g1191 ( 
.A(n_1136),
.B(n_1079),
.Y(n_1191)
);

INVx2_ASAP7_75t_L g1192 ( 
.A(n_1111),
.Y(n_1192)
);

CKINVDCx5p33_ASAP7_75t_R g1193 ( 
.A(n_1123),
.Y(n_1193)
);

BUFx6f_ASAP7_75t_L g1194 ( 
.A(n_1119),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_1135),
.Y(n_1195)
);

CKINVDCx5p33_ASAP7_75t_R g1196 ( 
.A(n_1138),
.Y(n_1196)
);

CKINVDCx20_ASAP7_75t_R g1197 ( 
.A(n_1160),
.Y(n_1197)
);

NOR2xp67_ASAP7_75t_L g1198 ( 
.A(n_1104),
.B(n_1074),
.Y(n_1198)
);

NOR2xp67_ASAP7_75t_L g1199 ( 
.A(n_1104),
.B(n_1077),
.Y(n_1199)
);

CKINVDCx5p33_ASAP7_75t_R g1200 ( 
.A(n_1145),
.Y(n_1200)
);

INVxp67_ASAP7_75t_SL g1201 ( 
.A(n_1132),
.Y(n_1201)
);

CKINVDCx20_ASAP7_75t_R g1202 ( 
.A(n_1145),
.Y(n_1202)
);

CKINVDCx20_ASAP7_75t_R g1203 ( 
.A(n_1136),
.Y(n_1203)
);

CKINVDCx20_ASAP7_75t_R g1204 ( 
.A(n_1117),
.Y(n_1204)
);

CKINVDCx5p33_ASAP7_75t_R g1205 ( 
.A(n_1157),
.Y(n_1205)
);

CKINVDCx5p33_ASAP7_75t_R g1206 ( 
.A(n_1157),
.Y(n_1206)
);

INVxp67_ASAP7_75t_L g1207 ( 
.A(n_1117),
.Y(n_1207)
);

CKINVDCx5p33_ASAP7_75t_R g1208 ( 
.A(n_1157),
.Y(n_1208)
);

CKINVDCx20_ASAP7_75t_R g1209 ( 
.A(n_1117),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1143),
.Y(n_1210)
);

INVx2_ASAP7_75t_L g1211 ( 
.A(n_1111),
.Y(n_1211)
);

NOR2xp33_ASAP7_75t_R g1212 ( 
.A(n_1132),
.B(n_1077),
.Y(n_1212)
);

HB1xp67_ASAP7_75t_L g1213 ( 
.A(n_1112),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_1143),
.Y(n_1214)
);

INVx3_ASAP7_75t_L g1215 ( 
.A(n_1132),
.Y(n_1215)
);

CKINVDCx5p33_ASAP7_75t_R g1216 ( 
.A(n_1157),
.Y(n_1216)
);

INVx1_ASAP7_75t_SL g1217 ( 
.A(n_1127),
.Y(n_1217)
);

CKINVDCx5p33_ASAP7_75t_R g1218 ( 
.A(n_1112),
.Y(n_1218)
);

INVx3_ASAP7_75t_L g1219 ( 
.A(n_1132),
.Y(n_1219)
);

CKINVDCx20_ASAP7_75t_R g1220 ( 
.A(n_1127),
.Y(n_1220)
);

NOR2xp33_ASAP7_75t_R g1221 ( 
.A(n_1134),
.B(n_1079),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1210),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1214),
.Y(n_1223)
);

BUFx3_ASAP7_75t_L g1224 ( 
.A(n_1169),
.Y(n_1224)
);

AND2x2_ASAP7_75t_L g1225 ( 
.A(n_1217),
.B(n_1112),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_1206),
.B(n_1104),
.Y(n_1226)
);

INVx2_ASAP7_75t_L g1227 ( 
.A(n_1177),
.Y(n_1227)
);

AND2x6_ASAP7_75t_L g1228 ( 
.A(n_1177),
.B(n_1127),
.Y(n_1228)
);

INVx2_ASAP7_75t_L g1229 ( 
.A(n_1192),
.Y(n_1229)
);

AND2x2_ASAP7_75t_L g1230 ( 
.A(n_1207),
.B(n_1112),
.Y(n_1230)
);

INVxp67_ASAP7_75t_L g1231 ( 
.A(n_1172),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1213),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1175),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1175),
.Y(n_1234)
);

BUFx6f_ASAP7_75t_L g1235 ( 
.A(n_1168),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_1206),
.B(n_1104),
.Y(n_1236)
);

AOI22xp33_ASAP7_75t_L g1237 ( 
.A1(n_1208),
.A2(n_1075),
.B1(n_1158),
.B2(n_1121),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1175),
.Y(n_1238)
);

INVx2_ASAP7_75t_L g1239 ( 
.A(n_1192),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1215),
.Y(n_1240)
);

INVx3_ASAP7_75t_L g1241 ( 
.A(n_1215),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_L g1242 ( 
.A(n_1208),
.B(n_1104),
.Y(n_1242)
);

NOR2xp33_ASAP7_75t_L g1243 ( 
.A(n_1191),
.B(n_1084),
.Y(n_1243)
);

BUFx6f_ASAP7_75t_L g1244 ( 
.A(n_1168),
.Y(n_1244)
);

CKINVDCx5p33_ASAP7_75t_R g1245 ( 
.A(n_1166),
.Y(n_1245)
);

INVx2_ASAP7_75t_L g1246 ( 
.A(n_1211),
.Y(n_1246)
);

INVxp67_ASAP7_75t_SL g1247 ( 
.A(n_1215),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1219),
.Y(n_1248)
);

INVx4_ASAP7_75t_L g1249 ( 
.A(n_1219),
.Y(n_1249)
);

BUFx8_ASAP7_75t_SL g1250 ( 
.A(n_1164),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1219),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1179),
.Y(n_1252)
);

INVx2_ASAP7_75t_L g1253 ( 
.A(n_1211),
.Y(n_1253)
);

BUFx6f_ASAP7_75t_L g1254 ( 
.A(n_1168),
.Y(n_1254)
);

AND2x6_ASAP7_75t_L g1255 ( 
.A(n_1186),
.B(n_1122),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1195),
.Y(n_1256)
);

INVx1_ASAP7_75t_SL g1257 ( 
.A(n_1189),
.Y(n_1257)
);

INVx1_ASAP7_75t_SL g1258 ( 
.A(n_1173),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1201),
.Y(n_1259)
);

OAI22xp33_ASAP7_75t_L g1260 ( 
.A1(n_1205),
.A2(n_983),
.B1(n_1085),
.B2(n_1084),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_L g1261 ( 
.A(n_1216),
.B(n_1112),
.Y(n_1261)
);

NOR2xp33_ASAP7_75t_L g1262 ( 
.A(n_1203),
.B(n_1085),
.Y(n_1262)
);

INVx5_ASAP7_75t_L g1263 ( 
.A(n_1168),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1218),
.Y(n_1264)
);

INVxp67_ASAP7_75t_L g1265 ( 
.A(n_1187),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_SL g1266 ( 
.A(n_1212),
.B(n_1100),
.Y(n_1266)
);

CKINVDCx20_ASAP7_75t_R g1267 ( 
.A(n_1167),
.Y(n_1267)
);

AND2x4_ASAP7_75t_L g1268 ( 
.A(n_1218),
.B(n_1122),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_SL g1269 ( 
.A(n_1221),
.B(n_1100),
.Y(n_1269)
);

INVx3_ASAP7_75t_L g1270 ( 
.A(n_1168),
.Y(n_1270)
);

INVx3_ASAP7_75t_L g1271 ( 
.A(n_1194),
.Y(n_1271)
);

CKINVDCx5p33_ASAP7_75t_R g1272 ( 
.A(n_1166),
.Y(n_1272)
);

BUFx3_ASAP7_75t_L g1273 ( 
.A(n_1169),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1194),
.Y(n_1274)
);

INVx2_ASAP7_75t_L g1275 ( 
.A(n_1194),
.Y(n_1275)
);

NAND2x1p5_ASAP7_75t_L g1276 ( 
.A(n_1194),
.B(n_1149),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1194),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1204),
.Y(n_1278)
);

INVx2_ASAP7_75t_L g1279 ( 
.A(n_1209),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_L g1280 ( 
.A(n_1198),
.B(n_1122),
.Y(n_1280)
);

NOR2xp33_ASAP7_75t_L g1281 ( 
.A(n_1188),
.B(n_1038),
.Y(n_1281)
);

CKINVDCx20_ASAP7_75t_R g1282 ( 
.A(n_1193),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1220),
.Y(n_1283)
);

INVx2_ASAP7_75t_L g1284 ( 
.A(n_1193),
.Y(n_1284)
);

INVx2_ASAP7_75t_SL g1285 ( 
.A(n_1184),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_SL g1286 ( 
.A(n_1176),
.B(n_1122),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1199),
.Y(n_1287)
);

INVx2_ASAP7_75t_L g1288 ( 
.A(n_1196),
.Y(n_1288)
);

INVx2_ASAP7_75t_L g1289 ( 
.A(n_1174),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1181),
.Y(n_1290)
);

NOR2xp33_ASAP7_75t_L g1291 ( 
.A(n_1178),
.B(n_1040),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1180),
.Y(n_1292)
);

AO22x2_ASAP7_75t_L g1293 ( 
.A1(n_1200),
.A2(n_1109),
.B1(n_594),
.B2(n_615),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_L g1294 ( 
.A(n_1190),
.B(n_1122),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_SL g1295 ( 
.A(n_1182),
.B(n_1131),
.Y(n_1295)
);

INVx2_ASAP7_75t_L g1296 ( 
.A(n_1183),
.Y(n_1296)
);

AND2x6_ASAP7_75t_L g1297 ( 
.A(n_1170),
.B(n_1131),
.Y(n_1297)
);

BUFx6f_ASAP7_75t_L g1298 ( 
.A(n_1170),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1171),
.Y(n_1299)
);

INVx2_ASAP7_75t_SL g1300 ( 
.A(n_1268),
.Y(n_1300)
);

NOR2xp33_ASAP7_75t_L g1301 ( 
.A(n_1243),
.B(n_1200),
.Y(n_1301)
);

AND2x2_ASAP7_75t_L g1302 ( 
.A(n_1288),
.B(n_1095),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1252),
.Y(n_1303)
);

INVxp67_ASAP7_75t_SL g1304 ( 
.A(n_1268),
.Y(n_1304)
);

INVx1_ASAP7_75t_SL g1305 ( 
.A(n_1257),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_SL g1306 ( 
.A(n_1249),
.B(n_1235),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1256),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_L g1308 ( 
.A(n_1225),
.B(n_1131),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_1225),
.B(n_1131),
.Y(n_1309)
);

CKINVDCx5p33_ASAP7_75t_R g1310 ( 
.A(n_1245),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_SL g1311 ( 
.A(n_1249),
.B(n_1134),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_L g1312 ( 
.A(n_1230),
.B(n_1131),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_L g1313 ( 
.A(n_1230),
.B(n_1147),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_L g1314 ( 
.A(n_1261),
.B(n_1147),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1232),
.Y(n_1315)
);

AOI22xp33_ASAP7_75t_L g1316 ( 
.A1(n_1293),
.A2(n_1197),
.B1(n_892),
.B2(n_906),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_L g1317 ( 
.A(n_1237),
.B(n_1147),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1222),
.Y(n_1318)
);

AND2x2_ASAP7_75t_L g1319 ( 
.A(n_1288),
.B(n_1185),
.Y(n_1319)
);

OAI221xp5_ASAP7_75t_L g1320 ( 
.A1(n_1284),
.A2(n_1087),
.B1(n_1069),
.B2(n_1088),
.C(n_1059),
.Y(n_1320)
);

NAND2xp5_ASAP7_75t_L g1321 ( 
.A(n_1259),
.B(n_1147),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_SL g1322 ( 
.A(n_1249),
.B(n_1134),
.Y(n_1322)
);

AOI22xp5_ASAP7_75t_L g1323 ( 
.A1(n_1264),
.A2(n_916),
.B1(n_919),
.B2(n_871),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_L g1324 ( 
.A(n_1268),
.B(n_1147),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_L g1325 ( 
.A(n_1290),
.B(n_1158),
.Y(n_1325)
);

INVxp67_ASAP7_75t_L g1326 ( 
.A(n_1291),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_SL g1327 ( 
.A(n_1235),
.B(n_1134),
.Y(n_1327)
);

NOR2x1p5_ASAP7_75t_L g1328 ( 
.A(n_1245),
.B(n_1165),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1222),
.Y(n_1329)
);

NAND2xp5_ASAP7_75t_SL g1330 ( 
.A(n_1235),
.B(n_1134),
.Y(n_1330)
);

NAND2xp5_ASAP7_75t_L g1331 ( 
.A(n_1290),
.B(n_1048),
.Y(n_1331)
);

NAND2xp5_ASAP7_75t_SL g1332 ( 
.A(n_1235),
.B(n_1142),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_SL g1333 ( 
.A(n_1235),
.B(n_1142),
.Y(n_1333)
);

NAND2xp5_ASAP7_75t_L g1334 ( 
.A(n_1294),
.B(n_1070),
.Y(n_1334)
);

CKINVDCx5p33_ASAP7_75t_R g1335 ( 
.A(n_1272),
.Y(n_1335)
);

INVx2_ASAP7_75t_L g1336 ( 
.A(n_1227),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_L g1337 ( 
.A(n_1286),
.B(n_1078),
.Y(n_1337)
);

INVx2_ASAP7_75t_L g1338 ( 
.A(n_1227),
.Y(n_1338)
);

NOR2xp33_ASAP7_75t_L g1339 ( 
.A(n_1265),
.B(n_1165),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_L g1340 ( 
.A(n_1255),
.B(n_1081),
.Y(n_1340)
);

NOR2xp33_ASAP7_75t_L g1341 ( 
.A(n_1284),
.B(n_1087),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1223),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_L g1343 ( 
.A(n_1255),
.B(n_1103),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1223),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1234),
.Y(n_1345)
);

NAND2xp5_ASAP7_75t_L g1346 ( 
.A(n_1255),
.B(n_1142),
.Y(n_1346)
);

INVxp67_ASAP7_75t_L g1347 ( 
.A(n_1262),
.Y(n_1347)
);

NOR2xp33_ASAP7_75t_L g1348 ( 
.A(n_1281),
.B(n_1260),
.Y(n_1348)
);

AND2x2_ASAP7_75t_SL g1349 ( 
.A(n_1298),
.B(n_1121),
.Y(n_1349)
);

O2A1O1Ixp33_ASAP7_75t_L g1350 ( 
.A1(n_1266),
.A2(n_1269),
.B(n_1238),
.C(n_1240),
.Y(n_1350)
);

AOI22xp33_ASAP7_75t_L g1351 ( 
.A1(n_1293),
.A2(n_936),
.B1(n_1015),
.B2(n_924),
.Y(n_1351)
);

AOI22xp5_ASAP7_75t_L g1352 ( 
.A1(n_1297),
.A2(n_1020),
.B1(n_620),
.B2(n_663),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_L g1353 ( 
.A(n_1255),
.B(n_1142),
.Y(n_1353)
);

NOR2xp33_ASAP7_75t_L g1354 ( 
.A(n_1231),
.B(n_1202),
.Y(n_1354)
);

NAND2x1p5_ASAP7_75t_L g1355 ( 
.A(n_1263),
.B(n_1121),
.Y(n_1355)
);

NAND2xp5_ASAP7_75t_L g1356 ( 
.A(n_1255),
.B(n_1142),
.Y(n_1356)
);

AOI22xp33_ASAP7_75t_L g1357 ( 
.A1(n_1293),
.A2(n_1121),
.B1(n_1109),
.B2(n_847),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_L g1358 ( 
.A(n_1255),
.B(n_1107),
.Y(n_1358)
);

INVx2_ASAP7_75t_L g1359 ( 
.A(n_1229),
.Y(n_1359)
);

NOR2xp33_ASAP7_75t_L g1360 ( 
.A(n_1282),
.B(n_1114),
.Y(n_1360)
);

INVx2_ASAP7_75t_SL g1361 ( 
.A(n_1255),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1234),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1238),
.Y(n_1363)
);

NOR2xp33_ASAP7_75t_L g1364 ( 
.A(n_1282),
.B(n_1114),
.Y(n_1364)
);

NAND2xp5_ASAP7_75t_SL g1365 ( 
.A(n_1244),
.B(n_1106),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_L g1366 ( 
.A(n_1247),
.B(n_1241),
.Y(n_1366)
);

NOR2xp33_ASAP7_75t_L g1367 ( 
.A(n_1285),
.B(n_1272),
.Y(n_1367)
);

NAND3xp33_ASAP7_75t_L g1368 ( 
.A(n_1278),
.B(n_647),
.C(n_789),
.Y(n_1368)
);

AND2x2_ASAP7_75t_L g1369 ( 
.A(n_1285),
.B(n_1056),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_SL g1370 ( 
.A(n_1244),
.B(n_1106),
.Y(n_1370)
);

CKINVDCx20_ASAP7_75t_R g1371 ( 
.A(n_1250),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_L g1372 ( 
.A(n_1241),
.B(n_1107),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_L g1373 ( 
.A(n_1241),
.B(n_1144),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1240),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_L g1375 ( 
.A(n_1297),
.B(n_1144),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_L g1376 ( 
.A(n_1297),
.B(n_1108),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_L g1377 ( 
.A(n_1297),
.B(n_1108),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1248),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1248),
.Y(n_1379)
);

INVx2_ASAP7_75t_L g1380 ( 
.A(n_1229),
.Y(n_1380)
);

INVx2_ASAP7_75t_L g1381 ( 
.A(n_1239),
.Y(n_1381)
);

INVx2_ASAP7_75t_SL g1382 ( 
.A(n_1228),
.Y(n_1382)
);

A2O1A1Ixp33_ASAP7_75t_L g1383 ( 
.A1(n_1233),
.A2(n_1151),
.B(n_1128),
.C(n_847),
.Y(n_1383)
);

AND2x2_ASAP7_75t_L g1384 ( 
.A(n_1279),
.B(n_1056),
.Y(n_1384)
);

NOR2xp33_ASAP7_75t_L g1385 ( 
.A(n_1298),
.B(n_1114),
.Y(n_1385)
);

NAND2xp5_ASAP7_75t_SL g1386 ( 
.A(n_1244),
.B(n_1129),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_SL g1387 ( 
.A(n_1244),
.B(n_1129),
.Y(n_1387)
);

INVx2_ASAP7_75t_L g1388 ( 
.A(n_1239),
.Y(n_1388)
);

NOR3xp33_ASAP7_75t_L g1389 ( 
.A(n_1278),
.B(n_1019),
.C(n_789),
.Y(n_1389)
);

INVxp67_ASAP7_75t_L g1390 ( 
.A(n_1283),
.Y(n_1390)
);

A2O1A1Ixp33_ASAP7_75t_L g1391 ( 
.A1(n_1251),
.A2(n_1128),
.B(n_1151),
.C(n_1019),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1297),
.B(n_1130),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1246),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_L g1394 ( 
.A(n_1297),
.B(n_1130),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_SL g1395 ( 
.A(n_1244),
.B(n_1133),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1246),
.Y(n_1396)
);

BUFx2_ASAP7_75t_R g1397 ( 
.A(n_1224),
.Y(n_1397)
);

NOR2xp33_ASAP7_75t_L g1398 ( 
.A(n_1298),
.B(n_1155),
.Y(n_1398)
);

NAND2xp33_ASAP7_75t_L g1399 ( 
.A(n_1228),
.B(n_1139),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1253),
.Y(n_1400)
);

CKINVDCx5p33_ASAP7_75t_R g1401 ( 
.A(n_1224),
.Y(n_1401)
);

INVx2_ASAP7_75t_SL g1402 ( 
.A(n_1228),
.Y(n_1402)
);

AND2x2_ASAP7_75t_SL g1403 ( 
.A(n_1301),
.B(n_1298),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_SL g1404 ( 
.A(n_1349),
.B(n_1254),
.Y(n_1404)
);

AOI21xp5_ASAP7_75t_L g1405 ( 
.A1(n_1399),
.A2(n_1253),
.B(n_1280),
.Y(n_1405)
);

NOR2xp33_ASAP7_75t_L g1406 ( 
.A(n_1348),
.B(n_1279),
.Y(n_1406)
);

AOI21xp5_ASAP7_75t_L g1407 ( 
.A1(n_1399),
.A2(n_1275),
.B(n_1274),
.Y(n_1407)
);

AND2x2_ASAP7_75t_L g1408 ( 
.A(n_1302),
.B(n_1283),
.Y(n_1408)
);

AOI21xp5_ASAP7_75t_L g1409 ( 
.A1(n_1385),
.A2(n_1275),
.B(n_1274),
.Y(n_1409)
);

NAND2xp5_ASAP7_75t_SL g1410 ( 
.A(n_1349),
.B(n_1254),
.Y(n_1410)
);

AOI21xp5_ASAP7_75t_L g1411 ( 
.A1(n_1398),
.A2(n_1277),
.B(n_1254),
.Y(n_1411)
);

CKINVDCx8_ASAP7_75t_R g1412 ( 
.A(n_1310),
.Y(n_1412)
);

CKINVDCx5p33_ASAP7_75t_R g1413 ( 
.A(n_1371),
.Y(n_1413)
);

NOR2xp33_ASAP7_75t_L g1414 ( 
.A(n_1347),
.B(n_1298),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_L g1415 ( 
.A(n_1304),
.B(n_1297),
.Y(n_1415)
);

AOI21xp5_ASAP7_75t_L g1416 ( 
.A1(n_1366),
.A2(n_1277),
.B(n_1254),
.Y(n_1416)
);

NAND2xp5_ASAP7_75t_L g1417 ( 
.A(n_1326),
.B(n_1289),
.Y(n_1417)
);

INVx2_ASAP7_75t_SL g1418 ( 
.A(n_1335),
.Y(n_1418)
);

AOI21xp5_ASAP7_75t_L g1419 ( 
.A1(n_1376),
.A2(n_1254),
.B(n_1270),
.Y(n_1419)
);

INVx2_ASAP7_75t_L g1420 ( 
.A(n_1336),
.Y(n_1420)
);

INVx2_ASAP7_75t_L g1421 ( 
.A(n_1336),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_L g1422 ( 
.A(n_1360),
.B(n_1364),
.Y(n_1422)
);

INVx3_ASAP7_75t_L g1423 ( 
.A(n_1361),
.Y(n_1423)
);

AND2x2_ASAP7_75t_L g1424 ( 
.A(n_1319),
.B(n_1341),
.Y(n_1424)
);

INVx1_ASAP7_75t_SL g1425 ( 
.A(n_1305),
.Y(n_1425)
);

INVx2_ASAP7_75t_L g1426 ( 
.A(n_1338),
.Y(n_1426)
);

AOI21xp5_ASAP7_75t_L g1427 ( 
.A1(n_1377),
.A2(n_1271),
.B(n_1270),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1315),
.Y(n_1428)
);

NAND2xp5_ASAP7_75t_L g1429 ( 
.A(n_1300),
.B(n_1289),
.Y(n_1429)
);

NAND2xp5_ASAP7_75t_L g1430 ( 
.A(n_1300),
.B(n_1296),
.Y(n_1430)
);

BUFx3_ASAP7_75t_L g1431 ( 
.A(n_1401),
.Y(n_1431)
);

AOI21xp5_ASAP7_75t_L g1432 ( 
.A1(n_1392),
.A2(n_1271),
.B(n_1270),
.Y(n_1432)
);

AOI21xp5_ASAP7_75t_L g1433 ( 
.A1(n_1394),
.A2(n_1271),
.B(n_1287),
.Y(n_1433)
);

AOI21x1_ASAP7_75t_L g1434 ( 
.A1(n_1306),
.A2(n_1287),
.B(n_1236),
.Y(n_1434)
);

OAI22xp5_ASAP7_75t_L g1435 ( 
.A1(n_1358),
.A2(n_1242),
.B1(n_1226),
.B2(n_1263),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1303),
.Y(n_1436)
);

BUFx6f_ASAP7_75t_L g1437 ( 
.A(n_1382),
.Y(n_1437)
);

AOI21xp5_ASAP7_75t_L g1438 ( 
.A1(n_1311),
.A2(n_1263),
.B(n_1276),
.Y(n_1438)
);

BUFx6f_ASAP7_75t_L g1439 ( 
.A(n_1382),
.Y(n_1439)
);

NOR2xp33_ASAP7_75t_L g1440 ( 
.A(n_1390),
.B(n_1273),
.Y(n_1440)
);

BUFx6f_ASAP7_75t_L g1441 ( 
.A(n_1402),
.Y(n_1441)
);

BUFx3_ASAP7_75t_L g1442 ( 
.A(n_1401),
.Y(n_1442)
);

AOI21xp5_ASAP7_75t_L g1443 ( 
.A1(n_1311),
.A2(n_1263),
.B(n_1276),
.Y(n_1443)
);

AOI21xp5_ASAP7_75t_L g1444 ( 
.A1(n_1322),
.A2(n_1263),
.B(n_1276),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1307),
.Y(n_1445)
);

AND2x2_ASAP7_75t_L g1446 ( 
.A(n_1354),
.B(n_1273),
.Y(n_1446)
);

NAND2xp5_ASAP7_75t_L g1447 ( 
.A(n_1334),
.B(n_1296),
.Y(n_1447)
);

AOI22xp5_ASAP7_75t_L g1448 ( 
.A1(n_1339),
.A2(n_1267),
.B1(n_1292),
.B2(n_1258),
.Y(n_1448)
);

HB1xp67_ASAP7_75t_L g1449 ( 
.A(n_1324),
.Y(n_1449)
);

NAND2xp5_ASAP7_75t_L g1450 ( 
.A(n_1367),
.B(n_1369),
.Y(n_1450)
);

NAND2xp5_ASAP7_75t_L g1451 ( 
.A(n_1384),
.B(n_1292),
.Y(n_1451)
);

NAND2x1_ASAP7_75t_L g1452 ( 
.A(n_1402),
.B(n_1228),
.Y(n_1452)
);

INVx2_ASAP7_75t_L g1453 ( 
.A(n_1338),
.Y(n_1453)
);

INVx2_ASAP7_75t_L g1454 ( 
.A(n_1359),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1318),
.Y(n_1455)
);

NAND2xp5_ASAP7_75t_L g1456 ( 
.A(n_1329),
.B(n_1293),
.Y(n_1456)
);

NAND2xp5_ASAP7_75t_L g1457 ( 
.A(n_1342),
.B(n_1228),
.Y(n_1457)
);

OAI21xp5_ASAP7_75t_L g1458 ( 
.A1(n_1375),
.A2(n_1373),
.B(n_1372),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_L g1459 ( 
.A(n_1344),
.B(n_1228),
.Y(n_1459)
);

AOI21x1_ASAP7_75t_L g1460 ( 
.A1(n_1306),
.A2(n_1295),
.B(n_1121),
.Y(n_1460)
);

AOI22xp33_ASAP7_75t_L g1461 ( 
.A1(n_1351),
.A2(n_1267),
.B1(n_1121),
.B2(n_998),
.Y(n_1461)
);

NAND2xp5_ASAP7_75t_SL g1462 ( 
.A(n_1361),
.B(n_1043),
.Y(n_1462)
);

A2O1A1Ixp33_ASAP7_75t_L g1463 ( 
.A1(n_1350),
.A2(n_619),
.B(n_699),
.C(n_608),
.Y(n_1463)
);

AOI21x1_ASAP7_75t_L g1464 ( 
.A1(n_1365),
.A2(n_1149),
.B(n_1128),
.Y(n_1464)
);

BUFx2_ASAP7_75t_L g1465 ( 
.A(n_1371),
.Y(n_1465)
);

INVx3_ASAP7_75t_L g1466 ( 
.A(n_1355),
.Y(n_1466)
);

INVx2_ASAP7_75t_L g1467 ( 
.A(n_1359),
.Y(n_1467)
);

NAND2x1p5_ASAP7_75t_L g1468 ( 
.A(n_1345),
.B(n_1149),
.Y(n_1468)
);

AND2x2_ASAP7_75t_L g1469 ( 
.A(n_1316),
.B(n_1299),
.Y(n_1469)
);

AOI21xp5_ASAP7_75t_L g1470 ( 
.A1(n_1322),
.A2(n_1155),
.B(n_1114),
.Y(n_1470)
);

OAI21xp5_ASAP7_75t_L g1471 ( 
.A1(n_1327),
.A2(n_1228),
.B(n_1153),
.Y(n_1471)
);

O2A1O1Ixp5_ASAP7_75t_L g1472 ( 
.A1(n_1365),
.A2(n_1152),
.B(n_1162),
.C(n_1143),
.Y(n_1472)
);

NAND2xp5_ASAP7_75t_L g1473 ( 
.A(n_1308),
.B(n_1299),
.Y(n_1473)
);

NAND2x1p5_ASAP7_75t_L g1474 ( 
.A(n_1362),
.B(n_1149),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_L g1475 ( 
.A(n_1309),
.B(n_1037),
.Y(n_1475)
);

A2O1A1Ixp33_ASAP7_75t_L g1476 ( 
.A1(n_1312),
.A2(n_619),
.B(n_699),
.C(n_608),
.Y(n_1476)
);

INVx3_ASAP7_75t_L g1477 ( 
.A(n_1355),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1363),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1374),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1378),
.Y(n_1480)
);

AOI21xp5_ASAP7_75t_L g1481 ( 
.A1(n_1327),
.A2(n_1155),
.B(n_1114),
.Y(n_1481)
);

OR2x2_ASAP7_75t_SL g1482 ( 
.A(n_1368),
.B(n_982),
.Y(n_1482)
);

AOI21xp5_ASAP7_75t_L g1483 ( 
.A1(n_1330),
.A2(n_1159),
.B(n_1155),
.Y(n_1483)
);

AND2x2_ASAP7_75t_L g1484 ( 
.A(n_1323),
.B(n_1389),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_SL g1485 ( 
.A(n_1346),
.B(n_1043),
.Y(n_1485)
);

O2A1O1Ixp33_ASAP7_75t_L g1486 ( 
.A1(n_1313),
.A2(n_798),
.B(n_820),
.C(n_714),
.Y(n_1486)
);

AOI21xp5_ASAP7_75t_L g1487 ( 
.A1(n_1330),
.A2(n_1159),
.B(n_1155),
.Y(n_1487)
);

AOI22xp5_ASAP7_75t_L g1488 ( 
.A1(n_1352),
.A2(n_668),
.B1(n_703),
.B2(n_598),
.Y(n_1488)
);

NOR2x1p5_ASAP7_75t_L g1489 ( 
.A(n_1397),
.B(n_1060),
.Y(n_1489)
);

NOR2xp33_ASAP7_75t_L g1490 ( 
.A(n_1331),
.B(n_1150),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_L g1491 ( 
.A(n_1340),
.B(n_1061),
.Y(n_1491)
);

OAI21xp5_ASAP7_75t_L g1492 ( 
.A1(n_1332),
.A2(n_1153),
.B(n_1151),
.Y(n_1492)
);

NOR2xp33_ASAP7_75t_L g1493 ( 
.A(n_1343),
.B(n_1154),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1379),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_1314),
.B(n_1064),
.Y(n_1495)
);

AOI21xp5_ASAP7_75t_L g1496 ( 
.A1(n_1332),
.A2(n_1159),
.B(n_1153),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1328),
.B(n_600),
.Y(n_1497)
);

AOI21xp5_ASAP7_75t_L g1498 ( 
.A1(n_1333),
.A2(n_1159),
.B(n_1140),
.Y(n_1498)
);

O2A1O1Ixp33_ASAP7_75t_L g1499 ( 
.A1(n_1320),
.A2(n_1325),
.B(n_798),
.C(n_820),
.Y(n_1499)
);

NAND2xp5_ASAP7_75t_L g1500 ( 
.A(n_1337),
.B(n_1067),
.Y(n_1500)
);

NOR2xp33_ASAP7_75t_L g1501 ( 
.A(n_1406),
.B(n_706),
.Y(n_1501)
);

O2A1O1Ixp33_ASAP7_75t_L g1502 ( 
.A1(n_1422),
.A2(n_714),
.B(n_1014),
.C(n_998),
.Y(n_1502)
);

CKINVDCx5p33_ASAP7_75t_R g1503 ( 
.A(n_1413),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1428),
.Y(n_1504)
);

OAI22x1_ASAP7_75t_L g1505 ( 
.A1(n_1406),
.A2(n_1484),
.B1(n_1448),
.B2(n_1488),
.Y(n_1505)
);

NOR2xp33_ASAP7_75t_L g1506 ( 
.A(n_1424),
.B(n_1414),
.Y(n_1506)
);

NAND2xp5_ASAP7_75t_L g1507 ( 
.A(n_1408),
.B(n_1414),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_L g1508 ( 
.A(n_1403),
.B(n_1357),
.Y(n_1508)
);

AOI21xp5_ASAP7_75t_L g1509 ( 
.A1(n_1405),
.A2(n_1411),
.B(n_1409),
.Y(n_1509)
);

INVx3_ASAP7_75t_SL g1510 ( 
.A(n_1418),
.Y(n_1510)
);

NOR2xp33_ASAP7_75t_SL g1511 ( 
.A(n_1403),
.B(n_1317),
.Y(n_1511)
);

AOI21xp5_ASAP7_75t_L g1512 ( 
.A1(n_1435),
.A2(n_1333),
.B(n_1370),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1436),
.Y(n_1513)
);

AOI21x1_ASAP7_75t_L g1514 ( 
.A1(n_1434),
.A2(n_1386),
.B(n_1370),
.Y(n_1514)
);

OAI22xp5_ASAP7_75t_L g1515 ( 
.A1(n_1450),
.A2(n_1356),
.B1(n_1353),
.B2(n_1321),
.Y(n_1515)
);

INVx5_ASAP7_75t_L g1516 ( 
.A(n_1437),
.Y(n_1516)
);

HB1xp67_ASAP7_75t_L g1517 ( 
.A(n_1425),
.Y(n_1517)
);

NAND2xp5_ASAP7_75t_SL g1518 ( 
.A(n_1440),
.B(n_1417),
.Y(n_1518)
);

AND2x4_ASAP7_75t_L g1519 ( 
.A(n_1431),
.B(n_1442),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_L g1520 ( 
.A(n_1473),
.B(n_1393),
.Y(n_1520)
);

AOI21xp5_ASAP7_75t_L g1521 ( 
.A1(n_1407),
.A2(n_1387),
.B(n_1386),
.Y(n_1521)
);

AOI21xp5_ASAP7_75t_L g1522 ( 
.A1(n_1404),
.A2(n_1395),
.B(n_1387),
.Y(n_1522)
);

NAND3xp33_ASAP7_75t_SL g1523 ( 
.A(n_1499),
.B(n_743),
.C(n_708),
.Y(n_1523)
);

O2A1O1Ixp5_ASAP7_75t_L g1524 ( 
.A1(n_1463),
.A2(n_1395),
.B(n_1391),
.C(n_1383),
.Y(n_1524)
);

AOI22x1_ASAP7_75t_L g1525 ( 
.A1(n_1458),
.A2(n_1396),
.B1(n_1400),
.B2(n_1014),
.Y(n_1525)
);

INVx3_ASAP7_75t_L g1526 ( 
.A(n_1437),
.Y(n_1526)
);

A2O1A1Ixp33_ASAP7_75t_SL g1527 ( 
.A1(n_1486),
.A2(n_1140),
.B(n_1141),
.C(n_1133),
.Y(n_1527)
);

NOR2xp33_ASAP7_75t_L g1528 ( 
.A(n_1446),
.B(n_794),
.Y(n_1528)
);

AOI21xp5_ASAP7_75t_L g1529 ( 
.A1(n_1404),
.A2(n_1391),
.B(n_1383),
.Y(n_1529)
);

OAI22xp5_ASAP7_75t_L g1530 ( 
.A1(n_1440),
.A2(n_591),
.B1(n_593),
.B2(n_592),
.Y(n_1530)
);

CKINVDCx14_ASAP7_75t_R g1531 ( 
.A(n_1465),
.Y(n_1531)
);

AND2x4_ASAP7_75t_SL g1532 ( 
.A(n_1449),
.B(n_1380),
.Y(n_1532)
);

AOI22xp33_ASAP7_75t_L g1533 ( 
.A1(n_1461),
.A2(n_626),
.B1(n_678),
.B2(n_600),
.Y(n_1533)
);

NOR2xp33_ASAP7_75t_L g1534 ( 
.A(n_1431),
.B(n_797),
.Y(n_1534)
);

BUFx3_ASAP7_75t_L g1535 ( 
.A(n_1442),
.Y(n_1535)
);

CKINVDCx8_ASAP7_75t_R g1536 ( 
.A(n_1412),
.Y(n_1536)
);

A2O1A1Ixp33_ASAP7_75t_L g1537 ( 
.A1(n_1490),
.A2(n_1381),
.B(n_1380),
.C(n_1388),
.Y(n_1537)
);

O2A1O1Ixp33_ASAP7_75t_L g1538 ( 
.A1(n_1476),
.A2(n_1463),
.B(n_1451),
.C(n_1455),
.Y(n_1538)
);

AOI21xp5_ASAP7_75t_L g1539 ( 
.A1(n_1410),
.A2(n_1388),
.B(n_1381),
.Y(n_1539)
);

AND2x2_ASAP7_75t_SL g1540 ( 
.A(n_1461),
.B(n_594),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1445),
.Y(n_1541)
);

OR2x6_ASAP7_75t_L g1542 ( 
.A(n_1489),
.B(n_1149),
.Y(n_1542)
);

AOI21xp5_ASAP7_75t_L g1543 ( 
.A1(n_1410),
.A2(n_1443),
.B(n_1438),
.Y(n_1543)
);

INVx4_ASAP7_75t_L g1544 ( 
.A(n_1437),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1478),
.Y(n_1545)
);

INVx3_ASAP7_75t_SL g1546 ( 
.A(n_1497),
.Y(n_1546)
);

NOR2xp33_ASAP7_75t_R g1547 ( 
.A(n_1429),
.B(n_600),
.Y(n_1547)
);

AOI21xp5_ASAP7_75t_L g1548 ( 
.A1(n_1444),
.A2(n_1150),
.B(n_1141),
.Y(n_1548)
);

AOI21xp5_ASAP7_75t_L g1549 ( 
.A1(n_1416),
.A2(n_1156),
.B(n_1154),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1479),
.Y(n_1550)
);

OAI22xp5_ASAP7_75t_L g1551 ( 
.A1(n_1415),
.A2(n_596),
.B1(n_599),
.B2(n_597),
.Y(n_1551)
);

O2A1O1Ixp5_ASAP7_75t_L g1552 ( 
.A1(n_1485),
.A2(n_604),
.B(n_616),
.C(n_590),
.Y(n_1552)
);

AOI21xp5_ASAP7_75t_L g1553 ( 
.A1(n_1471),
.A2(n_1156),
.B(n_1149),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1447),
.B(n_816),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_L g1555 ( 
.A(n_1449),
.B(n_883),
.Y(n_1555)
);

INVx2_ASAP7_75t_L g1556 ( 
.A(n_1420),
.Y(n_1556)
);

OAI22xp5_ASAP7_75t_L g1557 ( 
.A1(n_1457),
.A2(n_601),
.B1(n_605),
.B2(n_602),
.Y(n_1557)
);

AOI21xp5_ASAP7_75t_L g1558 ( 
.A1(n_1496),
.A2(n_1152),
.B(n_1143),
.Y(n_1558)
);

BUFx12f_ASAP7_75t_L g1559 ( 
.A(n_1482),
.Y(n_1559)
);

INVx2_ASAP7_75t_L g1560 ( 
.A(n_1421),
.Y(n_1560)
);

NAND2xp5_ASAP7_75t_SL g1561 ( 
.A(n_1437),
.B(n_1043),
.Y(n_1561)
);

OA22x2_ASAP7_75t_L g1562 ( 
.A1(n_1469),
.A2(n_1430),
.B1(n_1456),
.B2(n_1480),
.Y(n_1562)
);

AOI22xp33_ASAP7_75t_L g1563 ( 
.A1(n_1490),
.A2(n_626),
.B1(n_678),
.B2(n_600),
.Y(n_1563)
);

OAI22xp5_ASAP7_75t_L g1564 ( 
.A1(n_1459),
.A2(n_612),
.B1(n_614),
.B2(n_607),
.Y(n_1564)
);

BUFx6f_ASAP7_75t_L g1565 ( 
.A(n_1439),
.Y(n_1565)
);

NOR2xp33_ASAP7_75t_L g1566 ( 
.A(n_1494),
.B(n_1476),
.Y(n_1566)
);

OAI21xp5_ASAP7_75t_L g1567 ( 
.A1(n_1472),
.A2(n_1162),
.B(n_1152),
.Y(n_1567)
);

AOI21xp5_ASAP7_75t_L g1568 ( 
.A1(n_1419),
.A2(n_1162),
.B(n_1152),
.Y(n_1568)
);

AND2x2_ASAP7_75t_L g1569 ( 
.A(n_1475),
.B(n_626),
.Y(n_1569)
);

BUFx3_ASAP7_75t_L g1570 ( 
.A(n_1439),
.Y(n_1570)
);

NAND2xp5_ASAP7_75t_L g1571 ( 
.A(n_1500),
.B(n_971),
.Y(n_1571)
);

OAI22xp5_ASAP7_75t_L g1572 ( 
.A1(n_1493),
.A2(n_618),
.B1(n_623),
.B2(n_611),
.Y(n_1572)
);

OR2x2_ASAP7_75t_L g1573 ( 
.A(n_1426),
.B(n_1068),
.Y(n_1573)
);

OAI22xp5_ASAP7_75t_L g1574 ( 
.A1(n_1493),
.A2(n_627),
.B1(n_633),
.B2(n_625),
.Y(n_1574)
);

AOI21x1_ASAP7_75t_L g1575 ( 
.A1(n_1460),
.A2(n_1035),
.B(n_1034),
.Y(n_1575)
);

AOI21xp5_ASAP7_75t_L g1576 ( 
.A1(n_1492),
.A2(n_1163),
.B(n_1162),
.Y(n_1576)
);

OAI22xp5_ASAP7_75t_L g1577 ( 
.A1(n_1495),
.A2(n_636),
.B1(n_637),
.B2(n_635),
.Y(n_1577)
);

BUFx6f_ASAP7_75t_L g1578 ( 
.A(n_1439),
.Y(n_1578)
);

A2O1A1Ixp33_ASAP7_75t_L g1579 ( 
.A1(n_1433),
.A2(n_595),
.B(n_617),
.C(n_615),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_L g1580 ( 
.A(n_1453),
.B(n_1028),
.Y(n_1580)
);

INVx2_ASAP7_75t_L g1581 ( 
.A(n_1454),
.Y(n_1581)
);

INVx5_ASAP7_75t_L g1582 ( 
.A(n_1439),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_L g1583 ( 
.A(n_1467),
.B(n_1071),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1467),
.B(n_1082),
.Y(n_1584)
);

AO32x1_ASAP7_75t_L g1585 ( 
.A1(n_1472),
.A2(n_604),
.A3(n_621),
.B1(n_616),
.B2(n_590),
.Y(n_1585)
);

INVx2_ASAP7_75t_L g1586 ( 
.A(n_1468),
.Y(n_1586)
);

AND2x6_ASAP7_75t_L g1587 ( 
.A(n_1441),
.B(n_856),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1491),
.Y(n_1588)
);

HB1xp67_ASAP7_75t_L g1589 ( 
.A(n_1441),
.Y(n_1589)
);

AOI22x1_ASAP7_75t_L g1590 ( 
.A1(n_1427),
.A2(n_624),
.B1(n_628),
.B2(n_621),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1468),
.Y(n_1591)
);

A2O1A1Ixp33_ASAP7_75t_L g1592 ( 
.A1(n_1423),
.A2(n_615),
.B(n_617),
.C(n_595),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_L g1593 ( 
.A(n_1441),
.B(n_1086),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_L g1594 ( 
.A(n_1441),
.B(n_1090),
.Y(n_1594)
);

A2O1A1Ixp33_ASAP7_75t_L g1595 ( 
.A1(n_1423),
.A2(n_617),
.B(n_719),
.C(n_629),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_L g1596 ( 
.A(n_1466),
.B(n_645),
.Y(n_1596)
);

AOI21xp5_ASAP7_75t_L g1597 ( 
.A1(n_1485),
.A2(n_1163),
.B(n_1148),
.Y(n_1597)
);

AOI21xp5_ASAP7_75t_L g1598 ( 
.A1(n_1432),
.A2(n_1163),
.B(n_1148),
.Y(n_1598)
);

O2A1O1Ixp5_ASAP7_75t_L g1599 ( 
.A1(n_1452),
.A2(n_1462),
.B(n_1498),
.C(n_1464),
.Y(n_1599)
);

NOR2xp33_ASAP7_75t_L g1600 ( 
.A(n_1466),
.B(n_646),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_L g1601 ( 
.A(n_1477),
.B(n_648),
.Y(n_1601)
);

AOI22xp5_ASAP7_75t_L g1602 ( 
.A1(n_1477),
.A2(n_672),
.B1(n_684),
.B2(n_661),
.Y(n_1602)
);

AOI21xp5_ASAP7_75t_L g1603 ( 
.A1(n_1553),
.A2(n_1462),
.B(n_1474),
.Y(n_1603)
);

NAND3xp33_ASAP7_75t_L g1604 ( 
.A(n_1501),
.B(n_1502),
.C(n_1566),
.Y(n_1604)
);

HB1xp67_ASAP7_75t_L g1605 ( 
.A(n_1586),
.Y(n_1605)
);

AOI21xp33_ASAP7_75t_L g1606 ( 
.A1(n_1505),
.A2(n_1474),
.B(n_628),
.Y(n_1606)
);

AOI21x1_ASAP7_75t_L g1607 ( 
.A1(n_1575),
.A2(n_1483),
.B(n_1481),
.Y(n_1607)
);

OAI21x1_ASAP7_75t_L g1608 ( 
.A1(n_1509),
.A2(n_1487),
.B(n_1470),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1506),
.B(n_1043),
.Y(n_1609)
);

OAI21xp5_ASAP7_75t_L g1610 ( 
.A1(n_1518),
.A2(n_631),
.B(n_624),
.Y(n_1610)
);

INVx6_ASAP7_75t_SL g1611 ( 
.A(n_1519),
.Y(n_1611)
);

BUFx2_ASAP7_75t_L g1612 ( 
.A(n_1519),
.Y(n_1612)
);

AND2x2_ASAP7_75t_L g1613 ( 
.A(n_1528),
.B(n_626),
.Y(n_1613)
);

AOI21xp5_ASAP7_75t_L g1614 ( 
.A1(n_1512),
.A2(n_856),
.B(n_1163),
.Y(n_1614)
);

O2A1O1Ixp5_ASAP7_75t_L g1615 ( 
.A1(n_1543),
.A2(n_719),
.B(n_736),
.C(n_629),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_L g1616 ( 
.A(n_1507),
.B(n_631),
.Y(n_1616)
);

A2O1A1Ixp33_ASAP7_75t_L g1617 ( 
.A1(n_1538),
.A2(n_629),
.B(n_736),
.C(n_719),
.Y(n_1617)
);

NOR2xp33_ASAP7_75t_SL g1618 ( 
.A(n_1536),
.B(n_678),
.Y(n_1618)
);

OAI21x1_ASAP7_75t_L g1619 ( 
.A1(n_1599),
.A2(n_1124),
.B(n_1118),
.Y(n_1619)
);

BUFx2_ASAP7_75t_L g1620 ( 
.A(n_1535),
.Y(n_1620)
);

AOI21xp5_ASAP7_75t_L g1621 ( 
.A1(n_1515),
.A2(n_1148),
.B(n_1146),
.Y(n_1621)
);

AOI221x1_ASAP7_75t_L g1622 ( 
.A1(n_1529),
.A2(n_1523),
.B1(n_1551),
.B2(n_1595),
.C(n_1592),
.Y(n_1622)
);

AOI221xp5_ASAP7_75t_SL g1623 ( 
.A1(n_1572),
.A2(n_638),
.B1(n_639),
.B2(n_634),
.C(n_632),
.Y(n_1623)
);

HB1xp67_ASAP7_75t_L g1624 ( 
.A(n_1591),
.Y(n_1624)
);

AO31x2_ASAP7_75t_L g1625 ( 
.A1(n_1537),
.A2(n_1118),
.A3(n_1125),
.B(n_1124),
.Y(n_1625)
);

OAI22xp5_ASAP7_75t_L g1626 ( 
.A1(n_1602),
.A2(n_632),
.B1(n_638),
.B2(n_634),
.Y(n_1626)
);

AOI21xp5_ASAP7_75t_L g1627 ( 
.A1(n_1576),
.A2(n_1161),
.B(n_1146),
.Y(n_1627)
);

OR2x2_ASAP7_75t_L g1628 ( 
.A(n_1545),
.B(n_639),
.Y(n_1628)
);

AOI21xp5_ASAP7_75t_L g1629 ( 
.A1(n_1548),
.A2(n_1161),
.B(n_1146),
.Y(n_1629)
);

OAI21x1_ASAP7_75t_L g1630 ( 
.A1(n_1558),
.A2(n_1124),
.B(n_1118),
.Y(n_1630)
);

AOI21xp5_ASAP7_75t_L g1631 ( 
.A1(n_1521),
.A2(n_1161),
.B(n_800),
.Y(n_1631)
);

INVx2_ASAP7_75t_SL g1632 ( 
.A(n_1517),
.Y(n_1632)
);

OAI21xp5_ASAP7_75t_L g1633 ( 
.A1(n_1574),
.A2(n_650),
.B(n_649),
.Y(n_1633)
);

AND2x4_ASAP7_75t_L g1634 ( 
.A(n_1516),
.B(n_800),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_L g1635 ( 
.A(n_1554),
.B(n_649),
.Y(n_1635)
);

INVx3_ASAP7_75t_L g1636 ( 
.A(n_1516),
.Y(n_1636)
);

OAI21x1_ASAP7_75t_SL g1637 ( 
.A1(n_1522),
.A2(n_765),
.B(n_736),
.Y(n_1637)
);

OAI21x1_ASAP7_75t_L g1638 ( 
.A1(n_1539),
.A2(n_1124),
.B(n_1118),
.Y(n_1638)
);

NOR4xp25_ASAP7_75t_L g1639 ( 
.A(n_1563),
.B(n_651),
.C(n_654),
.D(n_650),
.Y(n_1639)
);

OAI21x1_ASAP7_75t_L g1640 ( 
.A1(n_1598),
.A2(n_1125),
.B(n_1083),
.Y(n_1640)
);

AOI21xp5_ASAP7_75t_L g1641 ( 
.A1(n_1549),
.A2(n_1567),
.B(n_1568),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1504),
.Y(n_1642)
);

AOI21x1_ASAP7_75t_L g1643 ( 
.A1(n_1514),
.A2(n_1597),
.B(n_1561),
.Y(n_1643)
);

AOI221x1_ASAP7_75t_L g1644 ( 
.A1(n_1579),
.A2(n_656),
.B1(n_660),
.B2(n_654),
.C(n_651),
.Y(n_1644)
);

AOI21xp5_ASAP7_75t_L g1645 ( 
.A1(n_1520),
.A2(n_786),
.B(n_765),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_L g1646 ( 
.A(n_1555),
.B(n_656),
.Y(n_1646)
);

A2O1A1Ixp33_ASAP7_75t_L g1647 ( 
.A1(n_1524),
.A2(n_786),
.B(n_808),
.C(n_765),
.Y(n_1647)
);

AOI21x1_ASAP7_75t_SL g1648 ( 
.A1(n_1596),
.A2(n_0),
.B(n_1),
.Y(n_1648)
);

AOI21xp5_ASAP7_75t_L g1649 ( 
.A1(n_1511),
.A2(n_808),
.B(n_786),
.Y(n_1649)
);

OAI21x1_ASAP7_75t_L g1650 ( 
.A1(n_1525),
.A2(n_1125),
.B(n_665),
.Y(n_1650)
);

AND2x2_ASAP7_75t_L g1651 ( 
.A(n_1534),
.B(n_678),
.Y(n_1651)
);

OAI21x1_ASAP7_75t_L g1652 ( 
.A1(n_1590),
.A2(n_1125),
.B(n_665),
.Y(n_1652)
);

NOR2xp33_ASAP7_75t_L g1653 ( 
.A(n_1511),
.B(n_729),
.Y(n_1653)
);

AOI221xp5_ASAP7_75t_SL g1654 ( 
.A1(n_1530),
.A2(n_670),
.B1(n_671),
.B2(n_669),
.C(n_660),
.Y(n_1654)
);

AOI21xp5_ASAP7_75t_L g1655 ( 
.A1(n_1527),
.A2(n_811),
.B(n_808),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1513),
.Y(n_1656)
);

OA21x2_ASAP7_75t_L g1657 ( 
.A1(n_1552),
.A2(n_1508),
.B(n_1550),
.Y(n_1657)
);

INVxp67_ASAP7_75t_SL g1658 ( 
.A(n_1593),
.Y(n_1658)
);

BUFx4f_ASAP7_75t_L g1659 ( 
.A(n_1510),
.Y(n_1659)
);

NOR2xp33_ASAP7_75t_SL g1660 ( 
.A(n_1503),
.B(n_729),
.Y(n_1660)
);

AOI22xp33_ASAP7_75t_L g1661 ( 
.A1(n_1540),
.A2(n_840),
.B1(n_868),
.B2(n_729),
.Y(n_1661)
);

OAI21x1_ASAP7_75t_L g1662 ( 
.A1(n_1526),
.A2(n_670),
.B(n_669),
.Y(n_1662)
);

OAI21x1_ASAP7_75t_L g1663 ( 
.A1(n_1526),
.A2(n_683),
.B(n_671),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1541),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_SL g1665 ( 
.A(n_1516),
.B(n_729),
.Y(n_1665)
);

OAI22xp5_ASAP7_75t_L g1666 ( 
.A1(n_1602),
.A2(n_686),
.B1(n_694),
.B2(n_683),
.Y(n_1666)
);

AND2x4_ASAP7_75t_L g1667 ( 
.A(n_1582),
.B(n_562),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_L g1668 ( 
.A(n_1588),
.B(n_686),
.Y(n_1668)
);

NAND2xp5_ASAP7_75t_L g1669 ( 
.A(n_1571),
.B(n_694),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_SL g1670 ( 
.A(n_1582),
.B(n_840),
.Y(n_1670)
);

BUFx2_ASAP7_75t_L g1671 ( 
.A(n_1570),
.Y(n_1671)
);

AND2x2_ASAP7_75t_L g1672 ( 
.A(n_1569),
.B(n_840),
.Y(n_1672)
);

NOR4xp25_ASAP7_75t_L g1673 ( 
.A(n_1533),
.B(n_704),
.C(n_705),
.D(n_696),
.Y(n_1673)
);

OAI21x1_ASAP7_75t_L g1674 ( 
.A1(n_1594),
.A2(n_704),
.B(n_696),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_L g1675 ( 
.A(n_1532),
.B(n_705),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_L g1676 ( 
.A(n_1547),
.B(n_713),
.Y(n_1676)
);

A2O1A1Ixp33_ASAP7_75t_L g1677 ( 
.A1(n_1600),
.A2(n_813),
.B(n_827),
.C(n_811),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1556),
.Y(n_1678)
);

INVx1_ASAP7_75t_SL g1679 ( 
.A(n_1546),
.Y(n_1679)
);

INVxp67_ASAP7_75t_L g1680 ( 
.A(n_1589),
.Y(n_1680)
);

O2A1O1Ixp33_ASAP7_75t_L g1681 ( 
.A1(n_1577),
.A2(n_721),
.B(n_726),
.C(n_713),
.Y(n_1681)
);

AOI21xp5_ASAP7_75t_L g1682 ( 
.A1(n_1582),
.A2(n_813),
.B(n_811),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1560),
.Y(n_1683)
);

INVx2_ASAP7_75t_L g1684 ( 
.A(n_1581),
.Y(n_1684)
);

INVx2_ASAP7_75t_L g1685 ( 
.A(n_1562),
.Y(n_1685)
);

OAI22xp5_ASAP7_75t_L g1686 ( 
.A1(n_1604),
.A2(n_1531),
.B1(n_1542),
.B2(n_1601),
.Y(n_1686)
);

OAI21x1_ASAP7_75t_L g1687 ( 
.A1(n_1608),
.A2(n_1584),
.B(n_1583),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_L g1688 ( 
.A(n_1632),
.B(n_1565),
.Y(n_1688)
);

OR2x2_ASAP7_75t_L g1689 ( 
.A(n_1624),
.B(n_1658),
.Y(n_1689)
);

AND2x4_ASAP7_75t_SL g1690 ( 
.A(n_1636),
.B(n_1565),
.Y(n_1690)
);

OAI21x1_ASAP7_75t_L g1691 ( 
.A1(n_1607),
.A2(n_1564),
.B(n_1557),
.Y(n_1691)
);

BUFx8_ASAP7_75t_SL g1692 ( 
.A(n_1659),
.Y(n_1692)
);

OAI21x1_ASAP7_75t_L g1693 ( 
.A1(n_1641),
.A2(n_1573),
.B(n_1580),
.Y(n_1693)
);

CKINVDCx5p33_ASAP7_75t_R g1694 ( 
.A(n_1659),
.Y(n_1694)
);

AOI22xp33_ASAP7_75t_L g1695 ( 
.A1(n_1685),
.A2(n_1542),
.B1(n_1559),
.B2(n_1587),
.Y(n_1695)
);

OAI21x1_ASAP7_75t_L g1696 ( 
.A1(n_1643),
.A2(n_1585),
.B(n_1587),
.Y(n_1696)
);

AND2x2_ASAP7_75t_L g1697 ( 
.A(n_1642),
.B(n_1565),
.Y(n_1697)
);

OAI21x1_ASAP7_75t_SL g1698 ( 
.A1(n_1637),
.A2(n_1603),
.B(n_1610),
.Y(n_1698)
);

AND2x2_ASAP7_75t_L g1699 ( 
.A(n_1656),
.B(n_1578),
.Y(n_1699)
);

OAI21x1_ASAP7_75t_L g1700 ( 
.A1(n_1615),
.A2(n_1585),
.B(n_1587),
.Y(n_1700)
);

AND2x4_ASAP7_75t_L g1701 ( 
.A(n_1624),
.B(n_1578),
.Y(n_1701)
);

INVx1_ASAP7_75t_SL g1702 ( 
.A(n_1612),
.Y(n_1702)
);

OAI21x1_ASAP7_75t_L g1703 ( 
.A1(n_1615),
.A2(n_1585),
.B(n_1587),
.Y(n_1703)
);

OA21x2_ASAP7_75t_L g1704 ( 
.A1(n_1617),
.A2(n_827),
.B(n_813),
.Y(n_1704)
);

OAI21xp5_ASAP7_75t_L g1705 ( 
.A1(n_1617),
.A2(n_726),
.B(n_721),
.Y(n_1705)
);

HB1xp67_ASAP7_75t_L g1706 ( 
.A(n_1680),
.Y(n_1706)
);

OAI21x1_ASAP7_75t_L g1707 ( 
.A1(n_1631),
.A2(n_740),
.B(n_738),
.Y(n_1707)
);

INVx3_ASAP7_75t_L g1708 ( 
.A(n_1625),
.Y(n_1708)
);

NAND2x1p5_ASAP7_75t_L g1709 ( 
.A(n_1657),
.B(n_1544),
.Y(n_1709)
);

INVx2_ASAP7_75t_L g1710 ( 
.A(n_1684),
.Y(n_1710)
);

AOI222xp33_ASAP7_75t_SL g1711 ( 
.A1(n_1626),
.A2(n_747),
.B1(n_740),
.B2(n_748),
.C1(n_746),
.C2(n_738),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1664),
.Y(n_1712)
);

NOR2xp33_ASAP7_75t_L g1713 ( 
.A(n_1660),
.B(n_1620),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1605),
.Y(n_1714)
);

OAI21x1_ASAP7_75t_L g1715 ( 
.A1(n_1619),
.A2(n_747),
.B(n_746),
.Y(n_1715)
);

NAND2x1p5_ASAP7_75t_L g1716 ( 
.A(n_1657),
.B(n_1544),
.Y(n_1716)
);

OAI21x1_ASAP7_75t_L g1717 ( 
.A1(n_1614),
.A2(n_749),
.B(n_748),
.Y(n_1717)
);

OAI21x1_ASAP7_75t_L g1718 ( 
.A1(n_1627),
.A2(n_756),
.B(n_749),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1605),
.Y(n_1719)
);

AOI21xp33_ASAP7_75t_L g1720 ( 
.A1(n_1653),
.A2(n_1542),
.B(n_1578),
.Y(n_1720)
);

AOI21xp5_ASAP7_75t_L g1721 ( 
.A1(n_1621),
.A2(n_896),
.B(n_827),
.Y(n_1721)
);

OA21x2_ASAP7_75t_L g1722 ( 
.A1(n_1647),
.A2(n_914),
.B(n_896),
.Y(n_1722)
);

A2O1A1Ixp33_ASAP7_75t_L g1723 ( 
.A1(n_1653),
.A2(n_897),
.B(n_958),
.C(n_943),
.Y(n_1723)
);

BUFx12f_ASAP7_75t_L g1724 ( 
.A(n_1671),
.Y(n_1724)
);

INVx3_ASAP7_75t_L g1725 ( 
.A(n_1625),
.Y(n_1725)
);

OAI21x1_ASAP7_75t_L g1726 ( 
.A1(n_1638),
.A2(n_759),
.B(n_756),
.Y(n_1726)
);

INVx2_ASAP7_75t_L g1727 ( 
.A(n_1684),
.Y(n_1727)
);

INVx2_ASAP7_75t_L g1728 ( 
.A(n_1678),
.Y(n_1728)
);

HB1xp67_ASAP7_75t_L g1729 ( 
.A(n_1680),
.Y(n_1729)
);

AO21x2_ASAP7_75t_L g1730 ( 
.A1(n_1606),
.A2(n_762),
.B(n_759),
.Y(n_1730)
);

NAND2x1p5_ASAP7_75t_L g1731 ( 
.A(n_1657),
.B(n_896),
.Y(n_1731)
);

OAI22xp5_ASAP7_75t_L g1732 ( 
.A1(n_1661),
.A2(n_764),
.B1(n_768),
.B2(n_762),
.Y(n_1732)
);

AO32x2_ASAP7_75t_L g1733 ( 
.A1(n_1666),
.A2(n_1008),
.A3(n_868),
.B1(n_840),
.B2(n_769),
.Y(n_1733)
);

INVx2_ASAP7_75t_L g1734 ( 
.A(n_1683),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1625),
.Y(n_1735)
);

OAI22xp5_ASAP7_75t_SL g1736 ( 
.A1(n_1661),
.A2(n_768),
.B1(n_769),
.B2(n_764),
.Y(n_1736)
);

OA21x2_ASAP7_75t_L g1737 ( 
.A1(n_1647),
.A2(n_956),
.B(n_914),
.Y(n_1737)
);

AOI21xp5_ASAP7_75t_L g1738 ( 
.A1(n_1609),
.A2(n_956),
.B(n_914),
.Y(n_1738)
);

HB1xp67_ASAP7_75t_L g1739 ( 
.A(n_1658),
.Y(n_1739)
);

INVx2_ASAP7_75t_L g1740 ( 
.A(n_1685),
.Y(n_1740)
);

CKINVDCx5p33_ASAP7_75t_R g1741 ( 
.A(n_1611),
.Y(n_1741)
);

AOI22xp33_ASAP7_75t_L g1742 ( 
.A1(n_1613),
.A2(n_868),
.B1(n_1008),
.B2(n_897),
.Y(n_1742)
);

OR2x2_ASAP7_75t_L g1743 ( 
.A(n_1628),
.B(n_864),
.Y(n_1743)
);

OAI21x1_ASAP7_75t_L g1744 ( 
.A1(n_1650),
.A2(n_775),
.B(n_771),
.Y(n_1744)
);

OAI221xp5_ASAP7_75t_L g1745 ( 
.A1(n_1639),
.A2(n_776),
.B1(n_778),
.B2(n_775),
.C(n_771),
.Y(n_1745)
);

AND2x4_ASAP7_75t_L g1746 ( 
.A(n_1701),
.B(n_1634),
.Y(n_1746)
);

OA21x2_ASAP7_75t_L g1747 ( 
.A1(n_1696),
.A2(n_1655),
.B(n_1677),
.Y(n_1747)
);

INVx6_ASAP7_75t_L g1748 ( 
.A(n_1724),
.Y(n_1748)
);

OAI21x1_ASAP7_75t_L g1749 ( 
.A1(n_1731),
.A2(n_1648),
.B(n_1630),
.Y(n_1749)
);

AO31x2_ASAP7_75t_L g1750 ( 
.A1(n_1735),
.A2(n_1644),
.A3(n_1677),
.B(n_1622),
.Y(n_1750)
);

AND2x2_ASAP7_75t_L g1751 ( 
.A(n_1702),
.B(n_1679),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1712),
.Y(n_1752)
);

NOR2x1_ASAP7_75t_SL g1753 ( 
.A(n_1724),
.B(n_1665),
.Y(n_1753)
);

AOI21xp5_ASAP7_75t_L g1754 ( 
.A1(n_1686),
.A2(n_1670),
.B(n_1665),
.Y(n_1754)
);

INVx1_ASAP7_75t_SL g1755 ( 
.A(n_1694),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1712),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1714),
.Y(n_1757)
);

AOI21xp5_ASAP7_75t_L g1758 ( 
.A1(n_1705),
.A2(n_1698),
.B(n_1670),
.Y(n_1758)
);

OAI21x1_ASAP7_75t_L g1759 ( 
.A1(n_1731),
.A2(n_1648),
.B(n_1674),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1714),
.Y(n_1760)
);

NAND2xp5_ASAP7_75t_L g1761 ( 
.A(n_1706),
.B(n_1616),
.Y(n_1761)
);

AOI21x1_ASAP7_75t_L g1762 ( 
.A1(n_1738),
.A2(n_1649),
.B(n_1645),
.Y(n_1762)
);

INVx2_ASAP7_75t_L g1763 ( 
.A(n_1710),
.Y(n_1763)
);

AO21x1_ASAP7_75t_L g1764 ( 
.A1(n_1705),
.A2(n_1676),
.B(n_1633),
.Y(n_1764)
);

AO21x2_ASAP7_75t_L g1765 ( 
.A1(n_1696),
.A2(n_1668),
.B(n_1675),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_L g1766 ( 
.A(n_1729),
.B(n_1651),
.Y(n_1766)
);

AO31x2_ASAP7_75t_L g1767 ( 
.A1(n_1735),
.A2(n_1682),
.A3(n_1629),
.B(n_1625),
.Y(n_1767)
);

OR2x6_ASAP7_75t_L g1768 ( 
.A(n_1689),
.B(n_1667),
.Y(n_1768)
);

NAND2x1p5_ASAP7_75t_L g1769 ( 
.A(n_1701),
.B(n_1667),
.Y(n_1769)
);

A2O1A1Ixp33_ASAP7_75t_L g1770 ( 
.A1(n_1723),
.A2(n_1623),
.B(n_1654),
.C(n_1681),
.Y(n_1770)
);

OAI21xp5_ASAP7_75t_L g1771 ( 
.A1(n_1721),
.A2(n_1634),
.B(n_1669),
.Y(n_1771)
);

OAI21x1_ASAP7_75t_L g1772 ( 
.A1(n_1731),
.A2(n_1640),
.B(n_1662),
.Y(n_1772)
);

OAI22xp5_ASAP7_75t_L g1773 ( 
.A1(n_1736),
.A2(n_1611),
.B1(n_1634),
.B2(n_1667),
.Y(n_1773)
);

OAI211xp5_ASAP7_75t_L g1774 ( 
.A1(n_1745),
.A2(n_1673),
.B(n_778),
.C(n_790),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_L g1775 ( 
.A(n_1702),
.B(n_1672),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1719),
.Y(n_1776)
);

AOI21xp5_ASAP7_75t_L g1777 ( 
.A1(n_1698),
.A2(n_1636),
.B(n_1663),
.Y(n_1777)
);

NAND2xp5_ASAP7_75t_L g1778 ( 
.A(n_1719),
.B(n_1635),
.Y(n_1778)
);

NAND2xp5_ASAP7_75t_L g1779 ( 
.A(n_1739),
.B(n_1646),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1689),
.Y(n_1780)
);

BUFx8_ASAP7_75t_SL g1781 ( 
.A(n_1692),
.Y(n_1781)
);

INVx2_ASAP7_75t_L g1782 ( 
.A(n_1710),
.Y(n_1782)
);

OR2x2_ASAP7_75t_L g1783 ( 
.A(n_1728),
.B(n_1734),
.Y(n_1783)
);

NAND2xp5_ASAP7_75t_SL g1784 ( 
.A(n_1701),
.B(n_1618),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1728),
.Y(n_1785)
);

HB1xp67_ASAP7_75t_L g1786 ( 
.A(n_1708),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1734),
.Y(n_1787)
);

INVx2_ASAP7_75t_SL g1788 ( 
.A(n_1741),
.Y(n_1788)
);

OAI21x1_ASAP7_75t_L g1789 ( 
.A1(n_1687),
.A2(n_1725),
.B(n_1708),
.Y(n_1789)
);

AO21x2_ASAP7_75t_L g1790 ( 
.A1(n_1720),
.A2(n_1652),
.B(n_790),
.Y(n_1790)
);

OAI21xp5_ASAP7_75t_L g1791 ( 
.A1(n_1693),
.A2(n_821),
.B(n_791),
.Y(n_1791)
);

OAI21xp5_ASAP7_75t_L g1792 ( 
.A1(n_1693),
.A2(n_821),
.B(n_791),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1740),
.Y(n_1793)
);

NAND2xp33_ASAP7_75t_R g1794 ( 
.A(n_1741),
.B(n_1611),
.Y(n_1794)
);

NAND2xp5_ASAP7_75t_L g1795 ( 
.A(n_1780),
.B(n_1709),
.Y(n_1795)
);

INVx2_ASAP7_75t_L g1796 ( 
.A(n_1789),
.Y(n_1796)
);

HB1xp67_ASAP7_75t_L g1797 ( 
.A(n_1757),
.Y(n_1797)
);

INVx2_ASAP7_75t_L g1798 ( 
.A(n_1789),
.Y(n_1798)
);

INVx3_ASAP7_75t_L g1799 ( 
.A(n_1749),
.Y(n_1799)
);

INVx2_ASAP7_75t_L g1800 ( 
.A(n_1763),
.Y(n_1800)
);

BUFx2_ASAP7_75t_L g1801 ( 
.A(n_1786),
.Y(n_1801)
);

OAI21x1_ASAP7_75t_L g1802 ( 
.A1(n_1749),
.A2(n_1725),
.B(n_1708),
.Y(n_1802)
);

INVx2_ASAP7_75t_L g1803 ( 
.A(n_1763),
.Y(n_1803)
);

INVx2_ASAP7_75t_L g1804 ( 
.A(n_1782),
.Y(n_1804)
);

INVx2_ASAP7_75t_L g1805 ( 
.A(n_1782),
.Y(n_1805)
);

NAND2xp5_ASAP7_75t_L g1806 ( 
.A(n_1760),
.B(n_1709),
.Y(n_1806)
);

OA21x2_ASAP7_75t_L g1807 ( 
.A1(n_1786),
.A2(n_1687),
.B(n_1691),
.Y(n_1807)
);

BUFx3_ASAP7_75t_L g1808 ( 
.A(n_1748),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1752),
.Y(n_1809)
);

AND2x2_ASAP7_75t_L g1810 ( 
.A(n_1756),
.B(n_1725),
.Y(n_1810)
);

OAI21xp5_ASAP7_75t_L g1811 ( 
.A1(n_1770),
.A2(n_1704),
.B(n_1722),
.Y(n_1811)
);

NAND3xp33_ASAP7_75t_L g1812 ( 
.A(n_1770),
.B(n_1711),
.C(n_1732),
.Y(n_1812)
);

OA21x2_ASAP7_75t_L g1813 ( 
.A1(n_1791),
.A2(n_1691),
.B(n_1700),
.Y(n_1813)
);

INVx2_ASAP7_75t_L g1814 ( 
.A(n_1785),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1776),
.Y(n_1815)
);

AO21x2_ASAP7_75t_L g1816 ( 
.A1(n_1764),
.A2(n_1703),
.B(n_1700),
.Y(n_1816)
);

HB1xp67_ASAP7_75t_L g1817 ( 
.A(n_1765),
.Y(n_1817)
);

OAI21x1_ASAP7_75t_L g1818 ( 
.A1(n_1777),
.A2(n_1716),
.B(n_1709),
.Y(n_1818)
);

AOI21xp5_ASAP7_75t_L g1819 ( 
.A1(n_1758),
.A2(n_1768),
.B(n_1754),
.Y(n_1819)
);

NAND2xp5_ASAP7_75t_L g1820 ( 
.A(n_1779),
.B(n_1716),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1787),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1793),
.Y(n_1822)
);

OR2x2_ASAP7_75t_L g1823 ( 
.A(n_1761),
.B(n_1768),
.Y(n_1823)
);

INVx2_ASAP7_75t_L g1824 ( 
.A(n_1783),
.Y(n_1824)
);

INVx2_ASAP7_75t_L g1825 ( 
.A(n_1767),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1778),
.Y(n_1826)
);

NAND2xp5_ASAP7_75t_L g1827 ( 
.A(n_1765),
.B(n_1716),
.Y(n_1827)
);

INVx2_ASAP7_75t_L g1828 ( 
.A(n_1767),
.Y(n_1828)
);

AND2x2_ASAP7_75t_L g1829 ( 
.A(n_1768),
.B(n_1697),
.Y(n_1829)
);

INVx1_ASAP7_75t_SL g1830 ( 
.A(n_1751),
.Y(n_1830)
);

INVx4_ASAP7_75t_L g1831 ( 
.A(n_1769),
.Y(n_1831)
);

AND2x2_ASAP7_75t_L g1832 ( 
.A(n_1747),
.B(n_1697),
.Y(n_1832)
);

INVx2_ASAP7_75t_L g1833 ( 
.A(n_1767),
.Y(n_1833)
);

AND2x2_ASAP7_75t_L g1834 ( 
.A(n_1747),
.B(n_1699),
.Y(n_1834)
);

AND2x2_ASAP7_75t_L g1835 ( 
.A(n_1747),
.B(n_1699),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1767),
.Y(n_1836)
);

BUFx2_ASAP7_75t_L g1837 ( 
.A(n_1746),
.Y(n_1837)
);

HB1xp67_ASAP7_75t_L g1838 ( 
.A(n_1766),
.Y(n_1838)
);

INVx5_ASAP7_75t_L g1839 ( 
.A(n_1746),
.Y(n_1839)
);

BUFx2_ASAP7_75t_L g1840 ( 
.A(n_1746),
.Y(n_1840)
);

INVx2_ASAP7_75t_L g1841 ( 
.A(n_1750),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1792),
.Y(n_1842)
);

INVx3_ASAP7_75t_L g1843 ( 
.A(n_1759),
.Y(n_1843)
);

INVx2_ASAP7_75t_L g1844 ( 
.A(n_1750),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1750),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1750),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1769),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_1772),
.Y(n_1848)
);

AOI22xp33_ASAP7_75t_L g1849 ( 
.A1(n_1812),
.A2(n_1736),
.B1(n_1730),
.B2(n_1771),
.Y(n_1849)
);

AOI22xp33_ASAP7_75t_L g1850 ( 
.A1(n_1812),
.A2(n_1730),
.B1(n_1711),
.B2(n_1784),
.Y(n_1850)
);

OAI22xp5_ASAP7_75t_L g1851 ( 
.A1(n_1812),
.A2(n_1784),
.B1(n_1748),
.B2(n_1775),
.Y(n_1851)
);

NAND4xp25_ASAP7_75t_L g1852 ( 
.A(n_1819),
.B(n_792),
.C(n_796),
.D(n_776),
.Y(n_1852)
);

OR2x2_ASAP7_75t_L g1853 ( 
.A(n_1838),
.B(n_1688),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1797),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1797),
.Y(n_1855)
);

AND2x2_ASAP7_75t_L g1856 ( 
.A(n_1830),
.B(n_1748),
.Y(n_1856)
);

OAI221xp5_ASAP7_75t_L g1857 ( 
.A1(n_1819),
.A2(n_1742),
.B1(n_1774),
.B2(n_1713),
.C(n_1695),
.Y(n_1857)
);

AOI21xp5_ASAP7_75t_L g1858 ( 
.A1(n_1811),
.A2(n_1753),
.B(n_1773),
.Y(n_1858)
);

AND2x2_ASAP7_75t_L g1859 ( 
.A(n_1830),
.B(n_1788),
.Y(n_1859)
);

AO31x2_ASAP7_75t_L g1860 ( 
.A1(n_1841),
.A2(n_1740),
.A3(n_1727),
.B(n_796),
.Y(n_1860)
);

OAI211xp5_ASAP7_75t_L g1861 ( 
.A1(n_1838),
.A2(n_804),
.B(n_805),
.C(n_792),
.Y(n_1861)
);

AOI221xp5_ASAP7_75t_L g1862 ( 
.A1(n_1845),
.A2(n_969),
.B1(n_994),
.B2(n_959),
.C(n_956),
.Y(n_1862)
);

OA211x2_ASAP7_75t_L g1863 ( 
.A1(n_1811),
.A2(n_1794),
.B(n_1781),
.C(n_1694),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1809),
.Y(n_1864)
);

OAI22xp5_ASAP7_75t_L g1865 ( 
.A1(n_1842),
.A2(n_1755),
.B1(n_1701),
.B2(n_1704),
.Y(n_1865)
);

OAI21xp33_ASAP7_75t_L g1866 ( 
.A1(n_1820),
.A2(n_805),
.B(n_804),
.Y(n_1866)
);

NOR2xp33_ASAP7_75t_L g1867 ( 
.A(n_1830),
.B(n_1781),
.Y(n_1867)
);

OAI211xp5_ASAP7_75t_L g1868 ( 
.A1(n_1801),
.A2(n_1806),
.B(n_1811),
.C(n_1820),
.Y(n_1868)
);

INVx2_ASAP7_75t_L g1869 ( 
.A(n_1800),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1809),
.Y(n_1870)
);

INVx2_ASAP7_75t_L g1871 ( 
.A(n_1814),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1809),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1815),
.Y(n_1873)
);

AOI221xp5_ASAP7_75t_L g1874 ( 
.A1(n_1845),
.A2(n_994),
.B1(n_969),
.B2(n_959),
.C(n_982),
.Y(n_1874)
);

INVx2_ASAP7_75t_SL g1875 ( 
.A(n_1808),
.Y(n_1875)
);

INVxp33_ASAP7_75t_L g1876 ( 
.A(n_1823),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_1815),
.Y(n_1877)
);

AOI22xp33_ASAP7_75t_L g1878 ( 
.A1(n_1842),
.A2(n_1730),
.B1(n_1704),
.B2(n_1722),
.Y(n_1878)
);

INVx1_ASAP7_75t_L g1879 ( 
.A(n_1815),
.Y(n_1879)
);

A2O1A1Ixp33_ASAP7_75t_L g1880 ( 
.A1(n_1842),
.A2(n_1743),
.B(n_1733),
.C(n_969),
.Y(n_1880)
);

INVx2_ASAP7_75t_L g1881 ( 
.A(n_1869),
.Y(n_1881)
);

INVx2_ASAP7_75t_L g1882 ( 
.A(n_1869),
.Y(n_1882)
);

OR2x2_ASAP7_75t_L g1883 ( 
.A(n_1854),
.B(n_1823),
.Y(n_1883)
);

OR2x2_ASAP7_75t_L g1884 ( 
.A(n_1855),
.B(n_1823),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_1864),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1870),
.Y(n_1886)
);

INVx2_ASAP7_75t_L g1887 ( 
.A(n_1871),
.Y(n_1887)
);

HB1xp67_ASAP7_75t_L g1888 ( 
.A(n_1872),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1873),
.Y(n_1889)
);

INVx2_ASAP7_75t_L g1890 ( 
.A(n_1860),
.Y(n_1890)
);

AOI22xp33_ASAP7_75t_L g1891 ( 
.A1(n_1849),
.A2(n_1844),
.B1(n_1841),
.B2(n_1845),
.Y(n_1891)
);

CKINVDCx20_ASAP7_75t_R g1892 ( 
.A(n_1867),
.Y(n_1892)
);

INVx2_ASAP7_75t_L g1893 ( 
.A(n_1860),
.Y(n_1893)
);

OR2x2_ASAP7_75t_L g1894 ( 
.A(n_1853),
.B(n_1823),
.Y(n_1894)
);

INVx2_ASAP7_75t_L g1895 ( 
.A(n_1877),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1879),
.Y(n_1896)
);

NAND2xp5_ASAP7_75t_L g1897 ( 
.A(n_1851),
.B(n_1826),
.Y(n_1897)
);

NAND2xp5_ASAP7_75t_L g1898 ( 
.A(n_1868),
.B(n_1826),
.Y(n_1898)
);

OR2x2_ASAP7_75t_L g1899 ( 
.A(n_1876),
.B(n_1826),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1876),
.Y(n_1900)
);

NAND2xp5_ASAP7_75t_L g1901 ( 
.A(n_1859),
.B(n_1810),
.Y(n_1901)
);

INVxp67_ASAP7_75t_L g1902 ( 
.A(n_1867),
.Y(n_1902)
);

NAND2xp5_ASAP7_75t_L g1903 ( 
.A(n_1856),
.B(n_1810),
.Y(n_1903)
);

AND2x2_ASAP7_75t_L g1904 ( 
.A(n_1875),
.B(n_1837),
.Y(n_1904)
);

AND2x4_ASAP7_75t_L g1905 ( 
.A(n_1858),
.B(n_1839),
.Y(n_1905)
);

INVx2_ASAP7_75t_L g1906 ( 
.A(n_1860),
.Y(n_1906)
);

NAND2xp5_ASAP7_75t_L g1907 ( 
.A(n_1865),
.B(n_1810),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1860),
.Y(n_1908)
);

HB1xp67_ASAP7_75t_L g1909 ( 
.A(n_1863),
.Y(n_1909)
);

INVx2_ASAP7_75t_L g1910 ( 
.A(n_1857),
.Y(n_1910)
);

AND2x2_ASAP7_75t_L g1911 ( 
.A(n_1850),
.B(n_1837),
.Y(n_1911)
);

AND2x2_ASAP7_75t_L g1912 ( 
.A(n_1905),
.B(n_1808),
.Y(n_1912)
);

AND2x2_ASAP7_75t_L g1913 ( 
.A(n_1905),
.B(n_1801),
.Y(n_1913)
);

AND2x4_ASAP7_75t_L g1914 ( 
.A(n_1905),
.B(n_1839),
.Y(n_1914)
);

INVx2_ASAP7_75t_L g1915 ( 
.A(n_1881),
.Y(n_1915)
);

INVx2_ASAP7_75t_L g1916 ( 
.A(n_1881),
.Y(n_1916)
);

AOI22xp33_ASAP7_75t_SL g1917 ( 
.A1(n_1911),
.A2(n_1861),
.B1(n_1817),
.B2(n_1844),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1888),
.Y(n_1918)
);

INVx1_ASAP7_75t_SL g1919 ( 
.A(n_1892),
.Y(n_1919)
);

INVx3_ASAP7_75t_L g1920 ( 
.A(n_1905),
.Y(n_1920)
);

AND2x2_ASAP7_75t_L g1921 ( 
.A(n_1904),
.B(n_1911),
.Y(n_1921)
);

INVx2_ASAP7_75t_L g1922 ( 
.A(n_1881),
.Y(n_1922)
);

INVx2_ASAP7_75t_SL g1923 ( 
.A(n_1895),
.Y(n_1923)
);

INVx1_ASAP7_75t_L g1924 ( 
.A(n_1885),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1885),
.Y(n_1925)
);

AND2x2_ASAP7_75t_L g1926 ( 
.A(n_1904),
.B(n_1801),
.Y(n_1926)
);

AOI22xp33_ASAP7_75t_L g1927 ( 
.A1(n_1910),
.A2(n_1849),
.B1(n_1852),
.B2(n_1844),
.Y(n_1927)
);

NOR2xp33_ASAP7_75t_L g1928 ( 
.A(n_1902),
.B(n_1808),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1886),
.Y(n_1929)
);

NAND2xp5_ASAP7_75t_L g1930 ( 
.A(n_1897),
.B(n_1846),
.Y(n_1930)
);

HB1xp67_ASAP7_75t_L g1931 ( 
.A(n_1895),
.Y(n_1931)
);

NAND2xp5_ASAP7_75t_L g1932 ( 
.A(n_1886),
.B(n_1846),
.Y(n_1932)
);

OR2x2_ASAP7_75t_L g1933 ( 
.A(n_1898),
.B(n_1846),
.Y(n_1933)
);

AND2x2_ASAP7_75t_L g1934 ( 
.A(n_1907),
.B(n_1837),
.Y(n_1934)
);

INVx1_ASAP7_75t_L g1935 ( 
.A(n_1889),
.Y(n_1935)
);

NAND2xp5_ASAP7_75t_L g1936 ( 
.A(n_1889),
.B(n_1896),
.Y(n_1936)
);

NAND2xp5_ASAP7_75t_L g1937 ( 
.A(n_1896),
.B(n_1821),
.Y(n_1937)
);

AND2x2_ASAP7_75t_L g1938 ( 
.A(n_1909),
.B(n_1808),
.Y(n_1938)
);

AND2x2_ASAP7_75t_L g1939 ( 
.A(n_1883),
.B(n_1840),
.Y(n_1939)
);

INVx1_ASAP7_75t_SL g1940 ( 
.A(n_1900),
.Y(n_1940)
);

INVx1_ASAP7_75t_SL g1941 ( 
.A(n_1900),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1899),
.Y(n_1942)
);

HB1xp67_ASAP7_75t_L g1943 ( 
.A(n_1883),
.Y(n_1943)
);

OR2x2_ASAP7_75t_L g1944 ( 
.A(n_1899),
.B(n_1841),
.Y(n_1944)
);

AND2x2_ASAP7_75t_L g1945 ( 
.A(n_1938),
.B(n_1884),
.Y(n_1945)
);

INVx1_ASAP7_75t_L g1946 ( 
.A(n_1924),
.Y(n_1946)
);

OAI22xp5_ASAP7_75t_L g1947 ( 
.A1(n_1917),
.A2(n_1891),
.B1(n_1910),
.B2(n_1850),
.Y(n_1947)
);

NOR3xp33_ASAP7_75t_L g1948 ( 
.A(n_1919),
.B(n_1910),
.C(n_1866),
.Y(n_1948)
);

INVx2_ASAP7_75t_L g1949 ( 
.A(n_1919),
.Y(n_1949)
);

OAI21xp5_ASAP7_75t_L g1950 ( 
.A1(n_1917),
.A2(n_1880),
.B(n_1884),
.Y(n_1950)
);

INVx1_ASAP7_75t_L g1951 ( 
.A(n_1924),
.Y(n_1951)
);

AND2x2_ASAP7_75t_SL g1952 ( 
.A(n_1938),
.B(n_1831),
.Y(n_1952)
);

AOI221xp5_ASAP7_75t_L g1953 ( 
.A1(n_1930),
.A2(n_1880),
.B1(n_1817),
.B2(n_1844),
.C(n_1841),
.Y(n_1953)
);

INVx1_ASAP7_75t_L g1954 ( 
.A(n_1925),
.Y(n_1954)
);

AND2x4_ASAP7_75t_SL g1955 ( 
.A(n_1928),
.B(n_1831),
.Y(n_1955)
);

HB1xp67_ASAP7_75t_L g1956 ( 
.A(n_1943),
.Y(n_1956)
);

AND2x2_ASAP7_75t_L g1957 ( 
.A(n_1921),
.B(n_1903),
.Y(n_1957)
);

OR2x2_ASAP7_75t_L g1958 ( 
.A(n_1943),
.B(n_1894),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_1925),
.Y(n_1959)
);

OAI211xp5_ASAP7_75t_L g1960 ( 
.A1(n_1940),
.A2(n_1843),
.B(n_1799),
.C(n_824),
.Y(n_1960)
);

NOR2xp33_ASAP7_75t_L g1961 ( 
.A(n_1940),
.B(n_1901),
.Y(n_1961)
);

NAND2xp5_ASAP7_75t_SL g1962 ( 
.A(n_1941),
.B(n_1839),
.Y(n_1962)
);

OR2x2_ASAP7_75t_L g1963 ( 
.A(n_1941),
.B(n_1894),
.Y(n_1963)
);

AND2x2_ASAP7_75t_L g1964 ( 
.A(n_1921),
.B(n_1840),
.Y(n_1964)
);

AND2x2_ASAP7_75t_L g1965 ( 
.A(n_1912),
.B(n_1840),
.Y(n_1965)
);

INVx1_ASAP7_75t_L g1966 ( 
.A(n_1929),
.Y(n_1966)
);

OAI22xp5_ASAP7_75t_L g1967 ( 
.A1(n_1927),
.A2(n_1839),
.B1(n_1831),
.B2(n_1829),
.Y(n_1967)
);

AND2x2_ASAP7_75t_L g1968 ( 
.A(n_1912),
.B(n_1843),
.Y(n_1968)
);

OAI22xp5_ASAP7_75t_L g1969 ( 
.A1(n_1930),
.A2(n_1839),
.B1(n_1831),
.B2(n_1829),
.Y(n_1969)
);

INVx1_ASAP7_75t_L g1970 ( 
.A(n_1929),
.Y(n_1970)
);

AOI22xp5_ASAP7_75t_L g1971 ( 
.A1(n_1933),
.A2(n_1908),
.B1(n_1834),
.B2(n_1835),
.Y(n_1971)
);

AO21x2_ASAP7_75t_L g1972 ( 
.A1(n_1942),
.A2(n_1882),
.B(n_1887),
.Y(n_1972)
);

INVx1_ASAP7_75t_L g1973 ( 
.A(n_1935),
.Y(n_1973)
);

AOI22xp33_ASAP7_75t_SL g1974 ( 
.A1(n_1933),
.A2(n_1832),
.B1(n_1835),
.B2(n_1834),
.Y(n_1974)
);

NOR2xp33_ASAP7_75t_L g1975 ( 
.A(n_1918),
.B(n_819),
.Y(n_1975)
);

HB1xp67_ASAP7_75t_L g1976 ( 
.A(n_1949),
.Y(n_1976)
);

NAND2xp5_ASAP7_75t_L g1977 ( 
.A(n_1949),
.B(n_1918),
.Y(n_1977)
);

INVx1_ASAP7_75t_L g1978 ( 
.A(n_1956),
.Y(n_1978)
);

NAND4xp25_ASAP7_75t_L g1979 ( 
.A(n_1961),
.B(n_1920),
.C(n_1934),
.D(n_1913),
.Y(n_1979)
);

INVx3_ASAP7_75t_L g1980 ( 
.A(n_1972),
.Y(n_1980)
);

OAI211xp5_ASAP7_75t_SL g1981 ( 
.A1(n_1962),
.A2(n_1920),
.B(n_1942),
.C(n_1936),
.Y(n_1981)
);

INVx1_ASAP7_75t_L g1982 ( 
.A(n_1946),
.Y(n_1982)
);

NAND2xp33_ASAP7_75t_SL g1983 ( 
.A(n_1945),
.B(n_1958),
.Y(n_1983)
);

AND2x2_ASAP7_75t_L g1984 ( 
.A(n_1945),
.B(n_1934),
.Y(n_1984)
);

NAND2xp5_ASAP7_75t_L g1985 ( 
.A(n_1948),
.B(n_1934),
.Y(n_1985)
);

NAND2xp5_ASAP7_75t_L g1986 ( 
.A(n_1957),
.B(n_1923),
.Y(n_1986)
);

AND2x2_ASAP7_75t_L g1987 ( 
.A(n_1952),
.B(n_1939),
.Y(n_1987)
);

OR2x2_ASAP7_75t_L g1988 ( 
.A(n_1963),
.B(n_1936),
.Y(n_1988)
);

NAND2xp5_ASAP7_75t_L g1989 ( 
.A(n_1957),
.B(n_1923),
.Y(n_1989)
);

AND2x2_ASAP7_75t_L g1990 ( 
.A(n_1952),
.B(n_1939),
.Y(n_1990)
);

AND2x2_ASAP7_75t_L g1991 ( 
.A(n_1964),
.B(n_1920),
.Y(n_1991)
);

AND2x2_ASAP7_75t_L g1992 ( 
.A(n_1964),
.B(n_1920),
.Y(n_1992)
);

OR2x2_ASAP7_75t_L g1993 ( 
.A(n_1951),
.B(n_1935),
.Y(n_1993)
);

INVx1_ASAP7_75t_L g1994 ( 
.A(n_1954),
.Y(n_1994)
);

INVx2_ASAP7_75t_L g1995 ( 
.A(n_1972),
.Y(n_1995)
);

AND2x2_ASAP7_75t_L g1996 ( 
.A(n_1955),
.B(n_1926),
.Y(n_1996)
);

AND2x2_ASAP7_75t_L g1997 ( 
.A(n_1955),
.B(n_1926),
.Y(n_1997)
);

NAND2xp5_ASAP7_75t_L g1998 ( 
.A(n_1975),
.B(n_1923),
.Y(n_1998)
);

AND2x2_ASAP7_75t_L g1999 ( 
.A(n_1965),
.B(n_1926),
.Y(n_1999)
);

NAND2xp5_ASAP7_75t_L g2000 ( 
.A(n_1975),
.B(n_1931),
.Y(n_2000)
);

AND2x2_ASAP7_75t_L g2001 ( 
.A(n_1965),
.B(n_1961),
.Y(n_2001)
);

INVx1_ASAP7_75t_L g2002 ( 
.A(n_1959),
.Y(n_2002)
);

AOI22xp33_ASAP7_75t_L g2003 ( 
.A1(n_1947),
.A2(n_1916),
.B1(n_1922),
.B2(n_1915),
.Y(n_2003)
);

INVx1_ASAP7_75t_L g2004 ( 
.A(n_1966),
.Y(n_2004)
);

NAND2xp5_ASAP7_75t_L g2005 ( 
.A(n_1960),
.B(n_1950),
.Y(n_2005)
);

INVx1_ASAP7_75t_L g2006 ( 
.A(n_1970),
.Y(n_2006)
);

INVx1_ASAP7_75t_L g2007 ( 
.A(n_1973),
.Y(n_2007)
);

AND2x2_ASAP7_75t_L g2008 ( 
.A(n_1968),
.B(n_1913),
.Y(n_2008)
);

INVx1_ASAP7_75t_L g2009 ( 
.A(n_1968),
.Y(n_2009)
);

OR2x2_ASAP7_75t_L g2010 ( 
.A(n_1971),
.B(n_1931),
.Y(n_2010)
);

AND2x2_ASAP7_75t_L g2011 ( 
.A(n_1974),
.B(n_1913),
.Y(n_2011)
);

NAND2xp5_ASAP7_75t_L g2012 ( 
.A(n_1953),
.B(n_1937),
.Y(n_2012)
);

NAND4xp25_ASAP7_75t_L g2013 ( 
.A(n_1962),
.B(n_1914),
.C(n_1937),
.D(n_1843),
.Y(n_2013)
);

AND2x4_ASAP7_75t_L g2014 ( 
.A(n_1969),
.B(n_1914),
.Y(n_2014)
);

AND2x2_ASAP7_75t_L g2015 ( 
.A(n_1967),
.B(n_1914),
.Y(n_2015)
);

NAND2xp5_ASAP7_75t_L g2016 ( 
.A(n_1949),
.B(n_1932),
.Y(n_2016)
);

NOR2xp33_ASAP7_75t_L g2017 ( 
.A(n_1949),
.B(n_1914),
.Y(n_2017)
);

NAND2xp5_ASAP7_75t_L g2018 ( 
.A(n_1949),
.B(n_1932),
.Y(n_2018)
);

HB1xp67_ASAP7_75t_L g2019 ( 
.A(n_1949),
.Y(n_2019)
);

INVx2_ASAP7_75t_L g2020 ( 
.A(n_1991),
.Y(n_2020)
);

NOR2xp33_ASAP7_75t_L g2021 ( 
.A(n_2000),
.B(n_1944),
.Y(n_2021)
);

AND2x2_ASAP7_75t_L g2022 ( 
.A(n_2001),
.B(n_1843),
.Y(n_2022)
);

AND2x2_ASAP7_75t_L g2023 ( 
.A(n_2001),
.B(n_1984),
.Y(n_2023)
);

OR2x2_ASAP7_75t_L g2024 ( 
.A(n_1976),
.B(n_1944),
.Y(n_2024)
);

OR2x2_ASAP7_75t_L g2025 ( 
.A(n_2019),
.B(n_1915),
.Y(n_2025)
);

INVx2_ASAP7_75t_L g2026 ( 
.A(n_1991),
.Y(n_2026)
);

INVx1_ASAP7_75t_SL g2027 ( 
.A(n_1983),
.Y(n_2027)
);

INVx2_ASAP7_75t_L g2028 ( 
.A(n_1992),
.Y(n_2028)
);

INVx1_ASAP7_75t_L g2029 ( 
.A(n_1993),
.Y(n_2029)
);

AND2x2_ASAP7_75t_L g2030 ( 
.A(n_1984),
.B(n_1843),
.Y(n_2030)
);

AND2x4_ASAP7_75t_L g2031 ( 
.A(n_1978),
.B(n_1915),
.Y(n_2031)
);

OR2x2_ASAP7_75t_L g2032 ( 
.A(n_1985),
.B(n_1916),
.Y(n_2032)
);

INVx1_ASAP7_75t_L g2033 ( 
.A(n_1993),
.Y(n_2033)
);

NAND2xp5_ASAP7_75t_L g2034 ( 
.A(n_1998),
.B(n_1916),
.Y(n_2034)
);

OR2x2_ASAP7_75t_L g2035 ( 
.A(n_1977),
.B(n_1986),
.Y(n_2035)
);

OR2x2_ASAP7_75t_L g2036 ( 
.A(n_1989),
.B(n_1922),
.Y(n_2036)
);

INVx1_ASAP7_75t_L g2037 ( 
.A(n_1994),
.Y(n_2037)
);

INVxp67_ASAP7_75t_SL g2038 ( 
.A(n_1980),
.Y(n_2038)
);

AND2x2_ASAP7_75t_L g2039 ( 
.A(n_1992),
.B(n_1843),
.Y(n_2039)
);

INVx2_ASAP7_75t_L g2040 ( 
.A(n_1999),
.Y(n_2040)
);

INVx1_ASAP7_75t_L g2041 ( 
.A(n_1994),
.Y(n_2041)
);

AND2x2_ASAP7_75t_L g2042 ( 
.A(n_1987),
.B(n_1829),
.Y(n_2042)
);

INVx1_ASAP7_75t_L g2043 ( 
.A(n_2002),
.Y(n_2043)
);

NAND2x1_ASAP7_75t_SL g2044 ( 
.A(n_1987),
.B(n_1922),
.Y(n_2044)
);

INVx1_ASAP7_75t_L g2045 ( 
.A(n_2002),
.Y(n_2045)
);

AND2x2_ASAP7_75t_L g2046 ( 
.A(n_1990),
.B(n_1829),
.Y(n_2046)
);

INVxp67_ASAP7_75t_SL g2047 ( 
.A(n_1980),
.Y(n_2047)
);

NAND3xp33_ASAP7_75t_L g2048 ( 
.A(n_1983),
.B(n_2003),
.C(n_1980),
.Y(n_2048)
);

AOI22xp5_ASAP7_75t_L g2049 ( 
.A1(n_2005),
.A2(n_1874),
.B1(n_1862),
.B2(n_1816),
.Y(n_2049)
);

INVx1_ASAP7_75t_L g2050 ( 
.A(n_1982),
.Y(n_2050)
);

BUFx2_ASAP7_75t_L g2051 ( 
.A(n_1988),
.Y(n_2051)
);

OR2x2_ASAP7_75t_L g2052 ( 
.A(n_1988),
.B(n_1979),
.Y(n_2052)
);

NAND2xp5_ASAP7_75t_L g2053 ( 
.A(n_2017),
.B(n_1887),
.Y(n_2053)
);

AOI22xp33_ASAP7_75t_L g2054 ( 
.A1(n_1995),
.A2(n_2012),
.B1(n_2010),
.B2(n_2011),
.Y(n_2054)
);

INVx2_ASAP7_75t_SL g2055 ( 
.A(n_1996),
.Y(n_2055)
);

NAND2xp5_ASAP7_75t_L g2056 ( 
.A(n_2004),
.B(n_819),
.Y(n_2056)
);

INVx1_ASAP7_75t_L g2057 ( 
.A(n_2006),
.Y(n_2057)
);

INVx1_ASAP7_75t_SL g2058 ( 
.A(n_1995),
.Y(n_2058)
);

INVx1_ASAP7_75t_SL g2059 ( 
.A(n_2016),
.Y(n_2059)
);

OR2x2_ASAP7_75t_L g2060 ( 
.A(n_2018),
.B(n_1887),
.Y(n_2060)
);

INVx1_ASAP7_75t_L g2061 ( 
.A(n_2007),
.Y(n_2061)
);

AND2x2_ASAP7_75t_L g2062 ( 
.A(n_1990),
.B(n_1799),
.Y(n_2062)
);

NAND2xp67_ASAP7_75t_L g2063 ( 
.A(n_2015),
.B(n_1882),
.Y(n_2063)
);

INVx1_ASAP7_75t_L g2064 ( 
.A(n_1999),
.Y(n_2064)
);

OR2x6_ASAP7_75t_L g2065 ( 
.A(n_2010),
.B(n_1743),
.Y(n_2065)
);

AND2x4_ASAP7_75t_L g2066 ( 
.A(n_1996),
.B(n_1839),
.Y(n_2066)
);

AND2x2_ASAP7_75t_L g2067 ( 
.A(n_1997),
.B(n_1799),
.Y(n_2067)
);

NOR2x1_ASAP7_75t_L g2068 ( 
.A(n_1981),
.B(n_2013),
.Y(n_2068)
);

NAND2xp5_ASAP7_75t_L g2069 ( 
.A(n_2009),
.B(n_824),
.Y(n_2069)
);

OR2x2_ASAP7_75t_L g2070 ( 
.A(n_2009),
.B(n_1882),
.Y(n_2070)
);

NAND2xp5_ASAP7_75t_L g2071 ( 
.A(n_2011),
.B(n_829),
.Y(n_2071)
);

INVx1_ASAP7_75t_SL g2072 ( 
.A(n_1997),
.Y(n_2072)
);

AND2x4_ASAP7_75t_L g2073 ( 
.A(n_2008),
.B(n_1839),
.Y(n_2073)
);

NAND2xp5_ASAP7_75t_L g2074 ( 
.A(n_2008),
.B(n_829),
.Y(n_2074)
);

INVx1_ASAP7_75t_L g2075 ( 
.A(n_2014),
.Y(n_2075)
);

OR2x2_ASAP7_75t_L g2076 ( 
.A(n_2014),
.B(n_1806),
.Y(n_2076)
);

NAND2xp5_ASAP7_75t_L g2077 ( 
.A(n_2014),
.B(n_830),
.Y(n_2077)
);

HB1xp67_ASAP7_75t_L g2078 ( 
.A(n_2015),
.Y(n_2078)
);

INVx1_ASAP7_75t_L g2079 ( 
.A(n_1976),
.Y(n_2079)
);

INVx1_ASAP7_75t_L g2080 ( 
.A(n_1976),
.Y(n_2080)
);

NAND2xp5_ASAP7_75t_L g2081 ( 
.A(n_1976),
.B(n_830),
.Y(n_2081)
);

HB1xp67_ASAP7_75t_L g2082 ( 
.A(n_1976),
.Y(n_2082)
);

INVx1_ASAP7_75t_L g2083 ( 
.A(n_1976),
.Y(n_2083)
);

INVx2_ASAP7_75t_L g2084 ( 
.A(n_2044),
.Y(n_2084)
);

OR2x2_ASAP7_75t_L g2085 ( 
.A(n_2051),
.B(n_832),
.Y(n_2085)
);

INVx2_ASAP7_75t_SL g2086 ( 
.A(n_2023),
.Y(n_2086)
);

NAND2xp5_ASAP7_75t_L g2087 ( 
.A(n_2059),
.B(n_832),
.Y(n_2087)
);

INVxp67_ASAP7_75t_SL g2088 ( 
.A(n_2082),
.Y(n_2088)
);

AOI211xp5_ASAP7_75t_L g2089 ( 
.A1(n_2048),
.A2(n_835),
.B(n_839),
.C(n_834),
.Y(n_2089)
);

INVx1_ASAP7_75t_L g2090 ( 
.A(n_2038),
.Y(n_2090)
);

A2O1A1Ixp33_ASAP7_75t_L g2091 ( 
.A1(n_2048),
.A2(n_835),
.B(n_839),
.C(n_834),
.Y(n_2091)
);

INVxp67_ASAP7_75t_L g2092 ( 
.A(n_2078),
.Y(n_2092)
);

HB1xp67_ASAP7_75t_L g2093 ( 
.A(n_2040),
.Y(n_2093)
);

AND2x2_ASAP7_75t_L g2094 ( 
.A(n_2072),
.B(n_1799),
.Y(n_2094)
);

OAI32xp33_ASAP7_75t_L g2095 ( 
.A1(n_2027),
.A2(n_2052),
.A3(n_2054),
.B1(n_2059),
.B2(n_2032),
.Y(n_2095)
);

INVxp67_ASAP7_75t_SL g2096 ( 
.A(n_2081),
.Y(n_2096)
);

INVx1_ASAP7_75t_L g2097 ( 
.A(n_2047),
.Y(n_2097)
);

INVx1_ASAP7_75t_L g2098 ( 
.A(n_2064),
.Y(n_2098)
);

NAND3xp33_ASAP7_75t_L g2099 ( 
.A(n_2079),
.B(n_994),
.C(n_959),
.Y(n_2099)
);

INVxp33_ASAP7_75t_L g2100 ( 
.A(n_2020),
.Y(n_2100)
);

INVx2_ASAP7_75t_L g2101 ( 
.A(n_2025),
.Y(n_2101)
);

INVx1_ASAP7_75t_L g2102 ( 
.A(n_2081),
.Y(n_2102)
);

OR2x2_ASAP7_75t_L g2103 ( 
.A(n_2072),
.B(n_845),
.Y(n_2103)
);

INVx2_ASAP7_75t_L g2104 ( 
.A(n_2026),
.Y(n_2104)
);

AOI32xp33_ASAP7_75t_L g2105 ( 
.A1(n_2068),
.A2(n_1834),
.A3(n_1835),
.B1(n_1832),
.B2(n_1799),
.Y(n_2105)
);

AND2x4_ASAP7_75t_L g2106 ( 
.A(n_2055),
.B(n_1839),
.Y(n_2106)
);

NAND2xp5_ASAP7_75t_L g2107 ( 
.A(n_2027),
.B(n_2028),
.Y(n_2107)
);

OAI322xp33_ASAP7_75t_L g2108 ( 
.A1(n_2080),
.A2(n_875),
.A3(n_953),
.B1(n_869),
.B2(n_861),
.C1(n_879),
.C2(n_867),
.Y(n_2108)
);

INVx1_ASAP7_75t_L g2109 ( 
.A(n_2074),
.Y(n_2109)
);

AOI22xp5_ASAP7_75t_L g2110 ( 
.A1(n_2049),
.A2(n_861),
.B1(n_867),
.B2(n_845),
.Y(n_2110)
);

A2O1A1Ixp33_ASAP7_75t_L g2111 ( 
.A1(n_2049),
.A2(n_869),
.B(n_879),
.C(n_875),
.Y(n_2111)
);

INVx2_ASAP7_75t_L g2112 ( 
.A(n_2065),
.Y(n_2112)
);

INVx1_ASAP7_75t_L g2113 ( 
.A(n_2083),
.Y(n_2113)
);

INVx1_ASAP7_75t_L g2114 ( 
.A(n_2056),
.Y(n_2114)
);

AOI21xp5_ASAP7_75t_L g2115 ( 
.A1(n_2071),
.A2(n_882),
.B(n_881),
.Y(n_2115)
);

INVx1_ASAP7_75t_L g2116 ( 
.A(n_2056),
.Y(n_2116)
);

NOR2xp33_ASAP7_75t_L g2117 ( 
.A(n_2035),
.B(n_881),
.Y(n_2117)
);

INVx1_ASAP7_75t_L g2118 ( 
.A(n_2077),
.Y(n_2118)
);

OAI22xp5_ASAP7_75t_L g2119 ( 
.A1(n_2075),
.A2(n_1839),
.B1(n_1799),
.B2(n_1831),
.Y(n_2119)
);

INVx1_ASAP7_75t_L g2120 ( 
.A(n_2029),
.Y(n_2120)
);

INVx1_ASAP7_75t_L g2121 ( 
.A(n_2033),
.Y(n_2121)
);

INVx1_ASAP7_75t_L g2122 ( 
.A(n_2069),
.Y(n_2122)
);

NOR2xp67_ASAP7_75t_L g2123 ( 
.A(n_2036),
.B(n_0),
.Y(n_2123)
);

AOI22xp5_ASAP7_75t_L g2124 ( 
.A1(n_2058),
.A2(n_882),
.B1(n_898),
.B2(n_890),
.Y(n_2124)
);

INVx2_ASAP7_75t_L g2125 ( 
.A(n_2065),
.Y(n_2125)
);

AND2x2_ASAP7_75t_L g2126 ( 
.A(n_2042),
.B(n_1839),
.Y(n_2126)
);

A2O1A1Ixp33_ASAP7_75t_L g2127 ( 
.A1(n_2021),
.A2(n_890),
.B(n_901),
.C(n_898),
.Y(n_2127)
);

AOI21xp33_ASAP7_75t_SL g2128 ( 
.A1(n_2071),
.A2(n_907),
.B(n_901),
.Y(n_2128)
);

NAND2xp5_ASAP7_75t_L g2129 ( 
.A(n_2031),
.B(n_907),
.Y(n_2129)
);

OR2x2_ASAP7_75t_L g2130 ( 
.A(n_2034),
.B(n_913),
.Y(n_2130)
);

INVx1_ASAP7_75t_L g2131 ( 
.A(n_2037),
.Y(n_2131)
);

AND2x2_ASAP7_75t_L g2132 ( 
.A(n_2046),
.B(n_913),
.Y(n_2132)
);

INVx3_ASAP7_75t_L g2133 ( 
.A(n_2066),
.Y(n_2133)
);

INVx1_ASAP7_75t_L g2134 ( 
.A(n_2041),
.Y(n_2134)
);

INVx1_ASAP7_75t_L g2135 ( 
.A(n_2043),
.Y(n_2135)
);

OAI21xp5_ASAP7_75t_SL g2136 ( 
.A1(n_2031),
.A2(n_2066),
.B(n_2057),
.Y(n_2136)
);

NOR2x1_ASAP7_75t_L g2137 ( 
.A(n_2045),
.B(n_917),
.Y(n_2137)
);

INVx1_ASAP7_75t_SL g2138 ( 
.A(n_2024),
.Y(n_2138)
);

NAND2xp5_ASAP7_75t_L g2139 ( 
.A(n_2050),
.B(n_917),
.Y(n_2139)
);

INVx1_ASAP7_75t_L g2140 ( 
.A(n_2058),
.Y(n_2140)
);

INVx1_ASAP7_75t_L g2141 ( 
.A(n_2061),
.Y(n_2141)
);

INVx1_ASAP7_75t_L g2142 ( 
.A(n_2065),
.Y(n_2142)
);

INVx1_ASAP7_75t_L g2143 ( 
.A(n_2060),
.Y(n_2143)
);

INVx1_ASAP7_75t_L g2144 ( 
.A(n_2070),
.Y(n_2144)
);

AOI22xp5_ASAP7_75t_L g2145 ( 
.A1(n_2053),
.A2(n_918),
.B1(n_921),
.B2(n_920),
.Y(n_2145)
);

OAI21xp5_ASAP7_75t_L g2146 ( 
.A1(n_2022),
.A2(n_920),
.B(n_918),
.Y(n_2146)
);

AOI32xp33_ASAP7_75t_L g2147 ( 
.A1(n_2062),
.A2(n_1835),
.A3(n_1834),
.B1(n_1832),
.B2(n_921),
.Y(n_2147)
);

INVx1_ASAP7_75t_L g2148 ( 
.A(n_2063),
.Y(n_2148)
);

AND2x2_ASAP7_75t_SL g2149 ( 
.A(n_2073),
.B(n_1831),
.Y(n_2149)
);

INVxp67_ASAP7_75t_SL g2150 ( 
.A(n_2076),
.Y(n_2150)
);

OR2x2_ASAP7_75t_L g2151 ( 
.A(n_2030),
.B(n_923),
.Y(n_2151)
);

INVx1_ASAP7_75t_L g2152 ( 
.A(n_2067),
.Y(n_2152)
);

INVx1_ASAP7_75t_L g2153 ( 
.A(n_2039),
.Y(n_2153)
);

NAND2xp5_ASAP7_75t_L g2154 ( 
.A(n_2073),
.B(n_923),
.Y(n_2154)
);

AND2x2_ASAP7_75t_L g2155 ( 
.A(n_2023),
.B(n_929),
.Y(n_2155)
);

NAND2xp5_ASAP7_75t_L g2156 ( 
.A(n_2023),
.B(n_929),
.Y(n_2156)
);

OAI21xp33_ASAP7_75t_L g2157 ( 
.A1(n_2054),
.A2(n_1798),
.B(n_1796),
.Y(n_2157)
);

INVx1_ASAP7_75t_L g2158 ( 
.A(n_2082),
.Y(n_2158)
);

INVx1_ASAP7_75t_L g2159 ( 
.A(n_2082),
.Y(n_2159)
);

INVx1_ASAP7_75t_L g2160 ( 
.A(n_2082),
.Y(n_2160)
);

AND2x2_ASAP7_75t_L g2161 ( 
.A(n_2023),
.B(n_932),
.Y(n_2161)
);

NAND2xp5_ASAP7_75t_L g2162 ( 
.A(n_2023),
.B(n_932),
.Y(n_2162)
);

INVxp67_ASAP7_75t_SL g2163 ( 
.A(n_2082),
.Y(n_2163)
);

INVx2_ASAP7_75t_L g2164 ( 
.A(n_2044),
.Y(n_2164)
);

INVx2_ASAP7_75t_L g2165 ( 
.A(n_2044),
.Y(n_2165)
);

INVx1_ASAP7_75t_L g2166 ( 
.A(n_2082),
.Y(n_2166)
);

OAI21xp33_ASAP7_75t_L g2167 ( 
.A1(n_2054),
.A2(n_938),
.B(n_937),
.Y(n_2167)
);

OAI21xp5_ASAP7_75t_L g2168 ( 
.A1(n_2048),
.A2(n_938),
.B(n_937),
.Y(n_2168)
);

INVx1_ASAP7_75t_L g2169 ( 
.A(n_2082),
.Y(n_2169)
);

OAI32xp33_ASAP7_75t_L g2170 ( 
.A1(n_2027),
.A2(n_1794),
.A3(n_940),
.B1(n_954),
.B2(n_953),
.Y(n_2170)
);

NAND2xp5_ASAP7_75t_L g2171 ( 
.A(n_2086),
.B(n_2155),
.Y(n_2171)
);

INVx1_ASAP7_75t_L g2172 ( 
.A(n_2093),
.Y(n_2172)
);

NAND2xp5_ASAP7_75t_L g2173 ( 
.A(n_2161),
.B(n_940),
.Y(n_2173)
);

NAND2xp5_ASAP7_75t_L g2174 ( 
.A(n_2088),
.B(n_945),
.Y(n_2174)
);

INVx2_ASAP7_75t_L g2175 ( 
.A(n_2103),
.Y(n_2175)
);

OAI21xp5_ASAP7_75t_L g2176 ( 
.A1(n_2091),
.A2(n_997),
.B(n_954),
.Y(n_2176)
);

AOI22xp33_ASAP7_75t_SL g2177 ( 
.A1(n_2095),
.A2(n_1893),
.B1(n_1906),
.B2(n_1890),
.Y(n_2177)
);

NAND2xp5_ASAP7_75t_SL g2178 ( 
.A(n_2092),
.B(n_1796),
.Y(n_2178)
);

OR2x2_ASAP7_75t_L g2179 ( 
.A(n_2138),
.B(n_945),
.Y(n_2179)
);

INVx1_ASAP7_75t_SL g2180 ( 
.A(n_2107),
.Y(n_2180)
);

NAND3xp33_ASAP7_75t_L g2181 ( 
.A(n_2089),
.B(n_2140),
.C(n_2168),
.Y(n_2181)
);

AOI22xp5_ASAP7_75t_L g2182 ( 
.A1(n_2084),
.A2(n_1893),
.B1(n_1906),
.B2(n_1890),
.Y(n_2182)
);

AOI22xp5_ASAP7_75t_L g2183 ( 
.A1(n_2164),
.A2(n_1893),
.B1(n_1906),
.B2(n_1890),
.Y(n_2183)
);

AOI21xp33_ASAP7_75t_L g2184 ( 
.A1(n_2165),
.A2(n_1908),
.B(n_957),
.Y(n_2184)
);

NAND2xp5_ASAP7_75t_L g2185 ( 
.A(n_2163),
.B(n_955),
.Y(n_2185)
);

OAI221xp5_ASAP7_75t_L g2186 ( 
.A1(n_2157),
.A2(n_968),
.B1(n_974),
.B2(n_957),
.C(n_955),
.Y(n_2186)
);

INVx1_ASAP7_75t_L g2187 ( 
.A(n_2085),
.Y(n_2187)
);

NOR2xp33_ASAP7_75t_L g2188 ( 
.A(n_2108),
.B(n_968),
.Y(n_2188)
);

A2O1A1Ixp33_ASAP7_75t_L g2189 ( 
.A1(n_2123),
.A2(n_978),
.B(n_981),
.C(n_974),
.Y(n_2189)
);

NAND2x1_ASAP7_75t_L g2190 ( 
.A(n_2133),
.B(n_978),
.Y(n_2190)
);

NAND2xp5_ASAP7_75t_SL g2191 ( 
.A(n_2158),
.B(n_1796),
.Y(n_2191)
);

OAI31xp33_ASAP7_75t_L g2192 ( 
.A1(n_2111),
.A2(n_1733),
.A3(n_984),
.B(n_997),
.Y(n_2192)
);

INVx1_ASAP7_75t_L g2193 ( 
.A(n_2137),
.Y(n_2193)
);

INVx3_ASAP7_75t_L g2194 ( 
.A(n_2133),
.Y(n_2194)
);

AOI211xp5_ASAP7_75t_L g2195 ( 
.A1(n_2100),
.A2(n_984),
.B(n_1003),
.C(n_981),
.Y(n_2195)
);

INVx2_ASAP7_75t_L g2196 ( 
.A(n_2132),
.Y(n_2196)
);

NAND2xp5_ASAP7_75t_L g2197 ( 
.A(n_2150),
.B(n_1003),
.Y(n_2197)
);

INVx2_ASAP7_75t_L g2198 ( 
.A(n_2101),
.Y(n_2198)
);

INVx2_ASAP7_75t_L g2199 ( 
.A(n_2130),
.Y(n_2199)
);

HB1xp67_ASAP7_75t_L g2200 ( 
.A(n_2159),
.Y(n_2200)
);

AND2x2_ASAP7_75t_L g2201 ( 
.A(n_2104),
.B(n_1013),
.Y(n_2201)
);

AOI22xp33_ASAP7_75t_L g2202 ( 
.A1(n_2148),
.A2(n_1828),
.B1(n_1833),
.B2(n_1825),
.Y(n_2202)
);

OR2x2_ASAP7_75t_L g2203 ( 
.A(n_2156),
.B(n_1013),
.Y(n_2203)
);

O2A1O1Ixp33_ASAP7_75t_L g2204 ( 
.A1(n_2170),
.A2(n_897),
.B(n_943),
.C(n_864),
.Y(n_2204)
);

NAND2xp5_ASAP7_75t_L g2205 ( 
.A(n_2117),
.B(n_653),
.Y(n_2205)
);

OAI21xp33_ASAP7_75t_SL g2206 ( 
.A1(n_2105),
.A2(n_1818),
.B(n_1798),
.Y(n_2206)
);

XOR2x2_ASAP7_75t_L g2207 ( 
.A(n_2123),
.B(n_2110),
.Y(n_2207)
);

NAND2xp5_ASAP7_75t_L g2208 ( 
.A(n_2143),
.B(n_655),
.Y(n_2208)
);

AOI22xp5_ASAP7_75t_L g2209 ( 
.A1(n_2110),
.A2(n_1832),
.B1(n_1816),
.B2(n_1827),
.Y(n_2209)
);

AOI21xp5_ASAP7_75t_L g2210 ( 
.A1(n_2167),
.A2(n_958),
.B(n_943),
.Y(n_2210)
);

A2O1A1Ixp33_ASAP7_75t_L g2211 ( 
.A1(n_2167),
.A2(n_958),
.B(n_659),
.C(n_662),
.Y(n_2211)
);

NOR2xp33_ASAP7_75t_L g2212 ( 
.A(n_2162),
.B(n_658),
.Y(n_2212)
);

NAND2xp5_ASAP7_75t_L g2213 ( 
.A(n_2147),
.B(n_666),
.Y(n_2213)
);

OAI21xp33_ASAP7_75t_SL g2214 ( 
.A1(n_2090),
.A2(n_1818),
.B(n_1798),
.Y(n_2214)
);

INVxp67_ASAP7_75t_L g2215 ( 
.A(n_2096),
.Y(n_2215)
);

AND2x4_ASAP7_75t_L g2216 ( 
.A(n_2160),
.B(n_1810),
.Y(n_2216)
);

O2A1O1Ixp33_ASAP7_75t_L g2217 ( 
.A1(n_2127),
.A2(n_1008),
.B(n_868),
.C(n_1733),
.Y(n_2217)
);

INVx1_ASAP7_75t_L g2218 ( 
.A(n_2087),
.Y(n_2218)
);

XOR2x2_ASAP7_75t_L g2219 ( 
.A(n_2099),
.B(n_1762),
.Y(n_2219)
);

AOI21xp5_ASAP7_75t_L g2220 ( 
.A1(n_2129),
.A2(n_674),
.B(n_667),
.Y(n_2220)
);

NAND2xp5_ASAP7_75t_SL g2221 ( 
.A(n_2166),
.B(n_2169),
.Y(n_2221)
);

OAI31xp33_ASAP7_75t_L g2222 ( 
.A1(n_2144),
.A2(n_1733),
.A3(n_1878),
.B(n_1827),
.Y(n_2222)
);

AND2x2_ASAP7_75t_L g2223 ( 
.A(n_2152),
.B(n_1816),
.Y(n_2223)
);

NOR4xp25_ASAP7_75t_L g2224 ( 
.A(n_2097),
.B(n_1008),
.C(n_1798),
.D(n_1796),
.Y(n_2224)
);

AOI21xp5_ASAP7_75t_L g2225 ( 
.A1(n_2136),
.A2(n_679),
.B(n_676),
.Y(n_2225)
);

OAI222xp33_ASAP7_75t_L g2226 ( 
.A1(n_2142),
.A2(n_1878),
.B1(n_1825),
.B2(n_1828),
.C1(n_1833),
.C2(n_1836),
.Y(n_2226)
);

INVx1_ASAP7_75t_L g2227 ( 
.A(n_2151),
.Y(n_2227)
);

INVx1_ASAP7_75t_L g2228 ( 
.A(n_2124),
.Y(n_2228)
);

INVx1_ASAP7_75t_L g2229 ( 
.A(n_2124),
.Y(n_2229)
);

AOI21xp5_ASAP7_75t_L g2230 ( 
.A1(n_2139),
.A2(n_682),
.B(n_680),
.Y(n_2230)
);

OAI32xp33_ASAP7_75t_L g2231 ( 
.A1(n_2113),
.A2(n_688),
.A3(n_691),
.B1(n_687),
.B2(n_685),
.Y(n_2231)
);

AOI21xp5_ASAP7_75t_L g2232 ( 
.A1(n_2115),
.A2(n_693),
.B(n_692),
.Y(n_2232)
);

AOI22xp33_ASAP7_75t_L g2233 ( 
.A1(n_2112),
.A2(n_1828),
.B1(n_1833),
.B2(n_1825),
.Y(n_2233)
);

INVx1_ASAP7_75t_SL g2234 ( 
.A(n_2098),
.Y(n_2234)
);

INVx1_ASAP7_75t_L g2235 ( 
.A(n_2102),
.Y(n_2235)
);

NOR4xp25_ASAP7_75t_L g2236 ( 
.A(n_2131),
.B(n_1848),
.C(n_1733),
.D(n_1795),
.Y(n_2236)
);

NAND2xp5_ASAP7_75t_L g2237 ( 
.A(n_2114),
.B(n_695),
.Y(n_2237)
);

INVx1_ASAP7_75t_L g2238 ( 
.A(n_2116),
.Y(n_2238)
);

NOR2xp33_ASAP7_75t_L g2239 ( 
.A(n_2109),
.B(n_697),
.Y(n_2239)
);

INVx1_ASAP7_75t_L g2240 ( 
.A(n_2154),
.Y(n_2240)
);

OAI21xp33_ASAP7_75t_L g2241 ( 
.A1(n_2153),
.A2(n_1848),
.B(n_1795),
.Y(n_2241)
);

NAND2xp5_ASAP7_75t_L g2242 ( 
.A(n_2145),
.B(n_2122),
.Y(n_2242)
);

INVx1_ASAP7_75t_L g2243 ( 
.A(n_2118),
.Y(n_2243)
);

INVx2_ASAP7_75t_L g2244 ( 
.A(n_2106),
.Y(n_2244)
);

A2O1A1Ixp33_ASAP7_75t_SL g2245 ( 
.A1(n_2141),
.A2(n_2121),
.B(n_2120),
.C(n_2134),
.Y(n_2245)
);

AOI22xp5_ASAP7_75t_L g2246 ( 
.A1(n_2145),
.A2(n_1816),
.B1(n_1813),
.B2(n_1848),
.Y(n_2246)
);

NOR2xp33_ASAP7_75t_SL g2247 ( 
.A(n_2125),
.B(n_1847),
.Y(n_2247)
);

OAI21xp33_ASAP7_75t_SL g2248 ( 
.A1(n_2135),
.A2(n_1818),
.B(n_1802),
.Y(n_2248)
);

AOI322xp5_ASAP7_75t_L g2249 ( 
.A1(n_2094),
.A2(n_1825),
.A3(n_1828),
.B1(n_1833),
.B2(n_1836),
.C1(n_1821),
.C2(n_1822),
.Y(n_2249)
);

NAND2xp5_ASAP7_75t_L g2250 ( 
.A(n_2146),
.B(n_698),
.Y(n_2250)
);

OAI32xp33_ASAP7_75t_L g2251 ( 
.A1(n_2119),
.A2(n_709),
.A3(n_710),
.B1(n_707),
.B2(n_700),
.Y(n_2251)
);

AOI222xp33_ASAP7_75t_L g2252 ( 
.A1(n_2149),
.A2(n_1836),
.B1(n_716),
.B2(n_712),
.C1(n_717),
.C2(n_715),
.Y(n_2252)
);

AOI22xp33_ASAP7_75t_L g2253 ( 
.A1(n_2126),
.A2(n_2106),
.B1(n_1816),
.B2(n_1813),
.Y(n_2253)
);

AOI21xp33_ASAP7_75t_L g2254 ( 
.A1(n_2128),
.A2(n_718),
.B(n_711),
.Y(n_2254)
);

INVx1_ASAP7_75t_L g2255 ( 
.A(n_2128),
.Y(n_2255)
);

INVx1_ASAP7_75t_L g2256 ( 
.A(n_2093),
.Y(n_2256)
);

INVx1_ASAP7_75t_L g2257 ( 
.A(n_2093),
.Y(n_2257)
);

INVx2_ASAP7_75t_L g2258 ( 
.A(n_2086),
.Y(n_2258)
);

INVx1_ASAP7_75t_SL g2259 ( 
.A(n_2138),
.Y(n_2259)
);

INVxp67_ASAP7_75t_L g2260 ( 
.A(n_2093),
.Y(n_2260)
);

INVx1_ASAP7_75t_L g2261 ( 
.A(n_2093),
.Y(n_2261)
);

INVxp67_ASAP7_75t_L g2262 ( 
.A(n_2093),
.Y(n_2262)
);

INVx1_ASAP7_75t_L g2263 ( 
.A(n_2093),
.Y(n_2263)
);

INVx1_ASAP7_75t_L g2264 ( 
.A(n_2093),
.Y(n_2264)
);

NAND2xp5_ASAP7_75t_L g2265 ( 
.A(n_2086),
.B(n_720),
.Y(n_2265)
);

AND2x2_ASAP7_75t_L g2266 ( 
.A(n_2086),
.B(n_1816),
.Y(n_2266)
);

NAND2xp5_ASAP7_75t_SL g2267 ( 
.A(n_2086),
.B(n_702),
.Y(n_2267)
);

INVx1_ASAP7_75t_L g2268 ( 
.A(n_2093),
.Y(n_2268)
);

NOR2xp67_ASAP7_75t_SL g2269 ( 
.A(n_2099),
.B(n_702),
.Y(n_2269)
);

O2A1O1Ixp33_ASAP7_75t_SL g2270 ( 
.A1(n_2092),
.A2(n_1847),
.B(n_4),
.C(n_2),
.Y(n_2270)
);

INVx1_ASAP7_75t_L g2271 ( 
.A(n_2093),
.Y(n_2271)
);

OR2x2_ASAP7_75t_L g2272 ( 
.A(n_2138),
.B(n_2),
.Y(n_2272)
);

AOI22xp5_ASAP7_75t_L g2273 ( 
.A1(n_2140),
.A2(n_1813),
.B1(n_1821),
.B2(n_1822),
.Y(n_2273)
);

INVx1_ASAP7_75t_L g2274 ( 
.A(n_2093),
.Y(n_2274)
);

NAND2xp5_ASAP7_75t_L g2275 ( 
.A(n_2086),
.B(n_722),
.Y(n_2275)
);

INVxp67_ASAP7_75t_L g2276 ( 
.A(n_2093),
.Y(n_2276)
);

NAND3xp33_ASAP7_75t_L g2277 ( 
.A(n_2089),
.B(n_725),
.C(n_723),
.Y(n_2277)
);

INVx2_ASAP7_75t_L g2278 ( 
.A(n_2086),
.Y(n_2278)
);

NAND2xp5_ASAP7_75t_L g2279 ( 
.A(n_2086),
.B(n_727),
.Y(n_2279)
);

INVx1_ASAP7_75t_L g2280 ( 
.A(n_2093),
.Y(n_2280)
);

AOI332xp33_ASAP7_75t_L g2281 ( 
.A1(n_2140),
.A2(n_9),
.A3(n_8),
.B1(n_5),
.B2(n_10),
.B3(n_3),
.C1(n_4),
.C2(n_6),
.Y(n_2281)
);

INVx1_ASAP7_75t_L g2282 ( 
.A(n_2093),
.Y(n_2282)
);

OAI22xp33_ASAP7_75t_L g2283 ( 
.A1(n_2084),
.A2(n_1813),
.B1(n_1847),
.B2(n_1822),
.Y(n_2283)
);

INVx2_ASAP7_75t_L g2284 ( 
.A(n_2086),
.Y(n_2284)
);

INVx1_ASAP7_75t_SL g2285 ( 
.A(n_2138),
.Y(n_2285)
);

AOI21xp33_ASAP7_75t_L g2286 ( 
.A1(n_2095),
.A2(n_730),
.B(n_728),
.Y(n_2286)
);

NAND2xp5_ASAP7_75t_L g2287 ( 
.A(n_2086),
.B(n_731),
.Y(n_2287)
);

NAND2xp5_ASAP7_75t_L g2288 ( 
.A(n_2086),
.B(n_732),
.Y(n_2288)
);

AOI322xp5_ASAP7_75t_L g2289 ( 
.A1(n_2140),
.A2(n_1814),
.A3(n_741),
.B1(n_742),
.B2(n_735),
.C1(n_745),
.C2(n_744),
.Y(n_2289)
);

AOI21xp5_ASAP7_75t_SL g2290 ( 
.A1(n_2091),
.A2(n_750),
.B(n_739),
.Y(n_2290)
);

NAND2xp5_ASAP7_75t_L g2291 ( 
.A(n_2086),
.B(n_751),
.Y(n_2291)
);

OR2x2_ASAP7_75t_L g2292 ( 
.A(n_2138),
.B(n_9),
.Y(n_2292)
);

NAND2xp5_ASAP7_75t_L g2293 ( 
.A(n_2086),
.B(n_752),
.Y(n_2293)
);

NAND2xp5_ASAP7_75t_L g2294 ( 
.A(n_2086),
.B(n_753),
.Y(n_2294)
);

NAND2x1p5_ASAP7_75t_L g2295 ( 
.A(n_2137),
.B(n_702),
.Y(n_2295)
);

OAI211xp5_ASAP7_75t_L g2296 ( 
.A1(n_2095),
.A2(n_754),
.B(n_757),
.C(n_755),
.Y(n_2296)
);

NAND3xp33_ASAP7_75t_L g2297 ( 
.A(n_2089),
.B(n_763),
.C(n_758),
.Y(n_2297)
);

AOI22xp33_ASAP7_75t_L g2298 ( 
.A1(n_2148),
.A2(n_1813),
.B1(n_1807),
.B2(n_1704),
.Y(n_2298)
);

AOI222xp33_ASAP7_75t_L g2299 ( 
.A1(n_2140),
.A2(n_774),
.B1(n_770),
.B2(n_780),
.C1(n_773),
.C2(n_766),
.Y(n_2299)
);

INVx1_ASAP7_75t_L g2300 ( 
.A(n_2093),
.Y(n_2300)
);

HB1xp67_ASAP7_75t_L g2301 ( 
.A(n_2086),
.Y(n_2301)
);

NAND2x1_ASAP7_75t_SL g2302 ( 
.A(n_2093),
.B(n_1807),
.Y(n_2302)
);

NOR2xp33_ASAP7_75t_L g2303 ( 
.A(n_2108),
.B(n_782),
.Y(n_2303)
);

INVx1_ASAP7_75t_L g2304 ( 
.A(n_2093),
.Y(n_2304)
);

NAND2xp5_ASAP7_75t_SL g2305 ( 
.A(n_2086),
.B(n_702),
.Y(n_2305)
);

AND2x4_ASAP7_75t_L g2306 ( 
.A(n_2086),
.B(n_1818),
.Y(n_2306)
);

INVx1_ASAP7_75t_L g2307 ( 
.A(n_2093),
.Y(n_2307)
);

NAND2xp5_ASAP7_75t_L g2308 ( 
.A(n_2086),
.B(n_783),
.Y(n_2308)
);

INVx1_ASAP7_75t_L g2309 ( 
.A(n_2093),
.Y(n_2309)
);

INVx1_ASAP7_75t_L g2310 ( 
.A(n_2093),
.Y(n_2310)
);

OAI22xp33_ASAP7_75t_L g2311 ( 
.A1(n_2084),
.A2(n_1813),
.B1(n_1814),
.B2(n_1807),
.Y(n_2311)
);

OR2x2_ASAP7_75t_L g2312 ( 
.A(n_2138),
.B(n_11),
.Y(n_2312)
);

AO21x2_ASAP7_75t_L g2313 ( 
.A1(n_2168),
.A2(n_12),
.B(n_13),
.Y(n_2313)
);

INVx1_ASAP7_75t_L g2314 ( 
.A(n_2093),
.Y(n_2314)
);

INVx1_ASAP7_75t_L g2315 ( 
.A(n_2093),
.Y(n_2315)
);

AOI22xp5_ASAP7_75t_L g2316 ( 
.A1(n_2140),
.A2(n_1813),
.B1(n_1807),
.B2(n_785),
.Y(n_2316)
);

NAND2xp5_ASAP7_75t_L g2317 ( 
.A(n_2086),
.B(n_788),
.Y(n_2317)
);

AOI21xp5_ASAP7_75t_L g2318 ( 
.A1(n_2095),
.A2(n_802),
.B(n_793),
.Y(n_2318)
);

OAI21xp5_ASAP7_75t_L g2319 ( 
.A1(n_2091),
.A2(n_809),
.B(n_803),
.Y(n_2319)
);

INVx1_ASAP7_75t_L g2320 ( 
.A(n_2093),
.Y(n_2320)
);

AND2x2_ASAP7_75t_L g2321 ( 
.A(n_2259),
.B(n_810),
.Y(n_2321)
);

NOR2xp33_ASAP7_75t_L g2322 ( 
.A(n_2285),
.B(n_812),
.Y(n_2322)
);

INVx1_ASAP7_75t_L g2323 ( 
.A(n_2301),
.Y(n_2323)
);

OAI21xp33_ASAP7_75t_SL g2324 ( 
.A1(n_2302),
.A2(n_2221),
.B(n_2180),
.Y(n_2324)
);

INVx1_ASAP7_75t_L g2325 ( 
.A(n_2272),
.Y(n_2325)
);

AOI22xp5_ASAP7_75t_L g2326 ( 
.A1(n_2198),
.A2(n_817),
.B1(n_818),
.B2(n_815),
.Y(n_2326)
);

AOI21xp5_ASAP7_75t_L g2327 ( 
.A1(n_2245),
.A2(n_825),
.B(n_823),
.Y(n_2327)
);

INVx2_ASAP7_75t_L g2328 ( 
.A(n_2295),
.Y(n_2328)
);

AOI321xp33_ASAP7_75t_L g2329 ( 
.A1(n_2236),
.A2(n_1814),
.A3(n_1824),
.B1(n_1804),
.B2(n_1805),
.C(n_1803),
.Y(n_2329)
);

INVx1_ASAP7_75t_L g2330 ( 
.A(n_2292),
.Y(n_2330)
);

OAI21xp33_ASAP7_75t_L g2331 ( 
.A1(n_2258),
.A2(n_831),
.B(n_826),
.Y(n_2331)
);

INVx1_ASAP7_75t_L g2332 ( 
.A(n_2312),
.Y(n_2332)
);

INVx2_ASAP7_75t_L g2333 ( 
.A(n_2194),
.Y(n_2333)
);

NAND2xp5_ASAP7_75t_L g2334 ( 
.A(n_2194),
.B(n_2260),
.Y(n_2334)
);

OAI21xp33_ASAP7_75t_L g2335 ( 
.A1(n_2278),
.A2(n_836),
.B(n_833),
.Y(n_2335)
);

INVx2_ASAP7_75t_L g2336 ( 
.A(n_2190),
.Y(n_2336)
);

OR2x2_ASAP7_75t_L g2337 ( 
.A(n_2172),
.B(n_13),
.Y(n_2337)
);

NAND2xp5_ASAP7_75t_L g2338 ( 
.A(n_2262),
.B(n_837),
.Y(n_2338)
);

OAI22xp5_ASAP7_75t_L g2339 ( 
.A1(n_2276),
.A2(n_1807),
.B1(n_841),
.B2(n_842),
.Y(n_2339)
);

INVx1_ASAP7_75t_L g2340 ( 
.A(n_2256),
.Y(n_2340)
);

INVx1_ASAP7_75t_L g2341 ( 
.A(n_2257),
.Y(n_2341)
);

NAND2xp5_ASAP7_75t_L g2342 ( 
.A(n_2299),
.B(n_838),
.Y(n_2342)
);

INVx1_ASAP7_75t_L g2343 ( 
.A(n_2261),
.Y(n_2343)
);

INVx1_ASAP7_75t_L g2344 ( 
.A(n_2263),
.Y(n_2344)
);

NAND2xp5_ASAP7_75t_L g2345 ( 
.A(n_2212),
.B(n_843),
.Y(n_2345)
);

OR2x2_ASAP7_75t_L g2346 ( 
.A(n_2264),
.B(n_14),
.Y(n_2346)
);

AOI221xp5_ASAP7_75t_L g2347 ( 
.A1(n_2186),
.A2(n_844),
.B1(n_850),
.B2(n_849),
.C(n_848),
.Y(n_2347)
);

INVx2_ASAP7_75t_L g2348 ( 
.A(n_2313),
.Y(n_2348)
);

NAND2xp5_ASAP7_75t_SL g2349 ( 
.A(n_2268),
.B(n_702),
.Y(n_2349)
);

AND2x2_ASAP7_75t_L g2350 ( 
.A(n_2284),
.B(n_2271),
.Y(n_2350)
);

OAI21xp5_ASAP7_75t_L g2351 ( 
.A1(n_2296),
.A2(n_852),
.B(n_851),
.Y(n_2351)
);

AOI31xp33_ASAP7_75t_SL g2352 ( 
.A1(n_2215),
.A2(n_2171),
.A3(n_2244),
.B(n_2252),
.Y(n_2352)
);

INVx1_ASAP7_75t_L g2353 ( 
.A(n_2274),
.Y(n_2353)
);

AOI221x1_ASAP7_75t_L g2354 ( 
.A1(n_2280),
.A2(n_865),
.B1(n_866),
.B2(n_858),
.C(n_806),
.Y(n_2354)
);

NOR2xp33_ASAP7_75t_L g2355 ( 
.A(n_2270),
.B(n_853),
.Y(n_2355)
);

NAND2xp5_ASAP7_75t_L g2356 ( 
.A(n_2303),
.B(n_855),
.Y(n_2356)
);

NOR2xp33_ASAP7_75t_L g2357 ( 
.A(n_2179),
.B(n_857),
.Y(n_2357)
);

AOI221xp5_ASAP7_75t_L g2358 ( 
.A1(n_2181),
.A2(n_859),
.B1(n_863),
.B2(n_862),
.C(n_860),
.Y(n_2358)
);

AND2x2_ASAP7_75t_L g2359 ( 
.A(n_2282),
.B(n_870),
.Y(n_2359)
);

INVx1_ASAP7_75t_L g2360 ( 
.A(n_2300),
.Y(n_2360)
);

XNOR2xp5_ASAP7_75t_L g2361 ( 
.A(n_2207),
.B(n_872),
.Y(n_2361)
);

INVx2_ASAP7_75t_L g2362 ( 
.A(n_2313),
.Y(n_2362)
);

NAND2xp5_ASAP7_75t_SL g2363 ( 
.A(n_2304),
.B(n_806),
.Y(n_2363)
);

AND2x4_ASAP7_75t_L g2364 ( 
.A(n_2307),
.B(n_14),
.Y(n_2364)
);

INVx1_ASAP7_75t_L g2365 ( 
.A(n_2309),
.Y(n_2365)
);

XOR2x2_ASAP7_75t_L g2366 ( 
.A(n_2277),
.B(n_15),
.Y(n_2366)
);

AND2x2_ASAP7_75t_L g2367 ( 
.A(n_2310),
.B(n_873),
.Y(n_2367)
);

AND2x2_ASAP7_75t_L g2368 ( 
.A(n_2314),
.B(n_874),
.Y(n_2368)
);

O2A1O1Ixp33_ASAP7_75t_L g2369 ( 
.A1(n_2286),
.A2(n_877),
.B(n_878),
.C(n_876),
.Y(n_2369)
);

OAI221xp5_ASAP7_75t_L g2370 ( 
.A1(n_2206),
.A2(n_887),
.B1(n_888),
.B2(n_886),
.C(n_880),
.Y(n_2370)
);

INVx3_ASAP7_75t_L g2371 ( 
.A(n_2315),
.Y(n_2371)
);

INVx1_ASAP7_75t_L g2372 ( 
.A(n_2320),
.Y(n_2372)
);

AOI21xp33_ASAP7_75t_SL g2373 ( 
.A1(n_2200),
.A2(n_18),
.B(n_17),
.Y(n_2373)
);

A2O1A1Ixp33_ASAP7_75t_L g2374 ( 
.A1(n_2281),
.A2(n_909),
.B(n_928),
.C(n_894),
.Y(n_2374)
);

O2A1O1Ixp33_ASAP7_75t_L g2375 ( 
.A1(n_2318),
.A2(n_893),
.B(n_899),
.C(n_891),
.Y(n_2375)
);

NAND2xp5_ASAP7_75t_L g2376 ( 
.A(n_2195),
.B(n_900),
.Y(n_2376)
);

NAND2xp5_ASAP7_75t_L g2377 ( 
.A(n_2234),
.B(n_902),
.Y(n_2377)
);

INVx2_ASAP7_75t_L g2378 ( 
.A(n_2175),
.Y(n_2378)
);

OAI22xp5_ASAP7_75t_L g2379 ( 
.A1(n_2316),
.A2(n_1807),
.B1(n_904),
.B2(n_905),
.Y(n_2379)
);

NAND2xp5_ASAP7_75t_L g2380 ( 
.A(n_2201),
.B(n_903),
.Y(n_2380)
);

INVx1_ASAP7_75t_L g2381 ( 
.A(n_2173),
.Y(n_2381)
);

AOI22xp33_ASAP7_75t_SL g2382 ( 
.A1(n_2206),
.A2(n_933),
.B1(n_947),
.B2(n_911),
.Y(n_2382)
);

NAND2xp5_ASAP7_75t_L g2383 ( 
.A(n_2193),
.B(n_2196),
.Y(n_2383)
);

OAI221xp5_ASAP7_75t_L g2384 ( 
.A1(n_2222),
.A2(n_2246),
.B1(n_2248),
.B2(n_2177),
.C(n_2209),
.Y(n_2384)
);

INVx1_ASAP7_75t_L g2385 ( 
.A(n_2187),
.Y(n_2385)
);

AOI211xp5_ASAP7_75t_L g2386 ( 
.A1(n_2251),
.A2(n_910),
.B(n_912),
.C(n_908),
.Y(n_2386)
);

INVxp33_ASAP7_75t_L g2387 ( 
.A(n_2188),
.Y(n_2387)
);

NAND2xp5_ASAP7_75t_L g2388 ( 
.A(n_2239),
.B(n_915),
.Y(n_2388)
);

NAND2xp5_ASAP7_75t_L g2389 ( 
.A(n_2289),
.B(n_2211),
.Y(n_2389)
);

AOI222xp33_ASAP7_75t_L g2390 ( 
.A1(n_2214),
.A2(n_934),
.B1(n_925),
.B2(n_935),
.C1(n_930),
.C2(n_922),
.Y(n_2390)
);

AOI22xp5_ASAP7_75t_L g2391 ( 
.A1(n_2228),
.A2(n_2229),
.B1(n_2227),
.B2(n_2250),
.Y(n_2391)
);

AOI222xp33_ASAP7_75t_L g2392 ( 
.A1(n_2214),
.A2(n_946),
.B1(n_941),
.B2(n_948),
.C1(n_944),
.C2(n_939),
.Y(n_2392)
);

NOR2xp33_ASAP7_75t_L g2393 ( 
.A(n_2205),
.B(n_949),
.Y(n_2393)
);

INVx1_ASAP7_75t_L g2394 ( 
.A(n_2203),
.Y(n_2394)
);

AOI22xp33_ASAP7_75t_L g2395 ( 
.A1(n_2218),
.A2(n_1807),
.B1(n_806),
.B2(n_865),
.Y(n_2395)
);

NAND2xp5_ASAP7_75t_L g2396 ( 
.A(n_2225),
.B(n_950),
.Y(n_2396)
);

OR2x2_ASAP7_75t_L g2397 ( 
.A(n_2265),
.B(n_2275),
.Y(n_2397)
);

NAND2xp5_ASAP7_75t_L g2398 ( 
.A(n_2235),
.B(n_2290),
.Y(n_2398)
);

AOI31xp33_ASAP7_75t_L g2399 ( 
.A1(n_2238),
.A2(n_961),
.A3(n_962),
.B(n_960),
.Y(n_2399)
);

INVx1_ASAP7_75t_L g2400 ( 
.A(n_2197),
.Y(n_2400)
);

NAND2xp5_ASAP7_75t_L g2401 ( 
.A(n_2230),
.B(n_963),
.Y(n_2401)
);

AOI311xp33_ASAP7_75t_L g2402 ( 
.A1(n_2243),
.A2(n_22),
.A3(n_15),
.B(n_19),
.C(n_23),
.Y(n_2402)
);

INVx1_ASAP7_75t_L g2403 ( 
.A(n_2279),
.Y(n_2403)
);

AOI21xp33_ASAP7_75t_L g2404 ( 
.A1(n_2204),
.A2(n_965),
.B(n_964),
.Y(n_2404)
);

INVx1_ASAP7_75t_L g2405 ( 
.A(n_2287),
.Y(n_2405)
);

OAI221xp5_ASAP7_75t_L g2406 ( 
.A1(n_2248),
.A2(n_973),
.B1(n_976),
.B2(n_970),
.C(n_966),
.Y(n_2406)
);

INVx1_ASAP7_75t_L g2407 ( 
.A(n_2288),
.Y(n_2407)
);

INVx1_ASAP7_75t_L g2408 ( 
.A(n_2291),
.Y(n_2408)
);

NOR3xp33_ASAP7_75t_L g2409 ( 
.A(n_2184),
.B(n_979),
.C(n_977),
.Y(n_2409)
);

AOI21xp5_ASAP7_75t_L g2410 ( 
.A1(n_2267),
.A2(n_985),
.B(n_980),
.Y(n_2410)
);

INVxp67_ASAP7_75t_SL g2411 ( 
.A(n_2213),
.Y(n_2411)
);

AOI31xp33_ASAP7_75t_L g2412 ( 
.A1(n_2174),
.A2(n_987),
.A3(n_988),
.B(n_986),
.Y(n_2412)
);

INVx2_ASAP7_75t_L g2413 ( 
.A(n_2199),
.Y(n_2413)
);

NAND2xp5_ASAP7_75t_L g2414 ( 
.A(n_2240),
.B(n_990),
.Y(n_2414)
);

INVx1_ASAP7_75t_L g2415 ( 
.A(n_2293),
.Y(n_2415)
);

OAI322xp33_ASAP7_75t_L g2416 ( 
.A1(n_2191),
.A2(n_989),
.A3(n_992),
.B1(n_1002),
.B2(n_1004),
.C1(n_996),
.C2(n_991),
.Y(n_2416)
);

AOI22xp5_ASAP7_75t_L g2417 ( 
.A1(n_2297),
.A2(n_1006),
.B1(n_1007),
.B2(n_1005),
.Y(n_2417)
);

OAI22xp5_ASAP7_75t_L g2418 ( 
.A1(n_2273),
.A2(n_1010),
.B1(n_1011),
.B2(n_1009),
.Y(n_2418)
);

INVx1_ASAP7_75t_L g2419 ( 
.A(n_2294),
.Y(n_2419)
);

OR2x2_ASAP7_75t_L g2420 ( 
.A(n_2308),
.B(n_19),
.Y(n_2420)
);

NAND2xp5_ASAP7_75t_L g2421 ( 
.A(n_2232),
.B(n_1016),
.Y(n_2421)
);

INVx1_ASAP7_75t_L g2422 ( 
.A(n_2317),
.Y(n_2422)
);

NAND2xp5_ASAP7_75t_L g2423 ( 
.A(n_2305),
.B(n_1017),
.Y(n_2423)
);

OAI21xp33_ASAP7_75t_L g2424 ( 
.A1(n_2216),
.A2(n_1021),
.B(n_1018),
.Y(n_2424)
);

O2A1O1Ixp33_ASAP7_75t_L g2425 ( 
.A1(n_2189),
.A2(n_1023),
.B(n_1024),
.C(n_1022),
.Y(n_2425)
);

OR2x2_ASAP7_75t_L g2426 ( 
.A(n_2208),
.B(n_2185),
.Y(n_2426)
);

NAND2xp5_ASAP7_75t_L g2427 ( 
.A(n_2220),
.B(n_2237),
.Y(n_2427)
);

AOI211xp5_ASAP7_75t_L g2428 ( 
.A1(n_2231),
.A2(n_1026),
.B(n_1027),
.C(n_1025),
.Y(n_2428)
);

AOI22xp33_ASAP7_75t_L g2429 ( 
.A1(n_2255),
.A2(n_806),
.B1(n_865),
.B2(n_858),
.Y(n_2429)
);

NAND2xp5_ASAP7_75t_L g2430 ( 
.A(n_2216),
.B(n_22),
.Y(n_2430)
);

NAND2xp5_ASAP7_75t_L g2431 ( 
.A(n_2176),
.B(n_24),
.Y(n_2431)
);

INVx2_ASAP7_75t_L g2432 ( 
.A(n_2306),
.Y(n_2432)
);

OAI22xp33_ASAP7_75t_L g2433 ( 
.A1(n_2247),
.A2(n_1737),
.B1(n_1722),
.B2(n_1800),
.Y(n_2433)
);

INVx1_ASAP7_75t_L g2434 ( 
.A(n_2242),
.Y(n_2434)
);

CKINVDCx14_ASAP7_75t_R g2435 ( 
.A(n_2266),
.Y(n_2435)
);

INVx1_ASAP7_75t_SL g2436 ( 
.A(n_2219),
.Y(n_2436)
);

AOI222xp33_ASAP7_75t_L g2437 ( 
.A1(n_2226),
.A2(n_866),
.B1(n_858),
.B2(n_999),
.C1(n_865),
.C2(n_806),
.Y(n_2437)
);

AOI22xp33_ASAP7_75t_SL g2438 ( 
.A1(n_2306),
.A2(n_806),
.B1(n_865),
.B2(n_858),
.Y(n_2438)
);

NOR2x1_ASAP7_75t_L g2439 ( 
.A(n_2319),
.B(n_2178),
.Y(n_2439)
);

NAND2xp5_ASAP7_75t_L g2440 ( 
.A(n_2355),
.B(n_2224),
.Y(n_2440)
);

AOI221xp5_ASAP7_75t_L g2441 ( 
.A1(n_2324),
.A2(n_2311),
.B1(n_2283),
.B2(n_2217),
.C(n_2253),
.Y(n_2441)
);

AOI211xp5_ASAP7_75t_L g2442 ( 
.A1(n_2324),
.A2(n_2223),
.B(n_2269),
.C(n_2192),
.Y(n_2442)
);

AOI22xp5_ASAP7_75t_SL g2443 ( 
.A1(n_2327),
.A2(n_2210),
.B1(n_2254),
.B2(n_2241),
.Y(n_2443)
);

AND2x2_ASAP7_75t_L g2444 ( 
.A(n_2350),
.B(n_2182),
.Y(n_2444)
);

OAI22xp5_ASAP7_75t_L g2445 ( 
.A1(n_2334),
.A2(n_2183),
.B1(n_2298),
.B2(n_2233),
.Y(n_2445)
);

A2O1A1Ixp33_ASAP7_75t_L g2446 ( 
.A1(n_2374),
.A2(n_2373),
.B(n_2435),
.C(n_2384),
.Y(n_2446)
);

AOI21xp5_ASAP7_75t_L g2447 ( 
.A1(n_2399),
.A2(n_2412),
.B(n_2406),
.Y(n_2447)
);

NAND2xp5_ASAP7_75t_L g2448 ( 
.A(n_2364),
.B(n_2249),
.Y(n_2448)
);

NOR2xp33_ASAP7_75t_L g2449 ( 
.A(n_2333),
.B(n_2202),
.Y(n_2449)
);

AOI21xp33_ASAP7_75t_L g2450 ( 
.A1(n_2387),
.A2(n_865),
.B(n_858),
.Y(n_2450)
);

NAND4xp25_ASAP7_75t_L g2451 ( 
.A(n_2323),
.B(n_28),
.C(n_25),
.D(n_27),
.Y(n_2451)
);

NAND2xp5_ASAP7_75t_L g2452 ( 
.A(n_2364),
.B(n_27),
.Y(n_2452)
);

NAND2xp5_ASAP7_75t_L g2453 ( 
.A(n_2321),
.B(n_28),
.Y(n_2453)
);

AOI21xp33_ASAP7_75t_L g2454 ( 
.A1(n_2390),
.A2(n_866),
.B(n_858),
.Y(n_2454)
);

OA22x2_ASAP7_75t_L g2455 ( 
.A1(n_2340),
.A2(n_1690),
.B1(n_1802),
.B2(n_1707),
.Y(n_2455)
);

NOR2x1_ASAP7_75t_SL g2456 ( 
.A(n_2337),
.B(n_866),
.Y(n_2456)
);

NOR2xp33_ASAP7_75t_L g2457 ( 
.A(n_2336),
.B(n_29),
.Y(n_2457)
);

AOI22xp5_ASAP7_75t_L g2458 ( 
.A1(n_2427),
.A2(n_1790),
.B1(n_1824),
.B2(n_999),
.Y(n_2458)
);

O2A1O1Ixp33_ASAP7_75t_L g2459 ( 
.A1(n_2352),
.A2(n_32),
.B(n_30),
.C(n_31),
.Y(n_2459)
);

OAI21xp5_ASAP7_75t_L g2460 ( 
.A1(n_2439),
.A2(n_1707),
.B(n_1802),
.Y(n_2460)
);

O2A1O1Ixp33_ASAP7_75t_L g2461 ( 
.A1(n_2371),
.A2(n_33),
.B(n_30),
.C(n_31),
.Y(n_2461)
);

NOR2xp33_ASAP7_75t_SL g2462 ( 
.A(n_2322),
.B(n_866),
.Y(n_2462)
);

OA22x2_ASAP7_75t_L g2463 ( 
.A1(n_2341),
.A2(n_1690),
.B1(n_1802),
.B2(n_1824),
.Y(n_2463)
);

NAND2xp5_ASAP7_75t_SL g2464 ( 
.A(n_2402),
.B(n_2371),
.Y(n_2464)
);

AOI22xp5_ASAP7_75t_L g2465 ( 
.A1(n_2325),
.A2(n_1790),
.B1(n_1824),
.B2(n_999),
.Y(n_2465)
);

NAND2xp5_ASAP7_75t_L g2466 ( 
.A(n_2330),
.B(n_2332),
.Y(n_2466)
);

AOI22xp33_ASAP7_75t_L g2467 ( 
.A1(n_2370),
.A2(n_2382),
.B1(n_2348),
.B2(n_2362),
.Y(n_2467)
);

AOI322xp5_ASAP7_75t_L g2468 ( 
.A1(n_2436),
.A2(n_1800),
.A3(n_1805),
.B1(n_1803),
.B2(n_1804),
.C1(n_999),
.C2(n_1000),
.Y(n_2468)
);

NAND2xp5_ASAP7_75t_L g2469 ( 
.A(n_2357),
.B(n_34),
.Y(n_2469)
);

AOI211xp5_ASAP7_75t_L g2470 ( 
.A1(n_2379),
.A2(n_999),
.B(n_1000),
.C(n_866),
.Y(n_2470)
);

NAND2xp5_ASAP7_75t_L g2471 ( 
.A(n_2434),
.B(n_35),
.Y(n_2471)
);

NOR3xp33_ASAP7_75t_L g2472 ( 
.A(n_2416),
.B(n_641),
.C(n_609),
.Y(n_2472)
);

NAND4xp25_ASAP7_75t_SL g2473 ( 
.A(n_2343),
.B(n_39),
.C(n_36),
.D(n_38),
.Y(n_2473)
);

NAND2xp5_ASAP7_75t_L g2474 ( 
.A(n_2359),
.B(n_36),
.Y(n_2474)
);

NAND2xp5_ASAP7_75t_SL g2475 ( 
.A(n_2358),
.B(n_999),
.Y(n_2475)
);

INVx1_ASAP7_75t_L g2476 ( 
.A(n_2346),
.Y(n_2476)
);

A2O1A1Ixp33_ASAP7_75t_L g2477 ( 
.A1(n_2432),
.A2(n_1000),
.B(n_1703),
.C(n_1800),
.Y(n_2477)
);

NAND4xp25_ASAP7_75t_L g2478 ( 
.A(n_2383),
.B(n_41),
.C(n_38),
.D(n_39),
.Y(n_2478)
);

OAI211xp5_ASAP7_75t_SL g2479 ( 
.A1(n_2385),
.A2(n_45),
.B(n_42),
.C(n_44),
.Y(n_2479)
);

NAND3xp33_ASAP7_75t_SL g2480 ( 
.A(n_2392),
.B(n_777),
.C(n_689),
.Y(n_2480)
);

NAND2xp5_ASAP7_75t_L g2481 ( 
.A(n_2367),
.B(n_42),
.Y(n_2481)
);

OAI221xp5_ASAP7_75t_L g2482 ( 
.A1(n_2329),
.A2(n_1000),
.B1(n_1737),
.B2(n_1722),
.C(n_1803),
.Y(n_2482)
);

OAI221xp5_ASAP7_75t_L g2483 ( 
.A1(n_2398),
.A2(n_1000),
.B1(n_1737),
.B2(n_1804),
.C(n_1803),
.Y(n_2483)
);

INVx1_ASAP7_75t_L g2484 ( 
.A(n_2380),
.Y(n_2484)
);

OAI21xp33_ASAP7_75t_L g2485 ( 
.A1(n_2389),
.A2(n_1000),
.B(n_1804),
.Y(n_2485)
);

OAI22xp5_ASAP7_75t_L g2486 ( 
.A1(n_2344),
.A2(n_1805),
.B1(n_1737),
.B2(n_1727),
.Y(n_2486)
);

OA22x2_ASAP7_75t_L g2487 ( 
.A1(n_2353),
.A2(n_1717),
.B1(n_1718),
.B2(n_1805),
.Y(n_2487)
);

AO22x2_ASAP7_75t_L g2488 ( 
.A1(n_2360),
.A2(n_46),
.B1(n_44),
.B2(n_45),
.Y(n_2488)
);

AOI221xp5_ASAP7_75t_L g2489 ( 
.A1(n_2418),
.A2(n_889),
.B1(n_927),
.B2(n_854),
.C(n_846),
.Y(n_2489)
);

NOR3xp33_ASAP7_75t_L g2490 ( 
.A(n_2377),
.B(n_942),
.C(n_931),
.Y(n_2490)
);

AOI221xp5_ASAP7_75t_L g2491 ( 
.A1(n_2339),
.A2(n_1001),
.B1(n_995),
.B2(n_952),
.C(n_50),
.Y(n_2491)
);

NOR2xp33_ASAP7_75t_SL g2492 ( 
.A(n_2413),
.B(n_734),
.Y(n_2492)
);

OAI21xp33_ASAP7_75t_L g2493 ( 
.A1(n_2403),
.A2(n_1718),
.B(n_1717),
.Y(n_2493)
);

NOR2x1_ASAP7_75t_L g2494 ( 
.A(n_2365),
.B(n_48),
.Y(n_2494)
);

NAND2xp5_ASAP7_75t_L g2495 ( 
.A(n_2368),
.B(n_48),
.Y(n_2495)
);

NOR2xp67_ASAP7_75t_L g2496 ( 
.A(n_2372),
.B(n_49),
.Y(n_2496)
);

NAND3x1_ASAP7_75t_L g2497 ( 
.A(n_2338),
.B(n_49),
.C(n_51),
.Y(n_2497)
);

AO21x1_ASAP7_75t_L g2498 ( 
.A1(n_2430),
.A2(n_52),
.B(n_53),
.Y(n_2498)
);

OAI22xp5_ASAP7_75t_L g2499 ( 
.A1(n_2397),
.A2(n_56),
.B1(n_54),
.B2(n_55),
.Y(n_2499)
);

NOR3xp33_ASAP7_75t_L g2500 ( 
.A(n_2425),
.B(n_55),
.C(n_57),
.Y(n_2500)
);

OAI211xp5_ASAP7_75t_L g2501 ( 
.A1(n_2331),
.A2(n_59),
.B(n_57),
.C(n_58),
.Y(n_2501)
);

OAI22xp5_ASAP7_75t_L g2502 ( 
.A1(n_2326),
.A2(n_62),
.B1(n_59),
.B2(n_61),
.Y(n_2502)
);

AOI21xp5_ASAP7_75t_L g2503 ( 
.A1(n_2342),
.A2(n_61),
.B(n_62),
.Y(n_2503)
);

NAND2xp5_ASAP7_75t_L g2504 ( 
.A(n_2393),
.B(n_65),
.Y(n_2504)
);

OA22x2_ASAP7_75t_L g2505 ( 
.A1(n_2361),
.A2(n_1772),
.B1(n_68),
.B2(n_66),
.Y(n_2505)
);

AOI21xp5_ASAP7_75t_L g2506 ( 
.A1(n_2375),
.A2(n_67),
.B(n_68),
.Y(n_2506)
);

AOI221x1_ASAP7_75t_L g2507 ( 
.A1(n_2424),
.A2(n_2335),
.B1(n_2409),
.B2(n_2408),
.C(n_2407),
.Y(n_2507)
);

OAI211xp5_ASAP7_75t_L g2508 ( 
.A1(n_2405),
.A2(n_2415),
.B(n_2422),
.C(n_2419),
.Y(n_2508)
);

AOI221xp5_ASAP7_75t_L g2509 ( 
.A1(n_2411),
.A2(n_2400),
.B1(n_2369),
.B2(n_2395),
.C(n_2426),
.Y(n_2509)
);

AND2x2_ASAP7_75t_L g2510 ( 
.A(n_2326),
.B(n_67),
.Y(n_2510)
);

INVxp67_ASAP7_75t_L g2511 ( 
.A(n_2431),
.Y(n_2511)
);

OAI221xp5_ASAP7_75t_L g2512 ( 
.A1(n_2378),
.A2(n_71),
.B1(n_69),
.B2(n_70),
.C(n_72),
.Y(n_2512)
);

AOI221xp5_ASAP7_75t_L g2513 ( 
.A1(n_2381),
.A2(n_75),
.B1(n_69),
.B2(n_74),
.C(n_76),
.Y(n_2513)
);

NAND2xp5_ASAP7_75t_SL g2514 ( 
.A(n_2428),
.B(n_734),
.Y(n_2514)
);

AOI21xp5_ASAP7_75t_SL g2515 ( 
.A1(n_2396),
.A2(n_74),
.B(n_75),
.Y(n_2515)
);

AOI32xp33_ASAP7_75t_L g2516 ( 
.A1(n_2328),
.A2(n_79),
.A3(n_77),
.B1(n_78),
.B2(n_80),
.Y(n_2516)
);

NAND3xp33_ASAP7_75t_SL g2517 ( 
.A(n_2391),
.B(n_77),
.C(n_78),
.Y(n_2517)
);

NOR2x1_ASAP7_75t_L g2518 ( 
.A(n_2420),
.B(n_79),
.Y(n_2518)
);

OAI21xp33_ASAP7_75t_L g2519 ( 
.A1(n_2366),
.A2(n_2414),
.B(n_2391),
.Y(n_2519)
);

OR2x2_ASAP7_75t_L g2520 ( 
.A(n_2388),
.B(n_80),
.Y(n_2520)
);

AOI21xp33_ASAP7_75t_SL g2521 ( 
.A1(n_2401),
.A2(n_81),
.B(n_82),
.Y(n_2521)
);

O2A1O1Ixp33_ASAP7_75t_L g2522 ( 
.A1(n_2421),
.A2(n_85),
.B(n_83),
.C(n_84),
.Y(n_2522)
);

OAI21xp33_ASAP7_75t_L g2523 ( 
.A1(n_2417),
.A2(n_1715),
.B(n_1744),
.Y(n_2523)
);

OAI321xp33_ASAP7_75t_L g2524 ( 
.A1(n_2394),
.A2(n_85),
.A3(n_87),
.B1(n_83),
.B2(n_84),
.C(n_86),
.Y(n_2524)
);

NOR2xp67_ASAP7_75t_L g2525 ( 
.A(n_2417),
.B(n_87),
.Y(n_2525)
);

AOI21xp5_ASAP7_75t_L g2526 ( 
.A1(n_2349),
.A2(n_88),
.B(n_89),
.Y(n_2526)
);

OAI211xp5_ASAP7_75t_L g2527 ( 
.A1(n_2363),
.A2(n_95),
.B(n_90),
.C(n_94),
.Y(n_2527)
);

AOI221xp5_ASAP7_75t_L g2528 ( 
.A1(n_2429),
.A2(n_99),
.B1(n_96),
.B2(n_97),
.C(n_101),
.Y(n_2528)
);

INVx1_ASAP7_75t_L g2529 ( 
.A(n_2376),
.Y(n_2529)
);

INVx1_ASAP7_75t_L g2530 ( 
.A(n_2356),
.Y(n_2530)
);

NAND2xp5_ASAP7_75t_L g2531 ( 
.A(n_2386),
.B(n_96),
.Y(n_2531)
);

OAI221xp5_ASAP7_75t_L g2532 ( 
.A1(n_2438),
.A2(n_2347),
.B1(n_2423),
.B2(n_2345),
.C(n_2351),
.Y(n_2532)
);

AOI211xp5_ASAP7_75t_L g2533 ( 
.A1(n_2404),
.A2(n_101),
.B(n_97),
.C(n_99),
.Y(n_2533)
);

AOI221xp5_ASAP7_75t_L g2534 ( 
.A1(n_2410),
.A2(n_104),
.B1(n_102),
.B2(n_103),
.C(n_105),
.Y(n_2534)
);

O2A1O1Ixp5_ASAP7_75t_L g2535 ( 
.A1(n_2433),
.A2(n_105),
.B(n_103),
.C(n_104),
.Y(n_2535)
);

NAND4xp25_ASAP7_75t_L g2536 ( 
.A(n_2354),
.B(n_108),
.C(n_106),
.D(n_107),
.Y(n_2536)
);

AOI22xp5_ASAP7_75t_L g2537 ( 
.A1(n_2437),
.A2(n_1744),
.B1(n_734),
.B2(n_1726),
.Y(n_2537)
);

INVx1_ASAP7_75t_L g2538 ( 
.A(n_2321),
.Y(n_2538)
);

AOI322xp5_ASAP7_75t_L g2539 ( 
.A1(n_2324),
.A2(n_112),
.A3(n_111),
.B1(n_109),
.B2(n_107),
.C1(n_108),
.C2(n_110),
.Y(n_2539)
);

AOI322xp5_ASAP7_75t_L g2540 ( 
.A1(n_2324),
.A2(n_117),
.A3(n_116),
.B1(n_113),
.B2(n_109),
.C1(n_112),
.C2(n_114),
.Y(n_2540)
);

OAI21x1_ASAP7_75t_L g2541 ( 
.A1(n_2371),
.A2(n_1726),
.B(n_1715),
.Y(n_2541)
);

AOI22xp5_ASAP7_75t_L g2542 ( 
.A1(n_2435),
.A2(n_734),
.B1(n_119),
.B2(n_114),
.Y(n_2542)
);

INVx1_ASAP7_75t_L g2543 ( 
.A(n_2321),
.Y(n_2543)
);

AOI221xp5_ASAP7_75t_L g2544 ( 
.A1(n_2324),
.A2(n_121),
.B1(n_117),
.B2(n_119),
.C(n_122),
.Y(n_2544)
);

NAND2xp5_ASAP7_75t_SL g2545 ( 
.A(n_2373),
.B(n_734),
.Y(n_2545)
);

AOI211xp5_ASAP7_75t_L g2546 ( 
.A1(n_2324),
.A2(n_123),
.B(n_121),
.C(n_122),
.Y(n_2546)
);

NOR3xp33_ASAP7_75t_L g2547 ( 
.A(n_2412),
.B(n_125),
.C(n_126),
.Y(n_2547)
);

AOI221x1_ASAP7_75t_L g2548 ( 
.A1(n_2323),
.A2(n_129),
.B1(n_126),
.B2(n_127),
.C(n_130),
.Y(n_2548)
);

AOI221xp5_ASAP7_75t_L g2549 ( 
.A1(n_2324),
.A2(n_131),
.B1(n_129),
.B2(n_130),
.C(n_132),
.Y(n_2549)
);

AND2x2_ASAP7_75t_SL g2550 ( 
.A(n_2350),
.B(n_132),
.Y(n_2550)
);

NAND2xp5_ASAP7_75t_L g2551 ( 
.A(n_2355),
.B(n_133),
.Y(n_2551)
);

NAND2xp5_ASAP7_75t_L g2552 ( 
.A(n_2355),
.B(n_133),
.Y(n_2552)
);

AOI21xp5_ASAP7_75t_L g2553 ( 
.A1(n_2324),
.A2(n_134),
.B(n_135),
.Y(n_2553)
);

OA22x2_ASAP7_75t_L g2554 ( 
.A1(n_2323),
.A2(n_137),
.B1(n_135),
.B2(n_136),
.Y(n_2554)
);

HB1xp67_ASAP7_75t_L g2555 ( 
.A(n_2333),
.Y(n_2555)
);

OAI21xp5_ASAP7_75t_SL g2556 ( 
.A1(n_2323),
.A2(n_136),
.B(n_138),
.Y(n_2556)
);

AOI221xp5_ASAP7_75t_L g2557 ( 
.A1(n_2324),
.A2(n_142),
.B1(n_140),
.B2(n_141),
.C(n_143),
.Y(n_2557)
);

INVx1_ASAP7_75t_L g2558 ( 
.A(n_2321),
.Y(n_2558)
);

NAND3xp33_ASAP7_75t_SL g2559 ( 
.A(n_2390),
.B(n_142),
.C(n_143),
.Y(n_2559)
);

AOI211xp5_ASAP7_75t_L g2560 ( 
.A1(n_2324),
.A2(n_146),
.B(n_144),
.C(n_145),
.Y(n_2560)
);

INVx1_ASAP7_75t_L g2561 ( 
.A(n_2321),
.Y(n_2561)
);

AOI21xp5_ASAP7_75t_L g2562 ( 
.A1(n_2324),
.A2(n_144),
.B(n_147),
.Y(n_2562)
);

AOI22xp5_ASAP7_75t_L g2563 ( 
.A1(n_2435),
.A2(n_734),
.B1(n_151),
.B2(n_149),
.Y(n_2563)
);

AOI221xp5_ASAP7_75t_L g2564 ( 
.A1(n_2324),
.A2(n_151),
.B1(n_149),
.B2(n_150),
.C(n_152),
.Y(n_2564)
);

OAI211xp5_ASAP7_75t_SL g2565 ( 
.A1(n_2324),
.A2(n_154),
.B(n_152),
.C(n_153),
.Y(n_2565)
);

NOR3x1_ASAP7_75t_L g2566 ( 
.A(n_2334),
.B(n_153),
.C(n_154),
.Y(n_2566)
);

NOR2x1_ASAP7_75t_L g2567 ( 
.A(n_2333),
.B(n_155),
.Y(n_2567)
);

AOI221xp5_ASAP7_75t_L g2568 ( 
.A1(n_2324),
.A2(n_157),
.B1(n_155),
.B2(n_156),
.C(n_158),
.Y(n_2568)
);

OAI21xp33_ASAP7_75t_L g2569 ( 
.A1(n_2436),
.A2(n_156),
.B(n_158),
.Y(n_2569)
);

AOI322xp5_ASAP7_75t_L g2570 ( 
.A1(n_2324),
.A2(n_165),
.A3(n_164),
.B1(n_162),
.B2(n_159),
.C1(n_160),
.C2(n_163),
.Y(n_2570)
);

AOI222xp33_ASAP7_75t_L g2571 ( 
.A1(n_2324),
.A2(n_163),
.B1(n_166),
.B2(n_159),
.C1(n_160),
.C2(n_164),
.Y(n_2571)
);

NOR3xp33_ASAP7_75t_L g2572 ( 
.A(n_2412),
.B(n_166),
.C(n_168),
.Y(n_2572)
);

NAND2xp5_ASAP7_75t_SL g2573 ( 
.A(n_2373),
.B(n_734),
.Y(n_2573)
);

INVx1_ASAP7_75t_L g2574 ( 
.A(n_2321),
.Y(n_2574)
);

OAI221xp5_ASAP7_75t_L g2575 ( 
.A1(n_2324),
.A2(n_171),
.B1(n_169),
.B2(n_170),
.C(n_172),
.Y(n_2575)
);

AOI221xp5_ASAP7_75t_L g2576 ( 
.A1(n_2324),
.A2(n_171),
.B1(n_169),
.B2(n_170),
.C(n_172),
.Y(n_2576)
);

AOI221xp5_ASAP7_75t_L g2577 ( 
.A1(n_2324),
.A2(n_178),
.B1(n_174),
.B2(n_175),
.C(n_179),
.Y(n_2577)
);

INVx1_ASAP7_75t_L g2578 ( 
.A(n_2321),
.Y(n_2578)
);

NAND3xp33_ASAP7_75t_L g2579 ( 
.A(n_2324),
.B(n_174),
.C(n_178),
.Y(n_2579)
);

A2O1A1O1Ixp25_ASAP7_75t_L g2580 ( 
.A1(n_2384),
.A2(n_182),
.B(n_179),
.C(n_181),
.D(n_183),
.Y(n_2580)
);

AOI221xp5_ASAP7_75t_L g2581 ( 
.A1(n_2324),
.A2(n_184),
.B1(n_181),
.B2(n_183),
.C(n_185),
.Y(n_2581)
);

OAI21xp5_ASAP7_75t_L g2582 ( 
.A1(n_2324),
.A2(n_184),
.B(n_186),
.Y(n_2582)
);

AOI221xp5_ASAP7_75t_L g2583 ( 
.A1(n_2324),
.A2(n_189),
.B1(n_187),
.B2(n_188),
.C(n_190),
.Y(n_2583)
);

NAND2xp5_ASAP7_75t_SL g2584 ( 
.A(n_2373),
.B(n_734),
.Y(n_2584)
);

INVx2_ASAP7_75t_L g2585 ( 
.A(n_2364),
.Y(n_2585)
);

AOI322xp5_ASAP7_75t_L g2586 ( 
.A1(n_2324),
.A2(n_187),
.A3(n_188),
.B1(n_189),
.B2(n_190),
.C1(n_191),
.C2(n_192),
.Y(n_2586)
);

AOI221xp5_ASAP7_75t_L g2587 ( 
.A1(n_2324),
.A2(n_194),
.B1(n_192),
.B2(n_193),
.C(n_195),
.Y(n_2587)
);

NOR2xp33_ASAP7_75t_L g2588 ( 
.A(n_2373),
.B(n_193),
.Y(n_2588)
);

OAI221xp5_ASAP7_75t_SL g2589 ( 
.A1(n_2570),
.A2(n_196),
.B1(n_194),
.B2(n_195),
.C(n_197),
.Y(n_2589)
);

OAI22xp5_ASAP7_75t_L g2590 ( 
.A1(n_2579),
.A2(n_199),
.B1(n_196),
.B2(n_197),
.Y(n_2590)
);

AOI22xp5_ASAP7_75t_L g2591 ( 
.A1(n_2449),
.A2(n_2444),
.B1(n_2529),
.B2(n_2441),
.Y(n_2591)
);

AOI221xp5_ASAP7_75t_L g2592 ( 
.A1(n_2553),
.A2(n_201),
.B1(n_199),
.B2(n_200),
.C(n_202),
.Y(n_2592)
);

OAI21xp5_ASAP7_75t_L g2593 ( 
.A1(n_2580),
.A2(n_200),
.B(n_201),
.Y(n_2593)
);

AOI22xp5_ASAP7_75t_L g2594 ( 
.A1(n_2445),
.A2(n_734),
.B1(n_205),
.B2(n_203),
.Y(n_2594)
);

INVx1_ASAP7_75t_L g2595 ( 
.A(n_2488),
.Y(n_2595)
);

AOI22xp33_ASAP7_75t_L g2596 ( 
.A1(n_2518),
.A2(n_1126),
.B1(n_1119),
.B2(n_206),
.Y(n_2596)
);

OAI321xp33_ASAP7_75t_L g2597 ( 
.A1(n_2565),
.A2(n_207),
.A3(n_209),
.B1(n_204),
.B2(n_205),
.C(n_208),
.Y(n_2597)
);

OAI31xp33_ASAP7_75t_L g2598 ( 
.A1(n_2575),
.A2(n_211),
.A3(n_209),
.B(n_210),
.Y(n_2598)
);

AOI21xp5_ASAP7_75t_L g2599 ( 
.A1(n_2562),
.A2(n_212),
.B(n_213),
.Y(n_2599)
);

INVx2_ASAP7_75t_L g2600 ( 
.A(n_2550),
.Y(n_2600)
);

AOI322xp5_ASAP7_75t_L g2601 ( 
.A1(n_2519),
.A2(n_214),
.A3(n_215),
.B1(n_216),
.B2(n_217),
.C1(n_218),
.C2(n_219),
.Y(n_2601)
);

AOI21xp5_ASAP7_75t_L g2602 ( 
.A1(n_2582),
.A2(n_214),
.B(n_216),
.Y(n_2602)
);

AND2x2_ASAP7_75t_L g2603 ( 
.A(n_2555),
.B(n_217),
.Y(n_2603)
);

INVx2_ASAP7_75t_L g2604 ( 
.A(n_2566),
.Y(n_2604)
);

AOI22xp5_ASAP7_75t_L g2605 ( 
.A1(n_2538),
.A2(n_221),
.B1(n_219),
.B2(n_220),
.Y(n_2605)
);

O2A1O1Ixp33_ASAP7_75t_L g2606 ( 
.A1(n_2546),
.A2(n_223),
.B(n_220),
.C(n_222),
.Y(n_2606)
);

INVx1_ASAP7_75t_L g2607 ( 
.A(n_2488),
.Y(n_2607)
);

NAND2xp5_ASAP7_75t_SL g2608 ( 
.A(n_2571),
.B(n_222),
.Y(n_2608)
);

AOI22xp5_ASAP7_75t_L g2609 ( 
.A1(n_2543),
.A2(n_2558),
.B1(n_2574),
.B2(n_2561),
.Y(n_2609)
);

OAI321xp33_ASAP7_75t_L g2610 ( 
.A1(n_2560),
.A2(n_227),
.A3(n_229),
.B1(n_224),
.B2(n_226),
.C(n_228),
.Y(n_2610)
);

AOI211xp5_ASAP7_75t_L g2611 ( 
.A1(n_2464),
.A2(n_2549),
.B(n_2557),
.C(n_2544),
.Y(n_2611)
);

INVx1_ASAP7_75t_L g2612 ( 
.A(n_2554),
.Y(n_2612)
);

OAI221xp5_ASAP7_75t_L g2613 ( 
.A1(n_2564),
.A2(n_2577),
.B1(n_2581),
.B2(n_2576),
.C(n_2568),
.Y(n_2613)
);

OAI22xp33_ASAP7_75t_L g2614 ( 
.A1(n_2448),
.A2(n_229),
.B1(n_227),
.B2(n_228),
.Y(n_2614)
);

NAND2xp33_ASAP7_75t_SL g2615 ( 
.A(n_2466),
.B(n_231),
.Y(n_2615)
);

AOI21xp33_ASAP7_75t_L g2616 ( 
.A1(n_2459),
.A2(n_232),
.B(n_233),
.Y(n_2616)
);

NOR2xp33_ASAP7_75t_L g2617 ( 
.A(n_2473),
.B(n_232),
.Y(n_2617)
);

INVxp67_ASAP7_75t_SL g2618 ( 
.A(n_2567),
.Y(n_2618)
);

NOR2xp67_ASAP7_75t_L g2619 ( 
.A(n_2451),
.B(n_2556),
.Y(n_2619)
);

OAI222xp33_ASAP7_75t_L g2620 ( 
.A1(n_2585),
.A2(n_2505),
.B1(n_2476),
.B2(n_2494),
.C1(n_2440),
.C2(n_2511),
.Y(n_2620)
);

NOR2x1_ASAP7_75t_L g2621 ( 
.A(n_2478),
.B(n_234),
.Y(n_2621)
);

OAI21xp5_ASAP7_75t_SL g2622 ( 
.A1(n_2583),
.A2(n_235),
.B(n_236),
.Y(n_2622)
);

OAI21xp5_ASAP7_75t_L g2623 ( 
.A1(n_2570),
.A2(n_235),
.B(n_236),
.Y(n_2623)
);

NAND2x1_ASAP7_75t_L g2624 ( 
.A(n_2578),
.B(n_237),
.Y(n_2624)
);

XNOR2xp5_ASAP7_75t_L g2625 ( 
.A(n_2497),
.B(n_237),
.Y(n_2625)
);

AOI22xp5_ASAP7_75t_L g2626 ( 
.A1(n_2530),
.A2(n_240),
.B1(n_238),
.B2(n_239),
.Y(n_2626)
);

A2O1A1Ixp33_ASAP7_75t_SL g2627 ( 
.A1(n_2508),
.A2(n_241),
.B(n_238),
.C(n_240),
.Y(n_2627)
);

AOI21xp5_ASAP7_75t_L g2628 ( 
.A1(n_2587),
.A2(n_242),
.B(n_243),
.Y(n_2628)
);

INVxp67_ASAP7_75t_SL g2629 ( 
.A(n_2496),
.Y(n_2629)
);

AOI21xp33_ASAP7_75t_L g2630 ( 
.A1(n_2442),
.A2(n_2443),
.B(n_2471),
.Y(n_2630)
);

AOI21xp5_ASAP7_75t_L g2631 ( 
.A1(n_2461),
.A2(n_245),
.B(n_246),
.Y(n_2631)
);

O2A1O1Ixp5_ASAP7_75t_SL g2632 ( 
.A1(n_2475),
.A2(n_248),
.B(n_245),
.C(n_247),
.Y(n_2632)
);

AOI222xp33_ASAP7_75t_L g2633 ( 
.A1(n_2467),
.A2(n_2446),
.B1(n_2559),
.B2(n_2517),
.C1(n_2482),
.C2(n_2545),
.Y(n_2633)
);

AOI21xp33_ASAP7_75t_SL g2634 ( 
.A1(n_2457),
.A2(n_247),
.B(n_249),
.Y(n_2634)
);

OAI22xp5_ASAP7_75t_L g2635 ( 
.A1(n_2453),
.A2(n_252),
.B1(n_250),
.B2(n_251),
.Y(n_2635)
);

AOI221xp5_ASAP7_75t_L g2636 ( 
.A1(n_2532),
.A2(n_2447),
.B1(n_2480),
.B2(n_2535),
.C(n_2484),
.Y(n_2636)
);

OAI322xp33_ASAP7_75t_SL g2637 ( 
.A1(n_2573),
.A2(n_252),
.A3(n_253),
.B1(n_254),
.B2(n_255),
.C1(n_257),
.C2(n_258),
.Y(n_2637)
);

INVx1_ASAP7_75t_L g2638 ( 
.A(n_2498),
.Y(n_2638)
);

AOI22xp33_ASAP7_75t_SL g2639 ( 
.A1(n_2443),
.A2(n_259),
.B1(n_253),
.B2(n_257),
.Y(n_2639)
);

AOI21xp33_ASAP7_75t_SL g2640 ( 
.A1(n_2588),
.A2(n_260),
.B(n_261),
.Y(n_2640)
);

NOR2xp33_ASAP7_75t_L g2641 ( 
.A(n_2479),
.B(n_260),
.Y(n_2641)
);

AOI22xp5_ASAP7_75t_L g2642 ( 
.A1(n_2490),
.A2(n_264),
.B1(n_261),
.B2(n_262),
.Y(n_2642)
);

AOI22xp5_ASAP7_75t_L g2643 ( 
.A1(n_2547),
.A2(n_267),
.B1(n_265),
.B2(n_266),
.Y(n_2643)
);

AOI22xp5_ASAP7_75t_SL g2644 ( 
.A1(n_2452),
.A2(n_268),
.B1(n_265),
.B2(n_266),
.Y(n_2644)
);

INVx1_ASAP7_75t_L g2645 ( 
.A(n_2474),
.Y(n_2645)
);

AOI221xp5_ASAP7_75t_L g2646 ( 
.A1(n_2522),
.A2(n_270),
.B1(n_268),
.B2(n_269),
.C(n_271),
.Y(n_2646)
);

OAI21xp33_ASAP7_75t_L g2647 ( 
.A1(n_2539),
.A2(n_272),
.B(n_273),
.Y(n_2647)
);

NOR2xp33_ASAP7_75t_L g2648 ( 
.A(n_2524),
.B(n_272),
.Y(n_2648)
);

OAI211xp5_ASAP7_75t_L g2649 ( 
.A1(n_2540),
.A2(n_277),
.B(n_275),
.C(n_276),
.Y(n_2649)
);

OAI221xp5_ASAP7_75t_L g2650 ( 
.A1(n_2586),
.A2(n_280),
.B1(n_275),
.B2(n_276),
.C(n_281),
.Y(n_2650)
);

O2A1O1Ixp33_ASAP7_75t_L g2651 ( 
.A1(n_2569),
.A2(n_287),
.B(n_281),
.C(n_283),
.Y(n_2651)
);

OAI322xp33_ASAP7_75t_L g2652 ( 
.A1(n_2542),
.A2(n_287),
.A3(n_288),
.B1(n_289),
.B2(n_290),
.C1(n_292),
.C2(n_293),
.Y(n_2652)
);

AOI22xp5_ASAP7_75t_L g2653 ( 
.A1(n_2572),
.A2(n_294),
.B1(n_288),
.B2(n_293),
.Y(n_2653)
);

AOI21x1_ASAP7_75t_L g2654 ( 
.A1(n_2548),
.A2(n_294),
.B(n_295),
.Y(n_2654)
);

NAND3xp33_ASAP7_75t_L g2655 ( 
.A(n_2509),
.B(n_296),
.C(n_297),
.Y(n_2655)
);

OAI21xp5_ASAP7_75t_L g2656 ( 
.A1(n_2526),
.A2(n_296),
.B(n_298),
.Y(n_2656)
);

AOI22xp5_ASAP7_75t_L g2657 ( 
.A1(n_2551),
.A2(n_300),
.B1(n_298),
.B2(n_299),
.Y(n_2657)
);

OAI222xp33_ASAP7_75t_L g2658 ( 
.A1(n_2455),
.A2(n_299),
.B1(n_302),
.B2(n_303),
.C1(n_304),
.C2(n_306),
.Y(n_2658)
);

O2A1O1Ixp33_ASAP7_75t_SL g2659 ( 
.A1(n_2481),
.A2(n_308),
.B(n_304),
.C(n_307),
.Y(n_2659)
);

OAI211xp5_ASAP7_75t_SL g2660 ( 
.A1(n_2468),
.A2(n_310),
.B(n_308),
.C(n_309),
.Y(n_2660)
);

NOR2x1_ASAP7_75t_L g2661 ( 
.A(n_2495),
.B(n_311),
.Y(n_2661)
);

OAI211xp5_ASAP7_75t_L g2662 ( 
.A1(n_2507),
.A2(n_313),
.B(n_311),
.C(n_312),
.Y(n_2662)
);

INVx1_ASAP7_75t_L g2663 ( 
.A(n_2510),
.Y(n_2663)
);

AOI22xp5_ASAP7_75t_L g2664 ( 
.A1(n_2552),
.A2(n_2525),
.B1(n_2563),
.B2(n_2504),
.Y(n_2664)
);

OAI21xp33_ASAP7_75t_L g2665 ( 
.A1(n_2460),
.A2(n_312),
.B(n_313),
.Y(n_2665)
);

AOI22xp5_ASAP7_75t_L g2666 ( 
.A1(n_2469),
.A2(n_316),
.B1(n_314),
.B2(n_315),
.Y(n_2666)
);

INVx1_ASAP7_75t_L g2667 ( 
.A(n_2520),
.Y(n_2667)
);

AOI221xp5_ASAP7_75t_SL g2668 ( 
.A1(n_2584),
.A2(n_319),
.B1(n_317),
.B2(n_318),
.C(n_320),
.Y(n_2668)
);

AOI21xp5_ASAP7_75t_L g2669 ( 
.A1(n_2531),
.A2(n_317),
.B(n_318),
.Y(n_2669)
);

INVx1_ASAP7_75t_L g2670 ( 
.A(n_2536),
.Y(n_2670)
);

NAND2xp5_ASAP7_75t_L g2671 ( 
.A(n_2516),
.B(n_319),
.Y(n_2671)
);

INVx1_ASAP7_75t_L g2672 ( 
.A(n_2499),
.Y(n_2672)
);

AOI211xp5_ASAP7_75t_SL g2673 ( 
.A1(n_2515),
.A2(n_322),
.B(n_320),
.C(n_321),
.Y(n_2673)
);

AOI21xp5_ASAP7_75t_L g2674 ( 
.A1(n_2506),
.A2(n_321),
.B(n_322),
.Y(n_2674)
);

INVxp67_ASAP7_75t_L g2675 ( 
.A(n_2456),
.Y(n_2675)
);

OAI21xp33_ASAP7_75t_L g2676 ( 
.A1(n_2477),
.A2(n_323),
.B(n_325),
.Y(n_2676)
);

AOI21xp5_ASAP7_75t_L g2677 ( 
.A1(n_2627),
.A2(n_2503),
.B(n_2527),
.Y(n_2677)
);

NAND2xp5_ASAP7_75t_L g2678 ( 
.A(n_2618),
.B(n_2521),
.Y(n_2678)
);

INVx1_ASAP7_75t_L g2679 ( 
.A(n_2603),
.Y(n_2679)
);

INVx1_ASAP7_75t_L g2680 ( 
.A(n_2625),
.Y(n_2680)
);

INVx1_ASAP7_75t_L g2681 ( 
.A(n_2654),
.Y(n_2681)
);

AOI211xp5_ASAP7_75t_SL g2682 ( 
.A1(n_2614),
.A2(n_2470),
.B(n_2450),
.C(n_2491),
.Y(n_2682)
);

OAI221xp5_ASAP7_75t_L g2683 ( 
.A1(n_2624),
.A2(n_2537),
.B1(n_2500),
.B2(n_2462),
.C(n_2501),
.Y(n_2683)
);

NOR3xp33_ASAP7_75t_L g2684 ( 
.A(n_2630),
.B(n_2514),
.C(n_2454),
.Y(n_2684)
);

NOR3x1_ASAP7_75t_L g2685 ( 
.A(n_2623),
.B(n_2512),
.C(n_2502),
.Y(n_2685)
);

INVx2_ASAP7_75t_L g2686 ( 
.A(n_2604),
.Y(n_2686)
);

AOI221xp5_ASAP7_75t_L g2687 ( 
.A1(n_2616),
.A2(n_2485),
.B1(n_2483),
.B2(n_2492),
.C(n_2534),
.Y(n_2687)
);

O2A1O1Ixp33_ASAP7_75t_L g2688 ( 
.A1(n_2638),
.A2(n_2472),
.B(n_2533),
.C(n_2513),
.Y(n_2688)
);

AOI322xp5_ASAP7_75t_L g2689 ( 
.A1(n_2612),
.A2(n_2528),
.A3(n_2465),
.B1(n_2458),
.B2(n_2493),
.C1(n_2523),
.C2(n_2489),
.Y(n_2689)
);

INVx1_ASAP7_75t_L g2690 ( 
.A(n_2661),
.Y(n_2690)
);

AOI222xp33_ASAP7_75t_L g2691 ( 
.A1(n_2595),
.A2(n_2486),
.B1(n_2487),
.B2(n_2463),
.C1(n_2541),
.C2(n_328),
.Y(n_2691)
);

INVx1_ASAP7_75t_L g2692 ( 
.A(n_2629),
.Y(n_2692)
);

AOI211xp5_ASAP7_75t_L g2693 ( 
.A1(n_2619),
.A2(n_2620),
.B(n_2613),
.C(n_2665),
.Y(n_2693)
);

OAI21xp5_ASAP7_75t_SL g2694 ( 
.A1(n_2658),
.A2(n_323),
.B(n_325),
.Y(n_2694)
);

NAND2xp5_ASAP7_75t_L g2695 ( 
.A(n_2673),
.B(n_326),
.Y(n_2695)
);

NAND2xp5_ASAP7_75t_L g2696 ( 
.A(n_2644),
.B(n_326),
.Y(n_2696)
);

AOI22xp5_ASAP7_75t_L g2697 ( 
.A1(n_2647),
.A2(n_329),
.B1(n_327),
.B2(n_328),
.Y(n_2697)
);

INVx1_ASAP7_75t_L g2698 ( 
.A(n_2607),
.Y(n_2698)
);

AOI211xp5_ASAP7_75t_L g2699 ( 
.A1(n_2662),
.A2(n_330),
.B(n_327),
.C(n_329),
.Y(n_2699)
);

INVx1_ASAP7_75t_L g2700 ( 
.A(n_2621),
.Y(n_2700)
);

INVx2_ASAP7_75t_L g2701 ( 
.A(n_2600),
.Y(n_2701)
);

AOI22xp5_ASAP7_75t_L g2702 ( 
.A1(n_2608),
.A2(n_333),
.B1(n_331),
.B2(n_332),
.Y(n_2702)
);

NAND2xp5_ASAP7_75t_L g2703 ( 
.A(n_2639),
.B(n_2668),
.Y(n_2703)
);

A2O1A1Ixp33_ASAP7_75t_L g2704 ( 
.A1(n_2602),
.A2(n_338),
.B(n_334),
.C(n_336),
.Y(n_2704)
);

AOI21xp5_ASAP7_75t_L g2705 ( 
.A1(n_2593),
.A2(n_334),
.B(n_336),
.Y(n_2705)
);

AOI211xp5_ASAP7_75t_L g2706 ( 
.A1(n_2617),
.A2(n_341),
.B(n_338),
.C(n_340),
.Y(n_2706)
);

NAND2xp5_ASAP7_75t_L g2707 ( 
.A(n_2668),
.B(n_340),
.Y(n_2707)
);

AOI22xp5_ASAP7_75t_L g2708 ( 
.A1(n_2645),
.A2(n_343),
.B1(n_341),
.B2(n_342),
.Y(n_2708)
);

INVx1_ASAP7_75t_L g2709 ( 
.A(n_2659),
.Y(n_2709)
);

OAI221xp5_ASAP7_75t_L g2710 ( 
.A1(n_2591),
.A2(n_344),
.B1(n_345),
.B2(n_346),
.C(n_347),
.Y(n_2710)
);

AOI22xp5_ASAP7_75t_L g2711 ( 
.A1(n_2615),
.A2(n_350),
.B1(n_344),
.B2(n_348),
.Y(n_2711)
);

OAI221xp5_ASAP7_75t_L g2712 ( 
.A1(n_2611),
.A2(n_348),
.B1(n_351),
.B2(n_352),
.C(n_353),
.Y(n_2712)
);

INVx1_ASAP7_75t_L g2713 ( 
.A(n_2667),
.Y(n_2713)
);

OAI211xp5_ASAP7_75t_L g2714 ( 
.A1(n_2609),
.A2(n_355),
.B(n_352),
.C(n_354),
.Y(n_2714)
);

AOI22xp5_ASAP7_75t_L g2715 ( 
.A1(n_2670),
.A2(n_2648),
.B1(n_2664),
.B2(n_2649),
.Y(n_2715)
);

AND2x2_ASAP7_75t_L g2716 ( 
.A(n_2656),
.B(n_354),
.Y(n_2716)
);

AOI221xp5_ASAP7_75t_L g2717 ( 
.A1(n_2596),
.A2(n_357),
.B1(n_358),
.B2(n_359),
.C(n_361),
.Y(n_2717)
);

NOR2xp33_ASAP7_75t_L g2718 ( 
.A(n_2597),
.B(n_357),
.Y(n_2718)
);

INVx2_ASAP7_75t_L g2719 ( 
.A(n_2663),
.Y(n_2719)
);

BUFx2_ASAP7_75t_L g2720 ( 
.A(n_2671),
.Y(n_2720)
);

INVx1_ASAP7_75t_L g2721 ( 
.A(n_2641),
.Y(n_2721)
);

INVx2_ASAP7_75t_L g2722 ( 
.A(n_2675),
.Y(n_2722)
);

INVx2_ASAP7_75t_L g2723 ( 
.A(n_2672),
.Y(n_2723)
);

A2O1A1Ixp33_ASAP7_75t_SL g2724 ( 
.A1(n_2594),
.A2(n_361),
.B(n_358),
.C(n_359),
.Y(n_2724)
);

AOI21xp5_ASAP7_75t_L g2725 ( 
.A1(n_2637),
.A2(n_362),
.B(n_363),
.Y(n_2725)
);

AOI22xp5_ASAP7_75t_L g2726 ( 
.A1(n_2590),
.A2(n_365),
.B1(n_362),
.B2(n_364),
.Y(n_2726)
);

HB1xp67_ASAP7_75t_L g2727 ( 
.A(n_2635),
.Y(n_2727)
);

OAI22xp5_ASAP7_75t_L g2728 ( 
.A1(n_2589),
.A2(n_366),
.B1(n_364),
.B2(n_365),
.Y(n_2728)
);

OAI21xp5_ASAP7_75t_L g2729 ( 
.A1(n_2655),
.A2(n_366),
.B(n_367),
.Y(n_2729)
);

NAND5xp2_ASAP7_75t_L g2730 ( 
.A(n_2633),
.B(n_367),
.C(n_368),
.D(n_369),
.E(n_371),
.Y(n_2730)
);

INVx1_ASAP7_75t_L g2731 ( 
.A(n_2643),
.Y(n_2731)
);

NAND3xp33_ASAP7_75t_L g2732 ( 
.A(n_2636),
.B(n_368),
.C(n_369),
.Y(n_2732)
);

INVx2_ASAP7_75t_L g2733 ( 
.A(n_2653),
.Y(n_2733)
);

INVx1_ASAP7_75t_L g2734 ( 
.A(n_2657),
.Y(n_2734)
);

INVxp67_ASAP7_75t_L g2735 ( 
.A(n_2730),
.Y(n_2735)
);

INVx1_ASAP7_75t_L g2736 ( 
.A(n_2681),
.Y(n_2736)
);

CKINVDCx5p33_ASAP7_75t_R g2737 ( 
.A(n_2701),
.Y(n_2737)
);

AOI211xp5_ASAP7_75t_L g2738 ( 
.A1(n_2692),
.A2(n_2622),
.B(n_2650),
.C(n_2640),
.Y(n_2738)
);

NOR3xp33_ASAP7_75t_L g2739 ( 
.A(n_2680),
.B(n_2610),
.C(n_2634),
.Y(n_2739)
);

AOI21xp5_ASAP7_75t_L g2740 ( 
.A1(n_2725),
.A2(n_2705),
.B(n_2677),
.Y(n_2740)
);

INVx1_ASAP7_75t_L g2741 ( 
.A(n_2690),
.Y(n_2741)
);

NOR2x1p5_ASAP7_75t_L g2742 ( 
.A(n_2719),
.B(n_2598),
.Y(n_2742)
);

NOR2x1_ASAP7_75t_L g2743 ( 
.A(n_2713),
.B(n_2652),
.Y(n_2743)
);

AOI221xp5_ASAP7_75t_L g2744 ( 
.A1(n_2698),
.A2(n_2676),
.B1(n_2669),
.B2(n_2651),
.C(n_2628),
.Y(n_2744)
);

INVx1_ASAP7_75t_L g2745 ( 
.A(n_2695),
.Y(n_2745)
);

O2A1O1Ixp33_ASAP7_75t_L g2746 ( 
.A1(n_2693),
.A2(n_2606),
.B(n_2597),
.C(n_2631),
.Y(n_2746)
);

OAI22xp33_ASAP7_75t_R g2747 ( 
.A1(n_2686),
.A2(n_2660),
.B1(n_2599),
.B2(n_2646),
.Y(n_2747)
);

AOI21xp5_ASAP7_75t_L g2748 ( 
.A1(n_2703),
.A2(n_2592),
.B(n_2674),
.Y(n_2748)
);

INVx1_ASAP7_75t_L g2749 ( 
.A(n_2709),
.Y(n_2749)
);

INVx1_ASAP7_75t_SL g2750 ( 
.A(n_2696),
.Y(n_2750)
);

OAI21xp33_ASAP7_75t_L g2751 ( 
.A1(n_2715),
.A2(n_2601),
.B(n_2642),
.Y(n_2751)
);

OR2x2_ASAP7_75t_L g2752 ( 
.A(n_2707),
.B(n_2605),
.Y(n_2752)
);

OAI21xp5_ASAP7_75t_L g2753 ( 
.A1(n_2732),
.A2(n_2632),
.B(n_2666),
.Y(n_2753)
);

HB1xp67_ASAP7_75t_L g2754 ( 
.A(n_2700),
.Y(n_2754)
);

AOI22xp5_ASAP7_75t_L g2755 ( 
.A1(n_2679),
.A2(n_2691),
.B1(n_2716),
.B2(n_2678),
.Y(n_2755)
);

INVx1_ASAP7_75t_L g2756 ( 
.A(n_2727),
.Y(n_2756)
);

NAND2xp5_ASAP7_75t_L g2757 ( 
.A(n_2699),
.B(n_2626),
.Y(n_2757)
);

INVxp67_ASAP7_75t_SL g2758 ( 
.A(n_2718),
.Y(n_2758)
);

AOI22xp5_ASAP7_75t_L g2759 ( 
.A1(n_2694),
.A2(n_374),
.B1(n_372),
.B2(n_373),
.Y(n_2759)
);

AOI21xp5_ASAP7_75t_L g2760 ( 
.A1(n_2714),
.A2(n_372),
.B(n_374),
.Y(n_2760)
);

AOI221xp5_ASAP7_75t_SL g2761 ( 
.A1(n_2688),
.A2(n_375),
.B1(n_377),
.B2(n_379),
.C(n_380),
.Y(n_2761)
);

AOI22xp33_ASAP7_75t_L g2762 ( 
.A1(n_2720),
.A2(n_1126),
.B1(n_1119),
.B2(n_1139),
.Y(n_2762)
);

OAI221xp5_ASAP7_75t_L g2763 ( 
.A1(n_2706),
.A2(n_375),
.B1(n_377),
.B2(n_381),
.C(n_382),
.Y(n_2763)
);

AOI21xp5_ASAP7_75t_L g2764 ( 
.A1(n_2712),
.A2(n_382),
.B(n_383),
.Y(n_2764)
);

AOI221xp5_ASAP7_75t_L g2765 ( 
.A1(n_2728),
.A2(n_383),
.B1(n_384),
.B2(n_385),
.C(n_386),
.Y(n_2765)
);

INVxp67_ASAP7_75t_L g2766 ( 
.A(n_2723),
.Y(n_2766)
);

OA22x2_ASAP7_75t_L g2767 ( 
.A1(n_2697),
.A2(n_388),
.B1(n_385),
.B2(n_387),
.Y(n_2767)
);

OAI21xp5_ASAP7_75t_L g2768 ( 
.A1(n_2704),
.A2(n_389),
.B(n_390),
.Y(n_2768)
);

INVx1_ASAP7_75t_L g2769 ( 
.A(n_2699),
.Y(n_2769)
);

AOI22xp33_ASAP7_75t_L g2770 ( 
.A1(n_2733),
.A2(n_1126),
.B1(n_1119),
.B2(n_1139),
.Y(n_2770)
);

NOR2x1_ASAP7_75t_L g2771 ( 
.A(n_2736),
.B(n_2722),
.Y(n_2771)
);

INVxp33_ASAP7_75t_L g2772 ( 
.A(n_2754),
.Y(n_2772)
);

INVxp33_ASAP7_75t_L g2773 ( 
.A(n_2743),
.Y(n_2773)
);

INVx1_ASAP7_75t_L g2774 ( 
.A(n_2737),
.Y(n_2774)
);

NOR2x1_ASAP7_75t_L g2775 ( 
.A(n_2749),
.B(n_2710),
.Y(n_2775)
);

AND2x2_ASAP7_75t_SL g2776 ( 
.A(n_2756),
.B(n_2685),
.Y(n_2776)
);

INVx1_ASAP7_75t_SL g2777 ( 
.A(n_2752),
.Y(n_2777)
);

INVx1_ASAP7_75t_L g2778 ( 
.A(n_2767),
.Y(n_2778)
);

INVx1_ASAP7_75t_L g2779 ( 
.A(n_2767),
.Y(n_2779)
);

AOI22xp5_ASAP7_75t_L g2780 ( 
.A1(n_2745),
.A2(n_2702),
.B1(n_2721),
.B2(n_2711),
.Y(n_2780)
);

NOR2x1_ASAP7_75t_L g2781 ( 
.A(n_2741),
.B(n_2729),
.Y(n_2781)
);

INVx1_ASAP7_75t_L g2782 ( 
.A(n_2766),
.Y(n_2782)
);

INVx1_ASAP7_75t_L g2783 ( 
.A(n_2735),
.Y(n_2783)
);

NOR2x1_ASAP7_75t_L g2784 ( 
.A(n_2740),
.B(n_2731),
.Y(n_2784)
);

OAI22x1_ASAP7_75t_L g2785 ( 
.A1(n_2759),
.A2(n_2726),
.B1(n_2708),
.B2(n_2734),
.Y(n_2785)
);

AOI22xp5_ASAP7_75t_L g2786 ( 
.A1(n_2758),
.A2(n_2706),
.B1(n_2717),
.B2(n_2684),
.Y(n_2786)
);

INVx1_ASAP7_75t_L g2787 ( 
.A(n_2742),
.Y(n_2787)
);

NOR2x1_ASAP7_75t_L g2788 ( 
.A(n_2763),
.B(n_2683),
.Y(n_2788)
);

AO22x2_ASAP7_75t_L g2789 ( 
.A1(n_2769),
.A2(n_2750),
.B1(n_2739),
.B2(n_2748),
.Y(n_2789)
);

NOR2x1_ASAP7_75t_L g2790 ( 
.A(n_2746),
.B(n_2724),
.Y(n_2790)
);

AND2x4_ASAP7_75t_L g2791 ( 
.A(n_2771),
.B(n_2774),
.Y(n_2791)
);

AOI22xp33_ASAP7_75t_SL g2792 ( 
.A1(n_2778),
.A2(n_2757),
.B1(n_2753),
.B2(n_2768),
.Y(n_2792)
);

NAND2xp5_ASAP7_75t_L g2793 ( 
.A(n_2779),
.B(n_2761),
.Y(n_2793)
);

INVx1_ASAP7_75t_L g2794 ( 
.A(n_2789),
.Y(n_2794)
);

NAND2x1p5_ASAP7_75t_SL g2795 ( 
.A(n_2784),
.B(n_2781),
.Y(n_2795)
);

XNOR2xp5_ASAP7_75t_L g2796 ( 
.A(n_2773),
.B(n_2755),
.Y(n_2796)
);

NAND2x1p5_ASAP7_75t_SL g2797 ( 
.A(n_2790),
.B(n_2747),
.Y(n_2797)
);

NAND2x1p5_ASAP7_75t_L g2798 ( 
.A(n_2776),
.B(n_2760),
.Y(n_2798)
);

AND3x4_ASAP7_75t_L g2799 ( 
.A(n_2775),
.B(n_2738),
.C(n_2751),
.Y(n_2799)
);

INVx1_ASAP7_75t_L g2800 ( 
.A(n_2789),
.Y(n_2800)
);

NAND2x1p5_ASAP7_75t_L g2801 ( 
.A(n_2782),
.B(n_2764),
.Y(n_2801)
);

AO22x2_ASAP7_75t_L g2802 ( 
.A1(n_2777),
.A2(n_2744),
.B1(n_2682),
.B2(n_2765),
.Y(n_2802)
);

HB1xp67_ASAP7_75t_L g2803 ( 
.A(n_2787),
.Y(n_2803)
);

NOR2x1_ASAP7_75t_L g2804 ( 
.A(n_2783),
.B(n_2689),
.Y(n_2804)
);

NOR2x1_ASAP7_75t_L g2805 ( 
.A(n_2788),
.B(n_2689),
.Y(n_2805)
);

INVx1_ASAP7_75t_L g2806 ( 
.A(n_2772),
.Y(n_2806)
);

NOR2xp33_ASAP7_75t_L g2807 ( 
.A(n_2786),
.B(n_2687),
.Y(n_2807)
);

AOI211xp5_ASAP7_75t_L g2808 ( 
.A1(n_2794),
.A2(n_2780),
.B(n_2785),
.C(n_2762),
.Y(n_2808)
);

AOI22xp33_ASAP7_75t_L g2809 ( 
.A1(n_2803),
.A2(n_2770),
.B1(n_1126),
.B2(n_1119),
.Y(n_2809)
);

OAI221xp5_ASAP7_75t_L g2810 ( 
.A1(n_2800),
.A2(n_390),
.B1(n_391),
.B2(n_392),
.C(n_393),
.Y(n_2810)
);

AO22x2_ASAP7_75t_L g2811 ( 
.A1(n_2799),
.A2(n_395),
.B1(n_392),
.B2(n_393),
.Y(n_2811)
);

NAND3xp33_ASAP7_75t_L g2812 ( 
.A(n_2805),
.B(n_395),
.C(n_399),
.Y(n_2812)
);

NOR3x2_ASAP7_75t_L g2813 ( 
.A(n_2795),
.B(n_399),
.C(n_400),
.Y(n_2813)
);

OAI22xp5_ASAP7_75t_L g2814 ( 
.A1(n_2806),
.A2(n_403),
.B1(n_401),
.B2(n_402),
.Y(n_2814)
);

CKINVDCx16_ASAP7_75t_R g2815 ( 
.A(n_2804),
.Y(n_2815)
);

INVx1_ASAP7_75t_L g2816 ( 
.A(n_2791),
.Y(n_2816)
);

OAI21xp33_ASAP7_75t_SL g2817 ( 
.A1(n_2793),
.A2(n_404),
.B(n_405),
.Y(n_2817)
);

OR2x2_ASAP7_75t_L g2818 ( 
.A(n_2797),
.B(n_2798),
.Y(n_2818)
);

NAND2xp5_ASAP7_75t_L g2819 ( 
.A(n_2796),
.B(n_404),
.Y(n_2819)
);

NOR2x1_ASAP7_75t_L g2820 ( 
.A(n_2807),
.B(n_406),
.Y(n_2820)
);

AND4x1_ASAP7_75t_L g2821 ( 
.A(n_2792),
.B(n_406),
.C(n_408),
.D(n_409),
.Y(n_2821)
);

OAI211xp5_ASAP7_75t_SL g2822 ( 
.A1(n_2802),
.A2(n_408),
.B(n_409),
.C(n_410),
.Y(n_2822)
);

OR2x2_ASAP7_75t_L g2823 ( 
.A(n_2801),
.B(n_412),
.Y(n_2823)
);

AOI322xp5_ASAP7_75t_L g2824 ( 
.A1(n_2804),
.A2(n_414),
.A3(n_415),
.B1(n_416),
.B2(n_417),
.C1(n_418),
.C2(n_419),
.Y(n_2824)
);

NAND3xp33_ASAP7_75t_L g2825 ( 
.A(n_2805),
.B(n_414),
.C(n_415),
.Y(n_2825)
);

NOR3xp33_ASAP7_75t_L g2826 ( 
.A(n_2794),
.B(n_416),
.C(n_417),
.Y(n_2826)
);

NAND2x1_ASAP7_75t_L g2827 ( 
.A(n_2816),
.B(n_420),
.Y(n_2827)
);

INVx1_ASAP7_75t_L g2828 ( 
.A(n_2811),
.Y(n_2828)
);

INVx2_ASAP7_75t_L g2829 ( 
.A(n_2811),
.Y(n_2829)
);

INVx1_ASAP7_75t_L g2830 ( 
.A(n_2815),
.Y(n_2830)
);

AND2x2_ASAP7_75t_L g2831 ( 
.A(n_2818),
.B(n_421),
.Y(n_2831)
);

INVx1_ASAP7_75t_L g2832 ( 
.A(n_2820),
.Y(n_2832)
);

XNOR2x1_ASAP7_75t_L g2833 ( 
.A(n_2823),
.B(n_422),
.Y(n_2833)
);

XNOR2x1_ASAP7_75t_L g2834 ( 
.A(n_2819),
.B(n_423),
.Y(n_2834)
);

NOR2xp67_ASAP7_75t_L g2835 ( 
.A(n_2812),
.B(n_423),
.Y(n_2835)
);

NOR3xp33_ASAP7_75t_L g2836 ( 
.A(n_2825),
.B(n_424),
.C(n_426),
.Y(n_2836)
);

NAND3xp33_ASAP7_75t_L g2837 ( 
.A(n_2824),
.B(n_424),
.C(n_426),
.Y(n_2837)
);

AND2x2_ASAP7_75t_SL g2838 ( 
.A(n_2821),
.B(n_427),
.Y(n_2838)
);

NAND2xp5_ASAP7_75t_L g2839 ( 
.A(n_2817),
.B(n_428),
.Y(n_2839)
);

OAI22xp5_ASAP7_75t_SL g2840 ( 
.A1(n_2810),
.A2(n_428),
.B1(n_431),
.B2(n_433),
.Y(n_2840)
);

AO22x1_ASAP7_75t_L g2841 ( 
.A1(n_2826),
.A2(n_431),
.B1(n_433),
.B2(n_434),
.Y(n_2841)
);

AOI21xp5_ASAP7_75t_L g2842 ( 
.A1(n_2814),
.A2(n_435),
.B(n_436),
.Y(n_2842)
);

INVx1_ASAP7_75t_L g2843 ( 
.A(n_2813),
.Y(n_2843)
);

INVx3_ASAP7_75t_L g2844 ( 
.A(n_2822),
.Y(n_2844)
);

INVx4_ASAP7_75t_L g2845 ( 
.A(n_2808),
.Y(n_2845)
);

NOR4xp75_ASAP7_75t_SL g2846 ( 
.A(n_2809),
.B(n_435),
.C(n_436),
.D(n_437),
.Y(n_2846)
);

XOR2x1_ASAP7_75t_L g2847 ( 
.A(n_2818),
.B(n_437),
.Y(n_2847)
);

AO22x2_ASAP7_75t_L g2848 ( 
.A1(n_2830),
.A2(n_2828),
.B1(n_2827),
.B2(n_2829),
.Y(n_2848)
);

INVx2_ASAP7_75t_L g2849 ( 
.A(n_2847),
.Y(n_2849)
);

INVxp67_ASAP7_75t_SL g2850 ( 
.A(n_2827),
.Y(n_2850)
);

INVx1_ASAP7_75t_L g2851 ( 
.A(n_2838),
.Y(n_2851)
);

INVx1_ASAP7_75t_SL g2852 ( 
.A(n_2831),
.Y(n_2852)
);

INVx2_ASAP7_75t_L g2853 ( 
.A(n_2833),
.Y(n_2853)
);

INVx2_ASAP7_75t_L g2854 ( 
.A(n_2845),
.Y(n_2854)
);

NAND2xp5_ASAP7_75t_L g2855 ( 
.A(n_2832),
.B(n_2843),
.Y(n_2855)
);

INVx2_ASAP7_75t_L g2856 ( 
.A(n_2834),
.Y(n_2856)
);

INVx1_ASAP7_75t_SL g2857 ( 
.A(n_2839),
.Y(n_2857)
);

INVx2_ASAP7_75t_L g2858 ( 
.A(n_2844),
.Y(n_2858)
);

AOI22xp5_ASAP7_75t_L g2859 ( 
.A1(n_2836),
.A2(n_438),
.B1(n_439),
.B2(n_442),
.Y(n_2859)
);

INVx2_ASAP7_75t_L g2860 ( 
.A(n_2841),
.Y(n_2860)
);

XOR2xp5_ASAP7_75t_L g2861 ( 
.A(n_2837),
.B(n_438),
.Y(n_2861)
);

INVx2_ASAP7_75t_L g2862 ( 
.A(n_2840),
.Y(n_2862)
);

NAND2xp5_ASAP7_75t_L g2863 ( 
.A(n_2850),
.B(n_2835),
.Y(n_2863)
);

OAI22xp5_ASAP7_75t_L g2864 ( 
.A1(n_2854),
.A2(n_2842),
.B1(n_2846),
.B2(n_444),
.Y(n_2864)
);

INVx1_ASAP7_75t_L g2865 ( 
.A(n_2848),
.Y(n_2865)
);

XNOR2x1_ASAP7_75t_L g2866 ( 
.A(n_2848),
.B(n_442),
.Y(n_2866)
);

AND2x2_ASAP7_75t_SL g2867 ( 
.A(n_2849),
.B(n_443),
.Y(n_2867)
);

NOR2x1_ASAP7_75t_L g2868 ( 
.A(n_2855),
.B(n_443),
.Y(n_2868)
);

INVx1_ASAP7_75t_L g2869 ( 
.A(n_2851),
.Y(n_2869)
);

NOR4xp25_ASAP7_75t_SL g2870 ( 
.A(n_2861),
.B(n_444),
.C(n_445),
.D(n_446),
.Y(n_2870)
);

CKINVDCx16_ASAP7_75t_R g2871 ( 
.A(n_2852),
.Y(n_2871)
);

INVx1_ASAP7_75t_L g2872 ( 
.A(n_2860),
.Y(n_2872)
);

AOI21xp33_ASAP7_75t_SL g2873 ( 
.A1(n_2858),
.A2(n_447),
.B(n_448),
.Y(n_2873)
);

NAND2xp5_ASAP7_75t_L g2874 ( 
.A(n_2857),
.B(n_450),
.Y(n_2874)
);

AOI22xp5_ASAP7_75t_L g2875 ( 
.A1(n_2853),
.A2(n_451),
.B1(n_452),
.B2(n_453),
.Y(n_2875)
);

XNOR2x2_ASAP7_75t_SL g2876 ( 
.A(n_2859),
.B(n_452),
.Y(n_2876)
);

XNOR2xp5_ASAP7_75t_L g2877 ( 
.A(n_2866),
.B(n_2856),
.Y(n_2877)
);

OAI22xp5_ASAP7_75t_L g2878 ( 
.A1(n_2871),
.A2(n_2862),
.B1(n_455),
.B2(n_456),
.Y(n_2878)
);

AOI22xp5_ASAP7_75t_L g2879 ( 
.A1(n_2865),
.A2(n_454),
.B1(n_455),
.B2(n_457),
.Y(n_2879)
);

NAND2xp5_ASAP7_75t_SL g2880 ( 
.A(n_2867),
.B(n_454),
.Y(n_2880)
);

HB1xp67_ASAP7_75t_L g2881 ( 
.A(n_2868),
.Y(n_2881)
);

OR2x2_ASAP7_75t_L g2882 ( 
.A(n_2863),
.B(n_457),
.Y(n_2882)
);

AO21x2_ASAP7_75t_L g2883 ( 
.A1(n_2872),
.A2(n_458),
.B(n_459),
.Y(n_2883)
);

OAI21x1_ASAP7_75t_L g2884 ( 
.A1(n_2864),
.A2(n_458),
.B(n_460),
.Y(n_2884)
);

INVx1_ASAP7_75t_L g2885 ( 
.A(n_2874),
.Y(n_2885)
);

INVx1_ASAP7_75t_L g2886 ( 
.A(n_2869),
.Y(n_2886)
);

INVx1_ASAP7_75t_L g2887 ( 
.A(n_2876),
.Y(n_2887)
);

OAI211xp5_ASAP7_75t_L g2888 ( 
.A1(n_2873),
.A2(n_460),
.B(n_462),
.C(n_463),
.Y(n_2888)
);

OAI22x1_ASAP7_75t_L g2889 ( 
.A1(n_2875),
.A2(n_465),
.B1(n_467),
.B2(n_468),
.Y(n_2889)
);

AO22x2_ASAP7_75t_L g2890 ( 
.A1(n_2870),
.A2(n_465),
.B1(n_467),
.B2(n_468),
.Y(n_2890)
);

OAI22xp5_ASAP7_75t_L g2891 ( 
.A1(n_2871),
.A2(n_470),
.B1(n_471),
.B2(n_473),
.Y(n_2891)
);

AOI22xp5_ASAP7_75t_L g2892 ( 
.A1(n_2886),
.A2(n_2887),
.B1(n_2877),
.B2(n_2878),
.Y(n_2892)
);

INVxp67_ASAP7_75t_SL g2893 ( 
.A(n_2881),
.Y(n_2893)
);

INVx5_ASAP7_75t_L g2894 ( 
.A(n_2884),
.Y(n_2894)
);

NAND4xp75_ASAP7_75t_L g2895 ( 
.A(n_2880),
.B(n_470),
.C(n_474),
.D(n_475),
.Y(n_2895)
);

NAND2xp5_ASAP7_75t_L g2896 ( 
.A(n_2885),
.B(n_474),
.Y(n_2896)
);

BUFx2_ASAP7_75t_L g2897 ( 
.A(n_2890),
.Y(n_2897)
);

NAND2xp5_ASAP7_75t_L g2898 ( 
.A(n_2890),
.B(n_475),
.Y(n_2898)
);

AO22x2_ASAP7_75t_L g2899 ( 
.A1(n_2882),
.A2(n_476),
.B1(n_477),
.B2(n_479),
.Y(n_2899)
);

XOR2xp5_ASAP7_75t_L g2900 ( 
.A(n_2889),
.B(n_476),
.Y(n_2900)
);

INVx1_ASAP7_75t_L g2901 ( 
.A(n_2883),
.Y(n_2901)
);

OAI22xp5_ASAP7_75t_L g2902 ( 
.A1(n_2879),
.A2(n_2891),
.B1(n_2888),
.B2(n_481),
.Y(n_2902)
);

OAI22xp5_ASAP7_75t_SL g2903 ( 
.A1(n_2886),
.A2(n_477),
.B1(n_480),
.B2(n_481),
.Y(n_2903)
);

NAND2xp5_ASAP7_75t_L g2904 ( 
.A(n_2893),
.B(n_483),
.Y(n_2904)
);

AOI21xp5_ASAP7_75t_L g2905 ( 
.A1(n_2897),
.A2(n_483),
.B(n_485),
.Y(n_2905)
);

AOI22xp5_ASAP7_75t_L g2906 ( 
.A1(n_2892),
.A2(n_486),
.B1(n_487),
.B2(n_488),
.Y(n_2906)
);

INVx1_ASAP7_75t_L g2907 ( 
.A(n_2894),
.Y(n_2907)
);

AND2x2_ASAP7_75t_L g2908 ( 
.A(n_2894),
.B(n_486),
.Y(n_2908)
);

OAI21xp5_ASAP7_75t_L g2909 ( 
.A1(n_2898),
.A2(n_2901),
.B(n_2900),
.Y(n_2909)
);

AOI21xp33_ASAP7_75t_L g2910 ( 
.A1(n_2896),
.A2(n_487),
.B(n_489),
.Y(n_2910)
);

AOI21xp33_ASAP7_75t_L g2911 ( 
.A1(n_2899),
.A2(n_489),
.B(n_490),
.Y(n_2911)
);

OAI22xp33_ASAP7_75t_L g2912 ( 
.A1(n_2902),
.A2(n_495),
.B1(n_496),
.B2(n_497),
.Y(n_2912)
);

AOI21xp5_ASAP7_75t_L g2913 ( 
.A1(n_2903),
.A2(n_498),
.B(n_499),
.Y(n_2913)
);

OAI22xp5_ASAP7_75t_L g2914 ( 
.A1(n_2895),
.A2(n_499),
.B1(n_500),
.B2(n_501),
.Y(n_2914)
);

AOI21xp5_ASAP7_75t_L g2915 ( 
.A1(n_2907),
.A2(n_501),
.B(n_502),
.Y(n_2915)
);

INVx1_ASAP7_75t_L g2916 ( 
.A(n_2908),
.Y(n_2916)
);

INVx1_ASAP7_75t_L g2917 ( 
.A(n_2904),
.Y(n_2917)
);

OAI21xp5_ASAP7_75t_L g2918 ( 
.A1(n_2909),
.A2(n_502),
.B(n_503),
.Y(n_2918)
);

AOI31xp33_ASAP7_75t_L g2919 ( 
.A1(n_2911),
.A2(n_504),
.A3(n_505),
.B(n_506),
.Y(n_2919)
);

AOI21xp5_ASAP7_75t_L g2920 ( 
.A1(n_2905),
.A2(n_504),
.B(n_506),
.Y(n_2920)
);

AOI21xp5_ASAP7_75t_L g2921 ( 
.A1(n_2910),
.A2(n_507),
.B(n_508),
.Y(n_2921)
);

A2O1A1Ixp33_ASAP7_75t_L g2922 ( 
.A1(n_2906),
.A2(n_508),
.B(n_509),
.C(n_510),
.Y(n_2922)
);

INVx1_ASAP7_75t_L g2923 ( 
.A(n_2914),
.Y(n_2923)
);

OAI22xp5_ASAP7_75t_SL g2924 ( 
.A1(n_2912),
.A2(n_510),
.B1(n_511),
.B2(n_512),
.Y(n_2924)
);

NOR2x1p5_ASAP7_75t_L g2925 ( 
.A(n_2916),
.B(n_2913),
.Y(n_2925)
);

OR2x6_ASAP7_75t_L g2926 ( 
.A(n_2917),
.B(n_513),
.Y(n_2926)
);

AOI222xp33_ASAP7_75t_SL g2927 ( 
.A1(n_2923),
.A2(n_513),
.B1(n_514),
.B2(n_515),
.C1(n_516),
.C2(n_517),
.Y(n_2927)
);

XNOR2xp5_ASAP7_75t_L g2928 ( 
.A(n_2921),
.B(n_514),
.Y(n_2928)
);

AOI21xp5_ASAP7_75t_L g2929 ( 
.A1(n_2919),
.A2(n_515),
.B(n_517),
.Y(n_2929)
);

AOI22xp5_ASAP7_75t_SL g2930 ( 
.A1(n_2928),
.A2(n_2920),
.B1(n_2918),
.B2(n_2915),
.Y(n_2930)
);

AOI22xp5_ASAP7_75t_SL g2931 ( 
.A1(n_2929),
.A2(n_2924),
.B1(n_2922),
.B2(n_520),
.Y(n_2931)
);

OA21x2_ASAP7_75t_L g2932 ( 
.A1(n_2930),
.A2(n_2925),
.B(n_2927),
.Y(n_2932)
);

XNOR2xp5_ASAP7_75t_L g2933 ( 
.A(n_2931),
.B(n_2926),
.Y(n_2933)
);

AOI221xp5_ASAP7_75t_L g2934 ( 
.A1(n_2933),
.A2(n_518),
.B1(n_519),
.B2(n_520),
.C(n_521),
.Y(n_2934)
);

AOI211xp5_ASAP7_75t_L g2935 ( 
.A1(n_2934),
.A2(n_2932),
.B(n_519),
.C(n_523),
.Y(n_2935)
);


endmodule