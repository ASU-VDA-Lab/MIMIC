module real_jpeg_12332_n_18 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_323, n_6, n_11, n_14, n_7, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_323;
input n_6;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_216;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx12f_ASAP7_75t_L g98 ( 
.A(n_0),
.Y(n_98)
);

BUFx16f_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

BUFx12_ASAP7_75t_L g60 ( 
.A(n_2),
.Y(n_60)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_3),
.Y(n_196)
);

AOI21xp33_ASAP7_75t_L g205 ( 
.A1(n_3),
.A2(n_58),
.B(n_206),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_3),
.B(n_81),
.Y(n_226)
);

OAI22xp33_ASAP7_75t_L g257 ( 
.A1(n_3),
.A2(n_34),
.B1(n_35),
.B2(n_196),
.Y(n_257)
);

O2A1O1Ixp33_ASAP7_75t_L g259 ( 
.A1(n_3),
.A2(n_35),
.B(n_46),
.C(n_260),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_3),
.B(n_72),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_3),
.B(n_98),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_3),
.B(n_41),
.Y(n_284)
);

A2O1A1Ixp33_ASAP7_75t_L g293 ( 
.A1(n_3),
.A2(n_27),
.B(n_29),
.C(n_294),
.Y(n_293)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_4),
.A2(n_58),
.B1(n_59),
.B2(n_143),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_4),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_4),
.A2(n_29),
.B1(n_30),
.B2(n_143),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_4),
.A2(n_34),
.B1(n_35),
.B2(n_143),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_4),
.A2(n_43),
.B1(n_47),
.B2(n_143),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_6),
.A2(n_58),
.B1(n_59),
.B2(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_6),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_6),
.A2(n_29),
.B1(n_30),
.B2(n_64),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_6),
.A2(n_34),
.B1(n_35),
.B2(n_64),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_6),
.A2(n_43),
.B1(n_47),
.B2(n_64),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_7),
.A2(n_58),
.B1(n_59),
.B2(n_171),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_7),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_7),
.A2(n_29),
.B1(n_30),
.B2(n_171),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_7),
.A2(n_34),
.B1(n_35),
.B2(n_171),
.Y(n_265)
);

OAI22xp33_ASAP7_75t_SL g272 ( 
.A1(n_7),
.A2(n_43),
.B1(n_47),
.B2(n_171),
.Y(n_272)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_8),
.A2(n_58),
.B1(n_59),
.B2(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_8),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_8),
.A2(n_29),
.B1(n_30),
.B2(n_106),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_8),
.A2(n_34),
.B1(n_35),
.B2(n_106),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_8),
.A2(n_43),
.B1(n_47),
.B2(n_106),
.Y(n_239)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

BUFx8_ASAP7_75t_L g56 ( 
.A(n_11),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_12),
.A2(n_58),
.B1(n_59),
.B2(n_67),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_12),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_12),
.A2(n_29),
.B1(n_30),
.B2(n_67),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_12),
.A2(n_34),
.B1(n_35),
.B2(n_67),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_12),
.A2(n_43),
.B1(n_47),
.B2(n_67),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_L g186 ( 
.A1(n_13),
.A2(n_58),
.B1(n_59),
.B2(n_187),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_13),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_13),
.A2(n_29),
.B1(n_30),
.B2(n_187),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_13),
.A2(n_34),
.B1(n_35),
.B2(n_187),
.Y(n_258)
);

OAI22xp33_ASAP7_75t_SL g279 ( 
.A1(n_13),
.A2(n_43),
.B1(n_47),
.B2(n_187),
.Y(n_279)
);

AOI22xp33_ASAP7_75t_L g36 ( 
.A1(n_14),
.A2(n_29),
.B1(n_30),
.B2(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_14),
.A2(n_37),
.B1(n_58),
.B2(n_59),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_14),
.A2(n_34),
.B1(n_35),
.B2(n_37),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g134 ( 
.A1(n_14),
.A2(n_37),
.B1(n_43),
.B2(n_47),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_15),
.A2(n_29),
.B1(n_30),
.B2(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_15),
.A2(n_34),
.B1(n_35),
.B2(n_39),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_15),
.A2(n_39),
.B1(n_43),
.B2(n_47),
.Y(n_99)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_17),
.A2(n_58),
.B1(n_59),
.B2(n_62),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_17),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_17),
.A2(n_29),
.B1(n_30),
.B2(n_62),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_17),
.A2(n_34),
.B1(n_35),
.B2(n_62),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_17),
.A2(n_43),
.B1(n_47),
.B2(n_62),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_87),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_85),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_73),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_21),
.B(n_73),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_65),
.C(n_68),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_22),
.A2(n_65),
.B1(n_114),
.B2(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_22),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_52),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_40),
.B2(n_51),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_25),
.B(n_40),
.C(n_52),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_26),
.A2(n_33),
.B1(n_36),
.B2(n_38),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_26),
.A2(n_33),
.B1(n_111),
.B2(n_140),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_26),
.A2(n_33),
.B1(n_140),
.B2(n_168),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_26),
.A2(n_33),
.B1(n_182),
.B2(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_27),
.A2(n_70),
.B1(n_71),
.B2(n_72),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_SL g75 ( 
.A1(n_27),
.A2(n_72),
.B(n_76),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_27),
.A2(n_70),
.B1(n_72),
.B2(n_110),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_27),
.A2(n_72),
.B1(n_181),
.B2(n_183),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_27),
.A2(n_72),
.B1(n_222),
.B2(n_224),
.Y(n_221)
);

AND2x2_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_33),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_29),
.A2(n_30),
.B1(n_31),
.B2(n_32),
.Y(n_28)
);

OA22x2_ASAP7_75t_L g54 ( 
.A1(n_29),
.A2(n_30),
.B1(n_55),
.B2(n_56),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_29),
.B(n_55),
.Y(n_194)
);

OAI32xp33_ASAP7_75t_L g235 ( 
.A1(n_29),
.A2(n_31),
.A3(n_34),
.B1(n_236),
.B2(n_237),
.Y(n_235)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

OAI32xp33_ASAP7_75t_L g193 ( 
.A1(n_30),
.A2(n_56),
.A3(n_58),
.B1(n_194),
.B2(n_195),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_30),
.B(n_196),
.Y(n_236)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_31),
.Y(n_32)
);

OA22x2_ASAP7_75t_L g33 ( 
.A1(n_31),
.A2(n_32),
.B1(n_34),
.B2(n_35),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_32),
.B(n_35),
.Y(n_237)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_33),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_L g292 ( 
.A1(n_33),
.A2(n_223),
.B(n_293),
.Y(n_292)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_34),
.Y(n_35)
);

OAI22xp33_ASAP7_75t_L g49 ( 
.A1(n_34),
.A2(n_35),
.B1(n_45),
.B2(n_46),
.Y(n_49)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_36),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_38),
.Y(n_76)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_40),
.B(n_65),
.C(n_69),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_40),
.A2(n_51),
.B1(n_69),
.B2(n_117),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_48),
.B(n_50),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_41),
.A2(n_48),
.B1(n_102),
.B2(n_103),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_41),
.A2(n_48),
.B1(n_50),
.B2(n_103),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_41),
.A2(n_48),
.B1(n_102),
.B2(n_137),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_41),
.A2(n_48),
.B1(n_165),
.B2(n_201),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_41),
.A2(n_48),
.B1(n_201),
.B2(n_230),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_41),
.A2(n_48),
.B1(n_257),
.B2(n_258),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_41),
.A2(n_48),
.B1(n_258),
.B2(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_42),
.B(n_49),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_42),
.A2(n_138),
.B1(n_164),
.B2(n_166),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_42),
.A2(n_166),
.B1(n_231),
.B2(n_296),
.Y(n_295)
);

OA22x2_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_45),
.B1(n_46),
.B2(n_47),
.Y(n_42)
);

INVx3_ASAP7_75t_SL g47 ( 
.A(n_43),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_43),
.B(n_97),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_43),
.B(n_281),
.Y(n_280)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

OAI21xp33_ASAP7_75t_L g260 ( 
.A1(n_45),
.A2(n_47),
.B(n_196),
.Y(n_260)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_48),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_53),
.A2(n_54),
.B1(n_61),
.B2(n_63),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_53),
.A2(n_54),
.B1(n_61),
.B2(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_53),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_53),
.A2(n_54),
.B1(n_66),
.B2(n_105),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_53),
.A2(n_54),
.B1(n_105),
.B2(n_142),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_53),
.A2(n_54),
.B1(n_142),
.B2(n_170),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_53),
.A2(n_54),
.B1(n_186),
.B2(n_205),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_54),
.B(n_57),
.Y(n_53)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_54),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_55),
.A2(n_56),
.B1(n_58),
.B2(n_59),
.Y(n_57)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_59),
.B(n_196),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_63),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_65),
.A2(n_114),
.B1(n_115),
.B2(n_116),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_65),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_68),
.B(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_69),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_84),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_77),
.B1(n_82),
.B2(n_83),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_75),
.Y(n_82)
);

CKINVDCx14_ASAP7_75t_R g83 ( 
.A(n_77),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_79),
.B1(n_80),
.B2(n_81),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_79),
.A2(n_81),
.B1(n_185),
.B2(n_188),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

AO21x1_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_149),
.B(n_319),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_144),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_90),
.B(n_120),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_90),
.B(n_120),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_107),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_91),
.B(n_113),
.C(n_118),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g91 ( 
.A1(n_92),
.A2(n_95),
.B(n_104),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_92),
.A2(n_93),
.B1(n_123),
.B2(n_124),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_100),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_94),
.A2(n_95),
.B1(n_104),
.B2(n_125),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_94),
.A2(n_95),
.B1(n_100),
.B2(n_101),
.Y(n_155)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_96),
.A2(n_98),
.B(n_99),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_96),
.A2(n_98),
.B1(n_99),
.B2(n_133),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_96),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_96),
.A2(n_98),
.B1(n_162),
.B2(n_192),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_96),
.A2(n_98),
.B1(n_192),
.B2(n_228),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_96),
.A2(n_98),
.B1(n_228),
.B2(n_239),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_96),
.A2(n_98),
.B1(n_239),
.B2(n_267),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_96),
.A2(n_98),
.B1(n_196),
.B2(n_279),
.Y(n_278)
);

AOI22xp33_ASAP7_75t_L g283 ( 
.A1(n_96),
.A2(n_98),
.B1(n_272),
.B2(n_279),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_97),
.A2(n_134),
.B1(n_160),
.B2(n_161),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_97),
.A2(n_160),
.B1(n_271),
.B2(n_273),
.Y(n_270)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

CKINVDCx14_ASAP7_75t_R g125 ( 
.A(n_104),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_113),
.B1(n_118),
.B2(n_119),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_108),
.Y(n_118)
);

OAI21xp33_ASAP7_75t_L g127 ( 
.A1(n_108),
.A2(n_109),
.B(n_112),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_112),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_113),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_116),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_126),
.C(n_128),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_121),
.A2(n_122),
.B1(n_126),
.B2(n_127),
.Y(n_173)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_128),
.B(n_173),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_139),
.C(n_141),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_129),
.A2(n_130),
.B1(n_153),
.B2(n_154),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_130),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_135),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_131),
.A2(n_132),
.B1(n_135),
.B2(n_136),
.Y(n_209)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_139),
.B(n_141),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g319 ( 
.A1(n_144),
.A2(n_320),
.B(n_321),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_146),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_145),
.B(n_146),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_150),
.A2(n_174),
.B(n_318),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_172),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_151),
.B(n_172),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_155),
.C(n_156),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_152),
.B(n_155),
.Y(n_316)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_156),
.B(n_316),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_167),
.C(n_169),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_157),
.A2(n_158),
.B1(n_211),
.B2(n_212),
.Y(n_210)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_163),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_159),
.B(n_163),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_162),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_165),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_167),
.B(n_169),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_168),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_170),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_175),
.A2(n_313),
.B(n_317),
.Y(n_174)
);

OAI221xp5_ASAP7_75t_L g175 ( 
.A1(n_176),
.A2(n_216),
.B1(n_311),
.B2(n_312),
.C(n_323),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_207),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_177),
.B(n_207),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_197),
.C(n_198),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_178),
.B(n_310),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_189),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_184),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_180),
.B(n_184),
.C(n_189),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_190),
.B(n_193),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_190),
.A2(n_191),
.B1(n_193),
.B2(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_193),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_195),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_197),
.B(n_198),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_202),
.C(n_204),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_199),
.A2(n_200),
.B1(n_202),
.B2(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_202),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_203),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_204),
.B(n_243),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_215),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_209),
.A2(n_210),
.B1(n_213),
.B2(n_214),
.Y(n_208)
);

CKINVDCx14_ASAP7_75t_R g213 ( 
.A(n_209),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_209),
.B(n_214),
.C(n_215),
.Y(n_314)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_210),
.Y(n_214)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_217),
.B(n_307),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_218),
.A2(n_250),
.B(n_306),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_240),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_219),
.B(n_240),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_229),
.C(n_232),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_220),
.B(n_303),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_SL g220 ( 
.A(n_221),
.B(n_225),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_221),
.B(n_226),
.C(n_227),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_227),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_229),
.A2(n_232),
.B1(n_233),
.B2(n_304),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_229),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_238),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_234),
.A2(n_235),
.B1(n_238),
.B2(n_298),
.Y(n_297)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

CKINVDCx16_ASAP7_75t_R g294 ( 
.A(n_236),
.Y(n_294)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_238),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_241),
.A2(n_242),
.B1(n_245),
.B2(n_249),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_241),
.B(n_246),
.C(n_248),
.Y(n_308)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_245),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_SL g245 ( 
.A(n_246),
.B(n_248),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_251),
.A2(n_300),
.B(n_305),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_252),
.A2(n_288),
.B(n_299),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_253),
.A2(n_268),
.B(n_287),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_261),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g287 ( 
.A(n_254),
.B(n_261),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_255),
.B(n_259),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_255),
.A2(n_256),
.B1(n_259),
.B2(n_275),
.Y(n_274)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_259),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_266),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_264),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_263),
.B(n_264),
.C(n_266),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_265),
.Y(n_296)
);

CKINVDCx14_ASAP7_75t_R g273 ( 
.A(n_267),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_269),
.A2(n_276),
.B(n_286),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_274),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_270),
.B(n_274),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_277),
.A2(n_282),
.B(n_285),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_278),
.B(n_280),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_284),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_283),
.B(n_284),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_290),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_289),
.B(n_290),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_297),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_295),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_292),
.B(n_295),
.C(n_297),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_302),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_SL g305 ( 
.A(n_301),
.B(n_302),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_309),
.Y(n_307)
);

OR2x2_ASAP7_75t_L g311 ( 
.A(n_308),
.B(n_309),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_315),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_314),
.B(n_315),
.Y(n_317)
);


endmodule