module fake_jpeg_558_n_389 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_389);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_389;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

BUFx16f_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx10_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx16_ASAP7_75t_R g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_3),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_8),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_1),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_5),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_9),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_48),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_49),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_22),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_50),
.Y(n_109)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_17),
.Y(n_51)
);

INVx2_ASAP7_75t_SL g102 ( 
.A(n_51),
.Y(n_102)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_52),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_22),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_53),
.Y(n_136)
);

INVx3_ASAP7_75t_SL g54 ( 
.A(n_17),
.Y(n_54)
);

HB1xp67_ASAP7_75t_L g140 ( 
.A(n_54),
.Y(n_140)
);

INVx4_ASAP7_75t_SL g55 ( 
.A(n_17),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_55),
.Y(n_128)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_56),
.Y(n_99)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_21),
.Y(n_57)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_57),
.Y(n_115)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_21),
.Y(n_58)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_58),
.Y(n_127)
);

INVx4_ASAP7_75t_SL g59 ( 
.A(n_46),
.Y(n_59)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_59),
.Y(n_100)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_23),
.Y(n_60)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_60),
.Y(n_122)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_29),
.Y(n_61)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_61),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_30),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_62),
.B(n_73),
.Y(n_130)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_29),
.Y(n_63)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_63),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_34),
.B(n_14),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_64),
.B(n_89),
.Y(n_105)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_25),
.Y(n_65)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_65),
.Y(n_108)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_26),
.Y(n_66)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_66),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_27),
.B(n_14),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_67),
.B(n_81),
.Y(n_112)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_16),
.Y(n_68)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_68),
.Y(n_111)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_16),
.Y(n_69)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_69),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_33),
.Y(n_70)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_70),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_33),
.Y(n_71)
);

INVx6_ASAP7_75t_L g138 ( 
.A(n_71),
.Y(n_138)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_23),
.Y(n_72)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_72),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_30),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_41),
.Y(n_74)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_74),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_39),
.Y(n_75)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_75),
.Y(n_118)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_34),
.Y(n_76)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_76),
.Y(n_132)
);

HB1xp67_ASAP7_75t_L g77 ( 
.A(n_46),
.Y(n_77)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_77),
.Y(n_133)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_16),
.Y(n_78)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_78),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_25),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_79),
.B(n_86),
.Y(n_134)
);

INVx11_ASAP7_75t_L g80 ( 
.A(n_46),
.Y(n_80)
);

INVx11_ASAP7_75t_L g101 ( 
.A(n_80),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_24),
.B(n_14),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_28),
.A2(n_13),
.B1(n_12),
.B2(n_9),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_82),
.A2(n_44),
.B1(n_40),
.B2(n_45),
.Y(n_119)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_19),
.Y(n_83)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_83),
.Y(n_141)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_19),
.Y(n_84)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_84),
.Y(n_143)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_32),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_85),
.B(n_90),
.Y(n_106)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_32),
.Y(n_86)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_28),
.Y(n_87)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_87),
.Y(n_124)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_38),
.Y(n_88)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_88),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_39),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_38),
.Y(n_90)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_46),
.Y(n_91)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_91),
.Y(n_142)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_16),
.Y(n_92)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_92),
.Y(n_144)
);

BUFx8_ASAP7_75t_L g93 ( 
.A(n_20),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_93),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_37),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_94),
.B(n_95),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_41),
.Y(n_95)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_18),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_96),
.B(n_97),
.Y(n_135)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_18),
.Y(n_97)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_18),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_98),
.B(n_35),
.Y(n_139)
);

AND2x2_ASAP7_75t_SL g113 ( 
.A(n_55),
.B(n_18),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_113),
.B(n_139),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_L g174 ( 
.A1(n_119),
.A2(n_129),
.B1(n_95),
.B2(n_49),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_59),
.A2(n_31),
.B1(n_37),
.B2(n_35),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_121),
.A2(n_145),
.B1(n_91),
.B2(n_71),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_L g125 ( 
.A1(n_48),
.A2(n_40),
.B1(n_44),
.B2(n_31),
.Y(n_125)
);

OAI22xp33_ASAP7_75t_L g153 ( 
.A1(n_125),
.A2(n_87),
.B1(n_65),
.B2(n_56),
.Y(n_153)
);

OAI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_50),
.A2(n_20),
.B1(n_35),
.B2(n_26),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_93),
.A2(n_35),
.B1(n_36),
.B2(n_47),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_67),
.A2(n_20),
.B(n_47),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_148),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_105),
.B(n_81),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_149),
.B(n_159),
.Y(n_192)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_137),
.Y(n_150)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_150),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_134),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_151),
.B(n_156),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_103),
.Y(n_152)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_152),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_153),
.A2(n_136),
.B1(n_109),
.B2(n_124),
.Y(n_205)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_133),
.Y(n_154)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_154),
.Y(n_197)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_106),
.Y(n_155)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_155),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_113),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_106),
.Y(n_157)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_157),
.Y(n_214)
);

O2A1O1Ixp33_ASAP7_75t_SL g158 ( 
.A1(n_125),
.A2(n_54),
.B(n_80),
.C(n_51),
.Y(n_158)
);

AO21x1_ASAP7_75t_L g198 ( 
.A1(n_158),
.A2(n_183),
.B(n_186),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_126),
.B(n_77),
.Y(n_159)
);

INVx6_ASAP7_75t_L g160 ( 
.A(n_103),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_160),
.Y(n_201)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_132),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_161),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_141),
.B(n_70),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_162),
.B(n_165),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_112),
.B(n_13),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_163),
.B(n_166),
.Y(n_194)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_142),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_164),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_143),
.B(n_122),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_131),
.B(n_9),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_130),
.B(n_51),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_167),
.B(n_168),
.Y(n_195)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_99),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_140),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_169),
.B(n_171),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_128),
.B(n_110),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_135),
.B(n_75),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_172),
.B(n_179),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_111),
.B(n_74),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_173),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_174),
.A2(n_188),
.B1(n_121),
.B2(n_145),
.Y(n_189)
);

OAI21xp33_ASAP7_75t_SL g204 ( 
.A1(n_175),
.A2(n_181),
.B(n_184),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_104),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_176),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_100),
.B(n_20),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_178),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_147),
.B(n_53),
.Y(n_179)
);

INVx6_ASAP7_75t_SL g180 ( 
.A(n_102),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g213 ( 
.A(n_180),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_129),
.A2(n_140),
.B1(n_114),
.B2(n_116),
.Y(n_181)
);

HB1xp67_ASAP7_75t_L g182 ( 
.A(n_123),
.Y(n_182)
);

BUFx12_ASAP7_75t_L g193 ( 
.A(n_182),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_104),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_144),
.B(n_1),
.Y(n_184)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_142),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_185),
.A2(n_187),
.B(n_180),
.Y(n_199)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_108),
.Y(n_186)
);

BUFx10_ASAP7_75t_L g187 ( 
.A(n_102),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_107),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_189),
.A2(n_202),
.B1(n_205),
.B2(n_206),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_159),
.B(n_177),
.C(n_165),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_191),
.B(n_157),
.C(n_161),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_199),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_170),
.A2(n_138),
.B1(n_107),
.B2(n_118),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_170),
.A2(n_138),
.B1(n_109),
.B2(n_136),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_172),
.A2(n_162),
.B1(n_179),
.B2(n_177),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_208),
.A2(n_219),
.B1(n_176),
.B2(n_152),
.Y(n_240)
);

AOI22x1_ASAP7_75t_L g215 ( 
.A1(n_177),
.A2(n_114),
.B1(n_120),
.B2(n_127),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_215),
.A2(n_158),
.B1(n_153),
.B2(n_116),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_155),
.A2(n_118),
.B1(n_124),
.B2(n_108),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_192),
.B(n_149),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_220),
.B(n_224),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_221),
.B(n_222),
.C(n_227),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_191),
.B(n_150),
.C(n_151),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_218),
.B(n_178),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_223),
.B(n_236),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_192),
.B(n_188),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_225),
.A2(n_243),
.B1(n_202),
.B2(n_242),
.Y(n_263)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_210),
.Y(n_226)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_226),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_200),
.B(n_146),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_208),
.B(n_154),
.C(n_115),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_228),
.B(n_229),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_200),
.B(n_209),
.Y(n_229)
);

O2A1O1Ixp33_ASAP7_75t_SL g231 ( 
.A1(n_198),
.A2(n_158),
.B(n_183),
.C(n_187),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g260 ( 
.A1(n_231),
.A2(n_244),
.B(n_204),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_218),
.A2(n_164),
.B(n_117),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_SL g257 ( 
.A1(n_232),
.A2(n_198),
.B(n_190),
.Y(n_257)
);

INVx4_ASAP7_75t_L g234 ( 
.A(n_196),
.Y(n_234)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_234),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_212),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_235),
.B(n_241),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_203),
.B(n_168),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_203),
.B(n_186),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_237),
.B(n_238),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_209),
.B(n_214),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_195),
.B(n_185),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_239),
.B(n_243),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_240),
.A2(n_242),
.B1(n_213),
.B2(n_206),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_217),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_205),
.A2(n_160),
.B1(n_36),
.B2(n_187),
.Y(n_242)
);

CKINVDCx14_ASAP7_75t_R g243 ( 
.A(n_215),
.Y(n_243)
);

OR2x2_ASAP7_75t_L g244 ( 
.A(n_190),
.B(n_187),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_195),
.B(n_2),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_245),
.B(n_213),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g246 ( 
.A(n_237),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_246),
.B(n_255),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_224),
.A2(n_215),
.B1(n_189),
.B2(n_214),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_249),
.A2(n_263),
.B1(n_230),
.B2(n_225),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_233),
.A2(n_199),
.B(n_198),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_250),
.A2(n_257),
.B(n_232),
.Y(n_268)
);

CKINVDCx16_ASAP7_75t_R g255 ( 
.A(n_236),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g272 ( 
.A(n_259),
.B(n_216),
.Y(n_272)
);

INVx1_ASAP7_75t_SL g275 ( 
.A(n_260),
.Y(n_275)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_226),
.Y(n_261)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_261),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_262),
.A2(n_230),
.B1(n_240),
.B2(n_235),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_239),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_264),
.B(n_266),
.Y(n_274)
);

BUFx24_ASAP7_75t_SL g266 ( 
.A(n_220),
.Y(n_266)
);

BUFx24_ASAP7_75t_SL g267 ( 
.A(n_223),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_267),
.B(n_194),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_268),
.B(n_280),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_248),
.B(n_238),
.Y(n_269)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_269),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_271),
.A2(n_246),
.B1(n_252),
.B2(n_253),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_272),
.B(n_287),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_248),
.B(n_229),
.Y(n_273)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_273),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_277),
.A2(n_285),
.B1(n_265),
.B2(n_250),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_278),
.B(n_194),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_247),
.B(n_222),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_279),
.B(n_253),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_254),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g281 ( 
.A1(n_260),
.A2(n_244),
.B(n_231),
.Y(n_281)
);

INVx1_ASAP7_75t_SL g291 ( 
.A(n_281),
.Y(n_291)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_256),
.Y(n_282)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_282),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_251),
.B(n_245),
.Y(n_283)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_283),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_254),
.B(n_227),
.Y(n_284)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_284),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_249),
.A2(n_204),
.B1(n_228),
.B2(n_231),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_256),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_286),
.B(n_201),
.Y(n_305)
);

OAI21xp33_ASAP7_75t_L g287 ( 
.A1(n_257),
.A2(n_244),
.B(n_221),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_279),
.B(n_247),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_290),
.B(n_270),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_292),
.B(n_270),
.C(n_269),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_285),
.A2(n_263),
.B1(n_265),
.B2(n_262),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_295),
.A2(n_296),
.B1(n_303),
.B2(n_276),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_277),
.A2(n_251),
.B1(n_252),
.B2(n_255),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_298),
.A2(n_299),
.B1(n_301),
.B2(n_302),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_SL g300 ( 
.A(n_273),
.B(n_247),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_SL g313 ( 
.A(n_300),
.B(n_268),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_271),
.A2(n_280),
.B1(n_283),
.B2(n_272),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_275),
.A2(n_261),
.B1(n_259),
.B2(n_258),
.Y(n_303)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_305),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_305),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g326 ( 
.A1(n_308),
.A2(n_321),
.B1(n_288),
.B2(n_297),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_292),
.B(n_284),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_309),
.B(n_310),
.Y(n_328)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_293),
.Y(n_311)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_311),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_312),
.B(n_314),
.C(n_315),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_SL g332 ( 
.A(n_313),
.B(n_317),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_290),
.B(n_275),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_300),
.B(n_274),
.C(n_281),
.Y(n_315)
);

BUFx6f_ASAP7_75t_L g316 ( 
.A(n_294),
.Y(n_316)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_316),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_SL g317 ( 
.A(n_297),
.B(n_274),
.Y(n_317)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_288),
.Y(n_319)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_319),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_301),
.B(n_286),
.C(n_282),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_320),
.B(n_323),
.Y(n_325)
);

AND3x1_ASAP7_75t_L g322 ( 
.A(n_289),
.B(n_276),
.C(n_258),
.Y(n_322)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_322),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_SL g323 ( 
.A(n_289),
.B(n_278),
.C(n_211),
.Y(n_323)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_326),
.Y(n_348)
);

INVx13_ASAP7_75t_L g327 ( 
.A(n_322),
.Y(n_327)
);

CKINVDCx16_ASAP7_75t_R g350 ( 
.A(n_327),
.Y(n_350)
);

BUFx12_ASAP7_75t_L g330 ( 
.A(n_314),
.Y(n_330)
);

HB1xp67_ASAP7_75t_L g340 ( 
.A(n_330),
.Y(n_340)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_307),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_335),
.A2(n_304),
.B1(n_241),
.B2(n_303),
.Y(n_339)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_316),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_SL g342 ( 
.A(n_336),
.B(n_304),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_L g337 ( 
.A1(n_318),
.A2(n_291),
.B(n_306),
.Y(n_337)
);

AOI21xp5_ASAP7_75t_L g346 ( 
.A1(n_337),
.A2(n_338),
.B(n_216),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_SL g338 ( 
.A1(n_313),
.A2(n_291),
.B(n_295),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_339),
.B(n_341),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_328),
.B(n_310),
.C(n_320),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_342),
.B(n_344),
.Y(n_353)
);

OAI21xp5_ASAP7_75t_L g343 ( 
.A1(n_329),
.A2(n_315),
.B(n_317),
.Y(n_343)
);

AOI21xp5_ASAP7_75t_L g361 ( 
.A1(n_343),
.A2(n_349),
.B(n_340),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_328),
.B(n_309),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_333),
.B(n_234),
.C(n_201),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_345),
.B(n_349),
.C(n_329),
.Y(n_354)
);

AOI21xp33_ASAP7_75t_L g358 ( 
.A1(n_346),
.A2(n_334),
.B(n_332),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_333),
.B(n_211),
.Y(n_347)
);

XOR2xp5_ASAP7_75t_L g359 ( 
.A(n_347),
.B(n_330),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_337),
.B(n_234),
.C(n_210),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_SL g351 ( 
.A(n_325),
.B(n_197),
.Y(n_351)
);

NOR2xp67_ASAP7_75t_L g355 ( 
.A(n_351),
.B(n_331),
.Y(n_355)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_354),
.Y(n_365)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_355),
.Y(n_369)
);

OAI21xp5_ASAP7_75t_SL g356 ( 
.A1(n_343),
.A2(n_325),
.B(n_338),
.Y(n_356)
);

AOI21xp5_ASAP7_75t_L g370 ( 
.A1(n_356),
.A2(n_358),
.B(n_361),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_341),
.B(n_332),
.C(n_335),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_357),
.B(n_360),
.Y(n_371)
);

AND2x2_ASAP7_75t_L g363 ( 
.A(n_359),
.B(n_344),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_L g360 ( 
.A1(n_348),
.A2(n_327),
.B1(n_324),
.B2(n_330),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_347),
.B(n_324),
.C(n_207),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_362),
.B(n_345),
.C(n_350),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_363),
.B(n_364),
.Y(n_373)
);

OAI21xp5_ASAP7_75t_SL g366 ( 
.A1(n_352),
.A2(n_207),
.B(n_196),
.Y(n_366)
);

AOI21xp5_ASAP7_75t_SL g377 ( 
.A1(n_366),
.A2(n_101),
.B(n_193),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_354),
.B(n_219),
.C(n_197),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_SL g376 ( 
.A(n_367),
.B(n_2),
.Y(n_376)
);

XOR2xp5_ASAP7_75t_L g368 ( 
.A(n_361),
.B(n_193),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_368),
.B(n_362),
.C(n_359),
.Y(n_374)
);

A2O1A1Ixp33_ASAP7_75t_L g372 ( 
.A1(n_370),
.A2(n_353),
.B(n_369),
.C(n_371),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_372),
.B(n_374),
.Y(n_381)
);

OAI21xp5_ASAP7_75t_SL g375 ( 
.A1(n_365),
.A2(n_363),
.B(n_357),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_SL g378 ( 
.A(n_375),
.B(n_376),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_377),
.B(n_368),
.C(n_367),
.Y(n_379)
);

OAI21xp5_ASAP7_75t_L g383 ( 
.A1(n_379),
.A2(n_193),
.B(n_3),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_373),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_380),
.A2(n_193),
.B1(n_101),
.B2(n_4),
.Y(n_382)
);

HB1xp67_ASAP7_75t_L g385 ( 
.A(n_382),
.Y(n_385)
);

OAI321xp33_ASAP7_75t_L g386 ( 
.A1(n_383),
.A2(n_384),
.A3(n_378),
.B1(n_6),
.B2(n_7),
.C(n_8),
.Y(n_386)
);

OAI311xp33_ASAP7_75t_L g384 ( 
.A1(n_381),
.A2(n_2),
.A3(n_3),
.B1(n_4),
.C1(n_5),
.Y(n_384)
);

OAI21xp5_ASAP7_75t_L g387 ( 
.A1(n_386),
.A2(n_5),
.B(n_6),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_387),
.B(n_385),
.C(n_7),
.Y(n_388)
);

OAI21xp5_ASAP7_75t_L g389 ( 
.A1(n_388),
.A2(n_6),
.B(n_8),
.Y(n_389)
);


endmodule