module fake_jpeg_245_n_230 (n_13, n_21, n_53, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_230);

input n_13;
input n_21;
input n_53;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_230;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_223;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_122;
wire n_75;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_91;
wire n_93;
wire n_54;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx3_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_51),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_25),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_21),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_37),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_3),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g62 ( 
.A(n_48),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_22),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_16),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_17),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_32),
.Y(n_66)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_31),
.Y(n_67)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_7),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_29),
.Y(n_70)
);

BUFx16f_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_10),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_47),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_6),
.Y(n_74)
);

BUFx5_ASAP7_75t_L g75 ( 
.A(n_42),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_11),
.Y(n_76)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_35),
.Y(n_77)
);

BUFx5_ASAP7_75t_L g78 ( 
.A(n_44),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_17),
.Y(n_79)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_55),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_80),
.Y(n_90)
);

INVx13_ASAP7_75t_L g81 ( 
.A(n_71),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_81),
.Y(n_88)
);

BUFx24_ASAP7_75t_L g82 ( 
.A(n_71),
.Y(n_82)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_82),
.Y(n_97)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_71),
.Y(n_83)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_83),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_65),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_84),
.B(n_80),
.Y(n_95)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_59),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_85),
.B(n_86),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_69),
.B(n_0),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_59),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_87),
.B(n_60),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_84),
.A2(n_64),
.B1(n_76),
.B2(n_65),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_89),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_85),
.A2(n_64),
.B1(n_76),
.B2(n_72),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_91),
.A2(n_74),
.B1(n_63),
.B2(n_62),
.Y(n_106)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_83),
.Y(n_92)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_92),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_95),
.Y(n_111)
);

OAI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_87),
.A2(n_67),
.B1(n_68),
.B2(n_77),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_96),
.A2(n_99),
.B1(n_68),
.B2(n_67),
.Y(n_114)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_80),
.Y(n_98)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_98),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_86),
.A2(n_70),
.B1(n_55),
.B2(n_57),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_100),
.B(n_77),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_82),
.B(n_61),
.Y(n_101)
);

OAI21xp33_ASAP7_75t_L g102 ( 
.A1(n_101),
.A2(n_82),
.B(n_79),
.Y(n_102)
);

CKINVDCx14_ASAP7_75t_R g138 ( 
.A(n_102),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_93),
.B(n_94),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_104),
.B(n_109),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_106),
.B(n_108),
.Y(n_132)
);

BUFx12f_ASAP7_75t_L g107 ( 
.A(n_94),
.Y(n_107)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_107),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_100),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_98),
.A2(n_70),
.B1(n_57),
.B2(n_58),
.Y(n_109)
);

INVx4_ASAP7_75t_SL g110 ( 
.A(n_88),
.Y(n_110)
);

INVxp67_ASAP7_75t_SL g140 ( 
.A(n_110),
.Y(n_140)
);

A2O1A1Ixp33_ASAP7_75t_L g112 ( 
.A1(n_93),
.A2(n_73),
.B(n_66),
.C(n_63),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_112),
.A2(n_116),
.B(n_119),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_114),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_115),
.B(n_117),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_92),
.B(n_81),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_101),
.B(n_88),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_99),
.B(n_54),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_118),
.B(n_120),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_90),
.A2(n_58),
.B1(n_56),
.B2(n_54),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_97),
.B(n_56),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_116),
.Y(n_121)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_121),
.Y(n_145)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_105),
.Y(n_122)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_122),
.Y(n_151)
);

INVx13_ASAP7_75t_L g124 ( 
.A(n_110),
.Y(n_124)
);

CKINVDCx14_ASAP7_75t_R g165 ( 
.A(n_124),
.Y(n_165)
);

INVx13_ASAP7_75t_L g125 ( 
.A(n_107),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_125),
.Y(n_154)
);

HB1xp67_ASAP7_75t_L g127 ( 
.A(n_103),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_127),
.B(n_131),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_113),
.A2(n_102),
.B(n_104),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_128),
.A2(n_82),
.B(n_78),
.Y(n_150)
);

INVx3_ASAP7_75t_SL g130 ( 
.A(n_103),
.Y(n_130)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_130),
.Y(n_149)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_111),
.Y(n_131)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_112),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_134),
.B(n_137),
.Y(n_153)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_107),
.Y(n_137)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_113),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_139),
.B(n_141),
.Y(n_156)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_114),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_109),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_142),
.B(n_0),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_133),
.B(n_90),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_143),
.B(n_147),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_138),
.B(n_90),
.C(n_81),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_144),
.B(n_36),
.C(n_34),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_129),
.A2(n_97),
.B1(n_78),
.B2(n_75),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_146),
.A2(n_158),
.B1(n_30),
.B2(n_28),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_136),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_150),
.A2(n_157),
.B(n_41),
.Y(n_171)
);

AO21x1_ASAP7_75t_L g152 ( 
.A1(n_135),
.A2(n_75),
.B(n_53),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_152),
.A2(n_164),
.B(n_8),
.Y(n_175)
);

CKINVDCx14_ASAP7_75t_R g184 ( 
.A(n_155),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_129),
.A2(n_52),
.B1(n_50),
.B2(n_49),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_132),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_126),
.B(n_43),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_159),
.B(n_160),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_123),
.B(n_1),
.Y(n_160)
);

INVx8_ASAP7_75t_L g161 ( 
.A(n_124),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_161),
.B(n_154),
.Y(n_174)
);

OR2x2_ASAP7_75t_L g162 ( 
.A(n_140),
.B(n_2),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_162),
.B(n_166),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_130),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_163)
);

OA21x2_ASAP7_75t_L g178 ( 
.A1(n_163),
.A2(n_9),
.B(n_10),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_140),
.A2(n_4),
.B(n_5),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_125),
.Y(n_166)
);

INVxp33_ASAP7_75t_L g167 ( 
.A(n_156),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_167),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_153),
.A2(n_137),
.B(n_136),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_169),
.B(n_170),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_150),
.A2(n_7),
.B(n_8),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_171),
.B(n_175),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_143),
.B(n_38),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_172),
.B(n_176),
.Y(n_189)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_148),
.Y(n_173)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_173),
.Y(n_192)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_174),
.Y(n_195)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_151),
.Y(n_177)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_177),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_178),
.A2(n_183),
.B1(n_163),
.B2(n_162),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_180),
.B(n_181),
.Y(n_190)
);

AOI322xp5_ASAP7_75t_L g181 ( 
.A1(n_145),
.A2(n_26),
.A3(n_24),
.B1(n_23),
.B2(n_27),
.C1(n_14),
.C2(n_15),
.Y(n_181)
);

MAJx2_ASAP7_75t_L g182 ( 
.A(n_144),
.B(n_9),
.C(n_11),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_182),
.B(n_186),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_157),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_159),
.B(n_12),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_151),
.Y(n_187)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_187),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_179),
.B(n_152),
.Y(n_193)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_193),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_169),
.Y(n_194)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_194),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_199),
.A2(n_178),
.B1(n_184),
.B2(n_175),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_189),
.B(n_176),
.C(n_182),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_201),
.B(n_202),
.C(n_205),
.Y(n_211)
);

NAND2x1_ASAP7_75t_L g202 ( 
.A(n_195),
.B(n_185),
.Y(n_202)
);

HB1xp67_ASAP7_75t_L g203 ( 
.A(n_196),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_203),
.B(n_206),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_204),
.A2(n_209),
.B1(n_197),
.B2(n_164),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_189),
.B(n_188),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_192),
.A2(n_167),
.B1(n_178),
.B2(n_170),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_200),
.A2(n_168),
.B1(n_165),
.B2(n_154),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_207),
.B(n_200),
.C(n_209),
.Y(n_212)
);

HB1xp67_ASAP7_75t_L g209 ( 
.A(n_198),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_212),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_210),
.B(n_191),
.C(n_190),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_213),
.B(n_214),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_208),
.B(n_172),
.C(n_199),
.Y(n_214)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_215),
.Y(n_221)
);

INVx11_ASAP7_75t_L g216 ( 
.A(n_203),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_216),
.B(n_147),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_219),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_218),
.B(n_211),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_223),
.B(n_220),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_224),
.B(n_220),
.C(n_221),
.Y(n_225)
);

AOI322xp5_ASAP7_75t_L g226 ( 
.A1(n_225),
.A2(n_222),
.A3(n_217),
.B1(n_197),
.B2(n_216),
.C1(n_149),
.C2(n_161),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_226),
.B(n_21),
.C(n_15),
.Y(n_227)
);

NOR3xp33_ASAP7_75t_L g228 ( 
.A(n_227),
.B(n_13),
.C(n_16),
.Y(n_228)
);

AOI321xp33_ASAP7_75t_L g229 ( 
.A1(n_228),
.A2(n_18),
.A3(n_19),
.B1(n_20),
.B2(n_158),
.C(n_134),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_229),
.B(n_20),
.Y(n_230)
);


endmodule