module fake_jpeg_31198_n_178 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_178);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_178;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_154;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx24_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_19),
.B(n_24),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_13),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_38),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_20),
.Y(n_56)
);

INVx2_ASAP7_75t_SL g57 ( 
.A(n_42),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_29),
.B(n_23),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_34),
.Y(n_59)
);

INVx1_ASAP7_75t_SL g60 ( 
.A(n_15),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_27),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_21),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_45),
.Y(n_63)
);

INVx13_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_13),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_14),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_16),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_30),
.Y(n_68)
);

INVx13_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_6),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_39),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_22),
.Y(n_72)
);

INVx13_ASAP7_75t_L g73 ( 
.A(n_1),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_33),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_18),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_64),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_77),
.Y(n_93)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_52),
.Y(n_78)
);

INVx11_ASAP7_75t_L g99 ( 
.A(n_78),
.Y(n_99)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_52),
.Y(n_79)
);

INVx5_ASAP7_75t_SL g98 ( 
.A(n_79),
.Y(n_98)
);

INVx2_ASAP7_75t_SL g80 ( 
.A(n_52),
.Y(n_80)
);

AO22x1_ASAP7_75t_L g95 ( 
.A1(n_80),
.A2(n_73),
.B1(n_74),
.B2(n_56),
.Y(n_95)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_66),
.Y(n_81)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_81),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_54),
.B(n_0),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_82),
.B(n_83),
.Y(n_86)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_61),
.Y(n_83)
);

A2O1A1Ixp33_ASAP7_75t_L g84 ( 
.A1(n_58),
.A2(n_51),
.B(n_17),
.C(n_25),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_84),
.B(n_44),
.Y(n_92)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_72),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_85),
.B(n_60),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_81),
.A2(n_66),
.B1(n_70),
.B2(n_74),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_87),
.A2(n_75),
.B1(n_71),
.B2(n_62),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_88),
.B(n_95),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_80),
.A2(n_70),
.B1(n_74),
.B2(n_56),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_89),
.A2(n_96),
.B1(n_71),
.B2(n_62),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_85),
.B(n_65),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_90),
.B(n_94),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_92),
.B(n_100),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_80),
.B(n_56),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_79),
.A2(n_78),
.B1(n_57),
.B2(n_76),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_77),
.B(n_53),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_97),
.B(n_3),
.Y(n_119)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_84),
.Y(n_100)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_100),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g122 ( 
.A1(n_101),
.A2(n_104),
.B1(n_111),
.B2(n_50),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_88),
.B(n_68),
.C(n_57),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_103),
.B(n_4),
.C(n_5),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_106),
.B(n_112),
.Y(n_123)
);

O2A1O1Ixp33_ASAP7_75t_SL g107 ( 
.A1(n_95),
.A2(n_94),
.B(n_98),
.C(n_88),
.Y(n_107)
);

A2O1A1Ixp33_ASAP7_75t_L g140 ( 
.A1(n_107),
.A2(n_31),
.B(n_28),
.C(n_10),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_95),
.A2(n_75),
.B1(n_55),
.B2(n_67),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_108),
.A2(n_113),
.B1(n_116),
.B2(n_120),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_92),
.B(n_59),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_109),
.B(n_110),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_86),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_91),
.A2(n_63),
.B1(n_69),
.B2(n_64),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_98),
.B(n_69),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_91),
.A2(n_73),
.B1(n_1),
.B2(n_2),
.Y(n_113)
);

BUFx2_ASAP7_75t_L g115 ( 
.A(n_93),
.Y(n_115)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_115),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_93),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_116)
);

BUFx6f_ASAP7_75t_SL g117 ( 
.A(n_93),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_117),
.Y(n_136)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_99),
.Y(n_118)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_118),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_119),
.B(n_102),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_99),
.A2(n_26),
.B1(n_49),
.B2(n_48),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_105),
.A2(n_4),
.B(n_5),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_121),
.B(n_129),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_122),
.A2(n_132),
.B1(n_11),
.B2(n_12),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_105),
.B(n_46),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_124),
.B(n_128),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_126),
.B(n_134),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_114),
.B(n_103),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_114),
.B(n_6),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_130),
.B(n_133),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_107),
.A2(n_41),
.B1(n_36),
.B2(n_35),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_115),
.B(n_7),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_117),
.B(n_7),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_113),
.Y(n_135)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_135),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_116),
.B(n_8),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_138),
.B(n_139),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_105),
.B(n_32),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_140),
.A2(n_12),
.B(n_139),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_106),
.B(n_8),
.Y(n_141)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_141),
.Y(n_146)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_118),
.Y(n_142)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_142),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_124),
.B(n_14),
.C(n_10),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_148),
.B(n_155),
.C(n_157),
.Y(n_161)
);

NOR3xp33_ASAP7_75t_SL g149 ( 
.A(n_131),
.B(n_9),
.C(n_11),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_149),
.B(n_153),
.Y(n_159)
);

NOR2x1_ASAP7_75t_L g150 ( 
.A(n_123),
.B(n_9),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_150),
.B(n_154),
.Y(n_163)
);

INVxp33_ASAP7_75t_L g152 ( 
.A(n_136),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_152),
.B(n_156),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_SL g155 ( 
.A(n_121),
.B(n_132),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_127),
.B(n_129),
.Y(n_157)
);

INVx2_ASAP7_75t_SL g160 ( 
.A(n_152),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_160),
.B(n_166),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_145),
.A2(n_125),
.B1(n_142),
.B2(n_137),
.Y(n_162)
);

CKINVDCx14_ASAP7_75t_R g170 ( 
.A(n_162),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_144),
.B(n_140),
.C(n_127),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_164),
.B(n_143),
.Y(n_167)
);

OAI32xp33_ASAP7_75t_L g165 ( 
.A1(n_158),
.A2(n_137),
.A3(n_147),
.B1(n_157),
.B2(n_155),
.Y(n_165)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_165),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_167),
.B(n_161),
.C(n_166),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_168),
.B(n_151),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_171),
.B(n_172),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_173),
.A2(n_169),
.B(n_163),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_174),
.Y(n_175)
);

NAND3xp33_ASAP7_75t_L g176 ( 
.A(n_175),
.B(n_163),
.C(n_146),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_176),
.B(n_159),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_177),
.A2(n_167),
.B(n_170),
.Y(n_178)
);


endmodule