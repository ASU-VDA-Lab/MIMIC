module real_jpeg_6869_n_13 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_13);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_13;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_215;
wire n_166;
wire n_176;
wire n_221;
wire n_104;
wire n_194;
wire n_153;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_184;
wire n_56;
wire n_164;
wire n_48;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_242;
wire n_141;
wire n_139;
wire n_33;
wire n_65;
wire n_188;
wire n_142;
wire n_175;
wire n_178;
wire n_76;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_195;
wire n_110;
wire n_61;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_150;
wire n_32;
wire n_20;
wire n_80;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_240;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_187;
wire n_75;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_167;
wire n_202;
wire n_128;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_253;
wire n_96;
wire n_89;
wire n_16;

INVx8_ASAP7_75t_L g55 ( 
.A(n_0),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_1),
.A2(n_67),
.B1(n_96),
.B2(n_97),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_1),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_1),
.A2(n_96),
.B1(n_162),
.B2(n_164),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_1),
.A2(n_96),
.B1(n_207),
.B2(n_211),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_2),
.A2(n_179),
.B1(n_182),
.B2(n_183),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_2),
.Y(n_183)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_4),
.A2(n_102),
.B1(n_104),
.B2(n_109),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_4),
.Y(n_109)
);

OAI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_4),
.A2(n_109),
.B1(n_207),
.B2(n_211),
.Y(n_206)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_5),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g36 ( 
.A1(n_6),
.A2(n_37),
.B1(n_43),
.B2(n_44),
.Y(n_36)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_6),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_6),
.A2(n_43),
.B1(n_143),
.B2(n_144),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_6),
.A2(n_43),
.B1(n_152),
.B2(n_155),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_7),
.Y(n_216)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_7),
.Y(n_230)
);

INVx8_ASAP7_75t_L g244 ( 
.A(n_7),
.Y(n_244)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_8),
.Y(n_172)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_8),
.Y(n_176)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_9),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_10),
.B(n_62),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_10),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_10),
.A2(n_139),
.B1(n_154),
.B2(n_195),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_10),
.B(n_202),
.C(n_203),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_10),
.B(n_127),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_10),
.B(n_229),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_10),
.B(n_100),
.Y(n_236)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_11),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_11),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g20 ( 
.A1(n_12),
.A2(n_21),
.B1(n_24),
.B2(n_25),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

XOR2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_189),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_187),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_146),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_16),
.B(n_146),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_73),
.C(n_110),
.Y(n_16)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_17),
.B(n_252),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_46),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_18),
.B(n_46),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_27),
.B(n_30),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_20),
.A2(n_31),
.B1(n_178),
.B2(n_184),
.Y(n_177)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

BUFx8_ASAP7_75t_L g92 ( 
.A(n_23),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_26),
.Y(n_91)
);

BUFx5_ASAP7_75t_L g203 ( 
.A(n_26),
.Y(n_203)
);

INVx3_ASAP7_75t_SL g27 ( 
.A(n_28),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_29),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_30),
.A2(n_234),
.B(n_235),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_36),
.Y(n_30)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_31),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_31),
.A2(n_240),
.B1(n_241),
.B2(n_242),
.Y(n_239)
);

OR2x2_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_33),
.Y(n_31)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_36),
.B(n_215),
.Y(n_214)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_41),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_42),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g181 ( 
.A(n_42),
.Y(n_181)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx8_ASAP7_75t_L g212 ( 
.A(n_45),
.Y(n_212)
);

AOI32xp33_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_51),
.A3(n_56),
.B1(n_61),
.B2(n_65),
.Y(n_46)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_49),
.Y(n_173)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

BUFx5_ASAP7_75t_L g126 ( 
.A(n_50),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_50),
.Y(n_138)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_54),
.Y(n_103)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_54),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_54),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_54),
.Y(n_154)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_55),
.Y(n_86)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_55),
.Y(n_108)
);

BUFx5_ASAP7_75t_L g157 ( 
.A(n_55),
.Y(n_157)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx2_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_59),
.Y(n_115)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_59),
.Y(n_129)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_60),
.Y(n_72)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_60),
.Y(n_123)
);

INVxp33_ASAP7_75t_L g140 ( 
.A(n_61),
.Y(n_140)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_64),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_64),
.Y(n_144)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_64),
.Y(n_165)
);

NAND2xp33_ASAP7_75t_SL g65 ( 
.A(n_66),
.B(n_70),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_69),
.Y(n_78)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_69),
.Y(n_200)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_73),
.A2(n_110),
.B1(n_111),
.B2(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_73),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_74),
.A2(n_95),
.B1(n_99),
.B2(n_101),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_74),
.A2(n_101),
.B(n_150),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_74),
.A2(n_150),
.B(n_194),
.Y(n_193)
);

INVx2_ASAP7_75t_SL g74 ( 
.A(n_75),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_75),
.B(n_151),
.Y(n_220)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_87),
.Y(n_75)
);

OAI22xp33_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_79),
.B1(n_82),
.B2(n_85),
.Y(n_76)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_81),
.Y(n_84)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_81),
.Y(n_94)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_86),
.Y(n_98)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_87),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_87),
.A2(n_95),
.B(n_220),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_91),
.B1(n_92),
.B2(n_93),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_89),
.Y(n_202)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

BUFx2_ASAP7_75t_L g182 ( 
.A(n_92),
.Y(n_182)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_100),
.B(n_151),
.Y(n_150)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx5_ASAP7_75t_SL g105 ( 
.A(n_106),
.Y(n_105)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_112),
.A2(n_134),
.B(n_141),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_112),
.B(n_167),
.Y(n_166)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

OR2x2_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_127),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_115),
.A2(n_116),
.B1(n_119),
.B2(n_124),
.Y(n_114)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx5_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_SL g119 ( 
.A(n_120),
.Y(n_119)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_125),
.A2(n_171),
.B1(n_173),
.B2(n_174),
.Y(n_170)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g143 ( 
.A(n_126),
.Y(n_143)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_127),
.Y(n_145)
);

AO22x2_ASAP7_75t_L g127 ( 
.A1(n_128),
.A2(n_129),
.B1(n_130),
.B2(n_133),
.Y(n_127)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx3_ASAP7_75t_SL g130 ( 
.A(n_131),
.Y(n_130)
);

INVx8_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g196 ( 
.A(n_133),
.Y(n_196)
);

OAI21xp33_ASAP7_75t_SL g134 ( 
.A1(n_135),
.A2(n_139),
.B(n_140),
.Y(n_134)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_138),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_139),
.B(n_170),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_139),
.A2(n_213),
.B(n_214),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_145),
.Y(n_141)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_142),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_145),
.A2(n_161),
.B(n_166),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_147),
.A2(n_148),
.B1(n_159),
.B2(n_186),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_SL g148 ( 
.A(n_149),
.B(n_158),
.Y(n_148)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx11_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx5_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_159),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_SL g159 ( 
.A(n_160),
.B(n_168),
.Y(n_159)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_177),
.Y(n_168)
);

INVx5_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx6_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_SL g179 ( 
.A(n_180),
.Y(n_179)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_190),
.A2(n_249),
.B(n_254),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_191),
.A2(n_223),
.B(n_248),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_204),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_192),
.B(n_204),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_193),
.B(n_197),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_193),
.A2(n_197),
.B1(n_198),
.B2(n_246),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_193),
.Y(n_246)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_201),
.Y(n_198)
);

HB1xp67_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_217),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_205),
.B(n_218),
.C(n_222),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_206),
.A2(n_213),
.B(n_214),
.Y(n_205)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_206),
.Y(n_241)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx6_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_211),
.Y(n_227)
);

INVx4_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx4_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_218),
.A2(n_219),
.B1(n_221),
.B2(n_222),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_224),
.A2(n_238),
.B(n_247),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_225),
.A2(n_232),
.B(n_237),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_231),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_228),
.Y(n_226)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_230),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_233),
.B(n_236),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_233),
.B(n_236),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_234),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_245),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_239),
.B(n_245),
.Y(n_247)
);

INVx4_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_251),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_250),
.B(n_251),
.Y(n_254)
);


endmodule