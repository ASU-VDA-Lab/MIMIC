module fake_jpeg_14430_n_350 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_350);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_350;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_16),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_SL g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_7),
.Y(n_25)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_13),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_3),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_10),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

INVx11_ASAP7_75t_SL g37 ( 
.A(n_15),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_17),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_11),
.Y(n_39)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_0),
.B(n_12),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_43),
.Y(n_82)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_45),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_46),
.Y(n_88)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_23),
.Y(n_47)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_47),
.Y(n_80)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_26),
.Y(n_48)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_48),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_24),
.A2(n_9),
.B1(n_16),
.B2(n_2),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_49),
.A2(n_24),
.B1(n_38),
.B2(n_35),
.Y(n_71)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_23),
.Y(n_50)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_50),
.Y(n_101)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_27),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_22),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_52),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_22),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_53),
.Y(n_110)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_54),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_22),
.Y(n_55)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_55),
.Y(n_75)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_32),
.Y(n_56)
);

HB1xp67_ASAP7_75t_L g78 ( 
.A(n_56),
.Y(n_78)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_27),
.Y(n_57)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_57),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_58),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_59),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_41),
.B(n_9),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_60),
.B(n_67),
.Y(n_74)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_27),
.Y(n_61)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_61),
.Y(n_94)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_27),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g103 ( 
.A(n_62),
.Y(n_103)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_27),
.Y(n_63)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_63),
.Y(n_72)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_64),
.Y(n_111)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_65),
.B(n_68),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_28),
.Y(n_66)
);

BUFx4f_ASAP7_75t_SL g106 ( 
.A(n_66),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_41),
.B(n_9),
.Y(n_67)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_29),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_28),
.Y(n_69)
);

BUFx12_ASAP7_75t_L g104 ( 
.A(n_69),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_71),
.A2(n_85),
.B1(n_87),
.B2(n_90),
.Y(n_130)
);

OR2x2_ASAP7_75t_L g79 ( 
.A(n_43),
.B(n_42),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_79),
.B(n_91),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_56),
.B(n_20),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_81),
.B(n_83),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_R g83 ( 
.A(n_44),
.B(n_20),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_45),
.B(n_19),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_84),
.B(n_95),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_57),
.A2(n_24),
.B1(n_28),
.B2(n_26),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_47),
.A2(n_36),
.B1(n_34),
.B2(n_29),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_86),
.A2(n_93),
.B1(n_97),
.B2(n_5),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_50),
.A2(n_36),
.B1(n_34),
.B2(n_29),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_68),
.A2(n_36),
.B1(n_34),
.B2(n_42),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_62),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_52),
.A2(n_18),
.B1(n_33),
.B2(n_35),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_54),
.B(n_38),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_65),
.A2(n_19),
.B1(n_31),
.B2(n_30),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_66),
.B(n_31),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_98),
.B(n_102),
.Y(n_125)
);

BUFx16f_ASAP7_75t_L g100 ( 
.A(n_63),
.Y(n_100)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_100),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_69),
.B(n_25),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_46),
.B(n_25),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_108),
.B(n_76),
.Y(n_131)
);

OR2x2_ASAP7_75t_L g109 ( 
.A(n_48),
.B(n_18),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_109),
.B(n_112),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_64),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_61),
.A2(n_26),
.B1(n_37),
.B2(n_30),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_113),
.A2(n_37),
.B1(n_55),
.B2(n_46),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_51),
.B(n_33),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_114),
.B(n_17),
.Y(n_148)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_78),
.Y(n_116)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_116),
.Y(n_160)
);

INVx5_ASAP7_75t_L g117 ( 
.A(n_73),
.Y(n_117)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_117),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_79),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_118),
.B(n_119),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_109),
.Y(n_119)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_82),
.Y(n_122)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_122),
.Y(n_190)
);

OAI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_71),
.A2(n_113),
.B1(n_85),
.B2(n_93),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_123),
.A2(n_141),
.B1(n_151),
.B2(n_75),
.Y(n_171)
);

AO22x1_ASAP7_75t_L g124 ( 
.A1(n_99),
.A2(n_59),
.B1(n_58),
.B2(n_53),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_124),
.A2(n_134),
.B(n_106),
.Y(n_163)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_70),
.Y(n_126)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_126),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_104),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_127),
.B(n_128),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_104),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_129),
.A2(n_73),
.B1(n_77),
.B2(n_110),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_131),
.B(n_132),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_104),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_89),
.A2(n_53),
.B1(n_10),
.B2(n_2),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_88),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g169 ( 
.A(n_135),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_111),
.A2(n_0),
.B1(n_1),
.B2(n_4),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_136),
.Y(n_157)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_80),
.Y(n_138)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_138),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_101),
.B(n_1),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_139),
.B(n_147),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_89),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_140),
.B(n_146),
.Y(n_170)
);

OAI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_90),
.A2(n_10),
.B1(n_4),
.B2(n_5),
.Y(n_141)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_107),
.Y(n_142)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_142),
.Y(n_174)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_107),
.Y(n_143)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_143),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_100),
.Y(n_144)
);

INVxp33_ASAP7_75t_L g166 ( 
.A(n_144),
.Y(n_166)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_111),
.Y(n_145)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_145),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_74),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_96),
.B(n_1),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_148),
.Y(n_159)
);

BUFx2_ASAP7_75t_L g149 ( 
.A(n_88),
.Y(n_149)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_149),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_106),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_150),
.Y(n_164)
);

OAI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_92),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_151)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_152),
.B(n_115),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_106),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_153),
.B(n_73),
.Y(n_177)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_77),
.Y(n_154)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_154),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_120),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_156),
.B(n_175),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_152),
.A2(n_105),
.B1(n_96),
.B2(n_75),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_162),
.A2(n_165),
.B1(n_167),
.B2(n_171),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_163),
.B(n_117),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_115),
.A2(n_131),
.B1(n_140),
.B2(n_119),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_122),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_137),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_176),
.B(n_180),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_177),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_116),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_125),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_183),
.B(n_126),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_130),
.A2(n_105),
.B1(n_110),
.B2(n_92),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_L g213 ( 
.A1(n_184),
.A2(n_186),
.B1(n_188),
.B2(n_149),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_185),
.A2(n_187),
.B1(n_149),
.B2(n_133),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_121),
.A2(n_94),
.B1(n_72),
.B2(n_103),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_L g187 ( 
.A1(n_118),
.A2(n_94),
.B1(n_72),
.B2(n_103),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_121),
.A2(n_103),
.B1(n_11),
.B2(n_13),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_158),
.A2(n_153),
.B(n_139),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g234 ( 
.A1(n_191),
.A2(n_201),
.B(n_202),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_170),
.B(n_146),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_192),
.B(n_200),
.Y(n_228)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_190),
.Y(n_193)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_193),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_168),
.B(n_178),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_194),
.B(n_197),
.Y(n_237)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_190),
.Y(n_195)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_195),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_165),
.B(n_145),
.C(n_128),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_196),
.B(n_214),
.C(n_220),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_168),
.B(n_147),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_170),
.B(n_134),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_158),
.A2(n_150),
.B(n_132),
.Y(n_201)
);

INVx8_ASAP7_75t_L g204 ( 
.A(n_166),
.Y(n_204)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_204),
.Y(n_236)
);

XOR2x1_ASAP7_75t_L g205 ( 
.A(n_178),
.B(n_124),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_SL g229 ( 
.A(n_205),
.B(n_171),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_156),
.B(n_138),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_206),
.B(n_207),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_176),
.B(n_154),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_208),
.B(n_216),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_173),
.A2(n_127),
.B(n_133),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_209),
.B(n_186),
.Y(n_226)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_160),
.Y(n_210)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_210),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_212),
.A2(n_217),
.B1(n_162),
.B2(n_164),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_213),
.A2(n_223),
.B1(n_157),
.B2(n_181),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_173),
.B(n_143),
.C(n_142),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_167),
.B(n_183),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_215),
.B(n_221),
.Y(n_238)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_160),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_167),
.A2(n_124),
.B1(n_135),
.B2(n_14),
.Y(n_217)
);

BUFx12f_ASAP7_75t_L g218 ( 
.A(n_169),
.Y(n_218)
);

BUFx5_ASAP7_75t_L g230 ( 
.A(n_218),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_159),
.B(n_8),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_219),
.B(n_188),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_167),
.B(n_8),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_177),
.B(n_13),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_189),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_222),
.B(n_179),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_L g223 ( 
.A1(n_184),
.A2(n_14),
.B1(n_15),
.B2(n_17),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_226),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_227),
.B(n_244),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_229),
.B(n_199),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_198),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_231),
.B(n_241),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_235),
.A2(n_248),
.B1(n_212),
.B2(n_195),
.Y(n_260)
);

OR2x2_ASAP7_75t_L g240 ( 
.A(n_215),
.B(n_163),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_240),
.A2(n_252),
.B(n_202),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_203),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_243),
.A2(n_211),
.B1(n_201),
.B2(n_191),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_192),
.B(n_189),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_194),
.B(n_182),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_245),
.B(n_247),
.C(n_225),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_204),
.B(n_161),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_246),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_196),
.B(n_182),
.C(n_155),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_199),
.A2(n_181),
.B1(n_179),
.B2(n_169),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_249),
.B(n_251),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_200),
.B(n_161),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_250),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_221),
.Y(n_251)
);

OR2x2_ASAP7_75t_L g252 ( 
.A(n_205),
.B(n_161),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_253),
.B(n_271),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_254),
.A2(n_238),
.B1(n_242),
.B2(n_224),
.Y(n_289)
);

AO21x1_ASAP7_75t_L g256 ( 
.A1(n_240),
.A2(n_202),
.B(n_209),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_256),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_243),
.A2(n_211),
.B1(n_197),
.B2(n_217),
.Y(n_259)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_259),
.Y(n_277)
);

AND2x2_ASAP7_75t_L g287 ( 
.A(n_260),
.B(n_270),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_245),
.B(n_220),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_261),
.B(n_268),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_L g281 ( 
.A1(n_262),
.A2(n_252),
.B(n_240),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_237),
.B(n_214),
.Y(n_263)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_263),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_248),
.A2(n_193),
.B1(n_216),
.B2(n_210),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_264),
.B(n_266),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_226),
.A2(n_222),
.B1(n_169),
.B2(n_174),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_235),
.A2(n_174),
.B1(n_155),
.B2(n_172),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_267),
.B(n_269),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_225),
.B(n_172),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_229),
.A2(n_14),
.B1(n_218),
.B2(n_251),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_247),
.A2(n_218),
.B1(n_228),
.B2(n_238),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_237),
.B(n_218),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_272),
.B(n_241),
.Y(n_279)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_232),
.Y(n_275)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_275),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_279),
.B(n_272),
.C(n_268),
.Y(n_294)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_281),
.Y(n_298)
);

AOI21xp33_ASAP7_75t_L g283 ( 
.A1(n_274),
.A2(n_228),
.B(n_265),
.Y(n_283)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_283),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_262),
.A2(n_252),
.B(n_234),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_285),
.B(n_288),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_255),
.B(n_231),
.Y(n_286)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_286),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_274),
.A2(n_234),
.B(n_224),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_289),
.A2(n_258),
.B1(n_266),
.B2(n_257),
.Y(n_299)
);

INVx1_ASAP7_75t_SL g290 ( 
.A(n_256),
.Y(n_290)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_290),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_SL g292 ( 
.A1(n_269),
.A2(n_236),
.B(n_232),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_292),
.B(n_264),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_294),
.B(n_280),
.C(n_288),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_282),
.B(n_270),
.C(n_263),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_297),
.B(n_301),
.C(n_277),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_299),
.B(n_307),
.Y(n_317)
);

OR2x2_ASAP7_75t_L g309 ( 
.A(n_300),
.B(n_308),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_282),
.B(n_261),
.C(n_271),
.Y(n_301)
);

XNOR2x1_ASAP7_75t_L g302 ( 
.A(n_280),
.B(n_253),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_302),
.B(n_289),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_284),
.B(n_258),
.Y(n_304)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_304),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_287),
.A2(n_260),
.B1(n_275),
.B2(n_242),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_305),
.A2(n_278),
.B1(n_290),
.B2(n_276),
.Y(n_310)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_293),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_278),
.B(n_292),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_310),
.B(n_319),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_311),
.B(n_313),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_312),
.B(n_318),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_294),
.B(n_273),
.C(n_287),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_314),
.B(n_305),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_306),
.B(n_249),
.Y(n_315)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_315),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_296),
.B(n_287),
.C(n_276),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_297),
.B(n_285),
.C(n_281),
.Y(n_319)
);

MAJx2_ASAP7_75t_L g320 ( 
.A(n_301),
.B(n_295),
.C(n_302),
.Y(n_320)
);

AOI21xp33_ASAP7_75t_L g327 ( 
.A1(n_320),
.A2(n_304),
.B(n_308),
.Y(n_327)
);

AO221x1_ASAP7_75t_L g322 ( 
.A1(n_315),
.A2(n_298),
.B1(n_233),
.B2(n_239),
.C(n_236),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_L g335 ( 
.A1(n_322),
.A2(n_325),
.B(n_327),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_323),
.B(n_309),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_L g325 ( 
.A1(n_309),
.A2(n_295),
.B(n_298),
.Y(n_325)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_317),
.Y(n_329)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_329),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_330),
.B(n_331),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_328),
.B(n_299),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_326),
.B(n_312),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_332),
.B(n_333),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_326),
.B(n_320),
.C(n_300),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_321),
.B(n_316),
.Y(n_336)
);

CKINVDCx14_ASAP7_75t_R g339 ( 
.A(n_336),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_333),
.B(n_324),
.C(n_323),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_338),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_335),
.A2(n_325),
.B1(n_303),
.B2(n_291),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_L g342 ( 
.A1(n_341),
.A2(n_303),
.B1(n_334),
.B2(n_291),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_342),
.A2(n_344),
.B1(n_341),
.B2(n_337),
.Y(n_346)
);

BUFx24_ASAP7_75t_SL g344 ( 
.A(n_339),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_343),
.B(n_340),
.C(n_338),
.Y(n_345)
);

AOI21xp5_ASAP7_75t_L g347 ( 
.A1(n_345),
.A2(n_346),
.B(n_330),
.Y(n_347)
);

AOI221xp5_ASAP7_75t_L g348 ( 
.A1(n_347),
.A2(n_324),
.B1(n_233),
.B2(n_239),
.C(n_267),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_348),
.B(n_230),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_349),
.B(n_230),
.Y(n_350)
);


endmodule