module real_jpeg_22681_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_64;
wire n_177;
wire n_131;
wire n_47;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_105;
wire n_40;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_126;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_148;
wire n_19;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_192;
wire n_203;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_202;
wire n_167;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_181;
wire n_85;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_0),
.A2(n_41),
.B1(n_42),
.B2(n_57),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_0),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_0),
.A2(n_57),
.B1(n_65),
.B2(n_66),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_0),
.A2(n_28),
.B1(n_29),
.B2(n_57),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g30 ( 
.A1(n_1),
.A2(n_28),
.B1(n_29),
.B2(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_2),
.A2(n_41),
.B1(n_42),
.B2(n_45),
.Y(n_40)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_2),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_2),
.A2(n_28),
.B1(n_29),
.B2(n_45),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_3),
.A2(n_65),
.B1(n_66),
.B2(n_72),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_3),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_3),
.A2(n_28),
.B1(n_29),
.B2(n_72),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_3),
.A2(n_41),
.B1(n_42),
.B2(n_72),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_4),
.A2(n_75),
.B1(n_82),
.B2(n_83),
.Y(n_81)
);

CKINVDCx14_ASAP7_75t_R g82 ( 
.A(n_4),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_4),
.A2(n_65),
.B1(n_66),
.B2(n_82),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_4),
.A2(n_41),
.B1(n_42),
.B2(n_82),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_4),
.A2(n_28),
.B1(n_29),
.B2(n_82),
.Y(n_148)
);

BUFx16f_ASAP7_75t_L g75 ( 
.A(n_5),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_6),
.A2(n_65),
.B1(n_66),
.B2(n_70),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_6),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_6),
.A2(n_70),
.B1(n_75),
.B2(n_83),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_6),
.A2(n_28),
.B1(n_29),
.B2(n_70),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_6),
.A2(n_41),
.B1(n_42),
.B2(n_70),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_7),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_7),
.B(n_80),
.Y(n_116)
);

AOI21xp33_ASAP7_75t_L g139 ( 
.A1(n_7),
.A2(n_14),
.B(n_29),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_7),
.A2(n_41),
.B1(n_42),
.B2(n_76),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_7),
.A2(n_26),
.B1(n_90),
.B2(n_148),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_7),
.B(n_120),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_7),
.B(n_65),
.Y(n_174)
);

AOI21xp33_ASAP7_75t_L g178 ( 
.A1(n_7),
.A2(n_65),
.B(n_174),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_8),
.B(n_28),
.Y(n_27)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_8),
.Y(n_90)
);

BUFx8_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_L g35 ( 
.A1(n_10),
.A2(n_28),
.B1(n_29),
.B2(n_36),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_10),
.Y(n_36)
);

OAI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_10),
.A2(n_36),
.B1(n_41),
.B2(n_42),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_11),
.Y(n_66)
);

INVx13_ASAP7_75t_L g64 ( 
.A(n_12),
.Y(n_64)
);

INVx13_ASAP7_75t_L g78 ( 
.A(n_13),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_13),
.A2(n_65),
.B1(n_66),
.B2(n_78),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_14),
.A2(n_28),
.B1(n_29),
.B2(n_39),
.Y(n_38)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

A2O1A1Ixp33_ASAP7_75t_L g49 ( 
.A1(n_14),
.A2(n_38),
.B(n_41),
.C(n_50),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_14),
.B(n_41),
.Y(n_50)
);

INVx11_ASAP7_75t_SL g44 ( 
.A(n_15),
.Y(n_44)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_124),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_122),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_19),
.Y(n_18)
);

AND2x2_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_105),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_20),
.B(n_105),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_84),
.B2(n_104),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_52),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_37),
.B2(n_51),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_30),
.B(n_32),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_26),
.A2(n_30),
.B1(n_89),
.B2(n_90),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_26),
.A2(n_34),
.B1(n_132),
.B2(n_148),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_26),
.A2(n_135),
.B(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_27),
.B(n_115),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_27),
.A2(n_131),
.B1(n_133),
.B2(n_134),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_27),
.A2(n_33),
.B(n_166),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_28),
.B(n_152),
.Y(n_151)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_35),
.Y(n_33)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_34),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_35),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_37),
.Y(n_51)
);

OAI21xp5_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_40),
.B(n_46),
.Y(n_37)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_38),
.A2(n_49),
.B1(n_142),
.B2(n_143),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_38),
.B(n_76),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_38),
.A2(n_49),
.B1(n_143),
.B2(n_163),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_38),
.A2(n_49),
.B1(n_163),
.B2(n_181),
.Y(n_180)
);

A2O1A1Ixp33_ASAP7_75t_L g138 ( 
.A1(n_39),
.A2(n_42),
.B(n_76),
.C(n_139),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_41),
.A2(n_42),
.B1(n_63),
.B2(n_64),
.Y(n_68)
);

AOI32xp33_ASAP7_75t_L g173 ( 
.A1(n_41),
.A2(n_64),
.A3(n_66),
.B1(n_174),
.B2(n_175),
.Y(n_173)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

NAND2xp33_ASAP7_75t_SL g175 ( 
.A(n_42),
.B(n_63),
.Y(n_175)
);

BUFx10_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_48),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_47),
.B(n_59),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_SL g54 ( 
.A1(n_49),
.A2(n_55),
.B(n_58),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_49),
.A2(n_181),
.B(n_197),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_60),
.C(n_73),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_53),
.A2(n_54),
.B1(n_60),
.B2(n_61),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g53 ( 
.A(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_56),
.B(n_59),
.Y(n_197)
);

CKINVDCx14_ASAP7_75t_R g60 ( 
.A(n_61),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_62),
.A2(n_68),
.B1(n_69),
.B2(n_71),
.Y(n_61)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_62),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_62),
.A2(n_68),
.B1(n_119),
.B2(n_178),
.Y(n_177)
);

A2O1A1Ixp33_ASAP7_75t_L g62 ( 
.A1(n_63),
.A2(n_65),
.B(n_67),
.C(n_68),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_63),
.B(n_65),
.Y(n_67)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_65),
.B(n_78),
.Y(n_87)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_66),
.A2(n_74),
.B1(n_79),
.B2(n_87),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_68),
.B(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_68),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_69),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_71),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_SL g106 ( 
.A(n_73),
.B(n_107),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_77),
.B1(n_80),
.B2(n_81),
.Y(n_73)
);

HAxp5_ASAP7_75t_SL g74 ( 
.A(n_75),
.B(n_76),
.CON(n_74),
.SN(n_74)
);

O2A1O1Ixp33_ASAP7_75t_L g77 ( 
.A1(n_75),
.A2(n_78),
.B(n_79),
.C(n_80),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_75),
.B(n_78),
.Y(n_79)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_75),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_76),
.B(n_90),
.Y(n_152)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_77),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_80),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_81),
.Y(n_95)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_84),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_91),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_88),
.Y(n_85)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_86),
.B(n_88),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_89),
.A2(n_90),
.B(n_114),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_92),
.A2(n_93),
.B1(n_98),
.B2(n_99),
.Y(n_91)
);

CKINVDCx14_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_94),
.A2(n_95),
.B1(n_96),
.B2(n_97),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_99),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_100),
.A2(n_101),
.B(n_102),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_100),
.A2(n_118),
.B1(n_120),
.B2(n_121),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_108),
.C(n_110),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_106),
.B(n_202),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_108),
.A2(n_109),
.B1(n_110),
.B2(n_111),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_109),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_111),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_116),
.C(n_117),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_112),
.A2(n_113),
.B1(n_116),
.B2(n_192),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_113),
.Y(n_112)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_116),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_SL g190 ( 
.A(n_117),
.B(n_191),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_125),
.A2(n_199),
.B(n_203),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_126),
.A2(n_186),
.B(n_198),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_168),
.B(n_185),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_128),
.A2(n_155),
.B(n_167),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_144),
.B(n_154),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_136),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_130),
.B(n_136),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_132),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_133),
.B(n_166),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_135),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_137),
.A2(n_138),
.B1(n_140),
.B2(n_141),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_138),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_138),
.B(n_140),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_141),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_145),
.A2(n_149),
.B(n_153),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_147),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_146),
.B(n_147),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_150),
.B(n_151),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_157),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_156),
.B(n_157),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_164),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_160),
.B1(n_161),
.B2(n_162),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_159),
.B(n_162),
.C(n_164),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_160),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_162),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_170),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_169),
.B(n_170),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_171),
.A2(n_176),
.B1(n_183),
.B2(n_184),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_171),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_173),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_172),
.B(n_173),
.Y(n_195)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_176),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_179),
.B1(n_180),
.B2(n_182),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_177),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_179),
.B(n_182),
.C(n_183),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_180),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_188),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_187),
.B(n_188),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_189),
.A2(n_190),
.B1(n_193),
.B2(n_194),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_189),
.B(n_195),
.C(n_196),
.Y(n_200)
);

CKINVDCx14_ASAP7_75t_R g189 ( 
.A(n_190),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_194),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_196),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_201),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_200),
.B(n_201),
.Y(n_203)
);


endmodule