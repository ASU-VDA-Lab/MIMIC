module fake_jpeg_13563_n_332 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_332);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_332;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_15),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

CKINVDCx14_ASAP7_75t_R g33 ( 
.A(n_14),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_1),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

BUFx16f_ASAP7_75t_L g39 ( 
.A(n_11),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

INVx13_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

BUFx4f_ASAP7_75t_SL g92 ( 
.A(n_41),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g97 ( 
.A(n_42),
.Y(n_97)
);

BUFx2_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_43),
.Y(n_87)
);

HAxp5_ASAP7_75t_SL g44 ( 
.A(n_33),
.B(n_8),
.CON(n_44),
.SN(n_44)
);

HAxp5_ASAP7_75t_SL g80 ( 
.A(n_44),
.B(n_54),
.CON(n_80),
.SN(n_80)
);

INVx13_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_33),
.B(n_8),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_46),
.B(n_21),
.Y(n_66)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_47),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g104 ( 
.A(n_48),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_26),
.B(n_0),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_49),
.B(n_58),
.Y(n_79)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_19),
.Y(n_50)
);

INVx11_ASAP7_75t_L g88 ( 
.A(n_50),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_26),
.B(n_32),
.Y(n_51)
);

A2O1A1Ixp33_ASAP7_75t_L g96 ( 
.A1(n_51),
.A2(n_24),
.B(n_16),
.C(n_27),
.Y(n_96)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_26),
.Y(n_52)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_52),
.Y(n_68)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_53),
.Y(n_108)
);

BUFx24_ASAP7_75t_L g54 ( 
.A(n_20),
.Y(n_54)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_54),
.Y(n_99)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_20),
.Y(n_55)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_32),
.Y(n_56)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_56),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_57),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_22),
.B(n_0),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_59),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_60),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_46),
.B(n_28),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_61),
.B(n_62),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_49),
.B(n_28),
.Y(n_62)
);

NAND2xp33_ASAP7_75t_SL g63 ( 
.A(n_51),
.B(n_20),
.Y(n_63)
);

NAND2x1_ASAP7_75t_SL g139 ( 
.A(n_63),
.B(n_66),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_54),
.A2(n_17),
.B1(n_22),
.B2(n_31),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_64),
.A2(n_67),
.B1(n_72),
.B2(n_100),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_51),
.A2(n_31),
.B1(n_22),
.B2(n_29),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_57),
.Y(n_70)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_70),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_40),
.B(n_21),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_71),
.B(n_81),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_43),
.A2(n_31),
.B1(n_29),
.B2(n_38),
.Y(n_72)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_57),
.Y(n_75)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_75),
.Y(n_113)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_77),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_80),
.A2(n_25),
.B1(n_36),
.B2(n_63),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_58),
.B(n_18),
.Y(n_81)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_55),
.Y(n_82)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_82),
.Y(n_130)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_47),
.Y(n_83)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_83),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_50),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_84),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_52),
.A2(n_29),
.B1(n_38),
.B2(n_17),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_85),
.A2(n_89),
.B1(n_23),
.B2(n_1),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_53),
.A2(n_29),
.B1(n_38),
.B2(n_17),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_56),
.B(n_30),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_91),
.B(n_94),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_48),
.Y(n_93)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_93),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_42),
.B(n_30),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_59),
.B(n_18),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_95),
.B(n_96),
.Y(n_126)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_54),
.Y(n_98)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_98),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_43),
.A2(n_35),
.B1(n_38),
.B2(n_24),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_60),
.B(n_37),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_101),
.B(n_103),
.Y(n_134)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_60),
.Y(n_102)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_102),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_48),
.B(n_37),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_41),
.B(n_39),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_105),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_41),
.B(n_36),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_106),
.A2(n_107),
.B1(n_39),
.B2(n_23),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_45),
.A2(n_35),
.B1(n_24),
.B2(n_27),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_109),
.Y(n_162)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_65),
.Y(n_111)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_111),
.Y(n_155)
);

A2O1A1Ixp33_ASAP7_75t_L g112 ( 
.A1(n_79),
.A2(n_39),
.B(n_25),
.C(n_45),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_112),
.B(n_92),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_114),
.Y(n_166)
);

BUFx4f_ASAP7_75t_L g115 ( 
.A(n_92),
.Y(n_115)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_115),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_64),
.A2(n_39),
.B1(n_9),
.B2(n_11),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_117),
.A2(n_118),
.B1(n_128),
.B2(n_141),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_100),
.A2(n_39),
.B1(n_23),
.B2(n_8),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_124),
.B(n_129),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_76),
.B(n_23),
.C(n_7),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_125),
.B(n_138),
.C(n_102),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_85),
.A2(n_23),
.B1(n_1),
.B2(n_2),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_127),
.A2(n_136),
.B(n_141),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_96),
.A2(n_7),
.B1(n_14),
.B2(n_13),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_68),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_129),
.A2(n_99),
.B1(n_98),
.B2(n_69),
.Y(n_146)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_86),
.Y(n_132)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_132),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_80),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_108),
.B(n_5),
.C(n_6),
.Y(n_138)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_87),
.Y(n_140)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_140),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_107),
.A2(n_5),
.B1(n_9),
.B2(n_12),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_75),
.A2(n_69),
.B1(n_70),
.B2(n_83),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_142),
.A2(n_110),
.B1(n_118),
.B2(n_113),
.Y(n_175)
);

OR2x2_ASAP7_75t_L g183 ( 
.A(n_144),
.B(n_130),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_120),
.B(n_78),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_145),
.B(n_149),
.Y(n_202)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_146),
.B(n_159),
.Y(n_210)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_111),
.Y(n_147)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_147),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_135),
.Y(n_148)
);

BUFx3_ASAP7_75t_L g194 ( 
.A(n_148),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_122),
.B(n_92),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_126),
.B(n_77),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_150),
.B(n_154),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_122),
.B(n_78),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_151),
.B(n_156),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_135),
.Y(n_152)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_152),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_153),
.B(n_143),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_126),
.B(n_73),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_131),
.B(n_97),
.Y(n_156)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_132),
.Y(n_161)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_161),
.Y(n_190)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_116),
.Y(n_163)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_163),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_134),
.B(n_119),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_165),
.B(n_172),
.Y(n_184)
);

INVx8_ASAP7_75t_L g167 ( 
.A(n_115),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_167),
.Y(n_201)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_115),
.Y(n_168)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_168),
.Y(n_205)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_116),
.Y(n_169)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_169),
.Y(n_208)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_113),
.Y(n_170)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_170),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_124),
.A2(n_90),
.B1(n_93),
.B2(n_87),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_171),
.B(n_146),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_123),
.B(n_13),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_134),
.B(n_97),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_173),
.B(n_174),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_120),
.B(n_97),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_175),
.A2(n_133),
.B1(n_142),
.B2(n_74),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_138),
.B(n_125),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_176),
.B(n_181),
.Y(n_213)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_121),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_177),
.Y(n_212)
);

NAND2x1p5_ASAP7_75t_L g178 ( 
.A(n_112),
.B(n_73),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_178),
.A2(n_158),
.B(n_160),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_139),
.B(n_88),
.C(n_104),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_179),
.B(n_130),
.C(n_143),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_180),
.A2(n_137),
.B(n_140),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_139),
.B(n_14),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_175),
.A2(n_121),
.B1(n_133),
.B2(n_90),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_182),
.A2(n_193),
.B1(n_199),
.B2(n_204),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_183),
.A2(n_200),
.B(n_185),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_185),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_186),
.B(n_187),
.C(n_163),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_154),
.B(n_137),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_191),
.B(n_195),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_150),
.B(n_15),
.Y(n_195)
);

BUFx4f_ASAP7_75t_SL g196 ( 
.A(n_167),
.Y(n_196)
);

INVx13_ASAP7_75t_L g219 ( 
.A(n_196),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_153),
.B(n_104),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_197),
.B(n_207),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_166),
.A2(n_74),
.B1(n_104),
.B2(n_88),
.Y(n_199)
);

OR2x2_ASAP7_75t_L g200 ( 
.A(n_144),
.B(n_82),
.Y(n_200)
);

A2O1A1Ixp33_ASAP7_75t_L g203 ( 
.A1(n_162),
.A2(n_178),
.B(n_179),
.C(n_180),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_203),
.B(n_211),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_157),
.A2(n_162),
.B1(n_180),
.B2(n_159),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_155),
.B(n_161),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_209),
.A2(n_216),
.B1(n_193),
.B2(n_182),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_178),
.B(n_155),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_157),
.A2(n_171),
.B1(n_158),
.B2(n_147),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_217),
.A2(n_177),
.B(n_168),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_192),
.B(n_160),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_218),
.B(n_223),
.C(n_225),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_202),
.B(n_189),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_220),
.B(n_227),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_222),
.A2(n_228),
.B(n_196),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_192),
.B(n_170),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_190),
.Y(n_226)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_226),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_189),
.B(n_164),
.Y(n_227)
);

AND2x6_ASAP7_75t_L g228 ( 
.A(n_203),
.B(n_169),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_209),
.A2(n_148),
.B1(n_152),
.B2(n_164),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_230),
.A2(n_237),
.B1(n_212),
.B2(n_201),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_183),
.B(n_211),
.Y(n_232)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_232),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_187),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_SL g257 ( 
.A1(n_233),
.A2(n_235),
.B1(n_238),
.B2(n_243),
.Y(n_257)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_190),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_183),
.B(n_217),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_SL g258 ( 
.A(n_236),
.B(n_239),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_200),
.A2(n_204),
.B1(n_216),
.B2(n_210),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_198),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_200),
.B(n_206),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_184),
.B(n_213),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_240),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_184),
.B(n_213),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_241),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_242),
.A2(n_214),
.B(n_196),
.Y(n_255)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_198),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_244),
.A2(n_210),
.B1(n_215),
.B2(n_208),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_245),
.A2(n_226),
.B1(n_243),
.B2(n_238),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_233),
.B(n_210),
.C(n_215),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_248),
.B(n_252),
.Y(n_280)
);

OAI32xp33_ASAP7_75t_L g250 ( 
.A1(n_224),
.A2(n_208),
.A3(n_188),
.B1(n_205),
.B2(n_199),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_250),
.B(n_256),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_251),
.A2(n_253),
.B1(n_259),
.B2(n_264),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_223),
.B(n_212),
.C(n_188),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_237),
.A2(n_201),
.B1(n_214),
.B2(n_205),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_255),
.A2(n_265),
.B(n_235),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_224),
.A2(n_236),
.B1(n_239),
.B2(n_242),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_218),
.B(n_196),
.C(n_194),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_SL g281 ( 
.A(n_260),
.B(n_266),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_232),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_262),
.B(n_261),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_230),
.A2(n_194),
.B1(n_229),
.B2(n_244),
.Y(n_264)
);

AND2x4_ASAP7_75t_L g265 ( 
.A(n_222),
.B(n_229),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_225),
.B(n_234),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_267),
.B(n_277),
.Y(n_286)
);

CKINVDCx16_ASAP7_75t_R g269 ( 
.A(n_257),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_269),
.B(n_272),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_270),
.A2(n_278),
.B1(n_255),
.B2(n_248),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_254),
.B(n_221),
.Y(n_271)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_271),
.Y(n_293)
);

CKINVDCx16_ASAP7_75t_R g272 ( 
.A(n_265),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_250),
.B(n_231),
.Y(n_273)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_273),
.Y(n_294)
);

AO22x1_ASAP7_75t_L g274 ( 
.A1(n_265),
.A2(n_228),
.B1(n_231),
.B2(n_219),
.Y(n_274)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_274),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_246),
.B(n_219),
.Y(n_275)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_275),
.Y(n_297)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_249),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_251),
.A2(n_240),
.B1(n_241),
.B2(n_253),
.Y(n_278)
);

CKINVDCx14_ASAP7_75t_R g296 ( 
.A(n_279),
.Y(n_296)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_245),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_282),
.Y(n_287)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_264),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_283),
.B(n_259),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_280),
.B(n_247),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_285),
.B(n_291),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_281),
.B(n_247),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_288),
.B(n_295),
.Y(n_298)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_289),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_290),
.B(n_276),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_280),
.B(n_281),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_278),
.B(n_252),
.Y(n_295)
);

HB1xp67_ASAP7_75t_L g299 ( 
.A(n_293),
.Y(n_299)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_299),
.Y(n_313)
);

OAI321xp33_ASAP7_75t_L g309 ( 
.A1(n_301),
.A2(n_294),
.A3(n_273),
.B1(n_268),
.B2(n_283),
.C(n_297),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_285),
.B(n_260),
.C(n_263),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_302),
.B(n_303),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_295),
.B(n_271),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_291),
.B(n_288),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_304),
.B(n_305),
.C(n_306),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_290),
.B(n_256),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_292),
.B(n_268),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_296),
.B(n_275),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_307),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_309),
.A2(n_265),
.B1(n_267),
.B2(n_277),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_306),
.B(n_279),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g320 ( 
.A1(n_311),
.A2(n_266),
.B(n_284),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_298),
.B(n_286),
.C(n_276),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_314),
.B(n_315),
.C(n_270),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_300),
.A2(n_287),
.B1(n_282),
.B2(n_284),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_316),
.B(n_308),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_317),
.B(n_319),
.Y(n_325)
);

OR2x2_ASAP7_75t_L g318 ( 
.A(n_312),
.B(n_286),
.Y(n_318)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_318),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_310),
.B(n_305),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_320),
.A2(n_321),
.B(n_322),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_SL g326 ( 
.A(n_325),
.B(n_324),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_326),
.B(n_327),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_323),
.B(n_318),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_L g329 ( 
.A1(n_328),
.A2(n_310),
.B(n_314),
.Y(n_329)
);

AOI221x1_ASAP7_75t_L g330 ( 
.A1(n_329),
.A2(n_319),
.B1(n_304),
.B2(n_298),
.C(n_274),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_330),
.A2(n_313),
.B1(n_274),
.B2(n_258),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_331),
.B(n_258),
.Y(n_332)
);


endmodule