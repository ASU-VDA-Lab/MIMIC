module fake_jpeg_29813_n_337 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_337);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_337;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_13),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx12_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

BUFx2_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_5),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_2),
.B(n_3),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_12),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx3_ASAP7_75t_SL g60 ( 
.A(n_36),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_37),
.Y(n_67)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_38),
.B(n_39),
.Y(n_52)
);

BUFx4f_ASAP7_75t_SL g39 ( 
.A(n_25),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_26),
.B(n_9),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_40),
.B(n_41),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_20),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_20),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_47),
.B(n_48),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_20),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_43),
.A2(n_34),
.B1(n_32),
.B2(n_18),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_49),
.A2(n_55),
.B1(n_59),
.B2(n_48),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_44),
.B(n_34),
.C(n_26),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_53),
.B(n_56),
.C(n_47),
.Y(n_88)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_54),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_43),
.A2(n_18),
.B1(n_29),
.B2(n_17),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_44),
.B(n_35),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_57),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_38),
.A2(n_18),
.B1(n_29),
.B2(n_35),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_41),
.A2(n_29),
.B1(n_35),
.B2(n_21),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_63),
.A2(n_24),
.B1(n_33),
.B2(n_37),
.Y(n_79)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_64),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g70 ( 
.A1(n_62),
.A2(n_39),
.B(n_40),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_70),
.A2(n_28),
.B(n_22),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_71),
.A2(n_49),
.B1(n_60),
.B2(n_65),
.Y(n_111)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_57),
.Y(n_72)
);

INVx1_ASAP7_75t_SL g100 ( 
.A(n_72),
.Y(n_100)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_73),
.Y(n_101)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_51),
.Y(n_74)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_74),
.Y(n_108)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_50),
.Y(n_75)
);

INVx1_ASAP7_75t_SL g113 ( 
.A(n_75),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_62),
.B(n_39),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_76),
.B(n_78),
.Y(n_103)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_65),
.Y(n_77)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_77),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_53),
.B(n_39),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_79),
.A2(n_37),
.B1(n_33),
.B2(n_24),
.Y(n_122)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_58),
.Y(n_80)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_80),
.Y(n_129)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_50),
.Y(n_81)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_81),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_52),
.B(n_39),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_83),
.B(n_86),
.Y(n_104)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_60),
.Y(n_84)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_84),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_52),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_85),
.B(n_89),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_56),
.B(n_30),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_64),
.Y(n_87)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_87),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_88),
.B(n_93),
.Y(n_119)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_61),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_61),
.Y(n_90)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_90),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_56),
.B(n_27),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_91),
.B(n_23),
.Y(n_105)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_61),
.Y(n_92)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_92),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_56),
.B(n_36),
.C(n_42),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_93),
.B(n_55),
.C(n_67),
.Y(n_102)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_60),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_94),
.B(n_95),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_59),
.B(n_16),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_67),
.B(n_16),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_96),
.B(n_28),
.Y(n_110)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_54),
.Y(n_97)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_97),
.Y(n_99)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_54),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_98),
.B(n_37),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_102),
.B(n_107),
.C(n_119),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_105),
.B(n_110),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_78),
.B(n_36),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_111),
.A2(n_117),
.B1(n_98),
.B2(n_97),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_83),
.Y(n_115)
);

CKINVDCx14_ASAP7_75t_R g140 ( 
.A(n_115),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_71),
.A2(n_66),
.B1(n_65),
.B2(n_58),
.Y(n_117)
);

NOR2x1_ASAP7_75t_R g118 ( 
.A(n_86),
.B(n_33),
.Y(n_118)
);

NOR2x1_ASAP7_75t_R g133 ( 
.A(n_118),
.B(n_70),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_73),
.B(n_74),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_121),
.B(n_127),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_122),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_123),
.A2(n_21),
.B(n_69),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_125),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_76),
.B(n_21),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_126),
.B(n_23),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_88),
.B(n_66),
.Y(n_127)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_109),
.Y(n_131)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_131),
.Y(n_160)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_99),
.Y(n_132)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_132),
.Y(n_164)
);

AO21x1_ASAP7_75t_L g176 ( 
.A1(n_133),
.A2(n_134),
.B(n_150),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_118),
.B(n_91),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_103),
.B(n_81),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_136),
.B(n_144),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_101),
.A2(n_108),
.B1(n_119),
.B2(n_115),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_137),
.A2(n_145),
.B1(n_153),
.B2(n_112),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_123),
.A2(n_84),
.B(n_22),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_138),
.A2(n_113),
.B(n_33),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_129),
.A2(n_80),
.B1(n_58),
.B2(n_66),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_141),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_142),
.A2(n_111),
.B1(n_113),
.B2(n_128),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_143),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_103),
.B(n_82),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_101),
.A2(n_68),
.B1(n_77),
.B2(n_82),
.Y(n_145)
);

BUFx24_ASAP7_75t_SL g146 ( 
.A(n_121),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_146),
.Y(n_156)
);

INVx6_ASAP7_75t_L g147 ( 
.A(n_106),
.Y(n_147)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_147),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_119),
.A2(n_92),
.B(n_90),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_148),
.A2(n_154),
.B(n_127),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_108),
.B(n_27),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_149),
.B(n_128),
.Y(n_169)
);

A2O1A1Ixp33_ASAP7_75t_SL g150 ( 
.A1(n_102),
.A2(n_68),
.B(n_37),
.C(n_67),
.Y(n_150)
);

INVx1_ASAP7_75t_SL g151 ( 
.A(n_124),
.Y(n_151)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_151),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_107),
.A2(n_69),
.B1(n_72),
.B2(n_46),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_157),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_155),
.B(n_104),
.C(n_114),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_159),
.B(n_165),
.C(n_167),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_145),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_161),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_133),
.A2(n_120),
.B(n_104),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_163),
.A2(n_179),
.B(n_8),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_155),
.B(n_109),
.C(n_124),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_135),
.B(n_105),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_169),
.B(n_10),
.Y(n_208)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_171),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_172),
.B(n_154),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_135),
.B(n_137),
.C(n_136),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_173),
.B(n_25),
.C(n_19),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_144),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_174),
.Y(n_204)
);

INVx13_ASAP7_75t_L g175 ( 
.A(n_132),
.Y(n_175)
);

INVx11_ASAP7_75t_L g194 ( 
.A(n_175),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_140),
.B(n_100),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_177),
.B(n_178),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_148),
.B(n_116),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_139),
.A2(n_100),
.B(n_116),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_142),
.A2(n_106),
.B1(n_129),
.B2(n_99),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_180),
.B(n_181),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_149),
.B(n_112),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_182),
.A2(n_150),
.B1(n_46),
.B2(n_42),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_139),
.A2(n_25),
.B(n_31),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_183),
.A2(n_138),
.B(n_151),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_134),
.B(n_153),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_SL g214 ( 
.A(n_184),
.B(n_19),
.Y(n_214)
);

INVx13_ASAP7_75t_L g185 ( 
.A(n_147),
.Y(n_185)
);

OAI21x1_ASAP7_75t_R g188 ( 
.A1(n_185),
.A2(n_150),
.B(n_152),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_186),
.A2(n_187),
.B(n_202),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_L g241 ( 
.A1(n_188),
.A2(n_19),
.B1(n_1),
.B2(n_4),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_167),
.B(n_152),
.Y(n_189)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_189),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_178),
.A2(n_134),
.B(n_150),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_192),
.A2(n_0),
.B(n_1),
.Y(n_238)
);

A2O1A1O1Ixp25_ASAP7_75t_L g195 ( 
.A1(n_162),
.A2(n_130),
.B(n_150),
.C(n_131),
.D(n_13),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_195),
.B(n_183),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_196),
.A2(n_213),
.B1(n_171),
.B2(n_180),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_166),
.B(n_10),
.Y(n_198)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_198),
.Y(n_235)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_160),
.Y(n_199)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_199),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_179),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_200),
.B(n_206),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_176),
.A2(n_25),
.B(n_1),
.Y(n_202)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_172),
.B(n_24),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_203),
.A2(n_216),
.B(n_7),
.Y(n_234)
);

BUFx5_ASAP7_75t_L g205 ( 
.A(n_185),
.Y(n_205)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_205),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_177),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_173),
.B(n_25),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_207),
.B(n_211),
.C(n_165),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_208),
.B(n_209),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_169),
.B(n_9),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_181),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_210),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_159),
.B(n_9),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_212),
.B(n_156),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_182),
.A2(n_161),
.B1(n_174),
.B2(n_184),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_214),
.B(n_176),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_217),
.B(n_192),
.C(n_203),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_218),
.B(n_199),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_220),
.A2(n_230),
.B1(n_231),
.B2(n_240),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_197),
.A2(n_158),
.B1(n_176),
.B2(n_157),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_221),
.A2(n_232),
.B1(n_233),
.B2(n_216),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_SL g249 ( 
.A(n_222),
.B(n_214),
.Y(n_249)
);

OAI21xp33_ASAP7_75t_L g223 ( 
.A1(n_204),
.A2(n_162),
.B(n_170),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_223),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_213),
.B(n_163),
.Y(n_224)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_224),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_226),
.B(n_234),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_190),
.B(n_170),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_229),
.B(n_237),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_197),
.A2(n_168),
.B1(n_160),
.B2(n_164),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_201),
.A2(n_168),
.B1(n_164),
.B2(n_185),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_201),
.A2(n_175),
.B1(n_156),
.B2(n_11),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_200),
.A2(n_175),
.B1(n_8),
.B2(n_12),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_190),
.B(n_19),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_238),
.B(n_241),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_204),
.A2(n_7),
.B1(n_15),
.B2(n_14),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_245),
.A2(n_234),
.B1(n_230),
.B2(n_195),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_225),
.B(n_206),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_246),
.B(n_252),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_229),
.B(n_207),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_247),
.B(n_249),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_222),
.B(n_211),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_250),
.B(n_253),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_240),
.B(n_210),
.Y(n_252)
);

XOR2x2_ASAP7_75t_L g253 ( 
.A(n_226),
.B(n_193),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_220),
.A2(n_193),
.B1(n_188),
.B2(n_203),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_255),
.A2(n_188),
.B1(n_231),
.B2(n_221),
.Y(n_267)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_256),
.Y(n_273)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_219),
.Y(n_257)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_257),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_258),
.B(n_261),
.C(n_263),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_235),
.B(n_205),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_259),
.B(n_264),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_217),
.B(n_191),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_236),
.B(n_191),
.Y(n_262)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_262),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_227),
.B(n_187),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_239),
.Y(n_264)
);

INVx13_ASAP7_75t_L g266 ( 
.A(n_262),
.Y(n_266)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_266),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_267),
.A2(n_269),
.B1(n_270),
.B2(n_275),
.Y(n_296)
);

BUFx2_ASAP7_75t_L g268 ( 
.A(n_254),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_268),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_260),
.A2(n_253),
.B1(n_255),
.B2(n_263),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_SL g271 ( 
.A1(n_248),
.A2(n_242),
.B1(n_233),
.B2(n_232),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_271),
.A2(n_243),
.B1(n_194),
.B2(n_261),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_260),
.B(n_215),
.Y(n_275)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_275),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_258),
.A2(n_228),
.B(n_215),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_278),
.A2(n_280),
.B(n_281),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_L g280 ( 
.A1(n_251),
.A2(n_228),
.B(n_223),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_243),
.A2(n_202),
.B(n_196),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_283),
.B(n_287),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_274),
.B(n_247),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_284),
.B(n_289),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_272),
.A2(n_194),
.B1(n_250),
.B2(n_249),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_274),
.B(n_244),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_279),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_290),
.B(n_292),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_265),
.B(n_244),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_291),
.B(n_296),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_277),
.B(n_237),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_278),
.A2(n_8),
.B(n_15),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_294),
.A2(n_276),
.B(n_269),
.Y(n_304)
);

FAx1_ASAP7_75t_L g295 ( 
.A(n_280),
.B(n_13),
.CI(n_4),
.CON(n_295),
.SN(n_295)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_295),
.B(n_270),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_282),
.B(n_19),
.C(n_4),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_297),
.B(n_273),
.Y(n_301)
);

CKINVDCx14_ASAP7_75t_R g312 ( 
.A(n_300),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_301),
.B(n_305),
.Y(n_313)
);

INVx6_ASAP7_75t_L g302 ( 
.A(n_293),
.Y(n_302)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_302),
.Y(n_311)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_304),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_286),
.B(n_268),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_288),
.A2(n_267),
.B1(n_285),
.B2(n_296),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_306),
.B(n_295),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_291),
.B(n_282),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_308),
.B(n_309),
.Y(n_318)
);

AOI21x1_ASAP7_75t_L g309 ( 
.A1(n_286),
.A2(n_266),
.B(n_281),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_303),
.A2(n_284),
.B(n_289),
.Y(n_310)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_310),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_302),
.B(n_297),
.Y(n_314)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_314),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_316),
.B(n_317),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_L g317 ( 
.A1(n_299),
.A2(n_295),
.B(n_265),
.Y(n_317)
);

AND2x2_ASAP7_75t_L g321 ( 
.A(n_318),
.B(n_306),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_321),
.B(n_324),
.Y(n_330)
);

AOI21xp33_ASAP7_75t_L g323 ( 
.A1(n_313),
.A2(n_307),
.B(n_298),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_SL g331 ( 
.A1(n_323),
.A2(n_0),
.B(n_5),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_314),
.B(n_298),
.Y(n_324)
);

AND2x2_ASAP7_75t_L g325 ( 
.A(n_315),
.B(n_308),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_325),
.B(n_326),
.Y(n_329)
);

AND2x2_ASAP7_75t_L g326 ( 
.A(n_312),
.B(n_0),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_322),
.B(n_311),
.C(n_4),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_327),
.B(n_328),
.Y(n_333)
);

AO221x1_ASAP7_75t_L g328 ( 
.A1(n_320),
.A2(n_0),
.B1(n_5),
.B2(n_6),
.C(n_319),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_331),
.B(n_329),
.C(n_320),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_SL g334 ( 
.A(n_332),
.B(n_330),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_SL g335 ( 
.A1(n_334),
.A2(n_333),
.B(n_5),
.Y(n_335)
);

BUFx24_ASAP7_75t_SL g336 ( 
.A(n_335),
.Y(n_336)
);

AOI21xp5_ASAP7_75t_L g337 ( 
.A1(n_336),
.A2(n_6),
.B(n_334),
.Y(n_337)
);


endmodule