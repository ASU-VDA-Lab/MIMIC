module real_jpeg_29475_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_255;
wire n_40;
wire n_105;
wire n_197;
wire n_173;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_150;
wire n_41;
wire n_74;
wire n_70;
wire n_32;
wire n_20;
wire n_80;
wire n_228;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_185;
wire n_125;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_167;
wire n_128;
wire n_202;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_206;
wire n_127;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_89;

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_0),
.A2(n_42),
.B1(n_43),
.B2(n_49),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_0),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_0),
.A2(n_49),
.B1(n_56),
.B2(n_58),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_0),
.A2(n_27),
.B1(n_28),
.B2(n_49),
.Y(n_126)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_1),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_2),
.A2(n_27),
.B1(n_28),
.B2(n_38),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_2),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_2),
.A2(n_38),
.B1(n_73),
.B2(n_74),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_2),
.A2(n_38),
.B1(n_56),
.B2(n_58),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_2),
.A2(n_38),
.B1(n_42),
.B2(n_43),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_L g34 ( 
.A1(n_3),
.A2(n_27),
.B1(n_28),
.B2(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_3),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_3),
.A2(n_35),
.B1(n_56),
.B2(n_58),
.Y(n_64)
);

OAI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_3),
.A2(n_35),
.B1(n_42),
.B2(n_43),
.Y(n_90)
);

BUFx12_ASAP7_75t_L g72 ( 
.A(n_4),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_5),
.A2(n_42),
.B1(n_43),
.B2(n_51),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_5),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_5),
.A2(n_27),
.B1(n_28),
.B2(n_51),
.Y(n_96)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

INVx13_ASAP7_75t_L g74 ( 
.A(n_7),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_8),
.A2(n_73),
.B1(n_74),
.B2(n_110),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_8),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_8),
.A2(n_56),
.B1(n_58),
.B2(n_110),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_8),
.A2(n_42),
.B1(n_43),
.B2(n_110),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_8),
.A2(n_27),
.B1(n_28),
.B2(n_110),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_9),
.A2(n_73),
.B1(n_74),
.B2(n_78),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_9),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_9),
.A2(n_56),
.B1(n_58),
.B2(n_78),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_9),
.A2(n_42),
.B1(n_43),
.B2(n_78),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_9),
.A2(n_27),
.B1(n_28),
.B2(n_78),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_10),
.A2(n_73),
.B1(n_74),
.B2(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_10),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_10),
.A2(n_56),
.B1(n_58),
.B2(n_135),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_10),
.A2(n_42),
.B1(n_43),
.B2(n_135),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_10),
.A2(n_27),
.B1(n_28),
.B2(n_135),
.Y(n_227)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_11),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_12),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_12),
.B(n_76),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_12),
.B(n_58),
.Y(n_178)
);

AOI21xp33_ASAP7_75t_L g182 ( 
.A1(n_12),
.A2(n_58),
.B(n_178),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_12),
.A2(n_42),
.B1(n_43),
.B2(n_124),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_12),
.A2(n_28),
.B(n_45),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_12),
.B(n_59),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_12),
.A2(n_85),
.B1(n_86),
.B2(n_227),
.Y(n_229)
);

BUFx24_ASAP7_75t_L g57 ( 
.A(n_13),
.Y(n_57)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_14),
.Y(n_62)
);

INVx11_ASAP7_75t_SL g30 ( 
.A(n_15),
.Y(n_30)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_138),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_136),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_112),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_19),
.B(n_112),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_93),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_81),
.B2(n_82),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_52),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_39),
.Y(n_23)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_24),
.B(n_39),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_36),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_25),
.A2(n_126),
.B(n_167),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_33),
.Y(n_25)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_26),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_26),
.A2(n_37),
.B(n_98),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_26),
.A2(n_31),
.B1(n_218),
.B2(n_220),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_31),
.Y(n_26)
);

OA22x2_ASAP7_75t_L g47 ( 
.A1(n_27),
.A2(n_28),
.B1(n_45),
.B2(n_46),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_27),
.B(n_231),
.Y(n_230)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx4f_ASAP7_75t_SL g28 ( 
.A(n_29),
.Y(n_28)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_31),
.B(n_37),
.Y(n_36)
);

INVx11_ASAP7_75t_L g167 ( 
.A(n_31),
.Y(n_167)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_32),
.A2(n_85),
.B1(n_96),
.B2(n_126),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_34),
.B(n_86),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_36),
.A2(n_85),
.B(n_214),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_37),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_40),
.A2(n_47),
.B1(n_48),
.B2(n_50),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_SL g88 ( 
.A1(n_40),
.A2(n_50),
.B(n_89),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_40),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_40),
.A2(n_89),
.B(n_146),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_40),
.A2(n_47),
.B1(n_185),
.B2(n_186),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_40),
.A2(n_186),
.B(n_196),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_40),
.A2(n_47),
.B1(n_203),
.B2(n_204),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_40),
.A2(n_47),
.B1(n_185),
.B2(n_204),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_47),
.Y(n_40)
);

OAI22xp33_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_43),
.B1(n_45),
.B2(n_46),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_42),
.A2(n_43),
.B1(n_61),
.B2(n_62),
.Y(n_60)
);

AOI32xp33_ASAP7_75t_L g176 ( 
.A1(n_42),
.A2(n_56),
.A3(n_177),
.B1(n_178),
.B2(n_179),
.Y(n_176)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

NAND2xp33_ASAP7_75t_SL g179 ( 
.A(n_43),
.B(n_61),
.Y(n_179)
);

A2O1A1Ixp33_ASAP7_75t_L g205 ( 
.A1(n_43),
.A2(n_46),
.B(n_124),
.C(n_206),
.Y(n_205)
);

BUFx10_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_47),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_47),
.A2(n_48),
.B(n_100),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_47),
.B(n_124),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_53),
.A2(n_54),
.B1(n_67),
.B2(n_68),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_54),
.Y(n_53)
);

AOI21xp5_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_59),
.B(n_63),
.Y(n_54)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_56),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_56),
.A2(n_58),
.B1(n_61),
.B2(n_62),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_56),
.A2(n_58),
.B1(n_71),
.B2(n_72),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_56),
.A2(n_75),
.B1(n_122),
.B2(n_123),
.Y(n_121)
);

BUFx4f_ASAP7_75t_SL g56 ( 
.A(n_57),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_58),
.B(n_71),
.Y(n_122)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_60),
.B(n_66),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_60),
.B(n_64),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_60),
.B(n_105),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_60),
.A2(n_65),
.B1(n_129),
.B2(n_150),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_60),
.A2(n_65),
.B1(n_150),
.B2(n_163),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_60),
.A2(n_65),
.B1(n_163),
.B2(n_182),
.Y(n_181)
);

INVx6_ASAP7_75t_L g177 ( 
.A(n_61),
.Y(n_177)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_65),
.Y(n_63)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_65),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_68),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_SL g68 ( 
.A1(n_69),
.A2(n_77),
.B(n_79),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_69),
.A2(n_77),
.B1(n_109),
.B2(n_111),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_69),
.A2(n_109),
.B1(n_111),
.B2(n_133),
.Y(n_132)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_70),
.A2(n_76),
.B1(n_123),
.B2(n_134),
.Y(n_151)
);

O2A1O1Ixp33_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_73),
.B(n_75),
.C(n_76),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_71),
.B(n_73),
.Y(n_75)
);

CKINVDCx14_ASAP7_75t_R g71 ( 
.A(n_72),
.Y(n_71)
);

HAxp5_ASAP7_75t_SL g123 ( 
.A(n_73),
.B(n_124),
.CON(n_123),
.SN(n_123)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_76),
.B(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_76),
.Y(n_111)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_84),
.B1(n_88),
.B2(n_92),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_84),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_86),
.B(n_87),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_L g95 ( 
.A1(n_85),
.A2(n_96),
.B(n_97),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_85),
.A2(n_167),
.B1(n_219),
.B2(n_227),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_86),
.B(n_124),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_88),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_90),
.B(n_91),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_90),
.B(n_101),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_91),
.B(n_147),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_102),
.C(n_107),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_94),
.B(n_114),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_99),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_95),
.B(n_99),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_98),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_102),
.A2(n_107),
.B1(n_108),
.B2(n_115),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_102),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_103),
.A2(n_104),
.B(n_106),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_103),
.A2(n_128),
.B(n_130),
.Y(n_127)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_108),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_116),
.C(n_118),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_113),
.A2(n_116),
.B1(n_117),
.B2(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_113),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_117),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_118),
.A2(n_119),
.B1(n_253),
.B2(n_254),
.Y(n_252)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_127),
.C(n_131),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_SL g152 ( 
.A(n_120),
.B(n_153),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_125),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_121),
.B(n_125),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_127),
.A2(n_131),
.B1(n_132),
.B2(n_154),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_127),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_132),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_134),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

O2A1O1Ixp33_ASAP7_75t_SL g138 ( 
.A1(n_139),
.A2(n_168),
.B(n_250),
.C(n_256),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_155),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_140),
.B(n_155),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_152),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_143),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_142),
.B(n_143),
.C(n_152),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_148),
.C(n_151),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_144),
.A2(n_145),
.B1(n_148),
.B2(n_149),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_149),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_SL g157 ( 
.A(n_151),
.B(n_158),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_159),
.C(n_161),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_156),
.A2(n_157),
.B1(n_245),
.B2(n_247),
.Y(n_244)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_159),
.A2(n_160),
.B1(n_161),
.B2(n_246),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_160),
.Y(n_159)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_161),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_164),
.C(n_166),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_162),
.B(n_190),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_164),
.A2(n_165),
.B1(n_166),
.B2(n_191),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_165),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_166),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_169),
.B(n_249),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_170),
.A2(n_242),
.B(n_248),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_171),
.A2(n_197),
.B(n_241),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_187),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_172),
.B(n_187),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_180),
.C(n_183),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_173),
.A2(n_174),
.B1(n_238),
.B2(n_239),
.Y(n_237)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_176),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_175),
.B(n_176),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_180),
.A2(n_181),
.B1(n_183),
.B2(n_184),
.Y(n_239)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_181),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_184),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_188),
.A2(n_189),
.B1(n_192),
.B2(n_193),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_188),
.B(n_194),
.C(n_195),
.Y(n_243)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_195),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_198),
.A2(n_235),
.B(n_240),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_199),
.A2(n_215),
.B(n_234),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_207),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_200),
.B(n_207),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_201),
.B(n_205),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_201),
.A2(n_202),
.B1(n_205),
.B2(n_222),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g201 ( 
.A(n_202),
.Y(n_201)
);

CKINVDCx16_ASAP7_75t_R g222 ( 
.A(n_205),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_213),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_209),
.A2(n_210),
.B1(n_211),
.B2(n_212),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_209),
.B(n_212),
.C(n_213),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_210),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g211 ( 
.A(n_212),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_214),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_216),
.A2(n_223),
.B(n_233),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_221),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_217),
.B(n_221),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_224),
.A2(n_228),
.B(n_232),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_226),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_225),
.B(n_226),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_229),
.B(n_230),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_237),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_236),
.B(n_237),
.Y(n_240)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_244),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_243),
.B(n_244),
.Y(n_248)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_245),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_252),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_251),
.B(n_252),
.Y(n_256)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);


endmodule