module fake_jpeg_20755_n_45 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_45);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_45;

wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_40;
wire n_19;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_32;

INVx11_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx5_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_7),
.B(n_3),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_20),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_25),
.B(n_26),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_24),
.B(n_0),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_23),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_27),
.B(n_28),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_21),
.B(n_0),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g29 ( 
.A(n_22),
.B(n_1),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_29),
.B(n_30),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_20),
.B(n_1),
.Y(n_30)
);

XNOR2xp5_ASAP7_75t_L g34 ( 
.A(n_28),
.B(n_22),
.Y(n_34)
);

XOR2xp5_ASAP7_75t_L g38 ( 
.A(n_34),
.B(n_19),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_25),
.A2(n_13),
.B1(n_18),
.B2(n_5),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_35),
.B(n_31),
.Y(n_37)
);

OR2x2_ASAP7_75t_L g36 ( 
.A(n_34),
.B(n_2),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_36),
.B(n_37),
.Y(n_40)
);

AO221x1_ASAP7_75t_L g41 ( 
.A1(n_38),
.A2(n_39),
.B1(n_33),
.B2(n_4),
.C(n_2),
.Y(n_41)
);

XOR2x2_ASAP7_75t_L g39 ( 
.A(n_32),
.B(n_19),
.Y(n_39)
);

OAI211xp5_ASAP7_75t_SL g42 ( 
.A1(n_41),
.A2(n_37),
.B(n_4),
.C(n_11),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_42),
.B(n_10),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_L g44 ( 
.A1(n_43),
.A2(n_41),
.B1(n_40),
.B2(n_16),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_44),
.A2(n_12),
.B1(n_14),
.B2(n_17),
.Y(n_45)
);


endmodule