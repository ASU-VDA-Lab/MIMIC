module fake_aes_8767_n_586 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_73, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_71, n_42, n_24, n_75, n_19, n_61, n_21, n_6, n_4, n_74, n_72, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_586);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_73;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_71;
input n_42;
input n_24;
input n_75;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_74;
input n_72;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_586;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_383;
wire n_288;
wire n_532;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_540;
wire n_563;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_554;
wire n_447;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_370;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_539;
wire n_197;
wire n_201;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_583;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_487;
wire n_451;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx20_ASAP7_75t_R g76 ( .A(n_28), .Y(n_76) );
INVx1_ASAP7_75t_L g77 ( .A(n_50), .Y(n_77) );
INVxp67_ASAP7_75t_SL g78 ( .A(n_0), .Y(n_78) );
CKINVDCx5p33_ASAP7_75t_R g79 ( .A(n_27), .Y(n_79) );
CKINVDCx5p33_ASAP7_75t_R g80 ( .A(n_36), .Y(n_80) );
INVxp67_ASAP7_75t_L g81 ( .A(n_5), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_38), .Y(n_82) );
INVx2_ASAP7_75t_L g83 ( .A(n_61), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_53), .Y(n_84) );
INVx1_ASAP7_75t_SL g85 ( .A(n_2), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_14), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_20), .Y(n_87) );
INVxp67_ASAP7_75t_L g88 ( .A(n_71), .Y(n_88) );
CKINVDCx20_ASAP7_75t_R g89 ( .A(n_51), .Y(n_89) );
INVxp67_ASAP7_75t_L g90 ( .A(n_32), .Y(n_90) );
NOR2xp67_ASAP7_75t_L g91 ( .A(n_33), .B(n_9), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_11), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_45), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_52), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_44), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_49), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_11), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_67), .Y(n_98) );
INVxp33_ASAP7_75t_L g99 ( .A(n_63), .Y(n_99) );
INVxp33_ASAP7_75t_SL g100 ( .A(n_21), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_35), .Y(n_101) );
INVxp33_ASAP7_75t_SL g102 ( .A(n_23), .Y(n_102) );
INVx2_ASAP7_75t_SL g103 ( .A(n_74), .Y(n_103) );
CKINVDCx20_ASAP7_75t_R g104 ( .A(n_70), .Y(n_104) );
CKINVDCx5p33_ASAP7_75t_R g105 ( .A(n_43), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_48), .Y(n_106) );
INVx2_ASAP7_75t_L g107 ( .A(n_10), .Y(n_107) );
INVx2_ASAP7_75t_L g108 ( .A(n_25), .Y(n_108) );
CKINVDCx5p33_ASAP7_75t_R g109 ( .A(n_47), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_34), .Y(n_110) );
CKINVDCx16_ASAP7_75t_R g111 ( .A(n_22), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_7), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_58), .Y(n_113) );
INVxp67_ASAP7_75t_SL g114 ( .A(n_20), .Y(n_114) );
INVxp67_ASAP7_75t_L g115 ( .A(n_29), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_31), .Y(n_116) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_26), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_6), .Y(n_118) );
CKINVDCx14_ASAP7_75t_R g119 ( .A(n_60), .Y(n_119) );
CKINVDCx5p33_ASAP7_75t_R g120 ( .A(n_40), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_1), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_65), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_57), .Y(n_123) );
INVxp67_ASAP7_75t_L g124 ( .A(n_64), .Y(n_124) );
INVx2_ASAP7_75t_L g125 ( .A(n_83), .Y(n_125) );
NAND2xp5_ASAP7_75t_SL g126 ( .A(n_103), .B(n_0), .Y(n_126) );
NAND2xp33_ASAP7_75t_R g127 ( .A(n_100), .B(n_1), .Y(n_127) );
INVx2_ASAP7_75t_L g128 ( .A(n_83), .Y(n_128) );
INVx2_ASAP7_75t_L g129 ( .A(n_108), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_77), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_77), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_82), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_82), .Y(n_133) );
INVx2_ASAP7_75t_L g134 ( .A(n_108), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_84), .Y(n_135) );
INVx3_ASAP7_75t_L g136 ( .A(n_107), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_84), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_93), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g139 ( .A(n_103), .B(n_2), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_86), .B(n_3), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_93), .Y(n_141) );
CKINVDCx20_ASAP7_75t_R g142 ( .A(n_111), .Y(n_142) );
NOR2xp33_ASAP7_75t_L g143 ( .A(n_99), .B(n_3), .Y(n_143) );
NOR2xp33_ASAP7_75t_R g144 ( .A(n_119), .B(n_30), .Y(n_144) );
CKINVDCx5p33_ASAP7_75t_R g145 ( .A(n_76), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_94), .Y(n_146) );
CKINVDCx5p33_ASAP7_75t_R g147 ( .A(n_89), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g148 ( .A(n_86), .B(n_4), .Y(n_148) );
INVx2_ASAP7_75t_L g149 ( .A(n_94), .Y(n_149) );
CKINVDCx20_ASAP7_75t_R g150 ( .A(n_104), .Y(n_150) );
NOR2xp33_ASAP7_75t_R g151 ( .A(n_79), .B(n_75), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_87), .B(n_4), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_95), .Y(n_153) );
NAND2xp33_ASAP7_75t_SL g154 ( .A(n_117), .B(n_5), .Y(n_154) );
HB1xp67_ASAP7_75t_L g155 ( .A(n_87), .Y(n_155) );
NOR2xp33_ASAP7_75t_R g156 ( .A(n_80), .B(n_37), .Y(n_156) );
OA21x2_ASAP7_75t_L g157 ( .A1(n_95), .A2(n_73), .B(n_72), .Y(n_157) );
INVx2_ASAP7_75t_L g158 ( .A(n_98), .Y(n_158) );
INVx3_ASAP7_75t_L g159 ( .A(n_107), .Y(n_159) );
CKINVDCx5p33_ASAP7_75t_R g160 ( .A(n_102), .Y(n_160) );
HB1xp67_ASAP7_75t_L g161 ( .A(n_92), .Y(n_161) );
HB1xp67_ASAP7_75t_L g162 ( .A(n_92), .Y(n_162) );
AND2x4_ASAP7_75t_L g163 ( .A(n_112), .B(n_6), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_112), .B(n_7), .Y(n_164) );
BUFx6f_ASAP7_75t_L g165 ( .A(n_98), .Y(n_165) );
INVx2_ASAP7_75t_SL g166 ( .A(n_101), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_101), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_165), .Y(n_168) );
BUFx6f_ASAP7_75t_L g169 ( .A(n_165), .Y(n_169) );
INVx8_ASAP7_75t_L g170 ( .A(n_163), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_130), .B(n_109), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_165), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_165), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_165), .Y(n_174) );
AND2x4_ASAP7_75t_L g175 ( .A(n_155), .B(n_118), .Y(n_175) );
NAND2xp5_ASAP7_75t_SL g176 ( .A(n_166), .B(n_124), .Y(n_176) );
AND2x4_ASAP7_75t_L g177 ( .A(n_155), .B(n_121), .Y(n_177) );
NOR2x1p5_ASAP7_75t_L g178 ( .A(n_145), .B(n_78), .Y(n_178) );
INVx2_ASAP7_75t_L g179 ( .A(n_165), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_163), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_130), .B(n_120), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_165), .Y(n_182) );
INVxp67_ASAP7_75t_L g183 ( .A(n_161), .Y(n_183) );
NOR2xp33_ASAP7_75t_L g184 ( .A(n_160), .B(n_88), .Y(n_184) );
AND2x2_ASAP7_75t_L g185 ( .A(n_161), .B(n_121), .Y(n_185) );
AND2x4_ASAP7_75t_L g186 ( .A(n_162), .B(n_118), .Y(n_186) );
INVx2_ASAP7_75t_L g187 ( .A(n_125), .Y(n_187) );
OR2x2_ASAP7_75t_L g188 ( .A(n_162), .B(n_81), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_149), .Y(n_189) );
NAND2xp5_ASAP7_75t_SL g190 ( .A(n_166), .B(n_90), .Y(n_190) );
BUFx2_ASAP7_75t_L g191 ( .A(n_144), .Y(n_191) );
AND2x2_ASAP7_75t_L g192 ( .A(n_131), .B(n_97), .Y(n_192) );
INVx2_ASAP7_75t_L g193 ( .A(n_125), .Y(n_193) );
INVx2_ASAP7_75t_L g194 ( .A(n_125), .Y(n_194) );
HB1xp67_ASAP7_75t_L g195 ( .A(n_147), .Y(n_195) );
INVx5_ASAP7_75t_L g196 ( .A(n_163), .Y(n_196) );
AND2x2_ASAP7_75t_L g197 ( .A(n_131), .B(n_132), .Y(n_197) );
CKINVDCx5p33_ASAP7_75t_R g198 ( .A(n_150), .Y(n_198) );
AO22x2_ASAP7_75t_L g199 ( .A1(n_163), .A2(n_123), .B1(n_122), .B2(n_116), .Y(n_199) );
AND2x2_ASAP7_75t_L g200 ( .A(n_132), .B(n_114), .Y(n_200) );
AOI22xp5_ASAP7_75t_L g201 ( .A1(n_163), .A2(n_85), .B1(n_122), .B2(n_116), .Y(n_201) );
OR2x2_ASAP7_75t_L g202 ( .A(n_133), .B(n_123), .Y(n_202) );
CKINVDCx5p33_ASAP7_75t_R g203 ( .A(n_142), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_133), .B(n_105), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_139), .Y(n_205) );
CKINVDCx20_ASAP7_75t_R g206 ( .A(n_154), .Y(n_206) );
NOR3xp33_ASAP7_75t_L g207 ( .A(n_143), .B(n_115), .C(n_113), .Y(n_207) );
NAND2xp5_ASAP7_75t_SL g208 ( .A(n_166), .B(n_96), .Y(n_208) );
BUFx6f_ASAP7_75t_L g209 ( .A(n_157), .Y(n_209) );
INVx3_ASAP7_75t_L g210 ( .A(n_128), .Y(n_210) );
INVx4_ASAP7_75t_L g211 ( .A(n_157), .Y(n_211) );
NOR3xp33_ASAP7_75t_L g212 ( .A(n_143), .B(n_110), .C(n_106), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_135), .B(n_113), .Y(n_213) );
BUFx4f_ASAP7_75t_L g214 ( .A(n_135), .Y(n_214) );
BUFx2_ASAP7_75t_L g215 ( .A(n_144), .Y(n_215) );
NAND2xp5_ASAP7_75t_SL g216 ( .A(n_137), .B(n_110), .Y(n_216) );
AND2x6_ASAP7_75t_L g217 ( .A(n_137), .B(n_106), .Y(n_217) );
NAND2xp5_ASAP7_75t_SL g218 ( .A(n_138), .B(n_91), .Y(n_218) );
AND2x4_ASAP7_75t_L g219 ( .A(n_138), .B(n_8), .Y(n_219) );
AOI22xp33_ASAP7_75t_L g220 ( .A1(n_141), .A2(n_8), .B1(n_9), .B2(n_10), .Y(n_220) );
BUFx6f_ASAP7_75t_L g221 ( .A(n_157), .Y(n_221) );
INVx1_ASAP7_75t_L g222 ( .A(n_139), .Y(n_222) );
INVxp67_ASAP7_75t_L g223 ( .A(n_127), .Y(n_223) );
AND2x4_ASAP7_75t_L g224 ( .A(n_141), .B(n_12), .Y(n_224) );
INVx2_ASAP7_75t_L g225 ( .A(n_128), .Y(n_225) );
INVx2_ASAP7_75t_L g226 ( .A(n_128), .Y(n_226) );
INVxp67_ASAP7_75t_SL g227 ( .A(n_146), .Y(n_227) );
AND2x2_ASAP7_75t_L g228 ( .A(n_146), .B(n_12), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_149), .Y(n_229) );
AND2x4_ASAP7_75t_L g230 ( .A(n_167), .B(n_13), .Y(n_230) );
AND2x4_ASAP7_75t_L g231 ( .A(n_167), .B(n_13), .Y(n_231) );
AND2x4_ASAP7_75t_L g232 ( .A(n_205), .B(n_164), .Y(n_232) );
AOI22xp5_ASAP7_75t_L g233 ( .A1(n_199), .A2(n_127), .B1(n_153), .B2(n_140), .Y(n_233) );
HB1xp67_ASAP7_75t_L g234 ( .A(n_183), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_222), .B(n_227), .Y(n_235) );
AOI22xp33_ASAP7_75t_L g236 ( .A1(n_199), .A2(n_153), .B1(n_164), .B2(n_148), .Y(n_236) );
CKINVDCx20_ASAP7_75t_R g237 ( .A(n_198), .Y(n_237) );
INVx2_ASAP7_75t_L g238 ( .A(n_189), .Y(n_238) );
INVx2_ASAP7_75t_SL g239 ( .A(n_170), .Y(n_239) );
NAND2xp5_ASAP7_75t_SL g240 ( .A(n_214), .B(n_151), .Y(n_240) );
NAND2xp5_ASAP7_75t_SL g241 ( .A(n_214), .B(n_151), .Y(n_241) );
NOR2xp33_ASAP7_75t_L g242 ( .A(n_184), .B(n_126), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_189), .Y(n_243) );
NOR2xp33_ASAP7_75t_L g244 ( .A(n_188), .B(n_148), .Y(n_244) );
OR2x6_ASAP7_75t_L g245 ( .A(n_170), .B(n_140), .Y(n_245) );
INVx2_ASAP7_75t_L g246 ( .A(n_229), .Y(n_246) );
NAND2x1p5_ASAP7_75t_L g247 ( .A(n_219), .B(n_157), .Y(n_247) );
AND2x4_ASAP7_75t_SL g248 ( .A(n_175), .B(n_149), .Y(n_248) );
AOI22xp33_ASAP7_75t_SL g249 ( .A1(n_175), .A2(n_152), .B1(n_159), .B2(n_136), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_180), .Y(n_250) );
BUFx6f_ASAP7_75t_L g251 ( .A(n_170), .Y(n_251) );
AOI221x1_ASAP7_75t_L g252 ( .A1(n_211), .A2(n_158), .B1(n_152), .B2(n_129), .C(n_134), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_197), .Y(n_253) );
BUFx6f_ASAP7_75t_L g254 ( .A(n_170), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_197), .Y(n_255) );
INVx2_ASAP7_75t_L g256 ( .A(n_179), .Y(n_256) );
OR2x2_ASAP7_75t_L g257 ( .A(n_188), .B(n_159), .Y(n_257) );
INVx3_ASAP7_75t_SL g258 ( .A(n_219), .Y(n_258) );
AOI22xp5_ASAP7_75t_L g259 ( .A1(n_199), .A2(n_158), .B1(n_134), .B2(n_129), .Y(n_259) );
O2A1O1Ixp5_ASAP7_75t_L g260 ( .A1(n_211), .A2(n_158), .B(n_134), .C(n_129), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_175), .B(n_159), .Y(n_261) );
INVx1_ASAP7_75t_SL g262 ( .A(n_177), .Y(n_262) );
BUFx2_ASAP7_75t_L g263 ( .A(n_199), .Y(n_263) );
AOI22xp33_ASAP7_75t_L g264 ( .A1(n_219), .A2(n_159), .B1(n_136), .B2(n_157), .Y(n_264) );
INVx2_ASAP7_75t_SL g265 ( .A(n_177), .Y(n_265) );
INVx4_ASAP7_75t_L g266 ( .A(n_196), .Y(n_266) );
INVx2_ASAP7_75t_L g267 ( .A(n_179), .Y(n_267) );
INVx1_ASAP7_75t_SL g268 ( .A(n_177), .Y(n_268) );
BUFx6f_ASAP7_75t_L g269 ( .A(n_209), .Y(n_269) );
INVx2_ASAP7_75t_L g270 ( .A(n_187), .Y(n_270) );
INVx4_ASAP7_75t_L g271 ( .A(n_196), .Y(n_271) );
BUFx3_ASAP7_75t_L g272 ( .A(n_217), .Y(n_272) );
AND2x4_ASAP7_75t_L g273 ( .A(n_186), .B(n_136), .Y(n_273) );
INVxp67_ASAP7_75t_SL g274 ( .A(n_224), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_187), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_186), .B(n_136), .Y(n_276) );
INVx2_ASAP7_75t_L g277 ( .A(n_193), .Y(n_277) );
INVx2_ASAP7_75t_L g278 ( .A(n_193), .Y(n_278) );
CKINVDCx5p33_ASAP7_75t_R g279 ( .A(n_203), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_186), .B(n_156), .Y(n_280) );
AND2x4_ASAP7_75t_L g281 ( .A(n_200), .B(n_14), .Y(n_281) );
INVx3_ASAP7_75t_L g282 ( .A(n_224), .Y(n_282) );
NAND2xp5_ASAP7_75t_SL g283 ( .A(n_214), .B(n_39), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_171), .B(n_15), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_194), .Y(n_285) );
INVx2_ASAP7_75t_L g286 ( .A(n_194), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_225), .Y(n_287) );
BUFx3_ASAP7_75t_L g288 ( .A(n_217), .Y(n_288) );
AO21x2_ASAP7_75t_L g289 ( .A1(n_212), .A2(n_15), .B(n_16), .Y(n_289) );
AND2x4_ASAP7_75t_L g290 ( .A(n_200), .B(n_16), .Y(n_290) );
AO21x2_ASAP7_75t_L g291 ( .A1(n_207), .A2(n_17), .B(n_18), .Y(n_291) );
AOI22xp33_ASAP7_75t_L g292 ( .A1(n_224), .A2(n_17), .B1(n_18), .B2(n_19), .Y(n_292) );
INVx3_ASAP7_75t_L g293 ( .A(n_230), .Y(n_293) );
OAI22xp5_ASAP7_75t_L g294 ( .A1(n_223), .A2(n_201), .B1(n_230), .B2(n_231), .Y(n_294) );
NOR2xp33_ASAP7_75t_L g295 ( .A(n_185), .B(n_46), .Y(n_295) );
BUFx3_ASAP7_75t_L g296 ( .A(n_217), .Y(n_296) );
BUFx6f_ASAP7_75t_L g297 ( .A(n_209), .Y(n_297) );
BUFx6f_ASAP7_75t_L g298 ( .A(n_209), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_181), .B(n_19), .Y(n_299) );
INVx2_ASAP7_75t_L g300 ( .A(n_238), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_243), .Y(n_301) );
INVxp67_ASAP7_75t_L g302 ( .A(n_234), .Y(n_302) );
HB1xp67_ASAP7_75t_L g303 ( .A(n_262), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_243), .Y(n_304) );
INVx4_ASAP7_75t_L g305 ( .A(n_251), .Y(n_305) );
AND2x4_ASAP7_75t_L g306 ( .A(n_232), .B(n_192), .Y(n_306) );
BUFx3_ASAP7_75t_L g307 ( .A(n_251), .Y(n_307) );
AOI21xp5_ASAP7_75t_L g308 ( .A1(n_274), .A2(n_235), .B(n_250), .Y(n_308) );
AND2x2_ASAP7_75t_L g309 ( .A(n_232), .B(n_185), .Y(n_309) );
OAI21x1_ASAP7_75t_SL g310 ( .A1(n_233), .A2(n_213), .B(n_211), .Y(n_310) );
OAI22xp33_ASAP7_75t_L g311 ( .A1(n_263), .A2(n_233), .B1(n_268), .B2(n_265), .Y(n_311) );
AND2x4_ASAP7_75t_L g312 ( .A(n_232), .B(n_192), .Y(n_312) );
INVx2_ASAP7_75t_L g313 ( .A(n_238), .Y(n_313) );
BUFx2_ASAP7_75t_L g314 ( .A(n_263), .Y(n_314) );
AOI22xp33_ASAP7_75t_L g315 ( .A1(n_290), .A2(n_231), .B1(n_230), .B2(n_217), .Y(n_315) );
AOI22xp33_ASAP7_75t_L g316 ( .A1(n_290), .A2(n_231), .B1(n_217), .B2(n_228), .Y(n_316) );
BUFx12f_ASAP7_75t_L g317 ( .A(n_279), .Y(n_317) );
AND2x2_ASAP7_75t_L g318 ( .A(n_244), .B(n_202), .Y(n_318) );
HB1xp67_ASAP7_75t_L g319 ( .A(n_248), .Y(n_319) );
OAI22xp33_ASAP7_75t_L g320 ( .A1(n_265), .A2(n_195), .B1(n_206), .B2(n_203), .Y(n_320) );
INVx2_ASAP7_75t_L g321 ( .A(n_270), .Y(n_321) );
AND2x4_ASAP7_75t_L g322 ( .A(n_245), .B(n_196), .Y(n_322) );
NAND2xp5_ASAP7_75t_SL g323 ( .A(n_251), .B(n_215), .Y(n_323) );
OR2x2_ASAP7_75t_L g324 ( .A(n_257), .B(n_198), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_275), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_275), .Y(n_326) );
AOI21xp5_ASAP7_75t_L g327 ( .A1(n_250), .A2(n_196), .B(n_209), .Y(n_327) );
AND2x2_ASAP7_75t_L g328 ( .A(n_248), .B(n_202), .Y(n_328) );
AOI22xp33_ASAP7_75t_L g329 ( .A1(n_290), .A2(n_217), .B1(n_228), .B2(n_196), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_282), .B(n_191), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_285), .Y(n_331) );
HB1xp67_ASAP7_75t_L g332 ( .A(n_245), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_285), .Y(n_333) );
NAND2xp5_ASAP7_75t_SL g334 ( .A(n_251), .B(n_215), .Y(n_334) );
BUFx2_ASAP7_75t_L g335 ( .A(n_258), .Y(n_335) );
NAND2x1p5_ASAP7_75t_L g336 ( .A(n_251), .B(n_210), .Y(n_336) );
AOI22xp5_ASAP7_75t_L g337 ( .A1(n_282), .A2(n_216), .B1(n_220), .B2(n_208), .Y(n_337) );
AND2x2_ASAP7_75t_SL g338 ( .A(n_236), .B(n_191), .Y(n_338) );
AND2x4_ASAP7_75t_L g339 ( .A(n_245), .B(n_178), .Y(n_339) );
BUFx3_ASAP7_75t_L g340 ( .A(n_254), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_293), .B(n_204), .Y(n_341) );
INVx2_ASAP7_75t_L g342 ( .A(n_270), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_287), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_293), .B(n_210), .Y(n_344) );
HB1xp67_ASAP7_75t_L g345 ( .A(n_245), .Y(n_345) );
AOI22x1_ASAP7_75t_L g346 ( .A1(n_247), .A2(n_209), .B1(n_221), .B2(n_172), .Y(n_346) );
NAND2x1p5_ASAP7_75t_L g347 ( .A(n_254), .B(n_226), .Y(n_347) );
BUFx2_ASAP7_75t_L g348 ( .A(n_258), .Y(n_348) );
NOR2xp67_ASAP7_75t_L g349 ( .A(n_293), .B(n_190), .Y(n_349) );
INVx2_ASAP7_75t_L g350 ( .A(n_321), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_301), .Y(n_351) );
AND2x2_ASAP7_75t_L g352 ( .A(n_306), .B(n_290), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_301), .Y(n_353) );
INVx8_ASAP7_75t_L g354 ( .A(n_306), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_304), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_304), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_325), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_325), .Y(n_358) );
INVx5_ASAP7_75t_L g359 ( .A(n_305), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_326), .Y(n_360) );
AOI22xp33_ASAP7_75t_L g361 ( .A1(n_338), .A2(n_306), .B1(n_312), .B2(n_309), .Y(n_361) );
INVx1_ASAP7_75t_SL g362 ( .A(n_324), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_306), .B(n_281), .Y(n_363) );
OAI21x1_ASAP7_75t_L g364 ( .A1(n_346), .A2(n_247), .B(n_252), .Y(n_364) );
OAI21xp5_ASAP7_75t_L g365 ( .A1(n_308), .A2(n_260), .B(n_252), .Y(n_365) );
INVx8_ASAP7_75t_L g366 ( .A(n_312), .Y(n_366) );
AOI22xp33_ASAP7_75t_L g367 ( .A1(n_338), .A2(n_281), .B1(n_206), .B2(n_294), .Y(n_367) );
BUFx2_ASAP7_75t_L g368 ( .A(n_314), .Y(n_368) );
INVx1_ASAP7_75t_SL g369 ( .A(n_324), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_326), .Y(n_370) );
AOI21xp33_ASAP7_75t_L g371 ( .A1(n_320), .A2(n_280), .B(n_242), .Y(n_371) );
OR2x6_ASAP7_75t_L g372 ( .A(n_312), .B(n_239), .Y(n_372) );
INVx2_ASAP7_75t_L g373 ( .A(n_321), .Y(n_373) );
OAI22xp5_ASAP7_75t_L g374 ( .A1(n_315), .A2(n_258), .B1(n_259), .B2(n_249), .Y(n_374) );
OR2x6_ASAP7_75t_L g375 ( .A(n_312), .B(n_239), .Y(n_375) );
INVx2_ASAP7_75t_L g376 ( .A(n_321), .Y(n_376) );
BUFx6f_ASAP7_75t_L g377 ( .A(n_307), .Y(n_377) );
AOI22xp33_ASAP7_75t_L g378 ( .A1(n_338), .A2(n_281), .B1(n_273), .B2(n_253), .Y(n_378) );
BUFx6f_ASAP7_75t_L g379 ( .A(n_307), .Y(n_379) );
OAI22xp5_ASAP7_75t_L g380 ( .A1(n_316), .A2(n_259), .B1(n_292), .B2(n_253), .Y(n_380) );
AOI22xp5_ASAP7_75t_SL g381 ( .A1(n_368), .A2(n_237), .B1(n_339), .B2(n_314), .Y(n_381) );
HB1xp67_ASAP7_75t_L g382 ( .A(n_362), .Y(n_382) );
AOI22xp33_ASAP7_75t_L g383 ( .A1(n_367), .A2(n_237), .B1(n_339), .B2(n_317), .Y(n_383) );
AOI22xp33_ASAP7_75t_L g384 ( .A1(n_378), .A2(n_339), .B1(n_317), .B2(n_318), .Y(n_384) );
AOI22xp33_ASAP7_75t_L g385 ( .A1(n_371), .A2(n_339), .B1(n_317), .B2(n_318), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_351), .Y(n_386) );
AOI22xp5_ASAP7_75t_L g387 ( .A1(n_380), .A2(n_311), .B1(n_369), .B2(n_361), .Y(n_387) );
BUFx6f_ASAP7_75t_L g388 ( .A(n_377), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_353), .Y(n_389) );
AND2x2_ASAP7_75t_L g390 ( .A(n_352), .B(n_309), .Y(n_390) );
HB1xp67_ASAP7_75t_L g391 ( .A(n_368), .Y(n_391) );
OAI22xp5_ASAP7_75t_L g392 ( .A1(n_363), .A2(n_329), .B1(n_333), .B2(n_343), .Y(n_392) );
AOI21x1_ASAP7_75t_L g393 ( .A1(n_364), .A2(n_310), .B(n_283), .Y(n_393) );
AOI22xp33_ASAP7_75t_L g394 ( .A1(n_374), .A2(n_352), .B1(n_310), .B2(n_354), .Y(n_394) );
AOI22xp5_ASAP7_75t_L g395 ( .A1(n_353), .A2(n_328), .B1(n_291), .B2(n_289), .Y(n_395) );
AOI22xp33_ASAP7_75t_L g396 ( .A1(n_354), .A2(n_328), .B1(n_345), .B2(n_332), .Y(n_396) );
AOI22xp33_ASAP7_75t_L g397 ( .A1(n_354), .A2(n_295), .B1(n_303), .B2(n_255), .Y(n_397) );
AOI22xp33_ASAP7_75t_L g398 ( .A1(n_354), .A2(n_255), .B1(n_291), .B2(n_273), .Y(n_398) );
INVx2_ASAP7_75t_L g399 ( .A(n_373), .Y(n_399) );
AOI221xp5_ASAP7_75t_L g400 ( .A1(n_357), .A2(n_302), .B1(n_218), .B2(n_273), .C(n_257), .Y(n_400) );
AOI221xp5_ASAP7_75t_L g401 ( .A1(n_357), .A2(n_273), .B1(n_261), .B2(n_276), .C(n_341), .Y(n_401) );
OAI22xp5_ASAP7_75t_L g402 ( .A1(n_355), .A2(n_331), .B1(n_333), .B2(n_343), .Y(n_402) );
HB1xp67_ASAP7_75t_L g403 ( .A(n_359), .Y(n_403) );
AOI221xp5_ASAP7_75t_L g404 ( .A1(n_358), .A2(n_341), .B1(n_284), .B2(n_299), .C(n_330), .Y(n_404) );
INVx2_ASAP7_75t_SL g405 ( .A(n_359), .Y(n_405) );
INVx5_ASAP7_75t_SL g406 ( .A(n_388), .Y(n_406) );
NAND2xp5_ASAP7_75t_SL g407 ( .A(n_381), .B(n_359), .Y(n_407) );
AOI221xp5_ASAP7_75t_L g408 ( .A1(n_400), .A2(n_358), .B1(n_370), .B2(n_360), .C(n_356), .Y(n_408) );
OAI221xp5_ASAP7_75t_L g409 ( .A1(n_383), .A2(n_319), .B1(n_375), .B2(n_372), .C(n_337), .Y(n_409) );
OR2x2_ASAP7_75t_L g410 ( .A(n_399), .B(n_391), .Y(n_410) );
AOI22xp33_ASAP7_75t_L g411 ( .A1(n_385), .A2(n_354), .B1(n_366), .B2(n_291), .Y(n_411) );
OAI221xp5_ASAP7_75t_SL g412 ( .A1(n_384), .A2(n_337), .B1(n_264), .B2(n_375), .C(n_372), .Y(n_412) );
AND2x2_ASAP7_75t_L g413 ( .A(n_399), .B(n_373), .Y(n_413) );
OAI221xp5_ASAP7_75t_L g414 ( .A1(n_397), .A2(n_372), .B1(n_375), .B2(n_330), .C(n_349), .Y(n_414) );
AOI221xp5_ASAP7_75t_L g415 ( .A1(n_404), .A2(n_370), .B1(n_360), .B2(n_356), .C(n_355), .Y(n_415) );
OAI21xp33_ASAP7_75t_L g416 ( .A1(n_395), .A2(n_365), .B(n_247), .Y(n_416) );
INVx2_ASAP7_75t_L g417 ( .A(n_399), .Y(n_417) );
OR2x2_ASAP7_75t_L g418 ( .A(n_386), .B(n_373), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_386), .Y(n_419) );
AOI22xp33_ASAP7_75t_L g420 ( .A1(n_394), .A2(n_366), .B1(n_289), .B2(n_375), .Y(n_420) );
NAND3xp33_ASAP7_75t_L g421 ( .A(n_395), .B(n_359), .C(n_169), .Y(n_421) );
AO21x2_ASAP7_75t_L g422 ( .A1(n_393), .A2(n_327), .B(n_376), .Y(n_422) );
OAI221xp5_ASAP7_75t_L g423 ( .A1(n_398), .A2(n_372), .B1(n_375), .B2(n_349), .C(n_335), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_389), .Y(n_424) );
OAI211xp5_ASAP7_75t_SL g425 ( .A1(n_382), .A2(n_176), .B(n_334), .C(n_323), .Y(n_425) );
OAI31xp33_ASAP7_75t_L g426 ( .A1(n_392), .A2(n_322), .A3(n_348), .B(n_335), .Y(n_426) );
AND2x2_ASAP7_75t_L g427 ( .A(n_390), .B(n_376), .Y(n_427) );
INVx2_ASAP7_75t_L g428 ( .A(n_388), .Y(n_428) );
NOR2xp33_ASAP7_75t_L g429 ( .A(n_381), .B(n_366), .Y(n_429) );
AND2x4_ASAP7_75t_L g430 ( .A(n_405), .B(n_403), .Y(n_430) );
AO21x2_ASAP7_75t_L g431 ( .A1(n_392), .A2(n_350), .B(n_289), .Y(n_431) );
NOR2x1_ASAP7_75t_L g432 ( .A(n_402), .B(n_305), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_402), .Y(n_433) );
AOI221xp5_ASAP7_75t_L g434 ( .A1(n_401), .A2(n_366), .B1(n_331), .B2(n_344), .C(n_246), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_405), .Y(n_435) );
NOR2xp67_ASAP7_75t_SL g436 ( .A(n_421), .B(n_359), .Y(n_436) );
AOI22xp5_ASAP7_75t_L g437 ( .A1(n_434), .A2(n_387), .B1(n_429), .B2(n_409), .Y(n_437) );
INVx3_ASAP7_75t_L g438 ( .A(n_406), .Y(n_438) );
AND2x2_ASAP7_75t_L g439 ( .A(n_413), .B(n_388), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_419), .Y(n_440) );
AND2x2_ASAP7_75t_L g441 ( .A(n_424), .B(n_388), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_424), .B(n_388), .Y(n_442) );
INVx2_ASAP7_75t_L g443 ( .A(n_417), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_433), .Y(n_444) );
INVx2_ASAP7_75t_L g445 ( .A(n_417), .Y(n_445) );
INVx4_ASAP7_75t_L g446 ( .A(n_430), .Y(n_446) );
NOR3xp33_ASAP7_75t_SL g447 ( .A(n_407), .B(n_241), .C(n_240), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_433), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_427), .B(n_396), .Y(n_449) );
AOI33xp33_ASAP7_75t_L g450 ( .A1(n_411), .A2(n_172), .A3(n_168), .B1(n_173), .B2(n_174), .B3(n_182), .Y(n_450) );
AND2x4_ASAP7_75t_L g451 ( .A(n_432), .B(n_359), .Y(n_451) );
OAI21xp5_ASAP7_75t_L g452 ( .A1(n_420), .A2(n_300), .B(n_313), .Y(n_452) );
AND2x2_ASAP7_75t_L g453 ( .A(n_427), .B(n_313), .Y(n_453) );
AND2x2_ASAP7_75t_L g454 ( .A(n_418), .B(n_300), .Y(n_454) );
OAI22xp5_ASAP7_75t_L g455 ( .A1(n_412), .A2(n_300), .B1(n_342), .B2(n_379), .Y(n_455) );
AND2x2_ASAP7_75t_L g456 ( .A(n_418), .B(n_342), .Y(n_456) );
AND2x2_ASAP7_75t_L g457 ( .A(n_410), .B(n_342), .Y(n_457) );
BUFx2_ASAP7_75t_L g458 ( .A(n_430), .Y(n_458) );
INVx2_ASAP7_75t_L g459 ( .A(n_428), .Y(n_459) );
A2O1A1Ixp33_ASAP7_75t_L g460 ( .A1(n_426), .A2(n_322), .B(n_348), .C(n_307), .Y(n_460) );
OAI33xp33_ASAP7_75t_L g461 ( .A1(n_425), .A2(n_173), .A3(n_182), .B1(n_174), .B2(n_168), .B3(n_21), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_415), .B(n_379), .Y(n_462) );
AO31x2_ASAP7_75t_L g463 ( .A1(n_428), .A2(n_344), .A3(n_246), .B(n_287), .Y(n_463) );
NAND4xp25_ASAP7_75t_L g464 ( .A(n_408), .B(n_322), .C(n_23), .D(n_24), .Y(n_464) );
AND2x2_ASAP7_75t_L g465 ( .A(n_431), .B(n_379), .Y(n_465) );
OR2x2_ASAP7_75t_L g466 ( .A(n_435), .B(n_379), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_431), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_431), .B(n_377), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_435), .Y(n_469) );
AOI221xp5_ASAP7_75t_L g470 ( .A1(n_414), .A2(n_322), .B1(n_221), .B2(n_169), .C(n_305), .Y(n_470) );
OAI211xp5_ASAP7_75t_L g471 ( .A1(n_423), .A2(n_305), .B(n_346), .C(n_340), .Y(n_471) );
AND2x4_ASAP7_75t_L g472 ( .A(n_422), .B(n_377), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_422), .Y(n_473) );
OA21x2_ASAP7_75t_L g474 ( .A1(n_416), .A2(n_278), .B(n_277), .Y(n_474) );
INVx2_ASAP7_75t_L g475 ( .A(n_443), .Y(n_475) );
INVx2_ASAP7_75t_L g476 ( .A(n_445), .Y(n_476) );
AOI22xp5_ASAP7_75t_L g477 ( .A1(n_464), .A2(n_377), .B1(n_406), .B2(n_340), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_457), .B(n_221), .Y(n_478) );
AND2x2_ASAP7_75t_L g479 ( .A(n_441), .B(n_221), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_454), .B(n_221), .Y(n_480) );
AND2x2_ASAP7_75t_L g481 ( .A(n_441), .B(n_41), .Y(n_481) );
AND2x2_ASAP7_75t_L g482 ( .A(n_442), .B(n_42), .Y(n_482) );
NOR3xp33_ASAP7_75t_L g483 ( .A(n_461), .B(n_266), .C(n_271), .Y(n_483) );
INVx2_ASAP7_75t_L g484 ( .A(n_445), .Y(n_484) );
OAI21x1_ASAP7_75t_L g485 ( .A1(n_473), .A2(n_347), .B(n_336), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_454), .B(n_286), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_440), .Y(n_487) );
AND2x2_ASAP7_75t_L g488 ( .A(n_442), .B(n_54), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_440), .B(n_286), .Y(n_489) );
OAI33xp33_ASAP7_75t_L g490 ( .A1(n_469), .A2(n_277), .A3(n_278), .B1(n_59), .B2(n_62), .B3(n_66), .Y(n_490) );
OR2x2_ASAP7_75t_L g491 ( .A(n_444), .B(n_347), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_444), .Y(n_492) );
BUFx2_ASAP7_75t_L g493 ( .A(n_446), .Y(n_493) );
OR2x2_ASAP7_75t_L g494 ( .A(n_448), .B(n_347), .Y(n_494) );
AND2x4_ASAP7_75t_L g495 ( .A(n_465), .B(n_55), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_448), .Y(n_496) );
AND2x2_ASAP7_75t_L g497 ( .A(n_439), .B(n_56), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_456), .B(n_453), .Y(n_498) );
NOR4xp25_ASAP7_75t_SL g499 ( .A(n_458), .B(n_68), .C(n_69), .D(n_336), .Y(n_499) );
AND2x2_ASAP7_75t_L g500 ( .A(n_439), .B(n_169), .Y(n_500) );
NAND2xp33_ASAP7_75t_SL g501 ( .A(n_446), .B(n_254), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_473), .Y(n_502) );
INVx2_ASAP7_75t_L g503 ( .A(n_459), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_459), .Y(n_504) );
A2O1A1Ixp33_ASAP7_75t_L g505 ( .A1(n_437), .A2(n_340), .B(n_296), .C(n_288), .Y(n_505) );
HB1xp67_ASAP7_75t_L g506 ( .A(n_463), .Y(n_506) );
NAND5xp2_ASAP7_75t_L g507 ( .A(n_437), .B(n_254), .C(n_296), .D(n_288), .E(n_272), .Y(n_507) );
NOR3xp33_ASAP7_75t_SL g508 ( .A(n_455), .B(n_266), .C(n_271), .Y(n_508) );
NOR2x1_ASAP7_75t_L g509 ( .A(n_446), .B(n_271), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_453), .B(n_169), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_467), .Y(n_511) );
OAI221xp5_ASAP7_75t_L g512 ( .A1(n_470), .A2(n_266), .B1(n_254), .B2(n_272), .C(n_269), .Y(n_512) );
AOI31xp33_ASAP7_75t_L g513 ( .A1(n_455), .A2(n_256), .A3(n_267), .B(n_269), .Y(n_513) );
INVx2_ASAP7_75t_L g514 ( .A(n_475), .Y(n_514) );
AND2x4_ASAP7_75t_SL g515 ( .A(n_497), .B(n_446), .Y(n_515) );
AOI21xp5_ASAP7_75t_L g516 ( .A1(n_501), .A2(n_513), .B(n_490), .Y(n_516) );
AND2x2_ASAP7_75t_L g517 ( .A(n_493), .B(n_468), .Y(n_517) );
INVxp67_ASAP7_75t_SL g518 ( .A(n_506), .Y(n_518) );
NAND2xp33_ASAP7_75t_SL g519 ( .A(n_508), .B(n_436), .Y(n_519) );
NAND3xp33_ASAP7_75t_SL g520 ( .A(n_477), .B(n_450), .C(n_460), .Y(n_520) );
OAI221xp5_ASAP7_75t_L g521 ( .A1(n_477), .A2(n_449), .B1(n_447), .B2(n_471), .C(n_462), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_487), .B(n_463), .Y(n_522) );
NOR2x1_ASAP7_75t_L g523 ( .A(n_509), .B(n_438), .Y(n_523) );
NOR2xp33_ASAP7_75t_SL g524 ( .A(n_495), .B(n_497), .Y(n_524) );
AOI21xp5_ASAP7_75t_L g525 ( .A1(n_507), .A2(n_474), .B(n_451), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_498), .B(n_463), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_492), .B(n_463), .Y(n_527) );
AOI221xp5_ASAP7_75t_L g528 ( .A1(n_511), .A2(n_452), .B1(n_472), .B2(n_438), .C(n_466), .Y(n_528) );
AOI22xp5_ASAP7_75t_L g529 ( .A1(n_495), .A2(n_472), .B1(n_452), .B2(n_474), .Y(n_529) );
OR2x6_ASAP7_75t_L g530 ( .A(n_495), .B(n_474), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_496), .Y(n_531) );
OAI21xp33_ASAP7_75t_L g532 ( .A1(n_511), .A2(n_269), .B(n_297), .Y(n_532) );
O2A1O1Ixp5_ASAP7_75t_L g533 ( .A1(n_502), .A2(n_298), .B(n_486), .C(n_488), .Y(n_533) );
NAND2xp33_ASAP7_75t_L g534 ( .A(n_481), .B(n_482), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_502), .Y(n_535) );
O2A1O1Ixp33_ASAP7_75t_SL g536 ( .A1(n_505), .A2(n_494), .B(n_491), .C(n_489), .Y(n_536) );
INVxp67_ASAP7_75t_L g537 ( .A(n_524), .Y(n_537) );
INVxp67_ASAP7_75t_L g538 ( .A(n_534), .Y(n_538) );
AOI21xp5_ASAP7_75t_L g539 ( .A1(n_519), .A2(n_510), .B(n_478), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_535), .Y(n_540) );
XNOR2x2_ASAP7_75t_L g541 ( .A(n_520), .B(n_481), .Y(n_541) );
INVx2_ASAP7_75t_L g542 ( .A(n_514), .Y(n_542) );
HB1xp67_ASAP7_75t_L g543 ( .A(n_517), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_526), .B(n_504), .Y(n_544) );
OR2x2_ASAP7_75t_L g545 ( .A(n_518), .B(n_503), .Y(n_545) );
XNOR2xp5_ASAP7_75t_L g546 ( .A(n_515), .B(n_500), .Y(n_546) );
INVx3_ASAP7_75t_L g547 ( .A(n_530), .Y(n_547) );
AOI21xp5_ASAP7_75t_L g548 ( .A1(n_516), .A2(n_480), .B(n_499), .Y(n_548) );
INVx3_ASAP7_75t_L g549 ( .A(n_530), .Y(n_549) );
AND2x2_ASAP7_75t_L g550 ( .A(n_530), .B(n_476), .Y(n_550) );
NOR3xp33_ASAP7_75t_SL g551 ( .A(n_521), .B(n_512), .C(n_483), .Y(n_551) );
NOR3xp33_ASAP7_75t_SL g552 ( .A(n_521), .B(n_479), .C(n_485), .Y(n_552) );
NAND3x1_ASAP7_75t_SL g553 ( .A(n_541), .B(n_523), .C(n_552), .Y(n_553) );
INVx1_ASAP7_75t_SL g554 ( .A(n_546), .Y(n_554) );
HB1xp67_ASAP7_75t_L g555 ( .A(n_545), .Y(n_555) );
INVx2_ASAP7_75t_L g556 ( .A(n_545), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_540), .Y(n_557) );
INVx2_ASAP7_75t_L g558 ( .A(n_542), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_544), .B(n_531), .Y(n_559) );
AOI221xp5_ASAP7_75t_L g560 ( .A1(n_538), .A2(n_528), .B1(n_536), .B2(n_527), .C(n_522), .Y(n_560) );
OR2x2_ASAP7_75t_L g561 ( .A(n_543), .B(n_476), .Y(n_561) );
INVx2_ASAP7_75t_L g562 ( .A(n_542), .Y(n_562) );
OA22x2_ASAP7_75t_L g563 ( .A1(n_547), .A2(n_529), .B1(n_532), .B2(n_484), .Y(n_563) );
NAND3xp33_ASAP7_75t_L g564 ( .A(n_551), .B(n_528), .C(n_533), .Y(n_564) );
OAI21xp5_ASAP7_75t_L g565 ( .A1(n_564), .A2(n_548), .B(n_525), .Y(n_565) );
HB1xp67_ASAP7_75t_L g566 ( .A(n_555), .Y(n_566) );
OAI221xp5_ASAP7_75t_SL g567 ( .A1(n_554), .A2(n_549), .B1(n_550), .B2(n_546), .C(n_539), .Y(n_567) );
NOR2xp33_ASAP7_75t_R g568 ( .A(n_553), .B(n_561), .Y(n_568) );
OAI211xp5_ASAP7_75t_L g569 ( .A1(n_553), .A2(n_559), .B(n_556), .C(n_557), .Y(n_569) );
OAI22xp5_ASAP7_75t_L g570 ( .A1(n_558), .A2(n_538), .B1(n_554), .B2(n_552), .Y(n_570) );
AOI31xp33_ASAP7_75t_SL g571 ( .A1(n_562), .A2(n_538), .A3(n_537), .B(n_560), .Y(n_571) );
OAI22xp5_ASAP7_75t_L g572 ( .A1(n_554), .A2(n_538), .B1(n_552), .B2(n_537), .Y(n_572) );
AOI21xp5_ASAP7_75t_L g573 ( .A1(n_564), .A2(n_563), .B(n_560), .Y(n_573) );
CKINVDCx5p33_ASAP7_75t_R g574 ( .A(n_568), .Y(n_574) );
CKINVDCx20_ASAP7_75t_R g575 ( .A(n_565), .Y(n_575) );
NOR2x1_ASAP7_75t_L g576 ( .A(n_571), .B(n_569), .Y(n_576) );
INVx2_ASAP7_75t_L g577 ( .A(n_566), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_577), .Y(n_578) );
XNOR2xp5_ASAP7_75t_L g579 ( .A(n_574), .B(n_572), .Y(n_579) );
HB1xp67_ASAP7_75t_L g580 ( .A(n_577), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_580), .Y(n_581) );
AOI22xp33_ASAP7_75t_L g582 ( .A1(n_579), .A2(n_576), .B1(n_575), .B2(n_573), .Y(n_582) );
XNOR2xp5_ASAP7_75t_L g583 ( .A(n_582), .B(n_579), .Y(n_583) );
HB1xp67_ASAP7_75t_L g584 ( .A(n_581), .Y(n_584) );
NAND3xp33_ASAP7_75t_L g585 ( .A(n_583), .B(n_578), .C(n_570), .Y(n_585) );
AOI21xp5_ASAP7_75t_L g586 ( .A1(n_585), .A2(n_584), .B(n_567), .Y(n_586) );
endmodule