module fake_jpeg_4085_n_49 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_49);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_49;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_43;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx3_ASAP7_75t_L g7 ( 
.A(n_3),
.Y(n_7)
);

BUFx6f_ASAP7_75t_L g8 ( 
.A(n_5),
.Y(n_8)
);

BUFx3_ASAP7_75t_L g9 ( 
.A(n_0),
.Y(n_9)
);

NOR2xp33_ASAP7_75t_L g10 ( 
.A(n_0),
.B(n_1),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

INVx13_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

BUFx3_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

INVx8_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_10),
.B(n_0),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_16),
.B(n_21),
.Y(n_34)
);

OAI21xp5_ASAP7_75t_L g17 ( 
.A1(n_12),
.A2(n_1),
.B(n_2),
.Y(n_17)
);

AOI21xp5_ASAP7_75t_L g31 ( 
.A1(n_17),
.A2(n_18),
.B(n_25),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g18 ( 
.A(n_11),
.B(n_2),
.C(n_4),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_SL g20 ( 
.A(n_7),
.B(n_6),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_20),
.Y(n_27)
);

AND2x2_ASAP7_75t_L g21 ( 
.A(n_12),
.B(n_8),
.Y(n_21)
);

OAI22xp33_ASAP7_75t_L g22 ( 
.A1(n_11),
.A2(n_8),
.B1(n_15),
.B2(n_9),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_22),
.A2(n_23),
.B1(n_19),
.B2(n_17),
.Y(n_26)
);

AO22x1_ASAP7_75t_SL g23 ( 
.A1(n_15),
.A2(n_9),
.B1(n_14),
.B2(n_13),
.Y(n_23)
);

CKINVDCx16_ASAP7_75t_R g24 ( 
.A(n_14),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_24),
.B(n_22),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g25 ( 
.A1(n_7),
.A2(n_14),
.B1(n_15),
.B2(n_8),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_26),
.B(n_30),
.C(n_35),
.Y(n_38)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_21),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_28),
.B(n_29),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_23),
.Y(n_32)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_18),
.Y(n_33)
);

CKINVDCx14_ASAP7_75t_R g37 ( 
.A(n_33),
.Y(n_37)
);

XOR2xp5_ASAP7_75t_L g39 ( 
.A(n_34),
.B(n_26),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_39),
.B(n_31),
.C(n_35),
.Y(n_42)
);

XOR2x1_ASAP7_75t_L g40 ( 
.A(n_34),
.B(n_29),
.Y(n_40)
);

XOR2xp5_ASAP7_75t_L g43 ( 
.A(n_40),
.B(n_39),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_42),
.B(n_43),
.C(n_38),
.Y(n_46)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_41),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_44),
.B(n_27),
.Y(n_45)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_45),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_47),
.A2(n_36),
.B1(n_37),
.B2(n_40),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_L g49 ( 
.A1(n_48),
.A2(n_31),
.B(n_46),
.Y(n_49)
);


endmodule