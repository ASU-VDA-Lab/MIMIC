module fake_jpeg_19415_n_124 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_124);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_124;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_49;
wire n_76;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_29),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_11),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_28),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_7),
.Y(n_48)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_41),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_1),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_13),
.Y(n_52)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_12),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_10),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_21),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_4),
.Y(n_57)
);

BUFx16f_ASAP7_75t_L g58 ( 
.A(n_22),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_5),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_19),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_48),
.B(n_0),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_62),
.B(n_57),
.Y(n_72)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_63),
.Y(n_70)
);

NAND3xp33_ASAP7_75t_L g64 ( 
.A(n_51),
.B(n_0),
.C(n_1),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_64),
.B(n_58),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_65),
.Y(n_76)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_58),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_66),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_67),
.Y(n_79)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_60),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_68),
.B(n_60),
.Y(n_71)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_69),
.Y(n_77)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_71),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_72),
.B(n_80),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_66),
.A2(n_49),
.B1(n_53),
.B2(n_43),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_73),
.A2(n_74),
.B1(n_56),
.B2(n_52),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_65),
.A2(n_61),
.B1(n_47),
.B2(n_50),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_67),
.Y(n_75)
);

INVx13_ASAP7_75t_L g82 ( 
.A(n_75),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_77),
.B(n_2),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_81),
.B(n_83),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_76),
.B(n_2),
.Y(n_83)
);

AND2x6_ASAP7_75t_L g84 ( 
.A(n_74),
.B(n_64),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_84),
.B(n_20),
.Y(n_96)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_78),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_86),
.Y(n_99)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_78),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_87),
.B(n_90),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_88),
.A2(n_89),
.B1(n_94),
.B2(n_90),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_73),
.A2(n_56),
.B1(n_55),
.B2(n_46),
.Y(n_89)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_76),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_70),
.A2(n_52),
.B1(n_55),
.B2(n_46),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_92),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_79),
.B(n_3),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_93),
.B(n_3),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_80),
.A2(n_44),
.B1(n_59),
.B2(n_23),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_85),
.B(n_84),
.C(n_91),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_95),
.B(n_8),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_96),
.B(n_98),
.Y(n_109)
);

OAI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_87),
.A2(n_18),
.B1(n_39),
.B2(n_38),
.Y(n_101)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_101),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_92),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_102),
.B(n_103),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_82),
.B(n_4),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_104),
.B(n_105),
.Y(n_111)
);

AND2x2_ASAP7_75t_SL g106 ( 
.A(n_82),
.B(n_26),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_SL g107 ( 
.A(n_106),
.B(n_6),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_107),
.B(n_108),
.C(n_106),
.Y(n_114)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_97),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_113),
.A2(n_99),
.B1(n_101),
.B2(n_100),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_114),
.B(n_115),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_110),
.A2(n_95),
.B(n_106),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_117),
.B(n_108),
.C(n_109),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_118),
.B(n_107),
.C(n_116),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_119),
.B(n_111),
.Y(n_120)
);

AOI322xp5_ASAP7_75t_L g121 ( 
.A1(n_120),
.A2(n_112),
.A3(n_9),
.B1(n_14),
.B2(n_15),
.C1(n_16),
.C2(n_17),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_121),
.A2(n_31),
.B(n_25),
.Y(n_122)
);

OAI21xp33_ASAP7_75t_R g123 ( 
.A1(n_122),
.A2(n_27),
.B(n_30),
.Y(n_123)
);

AOI221xp5_ASAP7_75t_L g124 ( 
.A1(n_123),
.A2(n_32),
.B1(n_34),
.B2(n_35),
.C(n_42),
.Y(n_124)
);


endmodule