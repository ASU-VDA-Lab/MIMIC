module real_jpeg_20360_n_11 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_10, n_9, n_11);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_11;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_104;
wire n_153;
wire n_64;
wire n_47;
wire n_131;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_140;
wire n_126;
wire n_13;
wire n_113;
wire n_155;
wire n_120;
wire n_93;
wire n_141;
wire n_95;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_134;
wire n_72;
wire n_159;
wire n_151;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

INVx13_ASAP7_75t_L g52 ( 
.A(n_0),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g21 ( 
.A1(n_1),
.A2(n_22),
.B1(n_23),
.B2(n_24),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_1),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_1),
.A2(n_24),
.B1(n_47),
.B2(n_48),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_1),
.A2(n_2),
.B1(n_24),
.B2(n_62),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_1),
.A2(n_24),
.B1(n_27),
.B2(n_29),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_2),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_2),
.A2(n_6),
.B1(n_32),
.B2(n_62),
.Y(n_68)
);

A2O1A1Ixp33_ASAP7_75t_L g82 ( 
.A1(n_2),
.A2(n_32),
.B(n_66),
.C(n_83),
.Y(n_82)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_3),
.A2(n_41),
.B(n_100),
.Y(n_99)
);

INVx8_ASAP7_75t_L g141 ( 
.A(n_3),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g47 ( 
.A(n_5),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_6),
.A2(n_22),
.B1(n_23),
.B2(n_32),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_6),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_6),
.A2(n_27),
.B1(n_29),
.B2(n_32),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_6),
.A2(n_32),
.B1(n_47),
.B2(n_48),
.Y(n_54)
);

AOI21xp33_ASAP7_75t_SL g83 ( 
.A1(n_6),
.A2(n_47),
.B(n_65),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_6),
.B(n_63),
.Y(n_97)
);

AOI21xp33_ASAP7_75t_L g112 ( 
.A1(n_6),
.A2(n_9),
.B(n_29),
.Y(n_112)
);

AOI21xp33_ASAP7_75t_SL g136 ( 
.A1(n_6),
.A2(n_23),
.B(n_51),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_7),
.A2(n_27),
.B1(n_29),
.B2(n_38),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_7),
.Y(n_38)
);

INVx13_ASAP7_75t_L g66 ( 
.A(n_8),
.Y(n_66)
);

A2O1A1Ixp33_ASAP7_75t_L g69 ( 
.A1(n_8),
.A2(n_62),
.B(n_64),
.C(n_70),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_8),
.B(n_62),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_9),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_26)
);

INVx6_ASAP7_75t_SL g28 ( 
.A(n_9),
.Y(n_28)
);

OAI22xp33_ASAP7_75t_L g34 ( 
.A1(n_9),
.A2(n_22),
.B1(n_23),
.B2(n_28),
.Y(n_34)
);

BUFx3_ASAP7_75t_SL g23 ( 
.A(n_10),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_103),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_101),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_14),
.Y(n_13)
);

AND2x2_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_86),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_15),
.B(n_86),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_71),
.Y(n_15)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_44),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_SL g17 ( 
.A1(n_18),
.A2(n_19),
.B1(n_35),
.B2(n_36),
.Y(n_17)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_18),
.A2(n_19),
.B1(n_110),
.B2(n_111),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_18),
.A2(n_19),
.B1(n_45),
.B2(n_91),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_19),
.B(n_111),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_19),
.B(n_45),
.C(n_134),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_25),
.B(n_30),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_21),
.A2(n_26),
.B1(n_31),
.B2(n_33),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_22),
.A2(n_23),
.B1(n_51),
.B2(n_52),
.Y(n_50)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

A2O1A1Ixp33_ASAP7_75t_L g111 ( 
.A1(n_23),
.A2(n_28),
.B(n_32),
.C(n_112),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_26),
.B(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_26),
.B(n_33),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_26),
.B(n_32),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_27),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_27),
.B(n_116),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_29),
.B(n_39),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_33),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g58 ( 
.A(n_31),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_32),
.B(n_39),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_32),
.B(n_50),
.Y(n_127)
);

A2O1A1Ixp33_ASAP7_75t_L g135 ( 
.A1(n_32),
.A2(n_47),
.B(n_52),
.C(n_136),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_36),
.Y(n_35)
);

OAI21xp5_ASAP7_75t_SL g36 ( 
.A1(n_37),
.A2(n_39),
.B(n_40),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_39),
.A2(n_42),
.B1(n_43),
.B2(n_85),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_43),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_42),
.B(n_141),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_43),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_57),
.C(n_60),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_45),
.A2(n_57),
.B1(n_90),
.B2(n_91),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_45),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g45 ( 
.A1(n_46),
.A2(n_49),
.B(n_53),
.Y(n_45)
);

CKINVDCx14_ASAP7_75t_R g74 ( 
.A(n_46),
.Y(n_74)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_47),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_47),
.A2(n_48),
.B1(n_65),
.B2(n_66),
.Y(n_64)
);

A2O1A1Ixp33_ASAP7_75t_L g55 ( 
.A1(n_48),
.A2(n_50),
.B(n_51),
.C(n_56),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_48),
.B(n_51),
.Y(n_56)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_50),
.A2(n_54),
.B1(n_55),
.B2(n_74),
.Y(n_73)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_55),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_57),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_59),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_60),
.A2(n_88),
.B1(n_89),
.B2(n_92),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_60),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_63),
.B(n_67),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_61),
.A2(n_63),
.B1(n_76),
.B2(n_77),
.Y(n_75)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_69),
.Y(n_67)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_68),
.Y(n_77)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_69),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_SL g71 ( 
.A(n_72),
.B(n_80),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_75),
.B1(n_78),
.B2(n_79),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_73),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_73),
.B(n_96),
.C(n_98),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_73),
.A2(n_79),
.B1(n_149),
.B2(n_150),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_75),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_84),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_81),
.A2(n_82),
.B1(n_84),
.B2(n_94),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_82),
.Y(n_81)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_84),
.Y(n_94)
);

NOR2x1_ASAP7_75t_R g117 ( 
.A(n_84),
.B(n_118),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_84),
.B(n_118),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_84),
.A2(n_94),
.B1(n_124),
.B2(n_129),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_84),
.B(n_125),
.C(n_127),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_85),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_93),
.C(n_95),
.Y(n_86)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_87),
.B(n_158),
.Y(n_157)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_89),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_93),
.B(n_95),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_96),
.A2(n_97),
.B1(n_98),
.B2(n_99),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_97),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_98),
.B(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_99),
.B(n_109),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_99),
.B(n_109),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_104),
.A2(n_155),
.B(n_159),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g104 ( 
.A1(n_105),
.A2(n_145),
.B(n_154),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_131),
.B(n_144),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_107),
.A2(n_121),
.B(n_130),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_113),
.B(n_120),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_111),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_114),
.A2(n_117),
.B(n_119),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_123),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_122),
.B(n_123),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_124),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_125),
.A2(n_126),
.B1(n_127),
.B2(n_128),
.Y(n_124)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_125),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_125),
.A2(n_128),
.B1(n_152),
.B2(n_153),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_125),
.B(n_148),
.C(n_153),
.Y(n_156)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_133),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_132),
.B(n_133),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_143),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_135),
.A2(n_137),
.B1(n_138),
.B2(n_142),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_135),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_137),
.B(n_142),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_138),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_140),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_147),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_146),
.B(n_147),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_151),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_150),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_152),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_157),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_156),
.B(n_157),
.Y(n_159)
);


endmodule