module fake_netlist_1_4113_n_46 (n_11, n_1, n_2, n_13, n_16, n_12, n_6, n_4, n_3, n_9, n_5, n_14, n_7, n_15, n_10, n_8, n_0, n_46);
input n_11;
input n_1;
input n_2;
input n_13;
input n_16;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_14;
input n_7;
input n_15;
input n_10;
input n_8;
input n_0;
output n_46;
wire n_45;
wire n_20;
wire n_38;
wire n_44;
wire n_36;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_25;
wire n_30;
wire n_33;
wire n_26;
wire n_18;
wire n_32;
wire n_41;
wire n_35;
wire n_17;
wire n_42;
wire n_24;
wire n_19;
wire n_27;
wire n_21;
wire n_43;
wire n_40;
wire n_29;
wire n_39;
NAND2xp5_ASAP7_75t_L g17 ( .A(n_6), .B(n_11), .Y(n_17) );
HB1xp67_ASAP7_75t_L g18 ( .A(n_14), .Y(n_18) );
INVx1_ASAP7_75t_L g19 ( .A(n_15), .Y(n_19) );
INVx1_ASAP7_75t_L g20 ( .A(n_10), .Y(n_20) );
CKINVDCx20_ASAP7_75t_R g21 ( .A(n_3), .Y(n_21) );
INVx1_ASAP7_75t_L g22 ( .A(n_5), .Y(n_22) );
OAI22xp5_ASAP7_75t_SL g23 ( .A1(n_16), .A2(n_7), .B1(n_12), .B2(n_13), .Y(n_23) );
OAI22xp5_ASAP7_75t_SL g24 ( .A1(n_8), .A2(n_4), .B1(n_5), .B2(n_2), .Y(n_24) );
INVx1_ASAP7_75t_L g25 ( .A(n_3), .Y(n_25) );
BUFx6f_ASAP7_75t_L g26 ( .A(n_19), .Y(n_26) );
INVx2_ASAP7_75t_L g27 ( .A(n_19), .Y(n_27) );
OR2x6_ASAP7_75t_L g28 ( .A(n_24), .B(n_0), .Y(n_28) );
NAND2xp5_ASAP7_75t_L g29 ( .A(n_18), .B(n_0), .Y(n_29) );
CKINVDCx6p67_ASAP7_75t_R g30 ( .A(n_29), .Y(n_30) );
OAI21x1_ASAP7_75t_L g31 ( .A1(n_27), .A2(n_20), .B(n_17), .Y(n_31) );
OAI21x1_ASAP7_75t_L g32 ( .A1(n_29), .A2(n_25), .B(n_22), .Y(n_32) );
INVx1_ASAP7_75t_L g33 ( .A(n_32), .Y(n_33) );
INVx1_ASAP7_75t_L g34 ( .A(n_32), .Y(n_34) );
OR2x2_ASAP7_75t_L g35 ( .A(n_33), .B(n_30), .Y(n_35) );
INVx2_ASAP7_75t_L g36 ( .A(n_34), .Y(n_36) );
INVx1_ASAP7_75t_L g37 ( .A(n_36), .Y(n_37) );
INVx2_ASAP7_75t_L g38 ( .A(n_35), .Y(n_38) );
AOI222xp33_ASAP7_75t_L g39 ( .A1(n_36), .A2(n_21), .B1(n_25), .B2(n_23), .C1(n_28), .C2(n_33), .Y(n_39) );
NAND2xp33_ASAP7_75t_SL g40 ( .A(n_37), .B(n_21), .Y(n_40) );
AOI211xp5_ASAP7_75t_L g41 ( .A1(n_38), .A2(n_31), .B(n_26), .C(n_30), .Y(n_41) );
OAI21xp33_ASAP7_75t_L g42 ( .A1(n_41), .A2(n_39), .B(n_28), .Y(n_42) );
AOI221xp5_ASAP7_75t_L g43 ( .A1(n_40), .A2(n_26), .B1(n_28), .B2(n_31), .C(n_6), .Y(n_43) );
BUFx2_ASAP7_75t_L g44 ( .A(n_43), .Y(n_44) );
AOI222xp33_ASAP7_75t_SL g45 ( .A1(n_44), .A2(n_42), .B1(n_7), .B2(n_8), .C1(n_9), .C2(n_1), .Y(n_45) );
INVxp67_ASAP7_75t_L g46 ( .A(n_45), .Y(n_46) );
endmodule