module real_jpeg_29411_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_131;
wire n_47;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_173;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_184;
wire n_200;
wire n_48;
wire n_56;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_178;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_44;
wire n_28;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_195;
wire n_110;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_167;
wire n_128;
wire n_202;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_206;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_0),
.B(n_52),
.Y(n_78)
);

INVx11_ASAP7_75t_L g82 ( 
.A(n_0),
.Y(n_82)
);

INVx5_ASAP7_75t_L g162 ( 
.A(n_0),
.Y(n_162)
);

BUFx12_ASAP7_75t_L g66 ( 
.A(n_1),
.Y(n_66)
);

OAI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_2),
.A2(n_63),
.B1(n_64),
.B2(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_2),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_2),
.A2(n_29),
.B1(n_30),
.B2(n_73),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_2),
.A2(n_36),
.B1(n_37),
.B2(n_73),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_2),
.A2(n_52),
.B1(n_54),
.B2(n_73),
.Y(n_158)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

OAI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_4),
.A2(n_63),
.B1(n_64),
.B2(n_71),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_4),
.Y(n_71)
);

AOI21xp33_ASAP7_75t_SL g76 ( 
.A1(n_4),
.A2(n_30),
.B(n_66),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_4),
.B(n_68),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_4),
.A2(n_36),
.B(n_131),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_4),
.B(n_36),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_4),
.B(n_91),
.Y(n_140)
);

OAI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_4),
.A2(n_102),
.B1(n_158),
.B2(n_162),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_4),
.A2(n_29),
.B(n_174),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_5),
.A2(n_52),
.B1(n_54),
.B2(n_80),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_5),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_5),
.A2(n_36),
.B1(n_37),
.B2(n_80),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_6),
.A2(n_52),
.B1(n_54),
.B2(n_106),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_6),
.Y(n_106)
);

INVx13_ASAP7_75t_L g65 ( 
.A(n_7),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_8),
.A2(n_52),
.B1(n_54),
.B2(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_8),
.Y(n_84)
);

OAI22xp33_ASAP7_75t_L g40 ( 
.A1(n_9),
.A2(n_29),
.B1(n_30),
.B2(n_41),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_9),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_9),
.A2(n_41),
.B1(n_63),
.B2(n_64),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_9),
.A2(n_36),
.B1(n_37),
.B2(n_41),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_9),
.A2(n_41),
.B1(n_52),
.B2(n_54),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_10),
.A2(n_29),
.B1(n_30),
.B2(n_43),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_10),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_L g145 ( 
.A1(n_10),
.A2(n_43),
.B1(n_52),
.B2(n_54),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_10),
.A2(n_36),
.B1(n_37),
.B2(n_43),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_11),
.A2(n_36),
.B1(n_37),
.B2(n_48),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_11),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_11),
.A2(n_29),
.B1(n_30),
.B2(n_48),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_11),
.A2(n_48),
.B1(n_52),
.B2(n_54),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_12),
.A2(n_52),
.B1(n_54),
.B2(n_55),
.Y(n_51)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_12),
.Y(n_55)
);

BUFx24_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

INVx11_ASAP7_75t_SL g53 ( 
.A(n_15),
.Y(n_53)
);

OAI22xp33_ASAP7_75t_L g58 ( 
.A1(n_16),
.A2(n_36),
.B1(n_37),
.B2(n_59),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_16),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_16),
.A2(n_52),
.B1(n_54),
.B2(n_59),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_122),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_120),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_95),
.Y(n_20)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_21),
.B(n_95),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_74),
.C(n_85),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_22),
.B(n_207),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_61),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_44),
.B2(n_45),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_24),
.B(n_45),
.C(n_61),
.Y(n_107)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_26),
.A2(n_33),
.B1(n_39),
.B2(n_42),
.Y(n_25)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_26),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_26),
.A2(n_33),
.B1(n_42),
.B2(n_117),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_26),
.A2(n_33),
.B1(n_89),
.B2(n_173),
.Y(n_172)
);

A2O1A1Ixp33_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_29),
.B(n_32),
.C(n_33),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_27),
.B(n_29),
.Y(n_32)
);

INVx1_ASAP7_75t_SL g27 ( 
.A(n_28),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_28),
.A2(n_34),
.B1(n_36),
.B2(n_37),
.Y(n_33)
);

AO22x1_ASAP7_75t_L g68 ( 
.A1(n_29),
.A2(n_30),
.B1(n_66),
.B2(n_69),
.Y(n_68)
);

OAI32xp33_ASAP7_75t_L g182 ( 
.A1(n_29),
.A2(n_34),
.A3(n_37),
.B1(n_175),
.B2(n_183),
.Y(n_182)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_30),
.B(n_71),
.Y(n_175)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_33),
.Y(n_91)
);

INVx6_ASAP7_75t_L g184 ( 
.A(n_34),
.Y(n_184)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

OAI22xp33_ASAP7_75t_L g56 ( 
.A1(n_36),
.A2(n_37),
.B1(n_55),
.B2(n_57),
.Y(n_56)
);

OAI32xp33_ASAP7_75t_L g134 ( 
.A1(n_36),
.A2(n_54),
.A3(n_57),
.B1(n_135),
.B2(n_136),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_36),
.B(n_184),
.Y(n_183)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_40),
.A2(n_88),
.B1(n_90),
.B2(n_91),
.Y(n_87)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_46),
.A2(n_49),
.B1(n_58),
.B2(n_60),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_47),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_47),
.A2(n_50),
.B1(n_51),
.B2(n_200),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_49),
.A2(n_60),
.B1(n_177),
.B2(n_178),
.Y(n_176)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_50),
.A2(n_51),
.B1(n_99),
.B2(n_100),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_50),
.A2(n_51),
.B1(n_130),
.B2(n_132),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_50),
.A2(n_51),
.B1(n_132),
.B2(n_143),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_51),
.B(n_56),
.Y(n_50)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_51),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_51),
.B(n_71),
.Y(n_159)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_52),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_52),
.B(n_55),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_52),
.B(n_164),
.Y(n_163)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_55),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_58),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_62),
.A2(n_68),
.B1(n_70),
.B2(n_72),
.Y(n_61)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_62),
.Y(n_111)
);

O2A1O1Ixp33_ASAP7_75t_L g62 ( 
.A1(n_63),
.A2(n_66),
.B(n_67),
.C(n_68),
.Y(n_62)
);

NAND2xp33_ASAP7_75t_SL g67 ( 
.A(n_63),
.B(n_66),
.Y(n_67)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

A2O1A1Ixp33_ASAP7_75t_L g75 ( 
.A1(n_64),
.A2(n_69),
.B(n_71),
.C(n_76),
.Y(n_75)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_66),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_68),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_71),
.B(n_82),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_72),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_74),
.A2(n_85),
.B1(n_86),
.B2(n_208),
.Y(n_207)
);

CKINVDCx16_ASAP7_75t_R g208 ( 
.A(n_74),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_77),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_75),
.B(n_77),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_79),
.B1(n_81),
.B2(n_83),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_78),
.A2(n_79),
.B1(n_81),
.B2(n_93),
.Y(n_92)
);

CKINVDCx14_ASAP7_75t_R g102 ( 
.A(n_78),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_78),
.A2(n_81),
.B1(n_151),
.B2(n_153),
.Y(n_150)
);

INVx11_ASAP7_75t_L g104 ( 
.A(n_81),
.Y(n_104)
);

INVx5_ASAP7_75t_SL g147 ( 
.A(n_81),
.Y(n_147)
);

INVx11_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_82),
.A2(n_102),
.B1(n_152),
.B2(n_158),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_83),
.Y(n_103)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_92),
.C(n_94),
.Y(n_86)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_87),
.B(n_195),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_89),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_92),
.B(n_94),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_93),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_108),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_107),
.Y(n_96)
);

XOR2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_101),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_102),
.A2(n_103),
.B1(n_104),
.B2(n_105),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_102),
.A2(n_145),
.B1(n_146),
.B2(n_147),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_102),
.A2(n_146),
.B1(n_147),
.B2(n_186),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_SL g108 ( 
.A(n_109),
.B(n_119),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_116),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_111),
.A2(n_112),
.B1(n_113),
.B2(n_114),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_115),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_118),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_121),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_204),
.B(n_209),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_124),
.A2(n_190),
.B(n_203),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_125),
.A2(n_168),
.B(n_189),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_126),
.A2(n_148),
.B(n_167),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_137),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_127),
.B(n_137),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_128),
.B(n_133),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_128),
.A2(n_129),
.B1(n_133),
.B2(n_134),
.Y(n_154)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_131),
.Y(n_135)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_144),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_139),
.A2(n_140),
.B1(n_141),
.B2(n_142),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_139),
.B(n_142),
.C(n_144),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_143),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_145),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_149),
.A2(n_155),
.B(n_166),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_154),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_150),
.B(n_154),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_152),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_156),
.A2(n_160),
.B(n_165),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_159),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_157),
.B(n_159),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_161),
.B(n_163),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_170),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_169),
.B(n_170),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_171),
.A2(n_181),
.B1(n_187),
.B2(n_188),
.Y(n_170)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_171),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_172),
.A2(n_176),
.B1(n_179),
.B2(n_180),
.Y(n_171)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_172),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_176),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_176),
.B(n_180),
.C(n_188),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_178),
.Y(n_200)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_181),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_185),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_182),
.B(n_185),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_192),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_191),
.B(n_192),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_193),
.A2(n_194),
.B1(n_196),
.B2(n_197),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_193),
.B(n_199),
.C(n_201),
.Y(n_205)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_198),
.A2(n_199),
.B1(n_201),
.B2(n_202),
.Y(n_197)
);

CKINVDCx14_ASAP7_75t_R g201 ( 
.A(n_198),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_199),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_206),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_205),
.B(n_206),
.Y(n_209)
);


endmodule