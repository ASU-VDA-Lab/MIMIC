module fake_ibex_2028_n_3977 (n_151, n_85, n_599, n_507, n_540, n_395, n_84, n_64, n_171, n_103, n_529, n_389, n_204, n_626, n_274, n_387, n_688, n_130, n_177, n_707, n_76, n_273, n_309, n_330, n_9, n_328, n_293, n_341, n_372, n_124, n_37, n_256, n_418, n_193, n_510, n_446, n_108, n_350, n_601, n_621, n_610, n_165, n_452, n_86, n_70, n_664, n_255, n_175, n_586, n_638, n_398, n_59, n_28, n_125, n_304, n_191, n_593, n_5, n_62, n_71, n_153, n_545, n_583, n_678, n_663, n_194, n_249, n_334, n_634, n_733, n_312, n_622, n_578, n_478, n_239, n_94, n_134, n_432, n_371, n_403, n_423, n_608, n_357, n_88, n_412, n_457, n_494, n_142, n_226, n_336, n_258, n_40, n_90, n_17, n_74, n_449, n_547, n_176, n_727, n_58, n_43, n_216, n_33, n_652, n_421, n_738, n_475, n_166, n_163, n_645, n_500, n_542, n_114, n_236, n_34, n_376, n_377, n_584, n_531, n_647, n_15, n_556, n_24, n_189, n_498, n_698, n_280, n_317, n_340, n_375, n_708, n_105, n_187, n_667, n_1, n_154, n_682, n_182, n_196, n_326, n_327, n_89, n_50, n_723, n_144, n_170, n_270, n_346, n_383, n_113, n_561, n_117, n_417, n_471, n_265, n_504, n_158, n_259, n_276, n_339, n_470, n_210, n_348, n_220, n_674, n_91, n_481, n_287, n_54, n_243, n_19, n_497, n_671, n_228, n_711, n_147, n_552, n_251, n_384, n_632, n_373, n_458, n_244, n_73, n_343, n_310, n_714, n_703, n_426, n_323, n_469, n_598, n_143, n_106, n_386, n_549, n_8, n_224, n_183, n_533, n_508, n_67, n_453, n_591, n_655, n_333, n_110, n_306, n_400, n_47, n_550, n_736, n_169, n_10, n_673, n_21, n_732, n_242, n_278, n_316, n_16, n_404, n_60, n_557, n_641, n_7, n_109, n_127, n_121, n_527, n_590, n_465, n_48, n_325, n_57, n_301, n_496, n_617, n_434, n_296, n_690, n_120, n_168, n_526, n_155, n_315, n_441, n_604, n_13, n_637, n_122, n_523, n_116, n_694, n_614, n_370, n_431, n_719, n_574, n_0, n_289, n_716, n_12, n_515, n_642, n_150, n_286, n_321, n_133, n_569, n_600, n_51, n_215, n_279, n_49, n_374, n_235, n_464, n_538, n_669, n_22, n_136, n_261, n_521, n_665, n_459, n_30, n_518, n_367, n_221, n_654, n_656, n_724, n_437, n_731, n_602, n_355, n_474, n_594, n_636, n_710, n_720, n_407, n_102, n_490, n_568, n_52, n_448, n_646, n_595, n_99, n_466, n_269, n_156, n_570, n_126, n_623, n_585, n_715, n_530, n_356, n_25, n_104, n_45, n_420, n_483, n_543, n_580, n_141, n_487, n_222, n_660, n_186, n_524, n_349, n_454, n_295, n_730, n_331, n_576, n_230, n_96, n_185, n_388, n_625, n_619, n_536, n_611, n_352, n_290, n_558, n_666, n_174, n_467, n_427, n_607, n_157, n_219, n_246, n_31, n_442, n_146, n_207, n_438, n_689, n_167, n_676, n_128, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_358, n_205, n_618, n_488, n_139, n_514, n_705, n_429, n_560, n_275, n_541, n_98, n_129, n_613, n_659, n_267, n_662, n_635, n_245, n_589, n_571, n_229, n_209, n_472, n_648, n_347, n_473, n_445, n_629, n_335, n_413, n_82, n_263, n_27, n_573, n_353, n_359, n_299, n_87, n_262, n_433, n_75, n_439, n_704, n_643, n_137, n_679, n_338, n_173, n_696, n_477, n_640, n_363, n_402, n_725, n_180, n_369, n_596, n_201, n_699, n_14, n_351, n_368, n_456, n_257, n_77, n_718, n_44, n_672, n_722, n_401, n_553, n_554, n_66, n_735, n_305, n_713, n_307, n_192, n_140, n_484, n_566, n_480, n_416, n_581, n_651, n_365, n_721, n_4, n_6, n_605, n_539, n_100, n_179, n_354, n_206, n_392, n_630, n_516, n_548, n_567, n_329, n_447, n_26, n_188, n_200, n_444, n_506, n_562, n_564, n_546, n_199, n_592, n_495, n_410, n_308, n_675, n_463, n_624, n_706, n_411, n_135, n_520, n_684, n_658, n_512, n_615, n_685, n_283, n_366, n_397, n_111, n_692, n_36, n_627, n_18, n_709, n_322, n_53, n_227, n_499, n_115, n_11, n_248, n_92, n_702, n_451, n_712, n_101, n_190, n_138, n_650, n_409, n_582, n_653, n_214, n_238, n_579, n_332, n_517, n_211, n_218, n_314, n_691, n_563, n_132, n_277, n_555, n_337, n_522, n_700, n_479, n_534, n_225, n_360, n_272, n_511, n_23, n_734, n_468, n_223, n_381, n_525, n_535, n_382, n_502, n_681, n_633, n_532, n_726, n_95, n_405, n_415, n_597, n_285, n_288, n_247, n_320, n_379, n_551, n_55, n_612, n_291, n_318, n_63, n_161, n_237, n_29, n_203, n_268, n_440, n_148, n_2, n_342, n_233, n_385, n_414, n_430, n_118, n_729, n_603, n_378, n_486, n_422, n_164, n_38, n_198, n_264, n_616, n_217, n_324, n_391, n_537, n_728, n_78, n_670, n_20, n_69, n_390, n_544, n_39, n_178, n_509, n_695, n_639, n_303, n_362, n_717, n_93, n_505, n_162, n_482, n_240, n_282, n_61, n_680, n_501, n_668, n_266, n_42, n_294, n_112, n_485, n_46, n_284, n_80, n_172, n_250, n_493, n_460, n_609, n_476, n_461, n_575, n_313, n_519, n_345, n_408, n_119, n_361, n_455, n_419, n_72, n_319, n_195, n_513, n_212, n_588, n_693, n_311, n_661, n_406, n_606, n_737, n_97, n_197, n_528, n_181, n_131, n_123, n_631, n_683, n_260, n_620, n_462, n_302, n_450, n_443, n_686, n_572, n_644, n_577, n_344, n_393, n_436, n_428, n_491, n_297, n_435, n_628, n_41, n_252, n_396, n_697, n_83, n_32, n_107, n_149, n_489, n_677, n_399, n_254, n_213, n_424, n_565, n_701, n_271, n_241, n_68, n_503, n_292, n_394, n_79, n_81, n_35, n_364, n_687, n_159, n_202, n_231, n_298, n_587, n_160, n_657, n_184, n_56, n_492, n_649, n_232, n_380, n_281, n_559, n_425, n_3977);

input n_151;
input n_85;
input n_599;
input n_507;
input n_540;
input n_395;
input n_84;
input n_64;
input n_171;
input n_103;
input n_529;
input n_389;
input n_204;
input n_626;
input n_274;
input n_387;
input n_688;
input n_130;
input n_177;
input n_707;
input n_76;
input n_273;
input n_309;
input n_330;
input n_9;
input n_328;
input n_293;
input n_341;
input n_372;
input n_124;
input n_37;
input n_256;
input n_418;
input n_193;
input n_510;
input n_446;
input n_108;
input n_350;
input n_601;
input n_621;
input n_610;
input n_165;
input n_452;
input n_86;
input n_70;
input n_664;
input n_255;
input n_175;
input n_586;
input n_638;
input n_398;
input n_59;
input n_28;
input n_125;
input n_304;
input n_191;
input n_593;
input n_5;
input n_62;
input n_71;
input n_153;
input n_545;
input n_583;
input n_678;
input n_663;
input n_194;
input n_249;
input n_334;
input n_634;
input n_733;
input n_312;
input n_622;
input n_578;
input n_478;
input n_239;
input n_94;
input n_134;
input n_432;
input n_371;
input n_403;
input n_423;
input n_608;
input n_357;
input n_88;
input n_412;
input n_457;
input n_494;
input n_142;
input n_226;
input n_336;
input n_258;
input n_40;
input n_90;
input n_17;
input n_74;
input n_449;
input n_547;
input n_176;
input n_727;
input n_58;
input n_43;
input n_216;
input n_33;
input n_652;
input n_421;
input n_738;
input n_475;
input n_166;
input n_163;
input n_645;
input n_500;
input n_542;
input n_114;
input n_236;
input n_34;
input n_376;
input n_377;
input n_584;
input n_531;
input n_647;
input n_15;
input n_556;
input n_24;
input n_189;
input n_498;
input n_698;
input n_280;
input n_317;
input n_340;
input n_375;
input n_708;
input n_105;
input n_187;
input n_667;
input n_1;
input n_154;
input n_682;
input n_182;
input n_196;
input n_326;
input n_327;
input n_89;
input n_50;
input n_723;
input n_144;
input n_170;
input n_270;
input n_346;
input n_383;
input n_113;
input n_561;
input n_117;
input n_417;
input n_471;
input n_265;
input n_504;
input n_158;
input n_259;
input n_276;
input n_339;
input n_470;
input n_210;
input n_348;
input n_220;
input n_674;
input n_91;
input n_481;
input n_287;
input n_54;
input n_243;
input n_19;
input n_497;
input n_671;
input n_228;
input n_711;
input n_147;
input n_552;
input n_251;
input n_384;
input n_632;
input n_373;
input n_458;
input n_244;
input n_73;
input n_343;
input n_310;
input n_714;
input n_703;
input n_426;
input n_323;
input n_469;
input n_598;
input n_143;
input n_106;
input n_386;
input n_549;
input n_8;
input n_224;
input n_183;
input n_533;
input n_508;
input n_67;
input n_453;
input n_591;
input n_655;
input n_333;
input n_110;
input n_306;
input n_400;
input n_47;
input n_550;
input n_736;
input n_169;
input n_10;
input n_673;
input n_21;
input n_732;
input n_242;
input n_278;
input n_316;
input n_16;
input n_404;
input n_60;
input n_557;
input n_641;
input n_7;
input n_109;
input n_127;
input n_121;
input n_527;
input n_590;
input n_465;
input n_48;
input n_325;
input n_57;
input n_301;
input n_496;
input n_617;
input n_434;
input n_296;
input n_690;
input n_120;
input n_168;
input n_526;
input n_155;
input n_315;
input n_441;
input n_604;
input n_13;
input n_637;
input n_122;
input n_523;
input n_116;
input n_694;
input n_614;
input n_370;
input n_431;
input n_719;
input n_574;
input n_0;
input n_289;
input n_716;
input n_12;
input n_515;
input n_642;
input n_150;
input n_286;
input n_321;
input n_133;
input n_569;
input n_600;
input n_51;
input n_215;
input n_279;
input n_49;
input n_374;
input n_235;
input n_464;
input n_538;
input n_669;
input n_22;
input n_136;
input n_261;
input n_521;
input n_665;
input n_459;
input n_30;
input n_518;
input n_367;
input n_221;
input n_654;
input n_656;
input n_724;
input n_437;
input n_731;
input n_602;
input n_355;
input n_474;
input n_594;
input n_636;
input n_710;
input n_720;
input n_407;
input n_102;
input n_490;
input n_568;
input n_52;
input n_448;
input n_646;
input n_595;
input n_99;
input n_466;
input n_269;
input n_156;
input n_570;
input n_126;
input n_623;
input n_585;
input n_715;
input n_530;
input n_356;
input n_25;
input n_104;
input n_45;
input n_420;
input n_483;
input n_543;
input n_580;
input n_141;
input n_487;
input n_222;
input n_660;
input n_186;
input n_524;
input n_349;
input n_454;
input n_295;
input n_730;
input n_331;
input n_576;
input n_230;
input n_96;
input n_185;
input n_388;
input n_625;
input n_619;
input n_536;
input n_611;
input n_352;
input n_290;
input n_558;
input n_666;
input n_174;
input n_467;
input n_427;
input n_607;
input n_157;
input n_219;
input n_246;
input n_31;
input n_442;
input n_146;
input n_207;
input n_438;
input n_689;
input n_167;
input n_676;
input n_128;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_358;
input n_205;
input n_618;
input n_488;
input n_139;
input n_514;
input n_705;
input n_429;
input n_560;
input n_275;
input n_541;
input n_98;
input n_129;
input n_613;
input n_659;
input n_267;
input n_662;
input n_635;
input n_245;
input n_589;
input n_571;
input n_229;
input n_209;
input n_472;
input n_648;
input n_347;
input n_473;
input n_445;
input n_629;
input n_335;
input n_413;
input n_82;
input n_263;
input n_27;
input n_573;
input n_353;
input n_359;
input n_299;
input n_87;
input n_262;
input n_433;
input n_75;
input n_439;
input n_704;
input n_643;
input n_137;
input n_679;
input n_338;
input n_173;
input n_696;
input n_477;
input n_640;
input n_363;
input n_402;
input n_725;
input n_180;
input n_369;
input n_596;
input n_201;
input n_699;
input n_14;
input n_351;
input n_368;
input n_456;
input n_257;
input n_77;
input n_718;
input n_44;
input n_672;
input n_722;
input n_401;
input n_553;
input n_554;
input n_66;
input n_735;
input n_305;
input n_713;
input n_307;
input n_192;
input n_140;
input n_484;
input n_566;
input n_480;
input n_416;
input n_581;
input n_651;
input n_365;
input n_721;
input n_4;
input n_6;
input n_605;
input n_539;
input n_100;
input n_179;
input n_354;
input n_206;
input n_392;
input n_630;
input n_516;
input n_548;
input n_567;
input n_329;
input n_447;
input n_26;
input n_188;
input n_200;
input n_444;
input n_506;
input n_562;
input n_564;
input n_546;
input n_199;
input n_592;
input n_495;
input n_410;
input n_308;
input n_675;
input n_463;
input n_624;
input n_706;
input n_411;
input n_135;
input n_520;
input n_684;
input n_658;
input n_512;
input n_615;
input n_685;
input n_283;
input n_366;
input n_397;
input n_111;
input n_692;
input n_36;
input n_627;
input n_18;
input n_709;
input n_322;
input n_53;
input n_227;
input n_499;
input n_115;
input n_11;
input n_248;
input n_92;
input n_702;
input n_451;
input n_712;
input n_101;
input n_190;
input n_138;
input n_650;
input n_409;
input n_582;
input n_653;
input n_214;
input n_238;
input n_579;
input n_332;
input n_517;
input n_211;
input n_218;
input n_314;
input n_691;
input n_563;
input n_132;
input n_277;
input n_555;
input n_337;
input n_522;
input n_700;
input n_479;
input n_534;
input n_225;
input n_360;
input n_272;
input n_511;
input n_23;
input n_734;
input n_468;
input n_223;
input n_381;
input n_525;
input n_535;
input n_382;
input n_502;
input n_681;
input n_633;
input n_532;
input n_726;
input n_95;
input n_405;
input n_415;
input n_597;
input n_285;
input n_288;
input n_247;
input n_320;
input n_379;
input n_551;
input n_55;
input n_612;
input n_291;
input n_318;
input n_63;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_440;
input n_148;
input n_2;
input n_342;
input n_233;
input n_385;
input n_414;
input n_430;
input n_118;
input n_729;
input n_603;
input n_378;
input n_486;
input n_422;
input n_164;
input n_38;
input n_198;
input n_264;
input n_616;
input n_217;
input n_324;
input n_391;
input n_537;
input n_728;
input n_78;
input n_670;
input n_20;
input n_69;
input n_390;
input n_544;
input n_39;
input n_178;
input n_509;
input n_695;
input n_639;
input n_303;
input n_362;
input n_717;
input n_93;
input n_505;
input n_162;
input n_482;
input n_240;
input n_282;
input n_61;
input n_680;
input n_501;
input n_668;
input n_266;
input n_42;
input n_294;
input n_112;
input n_485;
input n_46;
input n_284;
input n_80;
input n_172;
input n_250;
input n_493;
input n_460;
input n_609;
input n_476;
input n_461;
input n_575;
input n_313;
input n_519;
input n_345;
input n_408;
input n_119;
input n_361;
input n_455;
input n_419;
input n_72;
input n_319;
input n_195;
input n_513;
input n_212;
input n_588;
input n_693;
input n_311;
input n_661;
input n_406;
input n_606;
input n_737;
input n_97;
input n_197;
input n_528;
input n_181;
input n_131;
input n_123;
input n_631;
input n_683;
input n_260;
input n_620;
input n_462;
input n_302;
input n_450;
input n_443;
input n_686;
input n_572;
input n_644;
input n_577;
input n_344;
input n_393;
input n_436;
input n_428;
input n_491;
input n_297;
input n_435;
input n_628;
input n_41;
input n_252;
input n_396;
input n_697;
input n_83;
input n_32;
input n_107;
input n_149;
input n_489;
input n_677;
input n_399;
input n_254;
input n_213;
input n_424;
input n_565;
input n_701;
input n_271;
input n_241;
input n_68;
input n_503;
input n_292;
input n_394;
input n_79;
input n_81;
input n_35;
input n_364;
input n_687;
input n_159;
input n_202;
input n_231;
input n_298;
input n_587;
input n_160;
input n_657;
input n_184;
input n_56;
input n_492;
input n_649;
input n_232;
input n_380;
input n_281;
input n_559;
input n_425;

output n_3977;

wire n_1084;
wire n_2594;
wire n_1474;
wire n_1295;
wire n_1983;
wire n_2804;
wire n_3150;
wire n_992;
wire n_1582;
wire n_2201;
wire n_3853;
wire n_2512;
wire n_766;
wire n_3590;
wire n_2960;
wire n_2175;
wire n_2071;
wire n_2796;
wire n_1110;
wire n_3610;
wire n_2607;
wire n_1382;
wire n_3548;
wire n_3911;
wire n_3144;
wire n_2569;
wire n_2949;
wire n_1998;
wire n_2840;
wire n_1596;
wire n_926;
wire n_3319;
wire n_1079;
wire n_3077;
wire n_2835;
wire n_3915;
wire n_1100;
wire n_3559;
wire n_845;
wire n_2177;
wire n_1930;
wire n_2123;
wire n_1234;
wire n_3019;
wire n_2047;
wire n_1594;
wire n_1944;
wire n_2235;
wire n_1802;
wire n_2498;
wire n_3817;
wire n_773;
wire n_3755;
wire n_2038;
wire n_2504;
wire n_1469;
wire n_3812;
wire n_821;
wire n_2017;
wire n_873;
wire n_1227;
wire n_962;
wire n_1080;
wire n_862;
wire n_909;
wire n_2290;
wire n_3750;
wire n_3838;
wire n_957;
wire n_3272;
wire n_3255;
wire n_3674;
wire n_1652;
wire n_969;
wire n_1859;
wire n_1954;
wire n_2183;
wire n_2074;
wire n_2897;
wire n_1883;
wire n_1125;
wire n_2687;
wire n_3456;
wire n_2037;
wire n_1226;
wire n_1034;
wire n_2383;
wire n_3132;
wire n_1765;
wire n_872;
wire n_2392;
wire n_1873;
wire n_1619;
wire n_1666;
wire n_2682;
wire n_2640;
wire n_3605;
wire n_930;
wire n_1044;
wire n_3280;
wire n_3105;
wire n_3146;
wire n_1492;
wire n_1134;
wire n_1478;
wire n_1684;
wire n_1796;
wire n_3569;
wire n_1614;
wire n_2374;
wire n_3334;
wire n_3819;
wire n_2598;
wire n_1722;
wire n_3931;
wire n_911;
wire n_2023;
wire n_781;
wire n_2720;
wire n_3870;
wire n_802;
wire n_3340;
wire n_2322;
wire n_1233;
wire n_2335;
wire n_3025;
wire n_3411;
wire n_2955;
wire n_3458;
wire n_3653;
wire n_3519;
wire n_2276;
wire n_1045;
wire n_3235;
wire n_2989;
wire n_1856;
wire n_2230;
wire n_963;
wire n_1782;
wire n_2889;
wire n_3843;
wire n_2139;
wire n_2847;
wire n_3693;
wire n_3033;
wire n_1308;
wire n_1138;
wire n_2943;
wire n_1096;
wire n_2151;
wire n_2391;
wire n_1391;
wire n_3338;
wire n_3168;
wire n_884;
wire n_2396;
wire n_3440;
wire n_3135;
wire n_3904;
wire n_850;
wire n_3175;
wire n_3729;
wire n_3484;
wire n_1971;
wire n_2485;
wire n_2479;
wire n_3570;
wire n_879;
wire n_2179;
wire n_1957;
wire n_2188;
wire n_1144;
wire n_2360;
wire n_2359;
wire n_2506;
wire n_1392;
wire n_2158;
wire n_1268;
wire n_2571;
wire n_3187;
wire n_739;
wire n_3830;
wire n_3598;
wire n_2724;
wire n_3086;
wire n_2475;
wire n_853;
wire n_3721;
wire n_948;
wire n_2799;
wire n_1752;
wire n_1829;
wire n_1338;
wire n_3726;
wire n_1730;
wire n_1307;
wire n_875;
wire n_1327;
wire n_2644;
wire n_876;
wire n_3211;
wire n_1840;
wire n_2837;
wire n_3479;
wire n_3751;
wire n_989;
wire n_3262;
wire n_3407;
wire n_3804;
wire n_1908;
wire n_3315;
wire n_3537;
wire n_1668;
wire n_2343;
wire n_2605;
wire n_2887;
wire n_1641;
wire n_829;
wire n_2565;
wire n_825;
wire n_1480;
wire n_1463;
wire n_1823;
wire n_3251;
wire n_1681;
wire n_2921;
wire n_3724;
wire n_939;
wire n_1636;
wire n_1687;
wire n_3192;
wire n_3533;
wire n_3753;
wire n_3896;
wire n_2192;
wire n_1766;
wire n_3184;
wire n_3566;
wire n_3469;
wire n_3170;
wire n_1922;
wire n_3890;
wire n_2032;
wire n_2820;
wire n_3323;
wire n_1937;
wire n_2311;
wire n_3392;
wire n_3347;
wire n_893;
wire n_3242;
wire n_3395;
wire n_3839;
wire n_1654;
wire n_3577;
wire n_2995;
wire n_3330;
wire n_1258;
wire n_1344;
wire n_2208;
wire n_2198;
wire n_1929;
wire n_2707;
wire n_3472;
wire n_3509;
wire n_1749;
wire n_1680;
wire n_835;
wire n_1981;
wire n_1195;
wire n_2918;
wire n_3353;
wire n_3976;
wire n_824;
wire n_1945;
wire n_2638;
wire n_3939;
wire n_787;
wire n_2860;
wire n_2448;
wire n_3631;
wire n_2015;
wire n_3807;
wire n_2537;
wire n_1130;
wire n_2643;
wire n_1228;
wire n_2998;
wire n_2336;
wire n_3845;
wire n_3641;
wire n_2163;
wire n_3969;
wire n_1081;
wire n_2354;
wire n_3639;
wire n_3856;
wire n_1155;
wire n_1292;
wire n_2432;
wire n_2873;
wire n_3043;
wire n_1576;
wire n_1664;
wire n_2273;
wire n_3298;
wire n_1427;
wire n_852;
wire n_1133;
wire n_3049;
wire n_2421;
wire n_1926;
wire n_3208;
wire n_904;
wire n_2363;
wire n_2814;
wire n_3237;
wire n_3264;
wire n_3204;
wire n_2003;
wire n_1970;
wire n_3671;
wire n_3946;
wire n_3727;
wire n_2621;
wire n_3620;
wire n_3747;
wire n_1778;
wire n_2558;
wire n_2953;
wire n_2922;
wire n_2347;
wire n_3884;
wire n_3881;
wire n_3507;
wire n_3949;
wire n_3103;
wire n_2839;
wire n_3926;
wire n_1030;
wire n_1698;
wire n_3688;
wire n_1094;
wire n_2462;
wire n_3770;
wire n_1496;
wire n_1910;
wire n_2333;
wire n_1663;
wire n_2436;
wire n_1214;
wire n_1274;
wire n_2705;
wire n_2527;
wire n_1606;
wire n_769;
wire n_1595;
wire n_2164;
wire n_3711;
wire n_1509;
wire n_1618;
wire n_1648;
wire n_2944;
wire n_1886;
wire n_2269;
wire n_3748;
wire n_857;
wire n_765;
wire n_1070;
wire n_1841;
wire n_2472;
wire n_777;
wire n_2846;
wire n_2685;
wire n_3668;
wire n_3699;
wire n_1955;
wire n_3197;
wire n_917;
wire n_2413;
wire n_2249;
wire n_2362;
wire n_968;
wire n_3022;
wire n_3148;
wire n_2822;
wire n_3766;
wire n_1253;
wire n_3707;
wire n_1306;
wire n_1484;
wire n_2686;
wire n_1493;
wire n_2597;
wire n_3973;
wire n_1313;
wire n_2774;
wire n_3151;
wire n_2090;
wire n_2260;
wire n_3722;
wire n_3125;
wire n_2812;
wire n_3802;
wire n_3681;
wire n_2753;
wire n_3603;
wire n_1638;
wire n_2215;
wire n_1449;
wire n_1071;
wire n_1723;
wire n_1960;
wire n_2663;
wire n_3882;
wire n_793;
wire n_3129;
wire n_937;
wire n_2595;
wire n_2116;
wire n_3714;
wire n_3592;
wire n_1645;
wire n_3186;
wire n_973;
wire n_1038;
wire n_2280;
wire n_1943;
wire n_3541;
wire n_1863;
wire n_2844;
wire n_1269;
wire n_2393;
wire n_2773;
wire n_3565;
wire n_3883;
wire n_3030;
wire n_2906;
wire n_3097;
wire n_3943;
wire n_3809;
wire n_979;
wire n_1309;
wire n_1999;
wire n_3810;
wire n_3718;
wire n_1316;
wire n_1562;
wire n_3917;
wire n_1215;
wire n_3679;
wire n_3579;
wire n_2777;
wire n_2480;
wire n_3769;
wire n_1445;
wire n_2283;
wire n_2806;
wire n_3910;
wire n_2813;
wire n_2147;
wire n_1716;
wire n_1466;
wire n_1412;
wire n_3210;
wire n_3667;
wire n_3221;
wire n_1672;
wire n_1007;
wire n_2253;
wire n_1276;
wire n_3822;
wire n_1637;
wire n_3310;
wire n_841;
wire n_2900;
wire n_3858;
wire n_772;
wire n_810;
wire n_1401;
wire n_3764;
wire n_3795;
wire n_1817;
wire n_2951;
wire n_2145;
wire n_2122;
wire n_1588;
wire n_3765;
wire n_2216;
wire n_1301;
wire n_2579;
wire n_2876;
wire n_2242;
wire n_869;
wire n_1620;
wire n_1561;
wire n_3301;
wire n_2370;
wire n_2025;
wire n_1078;
wire n_2247;
wire n_3451;
wire n_1219;
wire n_1865;
wire n_3177;
wire n_3518;
wire n_3399;
wire n_1252;
wire n_2022;
wire n_2730;
wire n_3967;
wire n_1170;
wire n_1927;
wire n_2373;
wire n_1869;
wire n_3842;
wire n_1853;
wire n_2275;
wire n_2980;
wire n_2189;
wire n_2482;
wire n_745;
wire n_3799;
wire n_2767;
wire n_3676;
wire n_2899;
wire n_2826;
wire n_2112;
wire n_1753;
wire n_3351;
wire n_1322;
wire n_2008;
wire n_1305;
wire n_2088;
wire n_795;
wire n_1248;
wire n_2762;
wire n_2171;
wire n_3307;
wire n_762;
wire n_1388;
wire n_2859;
wire n_800;
wire n_2564;
wire n_3780;
wire n_3023;
wire n_784;
wire n_1653;
wire n_1375;
wire n_3224;
wire n_1356;
wire n_894;
wire n_1118;
wire n_2591;
wire n_1881;
wire n_3762;
wire n_3965;
wire n_1969;
wire n_3798;
wire n_1296;
wire n_3060;
wire n_971;
wire n_1326;
wire n_1350;
wire n_3627;
wire n_906;
wire n_2957;
wire n_2586;
wire n_3958;
wire n_1093;
wire n_1764;
wire n_2412;
wire n_2783;
wire n_978;
wire n_3777;
wire n_899;
wire n_1799;
wire n_3293;
wire n_1019;
wire n_902;
wire n_1689;
wire n_1250;
wire n_2550;
wire n_1190;
wire n_1304;
wire n_744;
wire n_2541;
wire n_1506;
wire n_881;
wire n_2987;
wire n_3259;
wire n_1702;
wire n_3916;
wire n_3381;
wire n_3630;
wire n_1558;
wire n_2750;
wire n_1650;
wire n_1520;
wire n_1073;
wire n_1453;
wire n_3961;
wire n_1108;
wire n_2722;
wire n_2509;
wire n_2727;
wire n_3618;
wire n_1794;
wire n_1423;
wire n_3836;
wire n_1239;
wire n_2399;
wire n_1370;
wire n_2719;
wire n_1209;
wire n_1708;
wire n_2213;
wire n_3038;
wire n_3732;
wire n_3779;
wire n_3521;
wire n_3203;
wire n_3295;
wire n_3923;
wire n_2723;
wire n_1616;
wire n_3199;
wire n_3808;
wire n_3093;
wire n_1569;
wire n_2664;
wire n_1434;
wire n_3716;
wire n_1649;
wire n_2389;
wire n_3450;
wire n_1936;
wire n_2114;
wire n_1717;
wire n_3567;
wire n_2107;
wire n_1609;
wire n_2257;
wire n_3435;
wire n_3530;
wire n_1613;
wire n_820;
wire n_805;
wire n_1988;
wire n_1132;
wire n_892;
wire n_1467;
wire n_1803;
wire n_2401;
wire n_1787;
wire n_2782;
wire n_2511;
wire n_3217;
wire n_1281;
wire n_3094;
wire n_3874;
wire n_1447;
wire n_2166;
wire n_2451;
wire n_2150;
wire n_1549;
wire n_2631;
wire n_1867;
wire n_1531;
wire n_2919;
wire n_3909;
wire n_3971;
wire n_1332;
wire n_2660;
wire n_2661;
wire n_2292;
wire n_3573;
wire n_3563;
wire n_3510;
wire n_3560;
wire n_2334;
wire n_1424;
wire n_3467;
wire n_2444;
wire n_2350;
wire n_1742;
wire n_2625;
wire n_3652;
wire n_1818;
wire n_870;
wire n_2199;
wire n_1709;
wire n_1610;
wire n_2219;
wire n_3847;
wire n_1298;
wire n_1844;
wire n_1387;
wire n_2649;
wire n_1040;
wire n_2203;
wire n_2693;
wire n_3194;
wire n_3607;
wire n_3371;
wire n_1159;
wire n_1368;
wire n_2281;
wire n_1154;
wire n_3202;
wire n_2539;
wire n_2431;
wire n_1701;
wire n_2084;
wire n_1243;
wire n_3572;
wire n_2387;
wire n_2646;
wire n_3375;
wire n_2397;
wire n_1121;
wire n_2746;
wire n_3241;
wire n_2256;
wire n_3317;
wire n_3800;
wire n_3887;
wire n_3963;
wire n_2445;
wire n_3461;
wire n_2729;
wire n_1571;
wire n_1980;
wire n_3951;
wire n_3355;
wire n_2529;
wire n_3583;
wire n_2019;
wire n_1407;
wire n_3282;
wire n_1235;
wire n_1821;
wire n_3832;
wire n_3508;
wire n_1003;
wire n_889;
wire n_3827;
wire n_2708;
wire n_3156;
wire n_3457;
wire n_2748;
wire n_816;
wire n_1058;
wire n_1835;
wire n_1862;
wire n_2224;
wire n_2697;
wire n_3531;
wire n_3415;
wire n_2470;
wire n_2355;
wire n_2890;
wire n_3698;
wire n_2731;
wire n_1543;
wire n_3466;
wire n_3386;
wire n_823;
wire n_2233;
wire n_2499;
wire n_3370;
wire n_1504;
wire n_3814;
wire n_1519;
wire n_1425;
wire n_1781;
wire n_3888;
wire n_2069;
wire n_2602;
wire n_1441;
wire n_2028;
wire n_3309;
wire n_3678;
wire n_1924;
wire n_2856;
wire n_1921;
wire n_3024;
wire n_1156;
wire n_2857;
wire n_1293;
wire n_1360;
wire n_749;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_3968;
wire n_819;
wire n_3950;
wire n_2070;
wire n_1042;
wire n_822;
wire n_1888;
wire n_3471;
wire n_743;
wire n_3117;
wire n_3320;
wire n_754;
wire n_1786;
wire n_2033;
wire n_3039;
wire n_3900;
wire n_1319;
wire n_1553;
wire n_3478;
wire n_3701;
wire n_3542;
wire n_1041;
wire n_2766;
wire n_3756;
wire n_2828;
wire n_3754;
wire n_1964;
wire n_1090;
wire n_3720;
wire n_3374;
wire n_1196;
wire n_3704;
wire n_1182;
wire n_1271;
wire n_3811;
wire n_2416;
wire n_3633;
wire n_2786;
wire n_1731;
wire n_1905;
wire n_2962;
wire n_1031;
wire n_3416;
wire n_2879;
wire n_2958;
wire n_3147;
wire n_3694;
wire n_2052;
wire n_3690;
wire n_981;
wire n_3628;
wire n_2425;
wire n_2800;
wire n_3514;
wire n_3091;
wire n_3006;
wire n_3348;
wire n_2118;
wire n_2259;
wire n_3859;
wire n_2162;
wire n_2236;
wire n_3455;
wire n_3957;
wire n_3660;
wire n_2377;
wire n_2718;
wire n_2577;
wire n_1591;
wire n_3426;
wire n_3165;
wire n_2289;
wire n_2288;
wire n_2841;
wire n_3075;
wire n_1671;
wire n_1795;
wire n_1409;
wire n_1015;
wire n_3448;
wire n_3788;
wire n_2744;
wire n_2101;
wire n_2795;
wire n_3524;
wire n_3634;
wire n_1377;
wire n_2473;
wire n_1583;
wire n_3520;
wire n_1521;
wire n_2632;
wire n_1152;
wire n_2456;
wire n_2924;
wire n_3054;
wire n_2264;
wire n_2076;
wire n_1036;
wire n_974;
wire n_2599;
wire n_1831;
wire n_3626;
wire n_3733;
wire n_864;
wire n_1987;
wire n_959;
wire n_1106;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_3171;
wire n_1733;
wire n_3365;
wire n_3684;
wire n_1634;
wire n_2853;
wire n_1932;
wire n_3775;
wire n_1452;
wire n_1552;
wire n_1318;
wire n_1508;
wire n_2217;
wire n_3741;
wire n_3854;
wire n_1217;
wire n_3594;
wire n_2866;
wire n_3970;
wire n_3153;
wire n_3291;
wire n_2655;
wire n_3487;
wire n_2454;
wire n_1715;
wire n_3966;
wire n_1189;
wire n_3300;
wire n_761;
wire n_748;
wire n_1713;
wire n_3621;
wire n_901;
wire n_1577;
wire n_2036;
wire n_1255;
wire n_2829;
wire n_2968;
wire n_2740;
wire n_3473;
wire n_1700;
wire n_2623;
wire n_2622;
wire n_3232;
wire n_2819;
wire n_1218;
wire n_2178;
wire n_1181;
wire n_3263;
wire n_3815;
wire n_1140;
wire n_1985;
wire n_1772;
wire n_2858;
wire n_3708;
wire n_1056;
wire n_2626;
wire n_1283;
wire n_3007;
wire n_3790;
wire n_1446;
wire n_2404;
wire n_1487;
wire n_3078;
wire n_2789;
wire n_2603;
wire n_840;
wire n_1203;
wire n_1421;
wire n_3640;
wire n_3218;
wire n_2821;
wire n_2424;
wire n_846;
wire n_1793;
wire n_1237;
wire n_2880;
wire n_2390;
wire n_2573;
wire n_2423;
wire n_859;
wire n_3849;
wire n_1109;
wire n_965;
wire n_2741;
wire n_2793;
wire n_3098;
wire n_3490;
wire n_3055;
wire n_1633;
wire n_3299;
wire n_2580;
wire n_3222;
wire n_1711;
wire n_3529;
wire n_3069;
wire n_3107;
wire n_3352;
wire n_3436;
wire n_1051;
wire n_1008;
wire n_2964;
wire n_3065;
wire n_2375;
wire n_1498;
wire n_2312;
wire n_2572;
wire n_2946;
wire n_1053;
wire n_1656;
wire n_1207;
wire n_1076;
wire n_1735;
wire n_2063;
wire n_1032;
wire n_936;
wire n_3082;
wire n_1884;
wire n_2176;
wire n_3813;
wire n_1825;
wire n_2805;
wire n_1589;
wire n_2717;
wire n_2204;
wire n_2863;
wire n_2575;
wire n_1210;
wire n_2319;
wire n_3757;
wire n_2877;
wire n_1933;
wire n_2522;
wire n_3357;
wire n_3855;
wire n_1996;
wire n_1510;
wire n_1201;
wire n_1842;
wire n_2852;
wire n_2132;
wire n_3964;
wire n_3110;
wire n_1246;
wire n_1677;
wire n_1236;
wire n_3364;
wire n_832;
wire n_2297;
wire n_3429;
wire n_3306;
wire n_3412;
wire n_3037;
wire n_3188;
wire n_2780;
wire n_3787;
wire n_1792;
wire n_1712;
wire n_3250;
wire n_1984;
wire n_1568;
wire n_2885;
wire n_1877;
wire n_3445;
wire n_1184;
wire n_1477;
wire n_2585;
wire n_2220;
wire n_2080;
wire n_1724;
wire n_2554;
wire n_3155;
wire n_2838;
wire n_1364;
wire n_3183;
wire n_1540;
wire n_1676;
wire n_1013;
wire n_3243;
wire n_2468;
wire n_929;
wire n_3248;
wire n_3214;
wire n_1136;
wire n_1890;
wire n_1075;
wire n_1249;
wire n_3128;
wire n_1918;
wire n_2606;
wire n_3642;
wire n_2549;
wire n_2461;
wire n_3468;
wire n_2006;
wire n_2440;
wire n_1229;
wire n_1440;
wire n_1490;
wire n_2152;
wire n_1179;
wire n_907;
wire n_1990;
wire n_3680;
wire n_1153;
wire n_3624;
wire n_1751;
wire n_2787;
wire n_3785;
wire n_2467;
wire n_2146;
wire n_2341;
wire n_3525;
wire n_1737;
wire n_3145;
wire n_2779;
wire n_1117;
wire n_1273;
wire n_3821;
wire n_2547;
wire n_2930;
wire n_2616;
wire n_1748;
wire n_2662;
wire n_1083;
wire n_3205;
wire n_3872;
wire n_1014;
wire n_3801;
wire n_2883;
wire n_938;
wire n_1178;
wire n_2935;
wire n_878;
wire n_2441;
wire n_3503;
wire n_2358;
wire n_2490;
wire n_3127;
wire n_3496;
wire n_2361;
wire n_1464;
wire n_1566;
wire n_3568;
wire n_944;
wire n_3312;
wire n_3003;
wire n_1848;
wire n_2062;
wire n_2277;
wire n_3841;
wire n_2650;
wire n_1982;
wire n_2252;
wire n_3932;
wire n_2888;
wire n_2339;
wire n_3614;
wire n_1334;
wire n_3879;
wire n_1963;
wire n_3394;
wire n_1695;
wire n_1418;
wire n_2999;
wire n_2402;
wire n_1137;
wire n_2910;
wire n_2552;
wire n_3331;
wire n_2590;
wire n_3119;
wire n_1977;
wire n_2294;
wire n_1200;
wire n_2295;
wire n_3345;
wire n_2530;
wire n_2379;
wire n_1120;
wire n_2300;
wire n_2792;
wire n_1602;
wire n_2965;
wire n_1776;
wire n_2372;
wire n_3341;
wire n_2382;
wire n_1852;
wire n_1522;
wire n_2523;
wire n_2557;
wire n_3544;
wire n_3868;
wire n_1279;
wire n_2505;
wire n_931;
wire n_3488;
wire n_827;
wire n_3554;
wire n_2481;
wire n_3692;
wire n_1064;
wire n_1408;
wire n_2832;
wire n_3913;
wire n_1028;
wire n_1264;
wire n_3535;
wire n_3730;
wire n_2808;
wire n_2287;
wire n_3597;
wire n_3396;
wire n_2954;
wire n_3526;
wire n_2102;
wire n_1935;
wire n_2046;
wire n_3367;
wire n_3492;
wire n_1146;
wire n_2785;
wire n_2751;
wire n_3558;
wire n_2142;
wire n_1548;
wire n_3703;
wire n_2977;
wire n_1682;
wire n_1608;
wire n_3776;
wire n_3599;
wire n_1009;
wire n_1260;
wire n_1896;
wire n_1704;
wire n_2160;
wire n_2699;
wire n_2234;
wire n_847;
wire n_2991;
wire n_1436;
wire n_3239;
wire n_2600;
wire n_1069;
wire n_1485;
wire n_2239;
wire n_1465;
wire n_3952;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_3826;
wire n_1232;
wire n_1979;
wire n_2328;
wire n_2715;
wire n_3781;
wire n_1345;
wire n_2434;
wire n_837;
wire n_1590;
wire n_2332;
wire n_2971;
wire n_954;
wire n_3578;
wire n_1628;
wire n_1773;
wire n_2133;
wire n_3553;
wire n_3072;
wire n_1545;
wire n_3249;
wire n_3580;
wire n_2369;
wire n_3470;
wire n_3584;
wire n_1471;
wire n_1738;
wire n_3441;
wire n_3797;
wire n_998;
wire n_1395;
wire n_1729;
wire n_1115;
wire n_2551;
wire n_3281;
wire n_801;
wire n_2823;
wire n_3274;
wire n_2094;
wire n_2613;
wire n_1479;
wire n_3505;
wire n_2306;
wire n_1046;
wire n_2419;
wire n_3397;
wire n_2934;
wire n_2807;
wire n_882;
wire n_942;
wire n_1627;
wire n_1431;
wire n_3956;
wire n_3880;
wire n_2525;
wire n_814;
wire n_3829;
wire n_1864;
wire n_943;
wire n_3087;
wire n_2568;
wire n_2629;
wire n_3587;
wire n_1086;
wire n_1523;
wire n_2197;
wire n_2010;
wire n_1756;
wire n_2097;
wire n_2733;
wire n_2241;
wire n_1470;
wire n_2098;
wire n_2109;
wire n_1761;
wire n_3796;
wire n_2648;
wire n_2458;
wire n_1836;
wire n_2398;
wire n_3401;
wire n_3032;
wire n_1593;
wire n_986;
wire n_1420;
wire n_2651;
wire n_1750;
wire n_1775;
wire n_2833;
wire n_1699;
wire n_3179;
wire n_927;
wire n_1563;
wire n_2905;
wire n_3460;
wire n_3954;
wire n_803;
wire n_2570;
wire n_3123;
wire n_1875;
wire n_3379;
wire n_1615;
wire n_2418;
wire n_2184;
wire n_1087;
wire n_3390;
wire n_3719;
wire n_757;
wire n_3948;
wire n_1400;
wire n_1539;
wire n_1599;
wire n_1806;
wire n_3070;
wire n_2842;
wire n_2711;
wire n_3477;
wire n_2635;
wire n_3646;
wire n_2469;
wire n_1575;
wire n_2209;
wire n_3074;
wire n_3897;
wire n_3020;
wire n_3142;
wire n_3975;
wire n_3164;
wire n_3475;
wire n_1448;
wire n_2077;
wire n_3136;
wire n_2520;
wire n_817;
wire n_2193;
wire n_3034;
wire n_2612;
wire n_2095;
wire n_3108;
wire n_2486;
wire n_2628;
wire n_2395;
wire n_951;
wire n_2521;
wire n_2908;
wire n_2053;
wire n_2752;
wire n_1580;
wire n_2124;
wire n_3974;
wire n_1574;
wire n_780;
wire n_2200;
wire n_1705;
wire n_3625;
wire n_2304;
wire n_1746;
wire n_1439;
wire n_2263;
wire n_2212;
wire n_2352;
wire n_2716;
wire n_3495;
wire n_863;
wire n_2185;
wire n_3169;
wire n_1832;
wire n_1128;
wire n_2476;
wire n_2376;
wire n_2979;
wire n_3398;
wire n_1266;
wire n_1300;
wire n_3759;
wire n_2781;
wire n_3419;
wire n_3629;
wire n_807;
wire n_741;
wire n_2460;
wire n_2170;
wire n_3600;
wire n_1785;
wire n_1870;
wire n_2484;
wire n_2721;
wire n_1405;
wire n_2884;
wire n_3383;
wire n_3167;
wire n_3687;
wire n_997;
wire n_2308;
wire n_3459;
wire n_3238;
wire n_2986;
wire n_3498;
wire n_1428;
wire n_2691;
wire n_2243;
wire n_2400;
wire n_3731;
wire n_3092;
wire n_3555;
wire n_2903;
wire n_891;
wire n_3659;
wire n_3254;
wire n_2507;
wire n_2759;
wire n_3434;
wire n_1528;
wire n_1495;
wire n_3131;
wire n_3682;
wire n_2654;
wire n_2463;
wire n_3840;
wire n_2975;
wire n_1357;
wire n_2503;
wire n_2478;
wire n_3178;
wire n_2794;
wire n_1512;
wire n_3672;
wire n_2496;
wire n_3378;
wire n_3481;
wire n_3885;
wire n_2974;
wire n_871;
wire n_2990;
wire n_2923;
wire n_1339;
wire n_1544;
wire n_1426;
wire n_2365;
wire n_3449;
wire n_3517;
wire n_3350;
wire n_2245;
wire n_1315;
wire n_1413;
wire n_2464;
wire n_811;
wire n_808;
wire n_3877;
wire n_945;
wire n_2925;
wire n_2270;
wire n_3260;
wire n_1706;
wire n_3936;
wire n_1560;
wire n_1592;
wire n_2776;
wire n_1461;
wire n_3166;
wire n_3953;
wire n_2695;
wire n_2630;
wire n_903;
wire n_1967;
wire n_2340;
wire n_3385;
wire n_2117;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_3834;
wire n_2488;
wire n_1378;
wire n_2042;
wire n_3656;
wire n_3257;
wire n_1048;
wire n_774;
wire n_2459;
wire n_3137;
wire n_3116;
wire n_1925;
wire n_2439;
wire n_3638;
wire n_2106;
wire n_1430;
wire n_2414;
wire n_1251;
wire n_3090;
wire n_1247;
wire n_3816;
wire n_2450;
wire n_836;
wire n_1475;
wire n_3337;
wire n_2465;
wire n_1263;
wire n_3316;
wire n_3925;
wire n_1185;
wire n_1683;
wire n_3575;
wire n_1122;
wire n_2765;
wire n_3387;
wire n_890;
wire n_874;
wire n_1505;
wire n_3010;
wire n_2941;
wire n_1163;
wire n_1514;
wire n_964;
wire n_2728;
wire n_3772;
wire n_2948;
wire n_916;
wire n_3428;
wire n_2298;
wire n_2771;
wire n_3219;
wire n_2936;
wire n_895;
wire n_3955;
wire n_3867;
wire n_1035;
wire n_2427;
wire n_2045;
wire n_2985;
wire n_1535;
wire n_3158;
wire n_3106;
wire n_751;
wire n_2190;
wire n_1127;
wire n_932;
wire n_3657;
wire n_1972;
wire n_3080;
wire n_2772;
wire n_2778;
wire n_947;
wire n_1004;
wire n_831;
wire n_3929;
wire n_778;
wire n_1898;
wire n_1254;
wire n_1148;
wire n_1667;
wire n_1845;
wire n_1104;
wire n_2205;
wire n_1011;
wire n_2684;
wire n_2875;
wire n_2524;
wire n_3284;
wire n_1437;
wire n_3835;
wire n_3723;
wire n_2747;
wire n_3389;
wire n_1707;
wire n_1941;
wire n_3902;
wire n_3927;
wire n_2422;
wire n_2064;
wire n_3088;
wire n_1679;
wire n_2342;
wire n_2755;
wire n_2301;
wire n_1497;
wire n_2002;
wire n_2055;
wire n_3564;
wire n_2385;
wire n_3095;
wire n_3864;
wire n_3026;
wire n_2545;
wire n_1578;
wire n_3294;
wire n_2050;
wire n_1143;
wire n_1783;
wire n_2712;
wire n_3695;
wire n_3279;
wire n_2584;
wire n_972;
wire n_1815;
wire n_2500;
wire n_3344;
wire n_1917;
wire n_1444;
wire n_920;
wire n_2442;
wire n_1067;
wire n_3328;
wire n_2763;
wire n_2788;
wire n_994;
wire n_2000;
wire n_2089;
wire n_1857;
wire n_2761;
wire n_1920;
wire n_2696;
wire n_3252;
wire n_887;
wire n_1162;
wire n_1997;
wire n_2578;
wire n_2745;
wire n_1894;
wire n_2110;
wire n_2904;
wire n_3064;
wire n_2896;
wire n_2997;
wire n_3314;
wire n_1349;
wire n_1331;
wire n_1223;
wire n_961;
wire n_991;
wire n_2127;
wire n_3735;
wire n_1323;
wire n_3891;
wire n_1739;
wire n_3130;
wire n_1777;
wire n_3028;
wire n_3228;
wire n_3710;
wire n_1353;
wire n_3409;
wire n_2386;
wire n_3706;
wire n_3324;
wire n_1429;
wire n_3073;
wire n_2029;
wire n_3209;
wire n_2026;
wire n_1546;
wire n_3588;
wire n_3420;
wire n_1432;
wire n_2103;
wire n_3322;
wire n_1950;
wire n_1320;
wire n_996;
wire n_3632;
wire n_3914;
wire n_915;
wire n_2238;
wire n_3289;
wire n_1174;
wire n_1874;
wire n_1834;
wire n_3372;
wire n_3499;
wire n_3552;
wire n_2862;
wire n_3850;
wire n_3100;
wire n_3405;
wire n_1727;
wire n_3377;
wire n_1286;
wire n_1657;
wire n_1741;
wire n_1294;
wire n_1601;
wire n_900;
wire n_3784;
wire n_3414;
wire n_1351;
wire n_2933;
wire n_2138;
wire n_1380;
wire n_1367;
wire n_3336;
wire n_3240;
wire n_3828;
wire n_1291;
wire n_2895;
wire n_3763;
wire n_1914;
wire n_3833;
wire n_1458;
wire n_1694;
wire n_1460;
wire n_2041;
wire n_3201;
wire n_2271;
wire n_2356;
wire n_3339;
wire n_1830;
wire n_2261;
wire n_3016;
wire n_1629;
wire n_3476;
wire n_3673;
wire n_2994;
wire n_2011;
wire n_2620;
wire n_1826;
wire n_1855;
wire n_1662;
wire n_2187;
wire n_2105;
wire n_3556;
wire n_1340;
wire n_2694;
wire n_3443;
wire n_2562;
wire n_2642;
wire n_3029;
wire n_3269;
wire n_3609;
wire n_3447;
wire n_3771;
wire n_2647;
wire n_1626;
wire n_2223;
wire n_1660;
wire n_1850;
wire n_1643;
wire n_1670;
wire n_1789;
wire n_2415;
wire n_3876;
wire n_3152;
wire n_3154;
wire n_2344;
wire n_3589;
wire n_2317;
wire n_2556;
wire n_1112;
wire n_1267;
wire n_2384;
wire n_2683;
wire n_1384;
wire n_1376;
wire n_1537;
wire n_1858;
wire n_3432;
wire n_3523;
wire n_2815;
wire n_1816;
wire n_2446;
wire n_3388;
wire n_1612;
wire n_2318;
wire n_1172;
wire n_2659;
wire n_3616;
wire n_3908;
wire n_1099;
wire n_2141;
wire n_3113;
wire n_3696;
wire n_2902;
wire n_2909;
wire n_1422;
wire n_1527;
wire n_3174;
wire n_3960;
wire n_3608;
wire n_3190;
wire n_1524;
wire n_1055;
wire n_3878;
wire n_798;
wire n_2849;
wire n_2947;
wire n_1754;
wire n_3048;
wire n_3686;
wire n_1177;
wire n_1025;
wire n_1991;
wire n_2566;
wire n_2679;
wire n_3292;
wire n_2210;
wire n_1517;
wire n_3940;
wire n_2502;
wire n_1225;
wire n_1962;
wire n_2346;
wire n_982;
wire n_3670;
wire n_1624;
wire n_785;
wire n_1952;
wire n_2180;
wire n_3002;
wire n_3376;
wire n_2087;
wire n_2920;
wire n_3290;
wire n_1598;
wire n_2952;
wire n_2617;
wire n_3585;
wire n_977;
wire n_2878;
wire n_1895;
wire n_2250;
wire n_1491;
wire n_1860;
wire n_2831;
wire n_1810;
wire n_1763;
wire n_923;
wire n_3778;
wire n_3912;
wire n_3818;
wire n_1607;
wire n_2865;
wire n_2075;
wire n_3047;
wire n_1625;
wire n_2959;
wire n_2610;
wire n_2380;
wire n_2420;
wire n_3335;
wire n_3265;
wire n_2240;
wire n_933;
wire n_2221;
wire n_1774;
wire n_1797;
wire n_2516;
wire n_2120;
wire n_1037;
wire n_1899;
wire n_2031;
wire n_3669;
wire n_3427;
wire n_1289;
wire n_1348;
wire n_838;
wire n_2892;
wire n_1021;
wire n_746;
wire n_1557;
wire n_1188;
wire n_1567;
wire n_2007;
wire n_742;
wire n_1191;
wire n_2004;
wire n_3356;
wire n_3431;
wire n_3220;
wire n_2024;
wire n_3783;
wire n_2086;
wire n_1503;
wire n_3422;
wire n_1052;
wire n_789;
wire n_1942;
wire n_3666;
wire n_3141;
wire n_2309;
wire n_842;
wire n_2274;
wire n_2698;
wire n_767;
wire n_1617;
wire n_1839;
wire n_3899;
wire n_3930;
wire n_1587;
wire n_2330;
wire n_2555;
wire n_2639;
wire n_1259;
wire n_2108;
wire n_3099;
wire n_3712;
wire n_2535;
wire n_1001;
wire n_2945;
wire n_3057;
wire n_2143;
wire n_2410;
wire n_3760;
wire n_1396;
wire n_2916;
wire n_1224;
wire n_1923;
wire n_3206;
wire n_3736;
wire n_2196;
wire n_2739;
wire n_2611;
wire n_1538;
wire n_2528;
wire n_3773;
wire n_2548;
wire n_3216;
wire n_2709;
wire n_3061;
wire n_3717;
wire n_2633;
wire n_1017;
wire n_2244;
wire n_2604;
wire n_3424;
wire n_3745;
wire n_3462;
wire n_2351;
wire n_2437;
wire n_3664;
wire n_2049;
wire n_1456;
wire n_3245;
wire n_1889;
wire n_3907;
wire n_2113;
wire n_2665;
wire n_1124;
wire n_1690;
wire n_3063;
wire n_2688;
wire n_2881;
wire n_3862;
wire n_3302;
wire n_1673;
wire n_3361;
wire n_2018;
wire n_3134;
wire n_922;
wire n_2817;
wire n_1790;
wire n_993;
wire n_851;
wire n_3196;
wire n_2085;
wire n_3304;
wire n_2581;
wire n_1725;
wire n_2809;
wire n_2149;
wire n_2268;
wire n_2320;
wire n_2237;
wire n_1135;
wire n_2255;
wire n_2001;
wire n_1820;
wire n_3921;
wire n_1800;
wire n_3277;
wire n_3480;
wire n_2758;
wire n_3746;
wire n_1494;
wire n_1550;
wire n_3906;
wire n_2060;
wire n_1066;
wire n_2214;
wire n_3474;
wire n_1169;
wire n_1726;
wire n_1946;
wire n_3111;
wire n_1938;
wire n_830;
wire n_3452;
wire n_1241;
wire n_3645;
wire n_2589;
wire n_1072;
wire n_2194;
wire n_1231;
wire n_1173;
wire n_2736;
wire n_1208;
wire n_1604;
wire n_1639;
wire n_2735;
wire n_2845;
wire n_3506;
wire n_826;
wire n_1976;
wire n_2154;
wire n_2035;
wire n_1337;
wire n_2732;
wire n_3162;
wire n_2984;
wire n_1906;
wire n_3004;
wire n_3886;
wire n_1647;
wire n_1901;
wire n_3096;
wire n_3333;
wire n_839;
wire n_768;
wire n_3705;
wire n_3031;
wire n_1278;
wire n_2059;
wire n_796;
wire n_797;
wire n_3276;
wire n_1006;
wire n_2956;
wire n_1238;
wire n_1415;
wire n_3959;
wire n_3743;
wire n_976;
wire n_1710;
wire n_3021;
wire n_1063;
wire n_2153;
wire n_2452;
wire n_1270;
wire n_2891;
wire n_834;
wire n_2457;
wire n_3825;
wire n_2144;
wire n_1476;
wire n_935;
wire n_1603;
wire n_925;
wire n_2592;
wire n_1054;
wire n_2027;
wire n_3404;
wire n_2072;
wire n_2737;
wire n_2012;
wire n_2251;
wire n_2963;
wire n_3512;
wire n_1644;
wire n_3892;
wire n_1406;
wire n_1489;
wire n_3591;
wire n_1880;
wire n_1993;
wire n_3860;
wire n_2137;
wire n_804;
wire n_1455;
wire n_1642;
wire n_1871;
wire n_2182;
wire n_2868;
wire n_3044;
wire n_2447;
wire n_3493;
wire n_2818;
wire n_3358;
wire n_3115;
wire n_1057;
wire n_1473;
wire n_3140;
wire n_3486;
wire n_2125;
wire n_2426;
wire n_2894;
wire n_1403;
wire n_2181;
wire n_3253;
wire n_2587;
wire n_1149;
wire n_1176;
wire n_1502;
wire n_1605;
wire n_868;
wire n_2099;
wire n_3920;
wire n_1202;
wire n_3848;
wire n_1065;
wire n_1897;
wire n_2477;
wire n_1457;
wire n_3172;
wire n_905;
wire n_2159;
wire n_3410;
wire n_975;
wire n_934;
wire n_775;
wire n_3273;
wire n_950;
wire n_2700;
wire n_1222;
wire n_3139;
wire n_1630;
wire n_3408;
wire n_2286;
wire n_3182;
wire n_1879;
wire n_1959;
wire n_2563;
wire n_1198;
wire n_2206;
wire n_3734;
wire n_3637;
wire n_1311;
wire n_3393;
wire n_1261;
wire n_2299;
wire n_3538;
wire n_2078;
wire n_3650;
wire n_3327;
wire n_2265;
wire n_776;
wire n_1114;
wire n_3513;
wire n_3709;
wire n_3011;
wire n_818;
wire n_1167;
wire n_3231;
wire n_2677;
wire n_2531;
wire n_2315;
wire n_3623;
wire n_3647;
wire n_3138;
wire n_2157;
wire n_3212;
wire n_1282;
wire n_2067;
wire n_2517;
wire n_1321;
wire n_1779;
wire n_3446;
wire n_3349;
wire n_3619;
wire n_3928;
wire n_2489;
wire n_1770;
wire n_1107;
wire n_3058;
wire n_3454;
wire n_1846;
wire n_2211;
wire n_1573;
wire n_2950;
wire n_815;
wire n_919;
wire n_2272;
wire n_1956;
wire n_3574;
wire n_2608;
wire n_3384;
wire n_2983;
wire n_1718;
wire n_2225;
wire n_3229;
wire n_2546;
wire n_3739;
wire n_1411;
wire n_2825;
wire n_1139;
wire n_1018;
wire n_858;
wire n_2345;
wire n_1324;
wire n_1669;
wire n_1501;
wire n_2742;
wire n_782;
wire n_1885;
wire n_1740;
wire n_1989;
wire n_3540;
wire n_1838;
wire n_3604;
wire n_833;
wire n_3649;
wire n_3824;
wire n_2680;
wire n_1343;
wire n_1801;
wire n_3439;
wire n_1371;
wire n_1513;
wire n_3740;
wire n_3001;
wire n_2861;
wire n_2976;
wire n_2161;
wire n_2191;
wire n_3611;
wire n_2329;
wire n_1788;
wire n_2093;
wire n_2348;
wire n_786;
wire n_2576;
wire n_2417;
wire n_2675;
wire n_2043;
wire n_3601;
wire n_2366;
wire n_1621;
wire n_2338;
wire n_3571;
wire n_1919;
wire n_1342;
wire n_752;
wire n_2756;
wire n_2893;
wire n_2009;
wire n_2248;
wire n_958;
wire n_1175;
wire n_3500;
wire n_1416;
wire n_1659;
wire n_2850;
wire n_3465;
wire n_1221;
wire n_3962;
wire n_3875;
wire n_1047;
wire n_1878;
wire n_1515;
wire n_1374;
wire n_3846;
wire n_2851;
wire n_2438;
wire n_1435;
wire n_1688;
wire n_792;
wire n_2973;
wire n_3651;
wire n_1314;
wire n_1433;
wire n_2567;
wire n_3085;
wire n_3059;
wire n_1242;
wire n_1119;
wire n_2229;
wire n_2867;
wire n_2810;
wire n_3871;
wire n_1085;
wire n_3027;
wire n_2388;
wire n_2981;
wire n_3438;
wire n_2222;
wire n_3112;
wire n_1907;
wire n_3464;
wire n_885;
wire n_1530;
wire n_3215;
wire n_3413;
wire n_877;
wire n_2871;
wire n_2135;
wire n_1088;
wire n_896;
wire n_2764;
wire n_2624;
wire n_1813;
wire n_1451;
wire n_1005;
wire n_1102;
wire n_3234;
wire n_794;
wire n_3648;
wire n_2471;
wire n_1288;
wire n_1275;
wire n_985;
wire n_1165;
wire n_897;
wire n_1622;
wire n_2757;
wire n_2714;
wire n_3066;
wire n_2669;
wire n_2869;
wire n_1105;
wire n_1459;
wire n_912;
wire n_2898;
wire n_2232;
wire n_3121;
wire n_2455;
wire n_2121;
wire n_1893;
wire n_2519;
wire n_1570;
wire n_2231;
wire n_2874;
wire n_995;
wire n_2278;
wire n_1000;
wire n_2284;
wire n_1931;
wire n_2433;
wire n_2803;
wire n_2816;
wire n_3402;
wire n_1256;
wire n_2798;
wire n_3425;
wire n_1303;
wire n_1994;
wire n_1771;
wire n_3308;
wire n_1526;
wire n_764;
wire n_1507;
wire n_1206;
wire n_1809;
wire n_855;
wire n_2367;
wire n_812;
wire n_2658;
wire n_3236;
wire n_3576;
wire n_3109;
wire n_1961;
wire n_3491;
wire n_3271;
wire n_3013;
wire n_2553;
wire n_1050;
wire n_2218;
wire n_2667;
wire n_3062;
wire n_3806;
wire n_1769;
wire n_2130;
wire n_3256;
wire n_1060;
wire n_3126;
wire n_1372;
wire n_1847;
wire n_756;
wire n_1565;
wire n_1257;
wire n_3805;
wire n_2325;
wire n_2406;
wire n_1632;
wire n_2864;
wire n_3346;
wire n_3104;
wire n_3391;
wire n_1542;
wire n_1586;
wire n_1547;
wire n_1362;
wire n_946;
wire n_3497;
wire n_1097;
wire n_3354;
wire n_3288;
wire n_3373;
wire n_3382;
wire n_3122;
wire n_2518;
wire n_2784;
wire n_3012;
wire n_3045;
wire n_1909;
wire n_2543;
wire n_3368;
wire n_2381;
wire n_2313;
wire n_3561;
wire n_956;
wire n_3586;
wire n_790;
wire n_2495;
wire n_2992;
wire n_1541;
wire n_2703;
wire n_1812;
wire n_3014;
wire n_1951;
wire n_1330;
wire n_1697;
wire n_2128;
wire n_2574;
wire n_1872;
wire n_1940;
wire n_2690;
wire n_1747;
wire n_3767;
wire n_1212;
wire n_1887;
wire n_1199;
wire n_3400;
wire n_3942;
wire n_2020;
wire n_3504;
wire n_1978;
wire n_2508;
wire n_3511;
wire n_2540;
wire n_1767;
wire n_1939;
wire n_2428;
wire n_3820;
wire n_3159;
wire n_1768;
wire n_1443;
wire n_3697;
wire n_2068;
wire n_2636;
wire n_2672;
wire n_3360;
wire n_1585;
wire n_1861;
wire n_2316;
wire n_3101;
wire n_1564;
wire n_1995;
wire n_1631;
wire n_2593;
wire n_1623;
wire n_2911;
wire n_861;
wire n_1828;
wire n_3937;
wire n_2364;
wire n_1389;
wire n_3303;
wire n_1131;
wire n_2641;
wire n_1798;
wire n_1077;
wire n_3120;
wire n_1554;
wire n_3549;
wire n_1481;
wire n_1584;
wire n_2021;
wire n_1928;
wire n_2713;
wire n_828;
wire n_2938;
wire n_3227;
wire n_1438;
wire n_3774;
wire n_3972;
wire n_3342;
wire n_1973;
wire n_2314;
wire n_2939;
wire n_2494;
wire n_2156;
wire n_753;
wire n_2126;
wire n_747;
wire n_1147;
wire n_3403;
wire n_1363;
wire n_3863;
wire n_2228;
wire n_1691;
wire n_1098;
wire n_1518;
wire n_1366;
wire n_1187;
wire n_1361;
wire n_2034;
wire n_1693;
wire n_2790;
wire n_2872;
wire n_3102;
wire n_3173;
wire n_2411;
wire n_2081;
wire n_1892;
wire n_1061;
wire n_3539;
wire n_2266;
wire n_2993;
wire n_3433;
wire n_2061;
wire n_3018;
wire n_1373;
wire n_2449;
wire n_1686;
wire n_2131;
wire n_3866;
wire n_3761;
wire n_2526;
wire n_2830;
wire n_1302;
wire n_3803;
wire n_3017;
wire n_3083;
wire n_2083;
wire n_886;
wire n_2119;
wire n_1010;
wire n_3844;
wire n_883;
wire n_2207;
wire n_2044;
wire n_2542;
wire n_755;
wire n_2091;
wire n_3918;
wire n_2843;
wire n_3362;
wire n_3035;
wire n_3191;
wire n_1029;
wire n_3485;
wire n_2394;
wire n_3051;
wire n_770;
wire n_1572;
wire n_1635;
wire n_3305;
wire n_3149;
wire n_2827;
wire n_941;
wire n_1245;
wire n_1317;
wire n_3643;
wire n_2615;
wire n_3278;
wire n_2487;
wire n_2701;
wire n_2929;
wire n_3163;
wire n_3343;
wire n_3752;
wire n_3786;
wire n_1329;
wire n_2409;
wire n_2637;
wire n_2337;
wire n_854;
wire n_2405;
wire n_2601;
wire n_2513;
wire n_3118;
wire n_1369;
wire n_1297;
wire n_1912;
wire n_3143;
wire n_1734;
wire n_3543;
wire n_3655;
wire n_3742;
wire n_3791;
wire n_1876;
wire n_2666;
wire n_3050;
wire n_2323;
wire n_3532;
wire n_740;
wire n_1811;
wire n_898;
wire n_928;
wire n_1285;
wire n_3042;
wire n_967;
wire n_2561;
wire n_3725;
wire n_2913;
wire n_2491;
wire n_1529;
wire n_1381;
wire n_1824;
wire n_2254;
wire n_1597;
wire n_1161;
wire n_1103;
wire n_3522;
wire n_1486;
wire n_1068;
wire n_1833;
wire n_2914;
wire n_3551;
wire n_2371;
wire n_914;
wire n_3444;
wire n_1986;
wire n_3898;
wire n_3366;
wire n_2882;
wire n_1024;
wire n_3009;
wire n_1141;
wire n_3453;
wire n_3297;
wire n_3176;
wire n_1949;
wire n_1197;
wire n_2493;
wire n_2408;
wire n_2429;
wire n_3326;
wire n_1168;
wire n_865;
wire n_3581;
wire n_3000;
wire n_2115;
wire n_2013;
wire n_2140;
wire n_2134;
wire n_2483;
wire n_2305;
wire n_1556;
wire n_3423;
wire n_3547;
wire n_1192;
wire n_1646;
wire n_1290;
wire n_3700;
wire n_2514;
wire n_2466;
wire n_3661;
wire n_1759;
wire n_2048;
wire n_2760;
wire n_987;
wire n_1299;
wire n_750;
wire n_2942;
wire n_3947;
wire n_2096;
wire n_3663;
wire n_2129;
wire n_3230;
wire n_3545;
wire n_1101;
wire n_2532;
wire n_3665;
wire n_2079;
wire n_2296;
wire n_3782;
wire n_1720;
wire n_880;
wire n_2671;
wire n_1911;
wire n_2293;
wire n_3296;
wire n_3831;
wire n_1336;
wire n_3068;
wire n_3071;
wire n_3683;
wire n_3919;
wire n_2734;
wire n_2870;
wire n_758;
wire n_1166;
wire n_1390;
wire n_2775;
wire n_1023;
wire n_1358;
wire n_813;
wire n_2310;
wire n_3223;
wire n_3318;
wire n_1211;
wire n_1397;
wire n_2674;
wire n_1284;
wire n_2005;
wire n_3794;
wire n_1359;
wire n_1116;
wire n_2811;
wire n_1758;
wire n_3226;
wire n_3702;
wire n_791;
wire n_1532;
wire n_2848;
wire n_1419;
wire n_2689;
wire n_1784;
wire n_1685;
wire n_1992;
wire n_1082;
wire n_3200;
wire n_3430;
wire n_1213;
wire n_2596;
wire n_2801;
wire n_980;
wire n_1193;
wire n_849;
wire n_1488;
wire n_2928;
wire n_3067;
wire n_2227;
wire n_2652;
wire n_3557;
wire n_1074;
wire n_3225;
wire n_3596;
wire n_3380;
wire n_3207;
wire n_1379;
wire n_759;
wire n_1721;
wire n_2972;
wire n_2627;
wire n_1827;
wire n_953;
wire n_1180;
wire n_1462;
wire n_3606;
wire n_3369;
wire n_3823;
wire n_3185;
wire n_2326;
wire n_3869;
wire n_1866;
wire n_3852;
wire n_1220;
wire n_1398;
wire n_2169;
wire n_2111;
wire n_1262;
wire n_1904;
wire n_2966;
wire n_3084;
wire n_3036;
wire n_1692;
wire n_2501;
wire n_2051;
wire n_1012;
wire n_1805;
wire n_960;
wire n_1022;
wire n_1760;
wire n_3737;
wire n_1240;
wire n_2173;
wire n_1183;
wire n_3285;
wire n_3160;
wire n_3483;
wire n_1204;
wire n_1151;
wire n_2824;
wire n_1814;
wire n_771;
wire n_2982;
wire n_999;
wire n_2634;
wire n_3286;
wire n_3124;
wire n_1092;
wire n_1808;
wire n_2768;
wire n_2668;
wire n_1658;
wire n_1386;
wire n_3015;
wire n_2588;
wire n_2931;
wire n_3321;
wire n_3081;
wire n_2492;
wire n_3636;
wire n_910;
wire n_2291;
wire n_3837;
wire n_3612;
wire n_3046;
wire n_844;
wire n_2172;
wire n_1728;
wire n_1020;
wire n_3076;
wire n_1142;
wire n_1385;
wire n_783;
wire n_2927;
wire n_1062;
wire n_1230;
wire n_1027;
wire n_1516;
wire n_3893;
wire n_3622;
wire n_3857;
wire n_2533;
wire n_1499;
wire n_1500;
wire n_2155;
wire n_2706;
wire n_1868;
wire n_966;
wire n_2303;
wire n_2104;
wire n_949;
wire n_2357;
wire n_2148;
wire n_2618;
wire n_2653;
wire n_2855;
wire n_3938;
wire n_924;
wire n_2937;
wire n_3728;
wire n_3359;
wire n_3114;
wire n_2331;
wire n_3332;
wire n_3905;
wire n_1600;
wire n_1661;
wire n_2967;
wire n_1965;
wire n_3005;
wire n_1757;
wire n_2136;
wire n_3617;
wire n_3602;
wire n_2403;
wire n_918;
wire n_3053;
wire n_2056;
wire n_1913;
wire n_2702;
wire n_3922;
wire n_2054;
wire n_1039;
wire n_2226;
wire n_3894;
wire n_2407;
wire n_2791;
wire n_1043;
wire n_1402;
wire n_2267;
wire n_1450;
wire n_2302;
wire n_2082;
wire n_2560;
wire n_2453;
wire n_3056;
wire n_3267;
wire n_2092;
wire n_3008;
wire n_1472;
wire n_1365;
wire n_2443;
wire n_2802;
wire n_3189;
wire n_3052;
wire n_2797;
wire n_2279;
wire n_1089;
wire n_1536;
wire n_1049;
wire n_1719;
wire n_1974;
wire n_1158;
wire n_2066;
wire n_2988;
wire n_3945;
wire n_763;
wire n_1882;
wire n_2770;
wire n_2961;
wire n_2704;
wire n_2996;
wire n_3924;
wire n_1915;
wire n_2836;
wire n_940;
wire n_1762;
wire n_2534;
wire n_1404;
wire n_3582;
wire n_3689;
wire n_788;
wire n_3283;
wire n_1736;
wire n_3421;
wire n_2907;
wire n_3311;
wire n_1160;
wire n_1442;
wire n_1948;
wire n_2168;
wire n_1216;
wire n_2681;
wire n_1891;
wire n_1026;
wire n_3247;
wire n_2886;
wire n_1454;
wire n_1033;
wire n_3613;
wire n_1383;
wire n_990;
wire n_3675;
wire n_1968;
wire n_2057;
wire n_2609;
wire n_2378;
wire n_888;
wire n_2749;
wire n_3658;
wire n_1325;
wire n_3133;
wire n_2754;
wire n_3527;
wire n_2014;
wire n_3901;
wire n_3041;
wire n_1483;
wire n_1703;
wire n_1205;
wire n_1822;
wire n_843;
wire n_1953;
wire n_3715;
wire n_1059;
wire n_2969;
wire n_799;
wire n_3713;
wire n_2692;
wire n_3261;
wire n_3550;
wire n_1804;
wire n_1581;
wire n_3287;
wire n_3534;
wire n_1837;
wire n_3889;
wire n_3325;
wire n_1744;
wire n_1975;
wire n_3437;
wire n_3744;
wire n_1414;
wire n_2246;
wire n_2324;
wire n_2738;
wire n_3861;
wire n_3161;
wire n_1002;
wire n_1851;
wire n_1755;
wire n_2195;
wire n_2940;
wire n_1111;
wire n_1819;
wire n_3313;
wire n_1341;
wire n_1807;
wire n_2670;
wire n_2645;
wire n_2202;
wire n_1310;
wire n_3275;
wire n_1745;
wire n_1714;
wire n_3198;
wire n_3463;
wire n_3941;
wire n_1958;
wire n_1611;
wire n_2559;
wire n_3516;
wire n_2262;
wire n_3562;
wire n_3933;
wire n_955;
wire n_1333;
wire n_1916;
wire n_2619;
wire n_2917;
wire n_2726;
wire n_3873;
wire n_3738;
wire n_2073;
wire n_952;
wire n_1675;
wire n_1947;
wire n_2165;
wire n_1640;
wire n_2016;
wire n_3157;
wire n_1551;
wire n_3793;
wire n_1145;
wire n_1533;
wire n_2307;
wire n_2515;
wire n_3792;
wire n_3546;
wire n_1511;
wire n_1791;
wire n_1113;
wire n_3089;
wire n_1651;
wire n_1966;
wire n_2058;
wire n_2678;
wire n_3406;
wire n_1468;
wire n_3442;
wire n_2327;
wire n_3758;
wire n_2656;
wire n_913;
wire n_2353;
wire n_1164;
wire n_2258;
wire n_3944;
wire n_3662;
wire n_3595;
wire n_1732;
wire n_3749;
wire n_2167;
wire n_3079;
wire n_1354;
wire n_3329;
wire n_2039;
wire n_1277;
wire n_1696;
wire n_1016;
wire n_3233;
wire n_1355;
wire n_809;
wire n_3691;
wire n_2544;
wire n_856;
wire n_779;
wire n_3193;
wire n_3635;
wire n_3501;
wire n_2538;
wire n_3270;
wire n_2582;
wire n_1559;
wire n_2321;
wire n_2915;
wire n_1579;
wire n_1280;
wire n_2854;
wire n_2932;
wire n_3258;
wire n_1335;
wire n_3266;
wire n_2285;
wire n_3213;
wire n_3789;
wire n_1934;
wire n_1900;
wire n_2040;
wire n_2174;
wire n_3246;
wire n_1843;
wire n_2186;
wire n_2510;
wire n_2030;
wire n_2614;
wire n_3418;
wire n_2435;
wire n_3934;
wire n_1665;
wire n_2583;
wire n_3417;
wire n_1678;
wire n_1091;
wire n_1780;
wire n_2725;
wire n_3865;
wire n_1287;
wire n_2769;
wire n_1482;
wire n_860;
wire n_1525;
wire n_848;
wire n_3244;
wire n_3195;
wire n_3593;
wire n_2100;
wire n_2349;
wire n_1902;
wire n_2536;
wire n_3903;
wire n_2474;
wire n_3895;
wire n_1194;
wire n_1150;
wire n_1399;
wire n_3685;
wire n_3851;
wire n_1903;
wire n_1674;
wire n_1849;
wire n_3768;
wire n_867;
wire n_983;
wire n_1417;
wire n_3482;
wire n_2282;
wire n_970;
wire n_3654;
wire n_2430;
wire n_2676;
wire n_921;
wire n_2673;
wire n_3515;
wire n_3489;
wire n_2926;
wire n_1534;
wire n_2912;
wire n_3181;
wire n_908;
wire n_3536;
wire n_1346;
wire n_2834;
wire n_3644;
wire n_3268;
wire n_1123;
wire n_2710;
wire n_1272;
wire n_2497;
wire n_1393;
wire n_2970;
wire n_984;
wire n_1655;
wire n_3040;
wire n_3494;
wire n_2978;
wire n_3615;
wire n_1410;
wire n_988;
wire n_2368;
wire n_3363;
wire n_760;
wire n_3528;
wire n_1157;
wire n_3502;
wire n_806;
wire n_3677;
wire n_2657;
wire n_3935;
wire n_1186;
wire n_2065;
wire n_2901;
wire n_3180;
wire n_1743;
wire n_2743;
wire n_1854;
wire n_866;

HB1xp67_ASAP7_75t_L g739 ( 
.A(n_168),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_333),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_578),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_445),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_672),
.Y(n_743)
);

INVx1_ASAP7_75t_SL g744 ( 
.A(n_717),
.Y(n_744)
);

INVxp67_ASAP7_75t_SL g745 ( 
.A(n_375),
.Y(n_745)
);

INVx2_ASAP7_75t_SL g746 ( 
.A(n_384),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_252),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_543),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_48),
.Y(n_749)
);

NOR2xp67_ASAP7_75t_L g750 ( 
.A(n_725),
.B(n_642),
.Y(n_750)
);

BUFx3_ASAP7_75t_L g751 ( 
.A(n_538),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_90),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_318),
.Y(n_753)
);

NOR2xp67_ASAP7_75t_L g754 ( 
.A(n_705),
.B(n_686),
.Y(n_754)
);

CKINVDCx5p33_ASAP7_75t_R g755 ( 
.A(n_420),
.Y(n_755)
);

CKINVDCx5p33_ASAP7_75t_R g756 ( 
.A(n_256),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_543),
.Y(n_757)
);

CKINVDCx20_ASAP7_75t_R g758 ( 
.A(n_675),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_479),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_80),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_568),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_732),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_1),
.Y(n_763)
);

CKINVDCx5p33_ASAP7_75t_R g764 ( 
.A(n_606),
.Y(n_764)
);

INVx1_ASAP7_75t_SL g765 ( 
.A(n_20),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_135),
.Y(n_766)
);

CKINVDCx16_ASAP7_75t_R g767 ( 
.A(n_233),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_318),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_198),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_577),
.Y(n_770)
);

NOR2xp67_ASAP7_75t_L g771 ( 
.A(n_626),
.B(n_339),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_730),
.Y(n_772)
);

CKINVDCx5p33_ASAP7_75t_R g773 ( 
.A(n_577),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_404),
.Y(n_774)
);

BUFx5_ASAP7_75t_L g775 ( 
.A(n_280),
.Y(n_775)
);

INVxp67_ASAP7_75t_L g776 ( 
.A(n_494),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_310),
.Y(n_777)
);

CKINVDCx5p33_ASAP7_75t_R g778 ( 
.A(n_501),
.Y(n_778)
);

CKINVDCx5p33_ASAP7_75t_R g779 ( 
.A(n_706),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_15),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_612),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_346),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_348),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_445),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_344),
.Y(n_785)
);

CKINVDCx5p33_ASAP7_75t_R g786 ( 
.A(n_502),
.Y(n_786)
);

CKINVDCx16_ASAP7_75t_R g787 ( 
.A(n_734),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_129),
.Y(n_788)
);

CKINVDCx5p33_ASAP7_75t_R g789 ( 
.A(n_85),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_606),
.Y(n_790)
);

CKINVDCx5p33_ASAP7_75t_R g791 ( 
.A(n_719),
.Y(n_791)
);

BUFx3_ASAP7_75t_L g792 ( 
.A(n_674),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_698),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_514),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_695),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_620),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_449),
.Y(n_797)
);

CKINVDCx20_ASAP7_75t_R g798 ( 
.A(n_283),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_49),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_296),
.Y(n_800)
);

BUFx6f_ASAP7_75t_L g801 ( 
.A(n_17),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_271),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_542),
.Y(n_803)
);

BUFx5_ASAP7_75t_L g804 ( 
.A(n_501),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_509),
.Y(n_805)
);

CKINVDCx5p33_ASAP7_75t_R g806 ( 
.A(n_151),
.Y(n_806)
);

BUFx2_ASAP7_75t_L g807 ( 
.A(n_192),
.Y(n_807)
);

BUFx2_ASAP7_75t_L g808 ( 
.A(n_43),
.Y(n_808)
);

BUFx6f_ASAP7_75t_L g809 ( 
.A(n_231),
.Y(n_809)
);

CKINVDCx5p33_ASAP7_75t_R g810 ( 
.A(n_198),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_91),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_143),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_224),
.Y(n_813)
);

CKINVDCx5p33_ASAP7_75t_R g814 ( 
.A(n_692),
.Y(n_814)
);

BUFx3_ASAP7_75t_L g815 ( 
.A(n_341),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_436),
.Y(n_816)
);

BUFx3_ASAP7_75t_L g817 ( 
.A(n_715),
.Y(n_817)
);

BUFx3_ASAP7_75t_L g818 ( 
.A(n_535),
.Y(n_818)
);

CKINVDCx20_ASAP7_75t_R g819 ( 
.A(n_448),
.Y(n_819)
);

CKINVDCx5p33_ASAP7_75t_R g820 ( 
.A(n_416),
.Y(n_820)
);

CKINVDCx5p33_ASAP7_75t_R g821 ( 
.A(n_284),
.Y(n_821)
);

CKINVDCx5p33_ASAP7_75t_R g822 ( 
.A(n_408),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_293),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_691),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_441),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_519),
.Y(n_826)
);

INVx1_ASAP7_75t_SL g827 ( 
.A(n_301),
.Y(n_827)
);

BUFx2_ASAP7_75t_L g828 ( 
.A(n_431),
.Y(n_828)
);

CKINVDCx20_ASAP7_75t_R g829 ( 
.A(n_597),
.Y(n_829)
);

CKINVDCx16_ASAP7_75t_R g830 ( 
.A(n_648),
.Y(n_830)
);

BUFx6f_ASAP7_75t_L g831 ( 
.A(n_71),
.Y(n_831)
);

CKINVDCx5p33_ASAP7_75t_R g832 ( 
.A(n_142),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_399),
.Y(n_833)
);

CKINVDCx5p33_ASAP7_75t_R g834 ( 
.A(n_712),
.Y(n_834)
);

CKINVDCx5p33_ASAP7_75t_R g835 ( 
.A(n_440),
.Y(n_835)
);

NOR2xp67_ASAP7_75t_L g836 ( 
.A(n_411),
.B(n_155),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_291),
.Y(n_837)
);

CKINVDCx5p33_ASAP7_75t_R g838 ( 
.A(n_452),
.Y(n_838)
);

INVx1_ASAP7_75t_SL g839 ( 
.A(n_16),
.Y(n_839)
);

CKINVDCx5p33_ASAP7_75t_R g840 ( 
.A(n_431),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_478),
.Y(n_841)
);

CKINVDCx5p33_ASAP7_75t_R g842 ( 
.A(n_29),
.Y(n_842)
);

CKINVDCx5p33_ASAP7_75t_R g843 ( 
.A(n_169),
.Y(n_843)
);

CKINVDCx5p33_ASAP7_75t_R g844 ( 
.A(n_491),
.Y(n_844)
);

XOR2xp5_ASAP7_75t_R g845 ( 
.A(n_145),
.B(n_701),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_268),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_216),
.Y(n_847)
);

BUFx6f_ASAP7_75t_L g848 ( 
.A(n_555),
.Y(n_848)
);

BUFx3_ASAP7_75t_L g849 ( 
.A(n_685),
.Y(n_849)
);

CKINVDCx16_ASAP7_75t_R g850 ( 
.A(n_713),
.Y(n_850)
);

CKINVDCx5p33_ASAP7_75t_R g851 ( 
.A(n_203),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_46),
.Y(n_852)
);

CKINVDCx5p33_ASAP7_75t_R g853 ( 
.A(n_53),
.Y(n_853)
);

CKINVDCx5p33_ASAP7_75t_R g854 ( 
.A(n_425),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_722),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_620),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_707),
.Y(n_857)
);

CKINVDCx5p33_ASAP7_75t_R g858 ( 
.A(n_278),
.Y(n_858)
);

CKINVDCx20_ASAP7_75t_R g859 ( 
.A(n_625),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_616),
.Y(n_860)
);

INVx1_ASAP7_75t_SL g861 ( 
.A(n_679),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_704),
.Y(n_862)
);

INVx1_ASAP7_75t_SL g863 ( 
.A(n_660),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_135),
.Y(n_864)
);

INVx2_ASAP7_75t_L g865 ( 
.A(n_633),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_221),
.Y(n_866)
);

CKINVDCx5p33_ASAP7_75t_R g867 ( 
.A(n_186),
.Y(n_867)
);

CKINVDCx5p33_ASAP7_75t_R g868 ( 
.A(n_64),
.Y(n_868)
);

BUFx5_ASAP7_75t_L g869 ( 
.A(n_345),
.Y(n_869)
);

CKINVDCx5p33_ASAP7_75t_R g870 ( 
.A(n_121),
.Y(n_870)
);

INVx1_ASAP7_75t_SL g871 ( 
.A(n_89),
.Y(n_871)
);

CKINVDCx5p33_ASAP7_75t_R g872 ( 
.A(n_335),
.Y(n_872)
);

CKINVDCx20_ASAP7_75t_R g873 ( 
.A(n_256),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_283),
.Y(n_874)
);

CKINVDCx5p33_ASAP7_75t_R g875 ( 
.A(n_33),
.Y(n_875)
);

CKINVDCx5p33_ASAP7_75t_R g876 ( 
.A(n_75),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_253),
.Y(n_877)
);

CKINVDCx5p33_ASAP7_75t_R g878 ( 
.A(n_735),
.Y(n_878)
);

CKINVDCx20_ASAP7_75t_R g879 ( 
.A(n_367),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_475),
.Y(n_880)
);

CKINVDCx5p33_ASAP7_75t_R g881 ( 
.A(n_23),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_80),
.Y(n_882)
);

CKINVDCx5p33_ASAP7_75t_R g883 ( 
.A(n_127),
.Y(n_883)
);

CKINVDCx5p33_ASAP7_75t_R g884 ( 
.A(n_693),
.Y(n_884)
);

CKINVDCx20_ASAP7_75t_R g885 ( 
.A(n_699),
.Y(n_885)
);

CKINVDCx5p33_ASAP7_75t_R g886 ( 
.A(n_723),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_626),
.Y(n_887)
);

CKINVDCx5p33_ASAP7_75t_R g888 ( 
.A(n_605),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_470),
.Y(n_889)
);

CKINVDCx5p33_ASAP7_75t_R g890 ( 
.A(n_636),
.Y(n_890)
);

BUFx2_ASAP7_75t_L g891 ( 
.A(n_10),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_670),
.Y(n_892)
);

NOR2xp33_ASAP7_75t_L g893 ( 
.A(n_437),
.B(n_435),
.Y(n_893)
);

BUFx6f_ASAP7_75t_L g894 ( 
.A(n_637),
.Y(n_894)
);

CKINVDCx5p33_ASAP7_75t_R g895 ( 
.A(n_264),
.Y(n_895)
);

CKINVDCx16_ASAP7_75t_R g896 ( 
.A(n_26),
.Y(n_896)
);

CKINVDCx5p33_ASAP7_75t_R g897 ( 
.A(n_522),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_530),
.Y(n_898)
);

CKINVDCx20_ASAP7_75t_R g899 ( 
.A(n_258),
.Y(n_899)
);

CKINVDCx5p33_ASAP7_75t_R g900 ( 
.A(n_624),
.Y(n_900)
);

CKINVDCx5p33_ASAP7_75t_R g901 ( 
.A(n_21),
.Y(n_901)
);

CKINVDCx5p33_ASAP7_75t_R g902 ( 
.A(n_167),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_79),
.Y(n_903)
);

CKINVDCx5p33_ASAP7_75t_R g904 ( 
.A(n_203),
.Y(n_904)
);

CKINVDCx5p33_ASAP7_75t_R g905 ( 
.A(n_523),
.Y(n_905)
);

CKINVDCx5p33_ASAP7_75t_R g906 ( 
.A(n_635),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_266),
.Y(n_907)
);

INVxp67_ASAP7_75t_L g908 ( 
.A(n_207),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_396),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_231),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_374),
.Y(n_911)
);

INVx2_ASAP7_75t_L g912 ( 
.A(n_623),
.Y(n_912)
);

CKINVDCx5p33_ASAP7_75t_R g913 ( 
.A(n_639),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_151),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_77),
.Y(n_915)
);

CKINVDCx5p33_ASAP7_75t_R g916 ( 
.A(n_557),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_112),
.Y(n_917)
);

CKINVDCx5p33_ASAP7_75t_R g918 ( 
.A(n_703),
.Y(n_918)
);

CKINVDCx5p33_ASAP7_75t_R g919 ( 
.A(n_627),
.Y(n_919)
);

CKINVDCx5p33_ASAP7_75t_R g920 ( 
.A(n_619),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_251),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_47),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_733),
.Y(n_923)
);

INVx1_ASAP7_75t_SL g924 ( 
.A(n_34),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_498),
.Y(n_925)
);

CKINVDCx5p33_ASAP7_75t_R g926 ( 
.A(n_381),
.Y(n_926)
);

CKINVDCx5p33_ASAP7_75t_R g927 ( 
.A(n_630),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_254),
.Y(n_928)
);

CKINVDCx5p33_ASAP7_75t_R g929 ( 
.A(n_138),
.Y(n_929)
);

INVx1_ASAP7_75t_SL g930 ( 
.A(n_50),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_121),
.Y(n_931)
);

CKINVDCx5p33_ASAP7_75t_R g932 ( 
.A(n_444),
.Y(n_932)
);

CKINVDCx5p33_ASAP7_75t_R g933 ( 
.A(n_322),
.Y(n_933)
);

CKINVDCx5p33_ASAP7_75t_R g934 ( 
.A(n_644),
.Y(n_934)
);

CKINVDCx5p33_ASAP7_75t_R g935 ( 
.A(n_60),
.Y(n_935)
);

CKINVDCx5p33_ASAP7_75t_R g936 ( 
.A(n_248),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_528),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_176),
.Y(n_938)
);

INVx1_ASAP7_75t_SL g939 ( 
.A(n_495),
.Y(n_939)
);

CKINVDCx5p33_ASAP7_75t_R g940 ( 
.A(n_49),
.Y(n_940)
);

CKINVDCx5p33_ASAP7_75t_R g941 ( 
.A(n_504),
.Y(n_941)
);

CKINVDCx5p33_ASAP7_75t_R g942 ( 
.A(n_456),
.Y(n_942)
);

CKINVDCx20_ASAP7_75t_R g943 ( 
.A(n_396),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_595),
.Y(n_944)
);

CKINVDCx5p33_ASAP7_75t_R g945 ( 
.A(n_684),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_403),
.Y(n_946)
);

CKINVDCx5p33_ASAP7_75t_R g947 ( 
.A(n_295),
.Y(n_947)
);

HB1xp67_ASAP7_75t_L g948 ( 
.A(n_204),
.Y(n_948)
);

INVx1_ASAP7_75t_SL g949 ( 
.A(n_622),
.Y(n_949)
);

CKINVDCx5p33_ASAP7_75t_R g950 ( 
.A(n_714),
.Y(n_950)
);

CKINVDCx5p33_ASAP7_75t_R g951 ( 
.A(n_430),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_548),
.Y(n_952)
);

BUFx6f_ASAP7_75t_L g953 ( 
.A(n_689),
.Y(n_953)
);

CKINVDCx20_ASAP7_75t_R g954 ( 
.A(n_224),
.Y(n_954)
);

CKINVDCx5p33_ASAP7_75t_R g955 ( 
.A(n_434),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_250),
.Y(n_956)
);

BUFx6f_ASAP7_75t_L g957 ( 
.A(n_164),
.Y(n_957)
);

CKINVDCx20_ASAP7_75t_R g958 ( 
.A(n_242),
.Y(n_958)
);

CKINVDCx5p33_ASAP7_75t_R g959 ( 
.A(n_456),
.Y(n_959)
);

CKINVDCx5p33_ASAP7_75t_R g960 ( 
.A(n_711),
.Y(n_960)
);

CKINVDCx5p33_ASAP7_75t_R g961 ( 
.A(n_47),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_708),
.Y(n_962)
);

CKINVDCx5p33_ASAP7_75t_R g963 ( 
.A(n_127),
.Y(n_963)
);

CKINVDCx5p33_ASAP7_75t_R g964 ( 
.A(n_716),
.Y(n_964)
);

NOR2xp33_ASAP7_75t_L g965 ( 
.A(n_186),
.B(n_568),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_355),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_126),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_358),
.Y(n_968)
);

CKINVDCx5p33_ASAP7_75t_R g969 ( 
.A(n_153),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_358),
.Y(n_970)
);

INVx2_ASAP7_75t_SL g971 ( 
.A(n_532),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_530),
.Y(n_972)
);

CKINVDCx5p33_ASAP7_75t_R g973 ( 
.A(n_175),
.Y(n_973)
);

INVx2_ASAP7_75t_L g974 ( 
.A(n_2),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_114),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_726),
.Y(n_976)
);

BUFx10_ASAP7_75t_L g977 ( 
.A(n_423),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_738),
.Y(n_978)
);

CKINVDCx5p33_ASAP7_75t_R g979 ( 
.A(n_649),
.Y(n_979)
);

HB1xp67_ASAP7_75t_L g980 ( 
.A(n_570),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_622),
.Y(n_981)
);

CKINVDCx5p33_ASAP7_75t_R g982 ( 
.A(n_190),
.Y(n_982)
);

BUFx10_ASAP7_75t_L g983 ( 
.A(n_226),
.Y(n_983)
);

CKINVDCx20_ASAP7_75t_R g984 ( 
.A(n_408),
.Y(n_984)
);

CKINVDCx5p33_ASAP7_75t_R g985 ( 
.A(n_140),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_123),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_329),
.Y(n_987)
);

INVx1_ASAP7_75t_SL g988 ( 
.A(n_539),
.Y(n_988)
);

CKINVDCx5p33_ASAP7_75t_R g989 ( 
.A(n_617),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_601),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_42),
.Y(n_991)
);

INVxp67_ASAP7_75t_L g992 ( 
.A(n_10),
.Y(n_992)
);

INVx1_ASAP7_75t_SL g993 ( 
.A(n_102),
.Y(n_993)
);

CKINVDCx5p33_ASAP7_75t_R g994 ( 
.A(n_138),
.Y(n_994)
);

INVx2_ASAP7_75t_SL g995 ( 
.A(n_434),
.Y(n_995)
);

CKINVDCx5p33_ASAP7_75t_R g996 ( 
.A(n_73),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_6),
.Y(n_997)
);

INVxp67_ASAP7_75t_L g998 ( 
.A(n_634),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_618),
.Y(n_999)
);

CKINVDCx5p33_ASAP7_75t_R g1000 ( 
.A(n_621),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_582),
.Y(n_1001)
);

CKINVDCx5p33_ASAP7_75t_R g1002 ( 
.A(n_404),
.Y(n_1002)
);

CKINVDCx20_ASAP7_75t_R g1003 ( 
.A(n_544),
.Y(n_1003)
);

CKINVDCx5p33_ASAP7_75t_R g1004 ( 
.A(n_9),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_223),
.Y(n_1005)
);

CKINVDCx5p33_ASAP7_75t_R g1006 ( 
.A(n_602),
.Y(n_1006)
);

BUFx10_ASAP7_75t_L g1007 ( 
.A(n_614),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_176),
.Y(n_1008)
);

CKINVDCx5p33_ASAP7_75t_R g1009 ( 
.A(n_61),
.Y(n_1009)
);

CKINVDCx5p33_ASAP7_75t_R g1010 ( 
.A(n_11),
.Y(n_1010)
);

CKINVDCx5p33_ASAP7_75t_R g1011 ( 
.A(n_90),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_350),
.Y(n_1012)
);

CKINVDCx5p33_ASAP7_75t_R g1013 ( 
.A(n_688),
.Y(n_1013)
);

CKINVDCx5p33_ASAP7_75t_R g1014 ( 
.A(n_457),
.Y(n_1014)
);

CKINVDCx5p33_ASAP7_75t_R g1015 ( 
.A(n_297),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_656),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_681),
.Y(n_1017)
);

CKINVDCx5p33_ASAP7_75t_R g1018 ( 
.A(n_463),
.Y(n_1018)
);

INVx2_ASAP7_75t_L g1019 ( 
.A(n_70),
.Y(n_1019)
);

INVx2_ASAP7_75t_L g1020 ( 
.A(n_143),
.Y(n_1020)
);

CKINVDCx5p33_ASAP7_75t_R g1021 ( 
.A(n_368),
.Y(n_1021)
);

HB1xp67_ASAP7_75t_L g1022 ( 
.A(n_357),
.Y(n_1022)
);

CKINVDCx5p33_ASAP7_75t_R g1023 ( 
.A(n_489),
.Y(n_1023)
);

INVx1_ASAP7_75t_SL g1024 ( 
.A(n_294),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_435),
.Y(n_1025)
);

CKINVDCx20_ASAP7_75t_R g1026 ( 
.A(n_228),
.Y(n_1026)
);

CKINVDCx5p33_ASAP7_75t_R g1027 ( 
.A(n_736),
.Y(n_1027)
);

INVx2_ASAP7_75t_SL g1028 ( 
.A(n_641),
.Y(n_1028)
);

CKINVDCx5p33_ASAP7_75t_R g1029 ( 
.A(n_665),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_690),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_682),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_250),
.Y(n_1032)
);

BUFx10_ASAP7_75t_L g1033 ( 
.A(n_220),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_406),
.Y(n_1034)
);

CKINVDCx5p33_ASAP7_75t_R g1035 ( 
.A(n_196),
.Y(n_1035)
);

BUFx3_ASAP7_75t_L g1036 ( 
.A(n_249),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_667),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_438),
.Y(n_1038)
);

CKINVDCx20_ASAP7_75t_R g1039 ( 
.A(n_152),
.Y(n_1039)
);

INVx2_ASAP7_75t_L g1040 ( 
.A(n_260),
.Y(n_1040)
);

CKINVDCx5p33_ASAP7_75t_R g1041 ( 
.A(n_7),
.Y(n_1041)
);

INVxp67_ASAP7_75t_L g1042 ( 
.A(n_167),
.Y(n_1042)
);

CKINVDCx5p33_ASAP7_75t_R g1043 ( 
.A(n_130),
.Y(n_1043)
);

CKINVDCx5p33_ASAP7_75t_R g1044 ( 
.A(n_59),
.Y(n_1044)
);

CKINVDCx5p33_ASAP7_75t_R g1045 ( 
.A(n_53),
.Y(n_1045)
);

INVx2_ASAP7_75t_L g1046 ( 
.A(n_702),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_361),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_628),
.Y(n_1048)
);

CKINVDCx20_ASAP7_75t_R g1049 ( 
.A(n_593),
.Y(n_1049)
);

BUFx10_ASAP7_75t_L g1050 ( 
.A(n_103),
.Y(n_1050)
);

BUFx3_ASAP7_75t_L g1051 ( 
.A(n_613),
.Y(n_1051)
);

BUFx6f_ASAP7_75t_L g1052 ( 
.A(n_375),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_16),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_472),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_238),
.Y(n_1055)
);

CKINVDCx5p33_ASAP7_75t_R g1056 ( 
.A(n_113),
.Y(n_1056)
);

BUFx3_ASAP7_75t_L g1057 ( 
.A(n_389),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_428),
.Y(n_1058)
);

INVx1_ASAP7_75t_SL g1059 ( 
.A(n_631),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_493),
.Y(n_1060)
);

CKINVDCx5p33_ASAP7_75t_R g1061 ( 
.A(n_291),
.Y(n_1061)
);

BUFx3_ASAP7_75t_L g1062 ( 
.A(n_134),
.Y(n_1062)
);

HB1xp67_ASAP7_75t_L g1063 ( 
.A(n_227),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_357),
.Y(n_1064)
);

CKINVDCx5p33_ASAP7_75t_R g1065 ( 
.A(n_300),
.Y(n_1065)
);

CKINVDCx5p33_ASAP7_75t_R g1066 ( 
.A(n_18),
.Y(n_1066)
);

CKINVDCx5p33_ASAP7_75t_R g1067 ( 
.A(n_687),
.Y(n_1067)
);

CKINVDCx5p33_ASAP7_75t_R g1068 ( 
.A(n_272),
.Y(n_1068)
);

INVx1_ASAP7_75t_SL g1069 ( 
.A(n_179),
.Y(n_1069)
);

CKINVDCx5p33_ASAP7_75t_R g1070 ( 
.A(n_413),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_523),
.Y(n_1071)
);

INVx1_ASAP7_75t_SL g1072 ( 
.A(n_181),
.Y(n_1072)
);

CKINVDCx5p33_ASAP7_75t_R g1073 ( 
.A(n_454),
.Y(n_1073)
);

CKINVDCx5p33_ASAP7_75t_R g1074 ( 
.A(n_328),
.Y(n_1074)
);

CKINVDCx5p33_ASAP7_75t_R g1075 ( 
.A(n_727),
.Y(n_1075)
);

CKINVDCx5p33_ASAP7_75t_R g1076 ( 
.A(n_700),
.Y(n_1076)
);

BUFx6f_ASAP7_75t_L g1077 ( 
.A(n_99),
.Y(n_1077)
);

INVx2_ASAP7_75t_L g1078 ( 
.A(n_473),
.Y(n_1078)
);

CKINVDCx5p33_ASAP7_75t_R g1079 ( 
.A(n_468),
.Y(n_1079)
);

CKINVDCx20_ASAP7_75t_R g1080 ( 
.A(n_611),
.Y(n_1080)
);

BUFx3_ASAP7_75t_L g1081 ( 
.A(n_643),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_14),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_55),
.Y(n_1083)
);

CKINVDCx5p33_ASAP7_75t_R g1084 ( 
.A(n_230),
.Y(n_1084)
);

CKINVDCx5p33_ASAP7_75t_R g1085 ( 
.A(n_632),
.Y(n_1085)
);

INVxp67_ASAP7_75t_L g1086 ( 
.A(n_8),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_201),
.Y(n_1087)
);

CKINVDCx20_ASAP7_75t_R g1088 ( 
.A(n_140),
.Y(n_1088)
);

CKINVDCx5p33_ASAP7_75t_R g1089 ( 
.A(n_219),
.Y(n_1089)
);

CKINVDCx5p33_ASAP7_75t_R g1090 ( 
.A(n_585),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_175),
.Y(n_1091)
);

INVx2_ASAP7_75t_SL g1092 ( 
.A(n_591),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_398),
.Y(n_1093)
);

CKINVDCx5p33_ASAP7_75t_R g1094 ( 
.A(n_655),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_553),
.Y(n_1095)
);

CKINVDCx5p33_ASAP7_75t_R g1096 ( 
.A(n_102),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_126),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_721),
.Y(n_1098)
);

CKINVDCx5p33_ASAP7_75t_R g1099 ( 
.A(n_156),
.Y(n_1099)
);

CKINVDCx5p33_ASAP7_75t_R g1100 ( 
.A(n_213),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_74),
.Y(n_1101)
);

CKINVDCx5p33_ASAP7_75t_R g1102 ( 
.A(n_234),
.Y(n_1102)
);

CKINVDCx5p33_ASAP7_75t_R g1103 ( 
.A(n_444),
.Y(n_1103)
);

BUFx2_ASAP7_75t_SL g1104 ( 
.A(n_516),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_93),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_100),
.Y(n_1106)
);

CKINVDCx5p33_ASAP7_75t_R g1107 ( 
.A(n_257),
.Y(n_1107)
);

INVxp33_ASAP7_75t_L g1108 ( 
.A(n_306),
.Y(n_1108)
);

CKINVDCx14_ASAP7_75t_R g1109 ( 
.A(n_737),
.Y(n_1109)
);

CKINVDCx5p33_ASAP7_75t_R g1110 ( 
.A(n_627),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_293),
.Y(n_1111)
);

CKINVDCx5p33_ASAP7_75t_R g1112 ( 
.A(n_413),
.Y(n_1112)
);

CKINVDCx20_ASAP7_75t_R g1113 ( 
.A(n_650),
.Y(n_1113)
);

BUFx3_ASAP7_75t_L g1114 ( 
.A(n_78),
.Y(n_1114)
);

CKINVDCx5p33_ASAP7_75t_R g1115 ( 
.A(n_544),
.Y(n_1115)
);

INVx1_ASAP7_75t_SL g1116 ( 
.A(n_308),
.Y(n_1116)
);

CKINVDCx20_ASAP7_75t_R g1117 ( 
.A(n_600),
.Y(n_1117)
);

CKINVDCx5p33_ASAP7_75t_R g1118 ( 
.A(n_221),
.Y(n_1118)
);

CKINVDCx5p33_ASAP7_75t_R g1119 ( 
.A(n_279),
.Y(n_1119)
);

CKINVDCx5p33_ASAP7_75t_R g1120 ( 
.A(n_7),
.Y(n_1120)
);

CKINVDCx5p33_ASAP7_75t_R g1121 ( 
.A(n_459),
.Y(n_1121)
);

CKINVDCx5p33_ASAP7_75t_R g1122 ( 
.A(n_210),
.Y(n_1122)
);

CKINVDCx5p33_ASAP7_75t_R g1123 ( 
.A(n_491),
.Y(n_1123)
);

CKINVDCx20_ASAP7_75t_R g1124 ( 
.A(n_683),
.Y(n_1124)
);

CKINVDCx5p33_ASAP7_75t_R g1125 ( 
.A(n_171),
.Y(n_1125)
);

CKINVDCx5p33_ASAP7_75t_R g1126 ( 
.A(n_220),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_338),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_82),
.Y(n_1128)
);

CKINVDCx5p33_ASAP7_75t_R g1129 ( 
.A(n_559),
.Y(n_1129)
);

CKINVDCx5p33_ASAP7_75t_R g1130 ( 
.A(n_60),
.Y(n_1130)
);

CKINVDCx5p33_ASAP7_75t_R g1131 ( 
.A(n_697),
.Y(n_1131)
);

CKINVDCx20_ASAP7_75t_R g1132 ( 
.A(n_374),
.Y(n_1132)
);

INVx1_ASAP7_75t_SL g1133 ( 
.A(n_14),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_729),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_181),
.Y(n_1135)
);

CKINVDCx5p33_ASAP7_75t_R g1136 ( 
.A(n_371),
.Y(n_1136)
);

CKINVDCx5p33_ASAP7_75t_R g1137 ( 
.A(n_629),
.Y(n_1137)
);

CKINVDCx5p33_ASAP7_75t_R g1138 ( 
.A(n_520),
.Y(n_1138)
);

BUFx10_ASAP7_75t_L g1139 ( 
.A(n_635),
.Y(n_1139)
);

CKINVDCx20_ASAP7_75t_R g1140 ( 
.A(n_402),
.Y(n_1140)
);

BUFx10_ASAP7_75t_L g1141 ( 
.A(n_614),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_671),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_332),
.Y(n_1143)
);

CKINVDCx5p33_ASAP7_75t_R g1144 ( 
.A(n_9),
.Y(n_1144)
);

BUFx3_ASAP7_75t_L g1145 ( 
.A(n_77),
.Y(n_1145)
);

BUFx6f_ASAP7_75t_L g1146 ( 
.A(n_382),
.Y(n_1146)
);

CKINVDCx5p33_ASAP7_75t_R g1147 ( 
.A(n_487),
.Y(n_1147)
);

INVx2_ASAP7_75t_SL g1148 ( 
.A(n_320),
.Y(n_1148)
);

CKINVDCx5p33_ASAP7_75t_R g1149 ( 
.A(n_465),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_300),
.Y(n_1150)
);

CKINVDCx20_ASAP7_75t_R g1151 ( 
.A(n_350),
.Y(n_1151)
);

HB1xp67_ASAP7_75t_L g1152 ( 
.A(n_673),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_678),
.Y(n_1153)
);

CKINVDCx5p33_ASAP7_75t_R g1154 ( 
.A(n_108),
.Y(n_1154)
);

CKINVDCx5p33_ASAP7_75t_R g1155 ( 
.A(n_170),
.Y(n_1155)
);

CKINVDCx5p33_ASAP7_75t_R g1156 ( 
.A(n_1),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_632),
.Y(n_1157)
);

INVx2_ASAP7_75t_L g1158 ( 
.A(n_647),
.Y(n_1158)
);

CKINVDCx5p33_ASAP7_75t_R g1159 ( 
.A(n_27),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_630),
.Y(n_1160)
);

CKINVDCx5p33_ASAP7_75t_R g1161 ( 
.A(n_248),
.Y(n_1161)
);

CKINVDCx5p33_ASAP7_75t_R g1162 ( 
.A(n_339),
.Y(n_1162)
);

CKINVDCx5p33_ASAP7_75t_R g1163 ( 
.A(n_302),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_128),
.Y(n_1164)
);

CKINVDCx5p33_ASAP7_75t_R g1165 ( 
.A(n_596),
.Y(n_1165)
);

CKINVDCx5p33_ASAP7_75t_R g1166 ( 
.A(n_378),
.Y(n_1166)
);

CKINVDCx5p33_ASAP7_75t_R g1167 ( 
.A(n_330),
.Y(n_1167)
);

CKINVDCx5p33_ASAP7_75t_R g1168 ( 
.A(n_482),
.Y(n_1168)
);

CKINVDCx5p33_ASAP7_75t_R g1169 ( 
.A(n_147),
.Y(n_1169)
);

CKINVDCx5p33_ASAP7_75t_R g1170 ( 
.A(n_131),
.Y(n_1170)
);

CKINVDCx5p33_ASAP7_75t_R g1171 ( 
.A(n_124),
.Y(n_1171)
);

CKINVDCx5p33_ASAP7_75t_R g1172 ( 
.A(n_133),
.Y(n_1172)
);

BUFx5_ASAP7_75t_L g1173 ( 
.A(n_50),
.Y(n_1173)
);

BUFx5_ASAP7_75t_L g1174 ( 
.A(n_615),
.Y(n_1174)
);

BUFx10_ASAP7_75t_L g1175 ( 
.A(n_97),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_142),
.Y(n_1176)
);

HB1xp67_ASAP7_75t_L g1177 ( 
.A(n_512),
.Y(n_1177)
);

CKINVDCx5p33_ASAP7_75t_R g1178 ( 
.A(n_680),
.Y(n_1178)
);

CKINVDCx5p33_ASAP7_75t_R g1179 ( 
.A(n_513),
.Y(n_1179)
);

CKINVDCx5p33_ASAP7_75t_R g1180 ( 
.A(n_316),
.Y(n_1180)
);

OAI22x1_ASAP7_75t_SL g1181 ( 
.A1(n_879),
.A2(n_943),
.B1(n_954),
.B2(n_899),
.Y(n_1181)
);

OA21x2_ASAP7_75t_L g1182 ( 
.A1(n_1046),
.A2(n_646),
.B(n_645),
.Y(n_1182)
);

BUFx3_ASAP7_75t_L g1183 ( 
.A(n_792),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_SL g1184 ( 
.A(n_1046),
.B(n_1158),
.Y(n_1184)
);

INVx2_ASAP7_75t_L g1185 ( 
.A(n_775),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_1152),
.Y(n_1186)
);

BUFx8_ASAP7_75t_SL g1187 ( 
.A(n_879),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_746),
.B(n_0),
.Y(n_1188)
);

OAI21x1_ASAP7_75t_L g1189 ( 
.A1(n_1158),
.A2(n_652),
.B(n_651),
.Y(n_1189)
);

AOI22xp5_ASAP7_75t_L g1190 ( 
.A1(n_767),
.A2(n_4),
.B1(n_2),
.B2(n_3),
.Y(n_1190)
);

AND2x2_ASAP7_75t_L g1191 ( 
.A(n_1108),
.B(n_3),
.Y(n_1191)
);

INVx2_ASAP7_75t_L g1192 ( 
.A(n_775),
.Y(n_1192)
);

BUFx12f_ASAP7_75t_L g1193 ( 
.A(n_977),
.Y(n_1193)
);

BUFx12f_ASAP7_75t_L g1194 ( 
.A(n_977),
.Y(n_1194)
);

BUFx6f_ASAP7_75t_L g1195 ( 
.A(n_953),
.Y(n_1195)
);

NOR2xp33_ASAP7_75t_SL g1196 ( 
.A(n_787),
.B(n_653),
.Y(n_1196)
);

AND2x4_ASAP7_75t_L g1197 ( 
.A(n_751),
.B(n_4),
.Y(n_1197)
);

OAI22x1_ASAP7_75t_L g1198 ( 
.A1(n_745),
.A2(n_8),
.B1(n_5),
.B2(n_6),
.Y(n_1198)
);

INVx3_ASAP7_75t_L g1199 ( 
.A(n_977),
.Y(n_1199)
);

INVx2_ASAP7_75t_L g1200 ( 
.A(n_775),
.Y(n_1200)
);

BUFx6f_ASAP7_75t_L g1201 ( 
.A(n_953),
.Y(n_1201)
);

BUFx8_ASAP7_75t_L g1202 ( 
.A(n_807),
.Y(n_1202)
);

OAI22xp5_ASAP7_75t_L g1203 ( 
.A1(n_896),
.A2(n_12),
.B1(n_5),
.B2(n_11),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_751),
.Y(n_1204)
);

INVx5_ASAP7_75t_L g1205 ( 
.A(n_953),
.Y(n_1205)
);

BUFx6f_ASAP7_75t_L g1206 ( 
.A(n_953),
.Y(n_1206)
);

BUFx6f_ASAP7_75t_L g1207 ( 
.A(n_801),
.Y(n_1207)
);

NOR2x1_ASAP7_75t_L g1208 ( 
.A(n_815),
.B(n_654),
.Y(n_1208)
);

AND2x2_ASAP7_75t_L g1209 ( 
.A(n_1108),
.B(n_12),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_815),
.Y(n_1210)
);

CKINVDCx5p33_ASAP7_75t_R g1211 ( 
.A(n_830),
.Y(n_1211)
);

AND2x2_ASAP7_75t_L g1212 ( 
.A(n_808),
.B(n_13),
.Y(n_1212)
);

INVx5_ASAP7_75t_L g1213 ( 
.A(n_1028),
.Y(n_1213)
);

INVx2_ASAP7_75t_L g1214 ( 
.A(n_775),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_971),
.B(n_13),
.Y(n_1215)
);

HB1xp67_ASAP7_75t_L g1216 ( 
.A(n_739),
.Y(n_1216)
);

INVx4_ASAP7_75t_L g1217 ( 
.A(n_743),
.Y(n_1217)
);

BUFx8_ASAP7_75t_SL g1218 ( 
.A(n_899),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_995),
.B(n_15),
.Y(n_1219)
);

BUFx12f_ASAP7_75t_L g1220 ( 
.A(n_983),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_818),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_SL g1222 ( 
.A(n_762),
.B(n_17),
.Y(n_1222)
);

OAI22x1_ASAP7_75t_SL g1223 ( 
.A1(n_943),
.A2(n_958),
.B1(n_984),
.B2(n_954),
.Y(n_1223)
);

NOR2xp33_ASAP7_75t_L g1224 ( 
.A(n_1092),
.B(n_18),
.Y(n_1224)
);

AND2x4_ASAP7_75t_L g1225 ( 
.A(n_818),
.B(n_19),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1036),
.Y(n_1226)
);

AND2x2_ASAP7_75t_L g1227 ( 
.A(n_828),
.B(n_19),
.Y(n_1227)
);

INVx2_ASAP7_75t_L g1228 ( 
.A(n_804),
.Y(n_1228)
);

AND2x2_ASAP7_75t_L g1229 ( 
.A(n_891),
.B(n_20),
.Y(n_1229)
);

NOR2x1_ASAP7_75t_L g1230 ( 
.A(n_1036),
.B(n_657),
.Y(n_1230)
);

OAI21x1_ASAP7_75t_L g1231 ( 
.A1(n_793),
.A2(n_659),
.B(n_658),
.Y(n_1231)
);

BUFx6f_ASAP7_75t_L g1232 ( 
.A(n_801),
.Y(n_1232)
);

OAI21x1_ASAP7_75t_L g1233 ( 
.A1(n_795),
.A2(n_662),
.B(n_661),
.Y(n_1233)
);

BUFx12f_ASAP7_75t_L g1234 ( 
.A(n_983),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1051),
.Y(n_1235)
);

HB1xp67_ASAP7_75t_L g1236 ( 
.A(n_948),
.Y(n_1236)
);

INVx2_ASAP7_75t_L g1237 ( 
.A(n_804),
.Y(n_1237)
);

AND2x4_ASAP7_75t_L g1238 ( 
.A(n_1057),
.B(n_21),
.Y(n_1238)
);

INVx4_ASAP7_75t_L g1239 ( 
.A(n_772),
.Y(n_1239)
);

INVx2_ASAP7_75t_L g1240 ( 
.A(n_804),
.Y(n_1240)
);

BUFx6f_ASAP7_75t_L g1241 ( 
.A(n_801),
.Y(n_1241)
);

OR2x2_ASAP7_75t_L g1242 ( 
.A(n_980),
.B(n_1022),
.Y(n_1242)
);

BUFx12f_ASAP7_75t_L g1243 ( 
.A(n_983),
.Y(n_1243)
);

BUFx3_ASAP7_75t_L g1244 ( 
.A(n_792),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1057),
.Y(n_1245)
);

INVx2_ASAP7_75t_L g1246 ( 
.A(n_804),
.Y(n_1246)
);

BUFx6f_ASAP7_75t_L g1247 ( 
.A(n_801),
.Y(n_1247)
);

BUFx8_ASAP7_75t_SL g1248 ( 
.A(n_958),
.Y(n_1248)
);

BUFx3_ASAP7_75t_L g1249 ( 
.A(n_817),
.Y(n_1249)
);

AND2x4_ASAP7_75t_L g1250 ( 
.A(n_1062),
.B(n_1114),
.Y(n_1250)
);

INVx5_ASAP7_75t_L g1251 ( 
.A(n_817),
.Y(n_1251)
);

BUFx6f_ASAP7_75t_L g1252 ( 
.A(n_809),
.Y(n_1252)
);

BUFx6f_ASAP7_75t_L g1253 ( 
.A(n_809),
.Y(n_1253)
);

AND2x2_ASAP7_75t_SL g1254 ( 
.A(n_850),
.B(n_663),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1062),
.Y(n_1255)
);

HB1xp67_ASAP7_75t_L g1256 ( 
.A(n_1063),
.Y(n_1256)
);

OA22x2_ASAP7_75t_SL g1257 ( 
.A1(n_845),
.A2(n_24),
.B1(n_22),
.B2(n_23),
.Y(n_1257)
);

INVx2_ASAP7_75t_L g1258 ( 
.A(n_804),
.Y(n_1258)
);

HB1xp67_ASAP7_75t_L g1259 ( 
.A(n_1177),
.Y(n_1259)
);

BUFx6f_ASAP7_75t_L g1260 ( 
.A(n_809),
.Y(n_1260)
);

BUFx6f_ASAP7_75t_L g1261 ( 
.A(n_809),
.Y(n_1261)
);

BUFx6f_ASAP7_75t_L g1262 ( 
.A(n_831),
.Y(n_1262)
);

INVx2_ASAP7_75t_L g1263 ( 
.A(n_869),
.Y(n_1263)
);

XNOR2x2_ASAP7_75t_L g1264 ( 
.A(n_765),
.B(n_22),
.Y(n_1264)
);

INVx2_ASAP7_75t_L g1265 ( 
.A(n_869),
.Y(n_1265)
);

INVx5_ASAP7_75t_L g1266 ( 
.A(n_849),
.Y(n_1266)
);

INVx3_ASAP7_75t_L g1267 ( 
.A(n_1007),
.Y(n_1267)
);

BUFx2_ASAP7_75t_L g1268 ( 
.A(n_1114),
.Y(n_1268)
);

BUFx3_ASAP7_75t_L g1269 ( 
.A(n_849),
.Y(n_1269)
);

INVx2_ASAP7_75t_L g1270 ( 
.A(n_869),
.Y(n_1270)
);

INVx3_ASAP7_75t_L g1271 ( 
.A(n_1007),
.Y(n_1271)
);

BUFx6f_ASAP7_75t_L g1272 ( 
.A(n_831),
.Y(n_1272)
);

INVx2_ASAP7_75t_L g1273 ( 
.A(n_869),
.Y(n_1273)
);

INVx2_ASAP7_75t_L g1274 ( 
.A(n_869),
.Y(n_1274)
);

BUFx12f_ASAP7_75t_L g1275 ( 
.A(n_1007),
.Y(n_1275)
);

INVx2_ASAP7_75t_L g1276 ( 
.A(n_869),
.Y(n_1276)
);

AND2x2_ASAP7_75t_L g1277 ( 
.A(n_1033),
.B(n_1050),
.Y(n_1277)
);

INVx2_ASAP7_75t_L g1278 ( 
.A(n_869),
.Y(n_1278)
);

OA21x2_ASAP7_75t_L g1279 ( 
.A1(n_824),
.A2(n_666),
.B(n_664),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_L g1280 ( 
.A(n_1148),
.B(n_25),
.Y(n_1280)
);

BUFx6f_ASAP7_75t_L g1281 ( 
.A(n_831),
.Y(n_1281)
);

INVx2_ASAP7_75t_L g1282 ( 
.A(n_1173),
.Y(n_1282)
);

AND2x4_ASAP7_75t_L g1283 ( 
.A(n_1145),
.B(n_25),
.Y(n_1283)
);

BUFx6f_ASAP7_75t_L g1284 ( 
.A(n_831),
.Y(n_1284)
);

INVx2_ASAP7_75t_L g1285 ( 
.A(n_1173),
.Y(n_1285)
);

AND2x2_ASAP7_75t_L g1286 ( 
.A(n_1033),
.B(n_26),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1145),
.Y(n_1287)
);

INVx4_ASAP7_75t_L g1288 ( 
.A(n_779),
.Y(n_1288)
);

BUFx8_ASAP7_75t_SL g1289 ( 
.A(n_984),
.Y(n_1289)
);

INVx6_ASAP7_75t_L g1290 ( 
.A(n_1033),
.Y(n_1290)
);

OAI21x1_ASAP7_75t_L g1291 ( 
.A1(n_855),
.A2(n_669),
.B(n_668),
.Y(n_1291)
);

BUFx8_ASAP7_75t_SL g1292 ( 
.A(n_1003),
.Y(n_1292)
);

BUFx12f_ASAP7_75t_L g1293 ( 
.A(n_1050),
.Y(n_1293)
);

AND2x4_ASAP7_75t_L g1294 ( 
.A(n_748),
.B(n_27),
.Y(n_1294)
);

CKINVDCx5p33_ASAP7_75t_R g1295 ( 
.A(n_1187),
.Y(n_1295)
);

CKINVDCx5p33_ASAP7_75t_R g1296 ( 
.A(n_1187),
.Y(n_1296)
);

CKINVDCx5p33_ASAP7_75t_R g1297 ( 
.A(n_1218),
.Y(n_1297)
);

CKINVDCx5p33_ASAP7_75t_R g1298 ( 
.A(n_1218),
.Y(n_1298)
);

CKINVDCx5p33_ASAP7_75t_R g1299 ( 
.A(n_1248),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1294),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_SL g1301 ( 
.A(n_1199),
.B(n_791),
.Y(n_1301)
);

CKINVDCx5p33_ASAP7_75t_R g1302 ( 
.A(n_1248),
.Y(n_1302)
);

CKINVDCx5p33_ASAP7_75t_R g1303 ( 
.A(n_1289),
.Y(n_1303)
);

CKINVDCx5p33_ASAP7_75t_R g1304 ( 
.A(n_1289),
.Y(n_1304)
);

CKINVDCx20_ASAP7_75t_R g1305 ( 
.A(n_1292),
.Y(n_1305)
);

AOI22xp5_ASAP7_75t_L g1306 ( 
.A1(n_1254),
.A2(n_885),
.B1(n_1113),
.B2(n_758),
.Y(n_1306)
);

AOI22xp5_ASAP7_75t_L g1307 ( 
.A1(n_1254),
.A2(n_885),
.B1(n_1113),
.B2(n_758),
.Y(n_1307)
);

CKINVDCx5p33_ASAP7_75t_R g1308 ( 
.A(n_1292),
.Y(n_1308)
);

CKINVDCx5p33_ASAP7_75t_R g1309 ( 
.A(n_1211),
.Y(n_1309)
);

CKINVDCx5p33_ASAP7_75t_R g1310 ( 
.A(n_1211),
.Y(n_1310)
);

HB1xp67_ASAP7_75t_L g1311 ( 
.A(n_1216),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1197),
.Y(n_1312)
);

CKINVDCx5p33_ASAP7_75t_R g1313 ( 
.A(n_1193),
.Y(n_1313)
);

CKINVDCx5p33_ASAP7_75t_R g1314 ( 
.A(n_1194),
.Y(n_1314)
);

CKINVDCx5p33_ASAP7_75t_R g1315 ( 
.A(n_1220),
.Y(n_1315)
);

AND3x2_ASAP7_75t_L g1316 ( 
.A(n_1196),
.B(n_908),
.C(n_776),
.Y(n_1316)
);

INVx2_ASAP7_75t_L g1317 ( 
.A(n_1250),
.Y(n_1317)
);

CKINVDCx5p33_ASAP7_75t_R g1318 ( 
.A(n_1234),
.Y(n_1318)
);

XNOR2xp5_ASAP7_75t_L g1319 ( 
.A(n_1181),
.B(n_1003),
.Y(n_1319)
);

INVx2_ASAP7_75t_L g1320 ( 
.A(n_1250),
.Y(n_1320)
);

CKINVDCx20_ASAP7_75t_R g1321 ( 
.A(n_1202),
.Y(n_1321)
);

CKINVDCx5p33_ASAP7_75t_R g1322 ( 
.A(n_1243),
.Y(n_1322)
);

CKINVDCx5p33_ASAP7_75t_R g1323 ( 
.A(n_1275),
.Y(n_1323)
);

NOR2xp33_ASAP7_75t_R g1324 ( 
.A(n_1293),
.B(n_1109),
.Y(n_1324)
);

CKINVDCx5p33_ASAP7_75t_R g1325 ( 
.A(n_1202),
.Y(n_1325)
);

AO21x2_ASAP7_75t_L g1326 ( 
.A1(n_1189),
.A2(n_862),
.B(n_857),
.Y(n_1326)
);

CKINVDCx5p33_ASAP7_75t_R g1327 ( 
.A(n_1217),
.Y(n_1327)
);

CKINVDCx5p33_ASAP7_75t_R g1328 ( 
.A(n_1217),
.Y(n_1328)
);

HB1xp67_ASAP7_75t_L g1329 ( 
.A(n_1216),
.Y(n_1329)
);

BUFx2_ASAP7_75t_L g1330 ( 
.A(n_1236),
.Y(n_1330)
);

CKINVDCx5p33_ASAP7_75t_R g1331 ( 
.A(n_1239),
.Y(n_1331)
);

CKINVDCx20_ASAP7_75t_R g1332 ( 
.A(n_1236),
.Y(n_1332)
);

NOR2xp33_ASAP7_75t_R g1333 ( 
.A(n_1199),
.B(n_1109),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1225),
.Y(n_1334)
);

AND2x2_ASAP7_75t_L g1335 ( 
.A(n_1256),
.B(n_1050),
.Y(n_1335)
);

BUFx6f_ASAP7_75t_L g1336 ( 
.A(n_1195),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1225),
.Y(n_1337)
);

CKINVDCx5p33_ASAP7_75t_R g1338 ( 
.A(n_1239),
.Y(n_1338)
);

CKINVDCx5p33_ASAP7_75t_R g1339 ( 
.A(n_1288),
.Y(n_1339)
);

HB1xp67_ASAP7_75t_L g1340 ( 
.A(n_1256),
.Y(n_1340)
);

OAI22xp5_ASAP7_75t_SL g1341 ( 
.A1(n_1190),
.A2(n_1039),
.B1(n_1049),
.B2(n_1026),
.Y(n_1341)
);

CKINVDCx20_ASAP7_75t_R g1342 ( 
.A(n_1259),
.Y(n_1342)
);

NOR2xp33_ASAP7_75t_R g1343 ( 
.A(n_1267),
.B(n_1124),
.Y(n_1343)
);

CKINVDCx5p33_ASAP7_75t_R g1344 ( 
.A(n_1288),
.Y(n_1344)
);

BUFx3_ASAP7_75t_L g1345 ( 
.A(n_1183),
.Y(n_1345)
);

CKINVDCx5p33_ASAP7_75t_R g1346 ( 
.A(n_1223),
.Y(n_1346)
);

CKINVDCx5p33_ASAP7_75t_R g1347 ( 
.A(n_1290),
.Y(n_1347)
);

CKINVDCx5p33_ASAP7_75t_R g1348 ( 
.A(n_1290),
.Y(n_1348)
);

BUFx6f_ASAP7_75t_L g1349 ( 
.A(n_1195),
.Y(n_1349)
);

CKINVDCx5p33_ASAP7_75t_R g1350 ( 
.A(n_1290),
.Y(n_1350)
);

CKINVDCx5p33_ASAP7_75t_R g1351 ( 
.A(n_1259),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_L g1352 ( 
.A(n_1277),
.B(n_1268),
.Y(n_1352)
);

HB1xp67_ASAP7_75t_L g1353 ( 
.A(n_1191),
.Y(n_1353)
);

XOR2x2_ASAP7_75t_L g1354 ( 
.A(n_1190),
.B(n_771),
.Y(n_1354)
);

INVx2_ASAP7_75t_L g1355 ( 
.A(n_1183),
.Y(n_1355)
);

CKINVDCx20_ASAP7_75t_R g1356 ( 
.A(n_1209),
.Y(n_1356)
);

NOR2xp67_ASAP7_75t_L g1357 ( 
.A(n_1267),
.B(n_1271),
.Y(n_1357)
);

CKINVDCx5p33_ASAP7_75t_R g1358 ( 
.A(n_1271),
.Y(n_1358)
);

OAI22xp33_ASAP7_75t_L g1359 ( 
.A1(n_1203),
.A2(n_1039),
.B1(n_1049),
.B2(n_1026),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1238),
.Y(n_1360)
);

CKINVDCx5p33_ASAP7_75t_R g1361 ( 
.A(n_1242),
.Y(n_1361)
);

CKINVDCx20_ASAP7_75t_R g1362 ( 
.A(n_1286),
.Y(n_1362)
);

INVx2_ASAP7_75t_L g1363 ( 
.A(n_1244),
.Y(n_1363)
);

CKINVDCx5p33_ASAP7_75t_R g1364 ( 
.A(n_1186),
.Y(n_1364)
);

CKINVDCx5p33_ASAP7_75t_R g1365 ( 
.A(n_1212),
.Y(n_1365)
);

CKINVDCx16_ASAP7_75t_R g1366 ( 
.A(n_1196),
.Y(n_1366)
);

CKINVDCx5p33_ASAP7_75t_R g1367 ( 
.A(n_1227),
.Y(n_1367)
);

CKINVDCx5p33_ASAP7_75t_R g1368 ( 
.A(n_1229),
.Y(n_1368)
);

CKINVDCx20_ASAP7_75t_R g1369 ( 
.A(n_1203),
.Y(n_1369)
);

INVx3_ASAP7_75t_L g1370 ( 
.A(n_1283),
.Y(n_1370)
);

CKINVDCx20_ASAP7_75t_R g1371 ( 
.A(n_1244),
.Y(n_1371)
);

CKINVDCx5p33_ASAP7_75t_R g1372 ( 
.A(n_1264),
.Y(n_1372)
);

INVx2_ASAP7_75t_L g1373 ( 
.A(n_1249),
.Y(n_1373)
);

CKINVDCx20_ASAP7_75t_R g1374 ( 
.A(n_1249),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1283),
.Y(n_1375)
);

NOR2xp33_ASAP7_75t_R g1376 ( 
.A(n_1269),
.B(n_1124),
.Y(n_1376)
);

CKINVDCx5p33_ASAP7_75t_R g1377 ( 
.A(n_1269),
.Y(n_1377)
);

NAND2xp5_ASAP7_75t_L g1378 ( 
.A(n_1213),
.B(n_1169),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1204),
.Y(n_1379)
);

NOR2xp33_ASAP7_75t_R g1380 ( 
.A(n_1210),
.B(n_814),
.Y(n_1380)
);

CKINVDCx20_ASAP7_75t_R g1381 ( 
.A(n_1222),
.Y(n_1381)
);

CKINVDCx5p33_ASAP7_75t_R g1382 ( 
.A(n_1213),
.Y(n_1382)
);

CKINVDCx5p33_ASAP7_75t_R g1383 ( 
.A(n_1213),
.Y(n_1383)
);

CKINVDCx5p33_ASAP7_75t_R g1384 ( 
.A(n_1213),
.Y(n_1384)
);

CKINVDCx5p33_ASAP7_75t_R g1385 ( 
.A(n_1224),
.Y(n_1385)
);

HB1xp67_ASAP7_75t_L g1386 ( 
.A(n_1188),
.Y(n_1386)
);

NOR2xp33_ASAP7_75t_R g1387 ( 
.A(n_1221),
.B(n_834),
.Y(n_1387)
);

INVx2_ASAP7_75t_L g1388 ( 
.A(n_1185),
.Y(n_1388)
);

CKINVDCx5p33_ASAP7_75t_R g1389 ( 
.A(n_1224),
.Y(n_1389)
);

CKINVDCx5p33_ASAP7_75t_R g1390 ( 
.A(n_1184),
.Y(n_1390)
);

CKINVDCx5p33_ASAP7_75t_R g1391 ( 
.A(n_1184),
.Y(n_1391)
);

CKINVDCx5p33_ASAP7_75t_R g1392 ( 
.A(n_1188),
.Y(n_1392)
);

CKINVDCx5p33_ASAP7_75t_R g1393 ( 
.A(n_1215),
.Y(n_1393)
);

CKINVDCx5p33_ASAP7_75t_R g1394 ( 
.A(n_1219),
.Y(n_1394)
);

CKINVDCx20_ASAP7_75t_R g1395 ( 
.A(n_1222),
.Y(n_1395)
);

CKINVDCx5p33_ASAP7_75t_R g1396 ( 
.A(n_1280),
.Y(n_1396)
);

NAND2xp33_ASAP7_75t_SL g1397 ( 
.A(n_1280),
.B(n_1080),
.Y(n_1397)
);

CKINVDCx5p33_ASAP7_75t_R g1398 ( 
.A(n_1226),
.Y(n_1398)
);

NOR2xp33_ASAP7_75t_R g1399 ( 
.A(n_1235),
.B(n_1245),
.Y(n_1399)
);

CKINVDCx5p33_ASAP7_75t_R g1400 ( 
.A(n_1255),
.Y(n_1400)
);

CKINVDCx5p33_ASAP7_75t_R g1401 ( 
.A(n_1287),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1192),
.Y(n_1402)
);

CKINVDCx5p33_ASAP7_75t_R g1403 ( 
.A(n_1198),
.Y(n_1403)
);

CKINVDCx5p33_ASAP7_75t_R g1404 ( 
.A(n_1228),
.Y(n_1404)
);

XOR2xp5_ASAP7_75t_L g1405 ( 
.A(n_1257),
.B(n_1080),
.Y(n_1405)
);

INVx2_ASAP7_75t_L g1406 ( 
.A(n_1237),
.Y(n_1406)
);

CKINVDCx5p33_ASAP7_75t_R g1407 ( 
.A(n_1246),
.Y(n_1407)
);

CKINVDCx5p33_ASAP7_75t_R g1408 ( 
.A(n_1263),
.Y(n_1408)
);

NOR2xp67_ASAP7_75t_L g1409 ( 
.A(n_1251),
.B(n_992),
.Y(n_1409)
);

CKINVDCx5p33_ASAP7_75t_R g1410 ( 
.A(n_1265),
.Y(n_1410)
);

CKINVDCx5p33_ASAP7_75t_R g1411 ( 
.A(n_1274),
.Y(n_1411)
);

CKINVDCx5p33_ASAP7_75t_R g1412 ( 
.A(n_1276),
.Y(n_1412)
);

CKINVDCx5p33_ASAP7_75t_R g1413 ( 
.A(n_1278),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1282),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1285),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_L g1416 ( 
.A(n_1251),
.B(n_1179),
.Y(n_1416)
);

NOR2xp67_ASAP7_75t_L g1417 ( 
.A(n_1251),
.B(n_998),
.Y(n_1417)
);

CKINVDCx20_ASAP7_75t_R g1418 ( 
.A(n_1257),
.Y(n_1418)
);

CKINVDCx5p33_ASAP7_75t_R g1419 ( 
.A(n_1200),
.Y(n_1419)
);

CKINVDCx5p33_ASAP7_75t_R g1420 ( 
.A(n_1200),
.Y(n_1420)
);

HB1xp67_ASAP7_75t_L g1421 ( 
.A(n_1214),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1240),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1240),
.Y(n_1423)
);

INVx2_ASAP7_75t_L g1424 ( 
.A(n_1258),
.Y(n_1424)
);

BUFx10_ASAP7_75t_L g1425 ( 
.A(n_1207),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1258),
.Y(n_1426)
);

CKINVDCx5p33_ASAP7_75t_R g1427 ( 
.A(n_1270),
.Y(n_1427)
);

NOR2xp33_ASAP7_75t_R g1428 ( 
.A(n_1251),
.B(n_878),
.Y(n_1428)
);

OA21x2_ASAP7_75t_L g1429 ( 
.A1(n_1231),
.A2(n_962),
.B(n_923),
.Y(n_1429)
);

CKINVDCx5p33_ASAP7_75t_R g1430 ( 
.A(n_1273),
.Y(n_1430)
);

BUFx6f_ASAP7_75t_L g1431 ( 
.A(n_1195),
.Y(n_1431)
);

NAND2xp33_ASAP7_75t_R g1432 ( 
.A(n_1279),
.B(n_740),
.Y(n_1432)
);

NOR2xp33_ASAP7_75t_R g1433 ( 
.A(n_1266),
.B(n_884),
.Y(n_1433)
);

CKINVDCx5p33_ASAP7_75t_R g1434 ( 
.A(n_1266),
.Y(n_1434)
);

CKINVDCx5p33_ASAP7_75t_R g1435 ( 
.A(n_1266),
.Y(n_1435)
);

NOR2xp33_ASAP7_75t_R g1436 ( 
.A(n_1205),
.B(n_886),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1208),
.Y(n_1437)
);

CKINVDCx5p33_ASAP7_75t_R g1438 ( 
.A(n_1205),
.Y(n_1438)
);

NAND2xp5_ASAP7_75t_L g1439 ( 
.A(n_1230),
.B(n_1166),
.Y(n_1439)
);

CKINVDCx5p33_ASAP7_75t_R g1440 ( 
.A(n_1207),
.Y(n_1440)
);

INVx2_ASAP7_75t_L g1441 ( 
.A(n_1207),
.Y(n_1441)
);

CKINVDCx5p33_ASAP7_75t_R g1442 ( 
.A(n_1232),
.Y(n_1442)
);

CKINVDCx5p33_ASAP7_75t_R g1443 ( 
.A(n_1232),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1233),
.Y(n_1444)
);

NOR2xp33_ASAP7_75t_R g1445 ( 
.A(n_1232),
.B(n_892),
.Y(n_1445)
);

INVx1_ASAP7_75t_SL g1446 ( 
.A(n_1182),
.Y(n_1446)
);

INVx2_ASAP7_75t_L g1447 ( 
.A(n_1241),
.Y(n_1447)
);

INVx2_ASAP7_75t_L g1448 ( 
.A(n_1241),
.Y(n_1448)
);

CKINVDCx5p33_ASAP7_75t_R g1449 ( 
.A(n_1241),
.Y(n_1449)
);

BUFx3_ASAP7_75t_L g1450 ( 
.A(n_1291),
.Y(n_1450)
);

NOR2xp33_ASAP7_75t_R g1451 ( 
.A(n_1247),
.B(n_918),
.Y(n_1451)
);

BUFx3_ASAP7_75t_L g1452 ( 
.A(n_1182),
.Y(n_1452)
);

CKINVDCx5p33_ASAP7_75t_R g1453 ( 
.A(n_1247),
.Y(n_1453)
);

CKINVDCx5p33_ASAP7_75t_R g1454 ( 
.A(n_1247),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1252),
.Y(n_1455)
);

CKINVDCx20_ASAP7_75t_R g1456 ( 
.A(n_1279),
.Y(n_1456)
);

CKINVDCx16_ASAP7_75t_R g1457 ( 
.A(n_1252),
.Y(n_1457)
);

CKINVDCx5p33_ASAP7_75t_R g1458 ( 
.A(n_1253),
.Y(n_1458)
);

CKINVDCx5p33_ASAP7_75t_R g1459 ( 
.A(n_1253),
.Y(n_1459)
);

CKINVDCx5p33_ASAP7_75t_R g1460 ( 
.A(n_1253),
.Y(n_1460)
);

CKINVDCx5p33_ASAP7_75t_R g1461 ( 
.A(n_1260),
.Y(n_1461)
);

CKINVDCx20_ASAP7_75t_R g1462 ( 
.A(n_1260),
.Y(n_1462)
);

NAND2x1_ASAP7_75t_L g1463 ( 
.A(n_1201),
.B(n_976),
.Y(n_1463)
);

OA21x2_ASAP7_75t_L g1464 ( 
.A1(n_1201),
.A2(n_1016),
.B(n_978),
.Y(n_1464)
);

INVx2_ASAP7_75t_L g1465 ( 
.A(n_1261),
.Y(n_1465)
);

CKINVDCx5p33_ASAP7_75t_R g1466 ( 
.A(n_1261),
.Y(n_1466)
);

CKINVDCx20_ASAP7_75t_R g1467 ( 
.A(n_1261),
.Y(n_1467)
);

NOR2xp33_ASAP7_75t_R g1468 ( 
.A(n_1262),
.B(n_934),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1262),
.Y(n_1469)
);

INVx2_ASAP7_75t_L g1470 ( 
.A(n_1262),
.Y(n_1470)
);

INVx2_ASAP7_75t_L g1471 ( 
.A(n_1272),
.Y(n_1471)
);

CKINVDCx5p33_ASAP7_75t_R g1472 ( 
.A(n_1272),
.Y(n_1472)
);

CKINVDCx20_ASAP7_75t_R g1473 ( 
.A(n_1272),
.Y(n_1473)
);

CKINVDCx5p33_ASAP7_75t_R g1474 ( 
.A(n_1281),
.Y(n_1474)
);

INVx4_ASAP7_75t_L g1475 ( 
.A(n_1201),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1284),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1284),
.B(n_1139),
.Y(n_1477)
);

BUFx6f_ASAP7_75t_SL g1478 ( 
.A(n_1206),
.Y(n_1478)
);

INVxp67_ASAP7_75t_SL g1479 ( 
.A(n_1206),
.Y(n_1479)
);

CKINVDCx5p33_ASAP7_75t_R g1480 ( 
.A(n_1206),
.Y(n_1480)
);

HB1xp67_ASAP7_75t_L g1481 ( 
.A(n_1216),
.Y(n_1481)
);

XNOR2xp5_ASAP7_75t_L g1482 ( 
.A(n_1306),
.B(n_1088),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1386),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1386),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_SL g1485 ( 
.A(n_1392),
.B(n_945),
.Y(n_1485)
);

NOR2xp33_ASAP7_75t_L g1486 ( 
.A(n_1352),
.B(n_1327),
.Y(n_1486)
);

BUFx6f_ASAP7_75t_L g1487 ( 
.A(n_1452),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_L g1488 ( 
.A(n_1393),
.B(n_950),
.Y(n_1488)
);

NAND2xp33_ASAP7_75t_L g1489 ( 
.A(n_1444),
.B(n_1394),
.Y(n_1489)
);

NOR2xp33_ASAP7_75t_L g1490 ( 
.A(n_1328),
.B(n_744),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_L g1491 ( 
.A(n_1396),
.B(n_960),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1317),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1320),
.Y(n_1493)
);

INVx2_ASAP7_75t_L g1494 ( 
.A(n_1355),
.Y(n_1494)
);

NOR3xp33_ASAP7_75t_L g1495 ( 
.A(n_1359),
.B(n_1086),
.C(n_1042),
.Y(n_1495)
);

NAND2xp5_ASAP7_75t_SL g1496 ( 
.A(n_1377),
.B(n_964),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1370),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_SL g1498 ( 
.A(n_1331),
.B(n_979),
.Y(n_1498)
);

BUFx8_ASAP7_75t_L g1499 ( 
.A(n_1330),
.Y(n_1499)
);

NOR2xp33_ASAP7_75t_L g1500 ( 
.A(n_1338),
.B(n_861),
.Y(n_1500)
);

NAND2xp5_ASAP7_75t_L g1501 ( 
.A(n_1353),
.B(n_1013),
.Y(n_1501)
);

INVx8_ASAP7_75t_L g1502 ( 
.A(n_1371),
.Y(n_1502)
);

NAND2xp5_ASAP7_75t_SL g1503 ( 
.A(n_1339),
.B(n_1027),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1477),
.Y(n_1504)
);

NOR3xp33_ASAP7_75t_L g1505 ( 
.A(n_1359),
.B(n_839),
.C(n_827),
.Y(n_1505)
);

NAND2xp5_ASAP7_75t_L g1506 ( 
.A(n_1353),
.B(n_1335),
.Y(n_1506)
);

NAND2xp5_ASAP7_75t_SL g1507 ( 
.A(n_1344),
.B(n_1029),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_L g1508 ( 
.A(n_1419),
.B(n_1067),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1379),
.Y(n_1509)
);

INVxp67_ASAP7_75t_L g1510 ( 
.A(n_1481),
.Y(n_1510)
);

NOR3xp33_ASAP7_75t_L g1511 ( 
.A(n_1341),
.B(n_924),
.C(n_871),
.Y(n_1511)
);

HB1xp67_ASAP7_75t_L g1512 ( 
.A(n_1332),
.Y(n_1512)
);

NAND2xp5_ASAP7_75t_SL g1513 ( 
.A(n_1385),
.B(n_1075),
.Y(n_1513)
);

AO221x1_ASAP7_75t_L g1514 ( 
.A1(n_1376),
.A2(n_1132),
.B1(n_1151),
.B2(n_1117),
.C(n_1088),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1312),
.Y(n_1515)
);

NOR2xp33_ASAP7_75t_SL g1516 ( 
.A(n_1366),
.B(n_1117),
.Y(n_1516)
);

NOR3xp33_ASAP7_75t_L g1517 ( 
.A(n_1397),
.B(n_1361),
.C(n_1372),
.Y(n_1517)
);

INVx2_ASAP7_75t_L g1518 ( 
.A(n_1363),
.Y(n_1518)
);

BUFx3_ASAP7_75t_L g1519 ( 
.A(n_1462),
.Y(n_1519)
);

INVx3_ASAP7_75t_L g1520 ( 
.A(n_1345),
.Y(n_1520)
);

NAND2xp5_ASAP7_75t_SL g1521 ( 
.A(n_1389),
.B(n_1076),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_L g1522 ( 
.A(n_1420),
.B(n_1094),
.Y(n_1522)
);

INVx2_ASAP7_75t_L g1523 ( 
.A(n_1373),
.Y(n_1523)
);

NOR2xp67_ASAP7_75t_L g1524 ( 
.A(n_1313),
.B(n_29),
.Y(n_1524)
);

NOR2xp33_ASAP7_75t_L g1525 ( 
.A(n_1358),
.B(n_863),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1334),
.Y(n_1526)
);

BUFx6f_ASAP7_75t_L g1527 ( 
.A(n_1450),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1427),
.B(n_1430),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_SL g1529 ( 
.A(n_1333),
.B(n_1131),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1337),
.Y(n_1530)
);

INVx2_ASAP7_75t_L g1531 ( 
.A(n_1421),
.Y(n_1531)
);

NOR3xp33_ASAP7_75t_L g1532 ( 
.A(n_1307),
.B(n_939),
.C(n_930),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1360),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1375),
.Y(n_1534)
);

INVx2_ASAP7_75t_L g1535 ( 
.A(n_1425),
.Y(n_1535)
);

XOR2xp5_ASAP7_75t_L g1536 ( 
.A(n_1342),
.B(n_1132),
.Y(n_1536)
);

INVx2_ASAP7_75t_L g1537 ( 
.A(n_1425),
.Y(n_1537)
);

NAND2xp33_ASAP7_75t_L g1538 ( 
.A(n_1456),
.B(n_1178),
.Y(n_1538)
);

NAND3xp33_ASAP7_75t_L g1539 ( 
.A(n_1365),
.B(n_747),
.C(n_741),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1300),
.Y(n_1540)
);

INVx2_ASAP7_75t_L g1541 ( 
.A(n_1429),
.Y(n_1541)
);

NOR2xp33_ASAP7_75t_L g1542 ( 
.A(n_1301),
.B(n_1017),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_L g1543 ( 
.A(n_1404),
.B(n_1173),
.Y(n_1543)
);

NOR2xp33_ASAP7_75t_L g1544 ( 
.A(n_1347),
.B(n_1030),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_SL g1545 ( 
.A(n_1348),
.B(n_1031),
.Y(n_1545)
);

INVx2_ASAP7_75t_L g1546 ( 
.A(n_1429),
.Y(n_1546)
);

NOR2xp33_ASAP7_75t_L g1547 ( 
.A(n_1350),
.B(n_1037),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_SL g1548 ( 
.A(n_1399),
.B(n_1098),
.Y(n_1548)
);

OR2x2_ASAP7_75t_L g1549 ( 
.A(n_1311),
.B(n_949),
.Y(n_1549)
);

NAND3xp33_ASAP7_75t_L g1550 ( 
.A(n_1367),
.B(n_1368),
.C(n_1364),
.Y(n_1550)
);

INVxp33_ASAP7_75t_L g1551 ( 
.A(n_1481),
.Y(n_1551)
);

INVx2_ASAP7_75t_L g1552 ( 
.A(n_1326),
.Y(n_1552)
);

NOR2xp33_ASAP7_75t_L g1553 ( 
.A(n_1398),
.B(n_1134),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1357),
.Y(n_1554)
);

NOR3xp33_ASAP7_75t_L g1555 ( 
.A(n_1403),
.B(n_993),
.C(n_988),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1407),
.B(n_1174),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_SL g1557 ( 
.A(n_1390),
.B(n_1142),
.Y(n_1557)
);

NOR2xp33_ASAP7_75t_L g1558 ( 
.A(n_1400),
.B(n_1153),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_L g1559 ( 
.A(n_1408),
.B(n_1174),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_L g1560 ( 
.A(n_1410),
.B(n_1174),
.Y(n_1560)
);

AND2x6_ASAP7_75t_L g1561 ( 
.A(n_1446),
.B(n_1081),
.Y(n_1561)
);

INVx1_ASAP7_75t_SL g1562 ( 
.A(n_1351),
.Y(n_1562)
);

NAND3xp33_ASAP7_75t_L g1563 ( 
.A(n_1311),
.B(n_755),
.C(n_752),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_L g1564 ( 
.A(n_1411),
.B(n_1174),
.Y(n_1564)
);

INVx2_ASAP7_75t_L g1565 ( 
.A(n_1326),
.Y(n_1565)
);

HB1xp67_ASAP7_75t_L g1566 ( 
.A(n_1329),
.Y(n_1566)
);

BUFx6f_ASAP7_75t_SL g1567 ( 
.A(n_1437),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_L g1568 ( 
.A(n_1412),
.B(n_1174),
.Y(n_1568)
);

NOR2xp33_ASAP7_75t_L g1569 ( 
.A(n_1401),
.B(n_756),
.Y(n_1569)
);

AOI22xp5_ASAP7_75t_L g1570 ( 
.A1(n_1329),
.A2(n_1180),
.B1(n_760),
.B2(n_763),
.Y(n_1570)
);

BUFx2_ASAP7_75t_R g1571 ( 
.A(n_1295),
.Y(n_1571)
);

INVx2_ASAP7_75t_L g1572 ( 
.A(n_1475),
.Y(n_1572)
);

NOR2xp33_ASAP7_75t_L g1573 ( 
.A(n_1391),
.B(n_759),
.Y(n_1573)
);

NOR3xp33_ASAP7_75t_L g1574 ( 
.A(n_1340),
.B(n_1059),
.C(n_1024),
.Y(n_1574)
);

BUFx8_ASAP7_75t_L g1575 ( 
.A(n_1478),
.Y(n_1575)
);

INVx3_ASAP7_75t_L g1576 ( 
.A(n_1457),
.Y(n_1576)
);

NOR2xp33_ASAP7_75t_L g1577 ( 
.A(n_1340),
.B(n_764),
.Y(n_1577)
);

INVx2_ASAP7_75t_L g1578 ( 
.A(n_1475),
.Y(n_1578)
);

BUFx6f_ASAP7_75t_L g1579 ( 
.A(n_1464),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_L g1580 ( 
.A(n_1413),
.B(n_1174),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_SL g1581 ( 
.A(n_1380),
.B(n_848),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1409),
.Y(n_1582)
);

BUFx8_ASAP7_75t_L g1583 ( 
.A(n_1478),
.Y(n_1583)
);

NOR2xp33_ASAP7_75t_L g1584 ( 
.A(n_1378),
.B(n_766),
.Y(n_1584)
);

INVx4_ASAP7_75t_L g1585 ( 
.A(n_1316),
.Y(n_1585)
);

NOR2x1p5_ASAP7_75t_L g1586 ( 
.A(n_1325),
.B(n_1314),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_L g1587 ( 
.A(n_1439),
.B(n_768),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_L g1588 ( 
.A(n_1387),
.B(n_770),
.Y(n_1588)
);

INVx2_ASAP7_75t_L g1589 ( 
.A(n_1424),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_SL g1590 ( 
.A(n_1324),
.B(n_848),
.Y(n_1590)
);

INVx2_ASAP7_75t_L g1591 ( 
.A(n_1480),
.Y(n_1591)
);

INVx2_ASAP7_75t_L g1592 ( 
.A(n_1388),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_L g1593 ( 
.A(n_1382),
.B(n_773),
.Y(n_1593)
);

INVx3_ASAP7_75t_L g1594 ( 
.A(n_1463),
.Y(n_1594)
);

INVx2_ASAP7_75t_L g1595 ( 
.A(n_1406),
.Y(n_1595)
);

INVx2_ASAP7_75t_L g1596 ( 
.A(n_1440),
.Y(n_1596)
);

INVxp67_ASAP7_75t_L g1597 ( 
.A(n_1315),
.Y(n_1597)
);

INVxp33_ASAP7_75t_L g1598 ( 
.A(n_1343),
.Y(n_1598)
);

INVx2_ASAP7_75t_L g1599 ( 
.A(n_1442),
.Y(n_1599)
);

INVx2_ASAP7_75t_L g1600 ( 
.A(n_1443),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_L g1601 ( 
.A(n_1383),
.B(n_778),
.Y(n_1601)
);

INVxp67_ASAP7_75t_SL g1602 ( 
.A(n_1374),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_SL g1603 ( 
.A(n_1428),
.B(n_848),
.Y(n_1603)
);

INVx2_ASAP7_75t_L g1604 ( 
.A(n_1449),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1417),
.Y(n_1605)
);

INVx2_ASAP7_75t_SL g1606 ( 
.A(n_1316),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1384),
.B(n_780),
.Y(n_1607)
);

NOR2xp67_ASAP7_75t_L g1608 ( 
.A(n_1318),
.B(n_30),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_SL g1609 ( 
.A(n_1433),
.B(n_848),
.Y(n_1609)
);

NOR2xp33_ASAP7_75t_L g1610 ( 
.A(n_1356),
.B(n_782),
.Y(n_1610)
);

NOR2xp33_ASAP7_75t_L g1611 ( 
.A(n_1362),
.B(n_783),
.Y(n_1611)
);

INVx2_ASAP7_75t_L g1612 ( 
.A(n_1453),
.Y(n_1612)
);

INVx2_ASAP7_75t_L g1613 ( 
.A(n_1454),
.Y(n_1613)
);

INVx2_ASAP7_75t_L g1614 ( 
.A(n_1458),
.Y(n_1614)
);

NOR2xp33_ASAP7_75t_SL g1615 ( 
.A(n_1309),
.B(n_1151),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_SL g1616 ( 
.A(n_1416),
.B(n_894),
.Y(n_1616)
);

NOR2xp33_ASAP7_75t_L g1617 ( 
.A(n_1310),
.B(n_786),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_SL g1618 ( 
.A(n_1436),
.B(n_1381),
.Y(n_1618)
);

OAI22xp5_ASAP7_75t_L g1619 ( 
.A1(n_1395),
.A2(n_789),
.B1(n_790),
.B2(n_788),
.Y(n_1619)
);

NOR2xp33_ASAP7_75t_L g1620 ( 
.A(n_1322),
.B(n_800),
.Y(n_1620)
);

BUFx5_ASAP7_75t_L g1621 ( 
.A(n_1422),
.Y(n_1621)
);

NAND2xp33_ASAP7_75t_L g1622 ( 
.A(n_1434),
.B(n_894),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_L g1623 ( 
.A(n_1423),
.B(n_802),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_SL g1624 ( 
.A(n_1323),
.B(n_894),
.Y(n_1624)
);

NAND2xp33_ASAP7_75t_L g1625 ( 
.A(n_1435),
.B(n_894),
.Y(n_1625)
);

NOR2xp33_ASAP7_75t_L g1626 ( 
.A(n_1402),
.B(n_805),
.Y(n_1626)
);

HAxp5_ASAP7_75t_SL g1627 ( 
.A(n_1319),
.B(n_798),
.CON(n_1627),
.SN(n_1627)
);

NOR2xp33_ASAP7_75t_R g1628 ( 
.A(n_1321),
.B(n_819),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_L g1629 ( 
.A(n_1426),
.B(n_806),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1354),
.B(n_1139),
.Y(n_1630)
);

NOR3xp33_ASAP7_75t_L g1631 ( 
.A(n_1346),
.B(n_1072),
.C(n_1069),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1414),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_L g1633 ( 
.A(n_1415),
.B(n_810),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1467),
.Y(n_1634)
);

BUFx6f_ASAP7_75t_L g1635 ( 
.A(n_1464),
.Y(n_1635)
);

AOI221xp5_ASAP7_75t_L g1636 ( 
.A1(n_1405),
.A2(n_753),
.B1(n_757),
.B2(n_749),
.C(n_742),
.Y(n_1636)
);

NOR2xp33_ASAP7_75t_L g1637 ( 
.A(n_1473),
.B(n_820),
.Y(n_1637)
);

NOR2xp33_ASAP7_75t_L g1638 ( 
.A(n_1438),
.B(n_821),
.Y(n_1638)
);

INVx2_ASAP7_75t_L g1639 ( 
.A(n_1459),
.Y(n_1639)
);

AND2x2_ASAP7_75t_L g1640 ( 
.A(n_1369),
.B(n_1139),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_SL g1641 ( 
.A(n_1445),
.B(n_957),
.Y(n_1641)
);

OR2x2_ASAP7_75t_L g1642 ( 
.A(n_1296),
.B(n_1116),
.Y(n_1642)
);

INVx2_ASAP7_75t_SL g1643 ( 
.A(n_1451),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_L g1644 ( 
.A(n_1468),
.B(n_822),
.Y(n_1644)
);

INVx3_ASAP7_75t_R g1645 ( 
.A(n_1305),
.Y(n_1645)
);

CKINVDCx5p33_ASAP7_75t_R g1646 ( 
.A(n_1297),
.Y(n_1646)
);

INVx2_ASAP7_75t_L g1647 ( 
.A(n_1460),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_L g1648 ( 
.A(n_1461),
.B(n_826),
.Y(n_1648)
);

INVxp67_ASAP7_75t_L g1649 ( 
.A(n_1298),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1466),
.Y(n_1650)
);

INVx2_ASAP7_75t_L g1651 ( 
.A(n_1472),
.Y(n_1651)
);

BUFx6f_ASAP7_75t_L g1652 ( 
.A(n_1474),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1479),
.Y(n_1653)
);

INVx2_ASAP7_75t_SL g1654 ( 
.A(n_1299),
.Y(n_1654)
);

BUFx6f_ASAP7_75t_L g1655 ( 
.A(n_1336),
.Y(n_1655)
);

NAND2x1_ASAP7_75t_L g1656 ( 
.A(n_1455),
.B(n_750),
.Y(n_1656)
);

INVx5_ASAP7_75t_L g1657 ( 
.A(n_1336),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_L g1658 ( 
.A(n_1469),
.B(n_832),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_SL g1659 ( 
.A(n_1418),
.B(n_957),
.Y(n_1659)
);

NOR2xp33_ASAP7_75t_L g1660 ( 
.A(n_1302),
.B(n_835),
.Y(n_1660)
);

NOR3xp33_ASAP7_75t_L g1661 ( 
.A(n_1303),
.B(n_1133),
.C(n_838),
.Y(n_1661)
);

NAND2xp33_ASAP7_75t_L g1662 ( 
.A(n_1432),
.B(n_957),
.Y(n_1662)
);

INVx2_ASAP7_75t_L g1663 ( 
.A(n_1476),
.Y(n_1663)
);

AOI221xp5_ASAP7_75t_L g1664 ( 
.A1(n_1304),
.A2(n_777),
.B1(n_781),
.B2(n_769),
.C(n_761),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_L g1665 ( 
.A(n_1441),
.B(n_840),
.Y(n_1665)
);

NOR2xp33_ASAP7_75t_L g1666 ( 
.A(n_1308),
.B(n_842),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_L g1667 ( 
.A(n_1447),
.B(n_843),
.Y(n_1667)
);

INVxp33_ASAP7_75t_L g1668 ( 
.A(n_1471),
.Y(n_1668)
);

INVx2_ASAP7_75t_L g1669 ( 
.A(n_1448),
.Y(n_1669)
);

INVxp67_ASAP7_75t_SL g1670 ( 
.A(n_1336),
.Y(n_1670)
);

NAND2xp5_ASAP7_75t_L g1671 ( 
.A(n_1470),
.B(n_844),
.Y(n_1671)
);

NOR2xp33_ASAP7_75t_L g1672 ( 
.A(n_1465),
.B(n_851),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_L g1673 ( 
.A(n_1336),
.B(n_853),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_L g1674 ( 
.A(n_1349),
.B(n_854),
.Y(n_1674)
);

INVxp67_ASAP7_75t_L g1675 ( 
.A(n_1349),
.Y(n_1675)
);

OR2x6_ASAP7_75t_L g1676 ( 
.A(n_1349),
.B(n_1104),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_SL g1677 ( 
.A(n_1349),
.B(n_957),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_SL g1678 ( 
.A(n_1431),
.B(n_1052),
.Y(n_1678)
);

BUFx6f_ASAP7_75t_SL g1679 ( 
.A(n_1431),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_L g1680 ( 
.A(n_1431),
.B(n_858),
.Y(n_1680)
);

BUFx6f_ASAP7_75t_L g1681 ( 
.A(n_1431),
.Y(n_1681)
);

NAND2xp5_ASAP7_75t_L g1682 ( 
.A(n_1386),
.B(n_867),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1386),
.Y(n_1683)
);

INVx2_ASAP7_75t_L g1684 ( 
.A(n_1355),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_SL g1685 ( 
.A(n_1392),
.B(n_1052),
.Y(n_1685)
);

NAND2xp5_ASAP7_75t_L g1686 ( 
.A(n_1386),
.B(n_868),
.Y(n_1686)
);

INVx2_ASAP7_75t_L g1687 ( 
.A(n_1355),
.Y(n_1687)
);

NAND2xp33_ASAP7_75t_L g1688 ( 
.A(n_1444),
.B(n_1052),
.Y(n_1688)
);

BUFx6f_ASAP7_75t_L g1689 ( 
.A(n_1452),
.Y(n_1689)
);

INVx2_ASAP7_75t_L g1690 ( 
.A(n_1355),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_L g1691 ( 
.A(n_1386),
.B(n_870),
.Y(n_1691)
);

INVx2_ASAP7_75t_L g1692 ( 
.A(n_1355),
.Y(n_1692)
);

AND2x2_ASAP7_75t_L g1693 ( 
.A(n_1330),
.B(n_1141),
.Y(n_1693)
);

INVx2_ASAP7_75t_L g1694 ( 
.A(n_1355),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_L g1695 ( 
.A(n_1386),
.B(n_872),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1386),
.Y(n_1696)
);

NOR3xp33_ASAP7_75t_L g1697 ( 
.A(n_1359),
.B(n_876),
.C(n_875),
.Y(n_1697)
);

BUFx6f_ASAP7_75t_L g1698 ( 
.A(n_1452),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1386),
.Y(n_1699)
);

NOR2xp33_ASAP7_75t_L g1700 ( 
.A(n_1386),
.B(n_881),
.Y(n_1700)
);

AND2x2_ASAP7_75t_L g1701 ( 
.A(n_1330),
.B(n_1141),
.Y(n_1701)
);

INVxp67_ASAP7_75t_L g1702 ( 
.A(n_1330),
.Y(n_1702)
);

NOR2xp33_ASAP7_75t_L g1703 ( 
.A(n_1386),
.B(n_883),
.Y(n_1703)
);

INVx2_ASAP7_75t_L g1704 ( 
.A(n_1355),
.Y(n_1704)
);

INVx2_ASAP7_75t_L g1705 ( 
.A(n_1355),
.Y(n_1705)
);

NAND2xp5_ASAP7_75t_SL g1706 ( 
.A(n_1392),
.B(n_1052),
.Y(n_1706)
);

INVx2_ASAP7_75t_SL g1707 ( 
.A(n_1386),
.Y(n_1707)
);

NOR2xp33_ASAP7_75t_L g1708 ( 
.A(n_1386),
.B(n_888),
.Y(n_1708)
);

CKINVDCx5p33_ASAP7_75t_R g1709 ( 
.A(n_1332),
.Y(n_1709)
);

INVx2_ASAP7_75t_L g1710 ( 
.A(n_1355),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1386),
.Y(n_1711)
);

AND2x2_ASAP7_75t_L g1712 ( 
.A(n_1330),
.B(n_1141),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_L g1713 ( 
.A(n_1386),
.B(n_890),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_L g1714 ( 
.A(n_1386),
.B(n_895),
.Y(n_1714)
);

HB1xp67_ASAP7_75t_L g1715 ( 
.A(n_1332),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_L g1716 ( 
.A(n_1386),
.B(n_897),
.Y(n_1716)
);

NAND2xp5_ASAP7_75t_SL g1717 ( 
.A(n_1392),
.B(n_1077),
.Y(n_1717)
);

AOI22xp5_ASAP7_75t_L g1718 ( 
.A1(n_1392),
.A2(n_1167),
.B1(n_1168),
.B2(n_1165),
.Y(n_1718)
);

NAND3xp33_ASAP7_75t_L g1719 ( 
.A(n_1392),
.B(n_901),
.C(n_900),
.Y(n_1719)
);

INVxp67_ASAP7_75t_L g1720 ( 
.A(n_1330),
.Y(n_1720)
);

INVx2_ASAP7_75t_SL g1721 ( 
.A(n_1386),
.Y(n_1721)
);

BUFx6f_ASAP7_75t_SL g1722 ( 
.A(n_1437),
.Y(n_1722)
);

INVx2_ASAP7_75t_SL g1723 ( 
.A(n_1386),
.Y(n_1723)
);

INVx2_ASAP7_75t_L g1724 ( 
.A(n_1355),
.Y(n_1724)
);

BUFx6f_ASAP7_75t_L g1725 ( 
.A(n_1452),
.Y(n_1725)
);

NAND2xp5_ASAP7_75t_L g1726 ( 
.A(n_1386),
.B(n_902),
.Y(n_1726)
);

NAND2xp5_ASAP7_75t_L g1727 ( 
.A(n_1386),
.B(n_904),
.Y(n_1727)
);

NAND2xp5_ASAP7_75t_L g1728 ( 
.A(n_1386),
.B(n_905),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1386),
.Y(n_1729)
);

NAND2xp33_ASAP7_75t_L g1730 ( 
.A(n_1444),
.B(n_1077),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_L g1731 ( 
.A(n_1386),
.B(n_906),
.Y(n_1731)
);

INVxp67_ASAP7_75t_L g1732 ( 
.A(n_1330),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1386),
.Y(n_1733)
);

NAND2xp5_ASAP7_75t_SL g1734 ( 
.A(n_1392),
.B(n_1077),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1707),
.Y(n_1735)
);

INVx3_ASAP7_75t_L g1736 ( 
.A(n_1575),
.Y(n_1736)
);

OR2x2_ASAP7_75t_L g1737 ( 
.A(n_1562),
.B(n_913),
.Y(n_1737)
);

INVx1_ASAP7_75t_SL g1738 ( 
.A(n_1709),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1721),
.Y(n_1739)
);

BUFx3_ASAP7_75t_L g1740 ( 
.A(n_1575),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1723),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1531),
.Y(n_1742)
);

NAND2xp5_ASAP7_75t_L g1743 ( 
.A(n_1483),
.B(n_916),
.Y(n_1743)
);

NOR2xp33_ASAP7_75t_L g1744 ( 
.A(n_1551),
.B(n_829),
.Y(n_1744)
);

NOR2xp33_ASAP7_75t_L g1745 ( 
.A(n_1510),
.B(n_859),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1497),
.Y(n_1746)
);

OAI21xp33_ASAP7_75t_L g1747 ( 
.A1(n_1700),
.A2(n_1162),
.B(n_1161),
.Y(n_1747)
);

BUFx3_ASAP7_75t_L g1748 ( 
.A(n_1583),
.Y(n_1748)
);

BUFx8_ASAP7_75t_L g1749 ( 
.A(n_1654),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_L g1750 ( 
.A(n_1484),
.B(n_919),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1683),
.Y(n_1751)
);

NOR2xp33_ASAP7_75t_L g1752 ( 
.A(n_1702),
.B(n_873),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1696),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1699),
.Y(n_1754)
);

AND2x4_ASAP7_75t_L g1755 ( 
.A(n_1711),
.B(n_836),
.Y(n_1755)
);

NAND2xp5_ASAP7_75t_L g1756 ( 
.A(n_1729),
.B(n_920),
.Y(n_1756)
);

OR2x6_ASAP7_75t_L g1757 ( 
.A(n_1502),
.B(n_774),
.Y(n_1757)
);

AND2x2_ASAP7_75t_L g1758 ( 
.A(n_1566),
.B(n_1175),
.Y(n_1758)
);

AOI22xp33_ASAP7_75t_L g1759 ( 
.A1(n_1697),
.A2(n_784),
.B1(n_794),
.B2(n_785),
.Y(n_1759)
);

NAND2xp5_ASAP7_75t_L g1760 ( 
.A(n_1733),
.B(n_926),
.Y(n_1760)
);

CKINVDCx5p33_ASAP7_75t_R g1761 ( 
.A(n_1499),
.Y(n_1761)
);

INVx4_ASAP7_75t_L g1762 ( 
.A(n_1576),
.Y(n_1762)
);

AOI22xp5_ASAP7_75t_L g1763 ( 
.A1(n_1720),
.A2(n_927),
.B1(n_932),
.B2(n_929),
.Y(n_1763)
);

NAND2xp5_ASAP7_75t_L g1764 ( 
.A(n_1703),
.B(n_933),
.Y(n_1764)
);

OR2x6_ASAP7_75t_L g1765 ( 
.A(n_1502),
.B(n_816),
.Y(n_1765)
);

AND2x4_ASAP7_75t_L g1766 ( 
.A(n_1504),
.B(n_796),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_L g1767 ( 
.A(n_1708),
.B(n_935),
.Y(n_1767)
);

NAND2xp5_ASAP7_75t_L g1768 ( 
.A(n_1506),
.B(n_936),
.Y(n_1768)
);

OAI22xp5_ASAP7_75t_L g1769 ( 
.A1(n_1528),
.A2(n_1140),
.B1(n_797),
.B2(n_803),
.Y(n_1769)
);

OAI21xp5_ASAP7_75t_L g1770 ( 
.A1(n_1552),
.A2(n_1565),
.B(n_1546),
.Y(n_1770)
);

HB1xp67_ASAP7_75t_L g1771 ( 
.A(n_1512),
.Y(n_1771)
);

INVx3_ASAP7_75t_L g1772 ( 
.A(n_1583),
.Y(n_1772)
);

NAND2xp5_ASAP7_75t_L g1773 ( 
.A(n_1682),
.B(n_940),
.Y(n_1773)
);

INVxp67_ASAP7_75t_L g1774 ( 
.A(n_1715),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1509),
.Y(n_1775)
);

BUFx6f_ASAP7_75t_L g1776 ( 
.A(n_1487),
.Y(n_1776)
);

AOI21xp5_ASAP7_75t_L g1777 ( 
.A1(n_1541),
.A2(n_754),
.B(n_1081),
.Y(n_1777)
);

AND2x2_ASAP7_75t_L g1778 ( 
.A(n_1732),
.B(n_1175),
.Y(n_1778)
);

AND2x6_ASAP7_75t_L g1779 ( 
.A(n_1487),
.B(n_816),
.Y(n_1779)
);

NOR2xp33_ASAP7_75t_L g1780 ( 
.A(n_1486),
.B(n_941),
.Y(n_1780)
);

AOI22xp33_ASAP7_75t_L g1781 ( 
.A1(n_1532),
.A2(n_811),
.B1(n_812),
.B2(n_799),
.Y(n_1781)
);

NAND3xp33_ASAP7_75t_L g1782 ( 
.A(n_1610),
.B(n_947),
.C(n_942),
.Y(n_1782)
);

INVx2_ASAP7_75t_L g1783 ( 
.A(n_1621),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1492),
.Y(n_1784)
);

BUFx3_ASAP7_75t_L g1785 ( 
.A(n_1499),
.Y(n_1785)
);

NAND2xp5_ASAP7_75t_L g1786 ( 
.A(n_1686),
.B(n_951),
.Y(n_1786)
);

NAND2xp5_ASAP7_75t_L g1787 ( 
.A(n_1691),
.B(n_955),
.Y(n_1787)
);

CKINVDCx11_ASAP7_75t_R g1788 ( 
.A(n_1519),
.Y(n_1788)
);

INVx5_ASAP7_75t_L g1789 ( 
.A(n_1576),
.Y(n_1789)
);

AOI22xp33_ASAP7_75t_L g1790 ( 
.A1(n_1505),
.A2(n_823),
.B1(n_825),
.B2(n_813),
.Y(n_1790)
);

NAND2xp5_ASAP7_75t_SL g1791 ( 
.A(n_1585),
.B(n_959),
.Y(n_1791)
);

BUFx6f_ASAP7_75t_L g1792 ( 
.A(n_1487),
.Y(n_1792)
);

INVx2_ASAP7_75t_SL g1793 ( 
.A(n_1549),
.Y(n_1793)
);

AND2x6_ASAP7_75t_L g1794 ( 
.A(n_1689),
.B(n_865),
.Y(n_1794)
);

AOI22xp33_ASAP7_75t_SL g1795 ( 
.A1(n_1516),
.A2(n_1175),
.B1(n_961),
.B2(n_969),
.Y(n_1795)
);

NOR2xp33_ASAP7_75t_L g1796 ( 
.A(n_1693),
.B(n_963),
.Y(n_1796)
);

NOR2xp33_ASAP7_75t_L g1797 ( 
.A(n_1701),
.B(n_1712),
.Y(n_1797)
);

AND2x4_ASAP7_75t_L g1798 ( 
.A(n_1515),
.B(n_833),
.Y(n_1798)
);

NAND2xp5_ASAP7_75t_L g1799 ( 
.A(n_1695),
.B(n_973),
.Y(n_1799)
);

BUFx3_ASAP7_75t_L g1800 ( 
.A(n_1652),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1493),
.Y(n_1801)
);

INVxp67_ASAP7_75t_L g1802 ( 
.A(n_1536),
.Y(n_1802)
);

BUFx6f_ASAP7_75t_L g1803 ( 
.A(n_1689),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1540),
.Y(n_1804)
);

NAND3xp33_ASAP7_75t_SL g1805 ( 
.A(n_1628),
.B(n_1170),
.C(n_1163),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1526),
.Y(n_1806)
);

BUFx2_ASAP7_75t_L g1807 ( 
.A(n_1602),
.Y(n_1807)
);

NOR2xp33_ASAP7_75t_L g1808 ( 
.A(n_1550),
.B(n_982),
.Y(n_1808)
);

AOI221xp5_ASAP7_75t_L g1809 ( 
.A1(n_1495),
.A2(n_846),
.B1(n_847),
.B2(n_841),
.C(n_837),
.Y(n_1809)
);

INVx3_ASAP7_75t_L g1810 ( 
.A(n_1520),
.Y(n_1810)
);

NOR2xp33_ASAP7_75t_R g1811 ( 
.A(n_1646),
.B(n_985),
.Y(n_1811)
);

NOR2xp33_ASAP7_75t_L g1812 ( 
.A(n_1573),
.B(n_989),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1530),
.Y(n_1813)
);

AOI22xp5_ASAP7_75t_L g1814 ( 
.A1(n_1577),
.A2(n_996),
.B1(n_1000),
.B2(n_994),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1533),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1534),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_L g1817 ( 
.A(n_1713),
.B(n_1714),
.Y(n_1817)
);

BUFx6f_ASAP7_75t_L g1818 ( 
.A(n_1689),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1632),
.Y(n_1819)
);

CKINVDCx5p33_ASAP7_75t_R g1820 ( 
.A(n_1571),
.Y(n_1820)
);

NAND2xp5_ASAP7_75t_SL g1821 ( 
.A(n_1606),
.B(n_1002),
.Y(n_1821)
);

NAND2xp5_ASAP7_75t_L g1822 ( 
.A(n_1716),
.B(n_1004),
.Y(n_1822)
);

CKINVDCx20_ASAP7_75t_R g1823 ( 
.A(n_1645),
.Y(n_1823)
);

INVx2_ASAP7_75t_L g1824 ( 
.A(n_1494),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1554),
.Y(n_1825)
);

HB1xp67_ASAP7_75t_L g1826 ( 
.A(n_1652),
.Y(n_1826)
);

NAND2xp5_ASAP7_75t_L g1827 ( 
.A(n_1726),
.B(n_1006),
.Y(n_1827)
);

INVxp67_ASAP7_75t_L g1828 ( 
.A(n_1615),
.Y(n_1828)
);

OA22x2_ASAP7_75t_L g1829 ( 
.A1(n_1482),
.A2(n_1010),
.B1(n_1011),
.B2(n_1009),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1518),
.Y(n_1830)
);

AND2x4_ASAP7_75t_L g1831 ( 
.A(n_1719),
.B(n_852),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1523),
.Y(n_1832)
);

NAND2xp5_ASAP7_75t_L g1833 ( 
.A(n_1727),
.B(n_1014),
.Y(n_1833)
);

NAND2xp5_ASAP7_75t_L g1834 ( 
.A(n_1728),
.B(n_1015),
.Y(n_1834)
);

AND2x6_ASAP7_75t_L g1835 ( 
.A(n_1698),
.B(n_865),
.Y(n_1835)
);

NOR3xp33_ASAP7_75t_SL g1836 ( 
.A(n_1636),
.B(n_1021),
.C(n_1018),
.Y(n_1836)
);

NAND2xp33_ASAP7_75t_SL g1837 ( 
.A(n_1598),
.B(n_1155),
.Y(n_1837)
);

NOR2xp33_ASAP7_75t_L g1838 ( 
.A(n_1731),
.B(n_1023),
.Y(n_1838)
);

BUFx3_ASAP7_75t_L g1839 ( 
.A(n_1652),
.Y(n_1839)
);

INVx2_ASAP7_75t_L g1840 ( 
.A(n_1684),
.Y(n_1840)
);

BUFx6f_ASAP7_75t_L g1841 ( 
.A(n_1698),
.Y(n_1841)
);

INVx3_ASAP7_75t_L g1842 ( 
.A(n_1520),
.Y(n_1842)
);

BUFx2_ASAP7_75t_L g1843 ( 
.A(n_1597),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1687),
.Y(n_1844)
);

AND2x4_ASAP7_75t_L g1845 ( 
.A(n_1563),
.B(n_856),
.Y(n_1845)
);

INVx2_ASAP7_75t_SL g1846 ( 
.A(n_1634),
.Y(n_1846)
);

NAND2xp5_ASAP7_75t_SL g1847 ( 
.A(n_1725),
.B(n_1035),
.Y(n_1847)
);

INVx2_ASAP7_75t_L g1848 ( 
.A(n_1690),
.Y(n_1848)
);

AOI22xp33_ASAP7_75t_L g1849 ( 
.A1(n_1517),
.A2(n_864),
.B1(n_866),
.B2(n_860),
.Y(n_1849)
);

INVx2_ASAP7_75t_L g1850 ( 
.A(n_1692),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1694),
.Y(n_1851)
);

INVx2_ASAP7_75t_L g1852 ( 
.A(n_1704),
.Y(n_1852)
);

AOI22xp33_ASAP7_75t_L g1853 ( 
.A1(n_1538),
.A2(n_877),
.B1(n_880),
.B2(n_874),
.Y(n_1853)
);

NAND2xp5_ASAP7_75t_L g1854 ( 
.A(n_1501),
.B(n_1488),
.Y(n_1854)
);

AND2x4_ASAP7_75t_L g1855 ( 
.A(n_1485),
.B(n_1582),
.Y(n_1855)
);

INVx3_ASAP7_75t_L g1856 ( 
.A(n_1535),
.Y(n_1856)
);

NAND2xp5_ASAP7_75t_SL g1857 ( 
.A(n_1725),
.B(n_1041),
.Y(n_1857)
);

INVx2_ASAP7_75t_L g1858 ( 
.A(n_1705),
.Y(n_1858)
);

AOI22xp5_ASAP7_75t_L g1859 ( 
.A1(n_1569),
.A2(n_1044),
.B1(n_1045),
.B2(n_1043),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1710),
.Y(n_1860)
);

INVx2_ASAP7_75t_L g1861 ( 
.A(n_1724),
.Y(n_1861)
);

BUFx2_ASAP7_75t_L g1862 ( 
.A(n_1640),
.Y(n_1862)
);

BUFx2_ASAP7_75t_L g1863 ( 
.A(n_1642),
.Y(n_1863)
);

NOR2xp67_ASAP7_75t_L g1864 ( 
.A(n_1649),
.B(n_28),
.Y(n_1864)
);

A2O1A1Ixp33_ASAP7_75t_L g1865 ( 
.A1(n_1542),
.A2(n_887),
.B(n_889),
.C(n_882),
.Y(n_1865)
);

AND2x2_ASAP7_75t_L g1866 ( 
.A(n_1570),
.B(n_1056),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1623),
.Y(n_1867)
);

AND2x6_ASAP7_75t_SL g1868 ( 
.A(n_1627),
.B(n_893),
.Y(n_1868)
);

CKINVDCx5p33_ASAP7_75t_R g1869 ( 
.A(n_1586),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1629),
.Y(n_1870)
);

BUFx12f_ASAP7_75t_L g1871 ( 
.A(n_1643),
.Y(n_1871)
);

NAND2xp5_ASAP7_75t_L g1872 ( 
.A(n_1491),
.B(n_1061),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1665),
.Y(n_1873)
);

AND2x2_ASAP7_75t_L g1874 ( 
.A(n_1611),
.B(n_1065),
.Y(n_1874)
);

AOI22xp5_ASAP7_75t_L g1875 ( 
.A1(n_1553),
.A2(n_1066),
.B1(n_1070),
.B2(n_1068),
.Y(n_1875)
);

INVx3_ASAP7_75t_L g1876 ( 
.A(n_1537),
.Y(n_1876)
);

INVx2_ASAP7_75t_L g1877 ( 
.A(n_1653),
.Y(n_1877)
);

INVx5_ASAP7_75t_L g1878 ( 
.A(n_1676),
.Y(n_1878)
);

INVx2_ASAP7_75t_L g1879 ( 
.A(n_1592),
.Y(n_1879)
);

INVx2_ASAP7_75t_L g1880 ( 
.A(n_1595),
.Y(n_1880)
);

INVxp67_ASAP7_75t_L g1881 ( 
.A(n_1637),
.Y(n_1881)
);

NAND2xp5_ASAP7_75t_L g1882 ( 
.A(n_1626),
.B(n_1073),
.Y(n_1882)
);

BUFx6f_ASAP7_75t_L g1883 ( 
.A(n_1725),
.Y(n_1883)
);

AOI22xp5_ASAP7_75t_L g1884 ( 
.A1(n_1558),
.A2(n_1074),
.B1(n_1084),
.B2(n_1079),
.Y(n_1884)
);

NAND2xp5_ASAP7_75t_SL g1885 ( 
.A(n_1527),
.B(n_1085),
.Y(n_1885)
);

OAI22xp5_ASAP7_75t_L g1886 ( 
.A1(n_1587),
.A2(n_907),
.B1(n_910),
.B2(n_898),
.Y(n_1886)
);

INVx3_ASAP7_75t_L g1887 ( 
.A(n_1676),
.Y(n_1887)
);

NOR2xp33_ASAP7_75t_L g1888 ( 
.A(n_1539),
.B(n_1089),
.Y(n_1888)
);

NOR2xp33_ASAP7_75t_L g1889 ( 
.A(n_1718),
.B(n_1090),
.Y(n_1889)
);

INVx5_ASAP7_75t_L g1890 ( 
.A(n_1527),
.Y(n_1890)
);

NAND2xp5_ASAP7_75t_L g1891 ( 
.A(n_1633),
.B(n_1096),
.Y(n_1891)
);

INVxp67_ASAP7_75t_L g1892 ( 
.A(n_1619),
.Y(n_1892)
);

O2A1O1Ixp33_ASAP7_75t_L g1893 ( 
.A1(n_1574),
.A2(n_914),
.B(n_915),
.C(n_911),
.Y(n_1893)
);

BUFx3_ASAP7_75t_L g1894 ( 
.A(n_1572),
.Y(n_1894)
);

NAND2x1p5_ASAP7_75t_L g1895 ( 
.A(n_1618),
.B(n_917),
.Y(n_1895)
);

INVx5_ASAP7_75t_L g1896 ( 
.A(n_1527),
.Y(n_1896)
);

BUFx4f_ASAP7_75t_L g1897 ( 
.A(n_1630),
.Y(n_1897)
);

INVxp67_ASAP7_75t_L g1898 ( 
.A(n_1617),
.Y(n_1898)
);

INVxp67_ASAP7_75t_L g1899 ( 
.A(n_1638),
.Y(n_1899)
);

NOR2xp33_ASAP7_75t_SL g1900 ( 
.A(n_1620),
.B(n_1099),
.Y(n_1900)
);

NAND2xp5_ASAP7_75t_L g1901 ( 
.A(n_1584),
.B(n_1100),
.Y(n_1901)
);

INVx3_ASAP7_75t_L g1902 ( 
.A(n_1591),
.Y(n_1902)
);

CKINVDCx5p33_ASAP7_75t_R g1903 ( 
.A(n_1567),
.Y(n_1903)
);

INVx2_ASAP7_75t_L g1904 ( 
.A(n_1589),
.Y(n_1904)
);

NAND2xp5_ASAP7_75t_L g1905 ( 
.A(n_1490),
.B(n_1500),
.Y(n_1905)
);

AND2x4_ASAP7_75t_L g1906 ( 
.A(n_1605),
.B(n_921),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1667),
.Y(n_1907)
);

A2O1A1Ixp33_ASAP7_75t_L g1908 ( 
.A1(n_1489),
.A2(n_925),
.B(n_928),
.C(n_922),
.Y(n_1908)
);

NOR2xp33_ASAP7_75t_L g1909 ( 
.A(n_1545),
.B(n_1102),
.Y(n_1909)
);

NAND2xp5_ASAP7_75t_L g1910 ( 
.A(n_1525),
.B(n_1103),
.Y(n_1910)
);

BUFx3_ASAP7_75t_L g1911 ( 
.A(n_1578),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1671),
.Y(n_1912)
);

NAND2xp5_ASAP7_75t_SL g1913 ( 
.A(n_1508),
.B(n_1107),
.Y(n_1913)
);

BUFx6f_ASAP7_75t_L g1914 ( 
.A(n_1579),
.Y(n_1914)
);

AND2x4_ASAP7_75t_L g1915 ( 
.A(n_1513),
.B(n_931),
.Y(n_1915)
);

NAND2xp5_ASAP7_75t_SL g1916 ( 
.A(n_1522),
.B(n_1110),
.Y(n_1916)
);

NOR2x1_ASAP7_75t_R g1917 ( 
.A(n_1588),
.B(n_1112),
.Y(n_1917)
);

AND2x4_ASAP7_75t_L g1918 ( 
.A(n_1521),
.B(n_937),
.Y(n_1918)
);

INVx1_ASAP7_75t_L g1919 ( 
.A(n_1658),
.Y(n_1919)
);

AND2x4_ASAP7_75t_L g1920 ( 
.A(n_1557),
.B(n_938),
.Y(n_1920)
);

AND2x2_ASAP7_75t_SL g1921 ( 
.A(n_1511),
.B(n_1661),
.Y(n_1921)
);

BUFx6f_ASAP7_75t_L g1922 ( 
.A(n_1579),
.Y(n_1922)
);

NAND3xp33_ASAP7_75t_SL g1923 ( 
.A(n_1664),
.B(n_1156),
.C(n_1154),
.Y(n_1923)
);

NAND2xp33_ASAP7_75t_SL g1924 ( 
.A(n_1567),
.B(n_1159),
.Y(n_1924)
);

BUFx2_ASAP7_75t_L g1925 ( 
.A(n_1648),
.Y(n_1925)
);

NAND3xp33_ASAP7_75t_SL g1926 ( 
.A(n_1631),
.B(n_1172),
.C(n_1171),
.Y(n_1926)
);

NOR2x1_ASAP7_75t_R g1927 ( 
.A(n_1659),
.B(n_1115),
.Y(n_1927)
);

OR2x6_ASAP7_75t_SL g1928 ( 
.A(n_1514),
.B(n_1118),
.Y(n_1928)
);

AND2x4_ASAP7_75t_L g1929 ( 
.A(n_1685),
.B(n_944),
.Y(n_1929)
);

AND2x4_ASAP7_75t_L g1930 ( 
.A(n_1706),
.B(n_952),
.Y(n_1930)
);

NAND2xp33_ASAP7_75t_L g1931 ( 
.A(n_1579),
.B(n_1119),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_1673),
.Y(n_1932)
);

BUFx4f_ASAP7_75t_L g1933 ( 
.A(n_1650),
.Y(n_1933)
);

CKINVDCx5p33_ASAP7_75t_R g1934 ( 
.A(n_1722),
.Y(n_1934)
);

INVx3_ASAP7_75t_L g1935 ( 
.A(n_1596),
.Y(n_1935)
);

NOR3xp33_ASAP7_75t_SL g1936 ( 
.A(n_1660),
.B(n_1121),
.C(n_1120),
.Y(n_1936)
);

NAND2xp5_ASAP7_75t_SL g1937 ( 
.A(n_1593),
.B(n_1122),
.Y(n_1937)
);

NAND2xp5_ASAP7_75t_L g1938 ( 
.A(n_1544),
.B(n_1547),
.Y(n_1938)
);

AND2x4_ASAP7_75t_L g1939 ( 
.A(n_1717),
.B(n_956),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1674),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1680),
.Y(n_1941)
);

CKINVDCx20_ASAP7_75t_R g1942 ( 
.A(n_1666),
.Y(n_1942)
);

NAND2xp5_ASAP7_75t_L g1943 ( 
.A(n_1548),
.B(n_1123),
.Y(n_1943)
);

NAND2xp5_ASAP7_75t_SL g1944 ( 
.A(n_1601),
.B(n_1125),
.Y(n_1944)
);

BUFx3_ASAP7_75t_L g1945 ( 
.A(n_1599),
.Y(n_1945)
);

NOR2xp33_ASAP7_75t_L g1946 ( 
.A(n_1607),
.B(n_1498),
.Y(n_1946)
);

CKINVDCx5p33_ASAP7_75t_R g1947 ( 
.A(n_1722),
.Y(n_1947)
);

INVx5_ASAP7_75t_L g1948 ( 
.A(n_1635),
.Y(n_1948)
);

OR2x6_ASAP7_75t_L g1949 ( 
.A(n_1524),
.B(n_903),
.Y(n_1949)
);

INVx1_ASAP7_75t_L g1950 ( 
.A(n_1734),
.Y(n_1950)
);

AND2x4_ASAP7_75t_SL g1951 ( 
.A(n_1600),
.B(n_903),
.Y(n_1951)
);

BUFx3_ASAP7_75t_L g1952 ( 
.A(n_1604),
.Y(n_1952)
);

INVx2_ASAP7_75t_SL g1953 ( 
.A(n_1612),
.Y(n_1953)
);

NOR2xp33_ASAP7_75t_R g1954 ( 
.A(n_1662),
.B(n_1126),
.Y(n_1954)
);

OR2x2_ASAP7_75t_L g1955 ( 
.A(n_1555),
.B(n_1129),
.Y(n_1955)
);

AND2x4_ASAP7_75t_L g1956 ( 
.A(n_1496),
.B(n_966),
.Y(n_1956)
);

INVx2_ASAP7_75t_L g1957 ( 
.A(n_1594),
.Y(n_1957)
);

A2O1A1Ixp33_ASAP7_75t_L g1958 ( 
.A1(n_1543),
.A2(n_967),
.B(n_970),
.C(n_968),
.Y(n_1958)
);

AND2x2_ASAP7_75t_L g1959 ( 
.A(n_1608),
.B(n_1130),
.Y(n_1959)
);

AOI22xp5_ASAP7_75t_L g1960 ( 
.A1(n_1529),
.A2(n_1559),
.B1(n_1560),
.B2(n_1556),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1656),
.Y(n_1961)
);

OAI21xp5_ASAP7_75t_L g1962 ( 
.A1(n_1564),
.A2(n_975),
.B(n_972),
.Y(n_1962)
);

AND2x2_ASAP7_75t_SL g1963 ( 
.A(n_1644),
.B(n_965),
.Y(n_1963)
);

AND2x2_ASAP7_75t_L g1964 ( 
.A(n_1503),
.B(n_1136),
.Y(n_1964)
);

NAND2xp5_ASAP7_75t_SL g1965 ( 
.A(n_1613),
.B(n_1137),
.Y(n_1965)
);

OR2x2_ASAP7_75t_L g1966 ( 
.A(n_1624),
.B(n_1138),
.Y(n_1966)
);

INVx1_ASAP7_75t_L g1967 ( 
.A(n_1614),
.Y(n_1967)
);

INVx1_ASAP7_75t_L g1968 ( 
.A(n_1639),
.Y(n_1968)
);

HB1xp67_ASAP7_75t_L g1969 ( 
.A(n_1647),
.Y(n_1969)
);

INVx3_ASAP7_75t_L g1970 ( 
.A(n_1651),
.Y(n_1970)
);

NAND2x1p5_ASAP7_75t_L g1971 ( 
.A(n_1590),
.B(n_981),
.Y(n_1971)
);

INVxp67_ASAP7_75t_L g1972 ( 
.A(n_1507),
.Y(n_1972)
);

INVx2_ASAP7_75t_L g1973 ( 
.A(n_1679),
.Y(n_1973)
);

INVxp67_ASAP7_75t_SL g1974 ( 
.A(n_1635),
.Y(n_1974)
);

NAND2xp5_ASAP7_75t_L g1975 ( 
.A(n_1568),
.B(n_1580),
.Y(n_1975)
);

INVx1_ASAP7_75t_L g1976 ( 
.A(n_1672),
.Y(n_1976)
);

INVx1_ASAP7_75t_L g1977 ( 
.A(n_1581),
.Y(n_1977)
);

INVx1_ASAP7_75t_L g1978 ( 
.A(n_1616),
.Y(n_1978)
);

INVx2_ASAP7_75t_L g1979 ( 
.A(n_1679),
.Y(n_1979)
);

AND2x2_ASAP7_75t_SL g1980 ( 
.A(n_1622),
.B(n_909),
.Y(n_1980)
);

INVx1_ASAP7_75t_L g1981 ( 
.A(n_1603),
.Y(n_1981)
);

AND2x4_ASAP7_75t_L g1982 ( 
.A(n_1609),
.B(n_986),
.Y(n_1982)
);

INVx1_ASAP7_75t_L g1983 ( 
.A(n_1641),
.Y(n_1983)
);

INVx1_ASAP7_75t_L g1984 ( 
.A(n_1625),
.Y(n_1984)
);

AND2x4_ASAP7_75t_L g1985 ( 
.A(n_1561),
.B(n_987),
.Y(n_1985)
);

AND2x2_ASAP7_75t_L g1986 ( 
.A(n_1561),
.B(n_1144),
.Y(n_1986)
);

AND2x2_ASAP7_75t_L g1987 ( 
.A(n_1668),
.B(n_1147),
.Y(n_1987)
);

NAND2xp5_ASAP7_75t_L g1988 ( 
.A(n_1688),
.B(n_1149),
.Y(n_1988)
);

AOI22xp33_ASAP7_75t_L g1989 ( 
.A1(n_1730),
.A2(n_991),
.B1(n_997),
.B2(n_990),
.Y(n_1989)
);

A2O1A1Ixp33_ASAP7_75t_L g1990 ( 
.A1(n_1670),
.A2(n_1001),
.B(n_1005),
.C(n_999),
.Y(n_1990)
);

AND2x2_ASAP7_75t_L g1991 ( 
.A(n_1657),
.B(n_1008),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1677),
.Y(n_1992)
);

NAND3xp33_ASAP7_75t_SL g1993 ( 
.A(n_1678),
.B(n_1025),
.C(n_1012),
.Y(n_1993)
);

OR2x6_ASAP7_75t_L g1994 ( 
.A(n_1675),
.B(n_909),
.Y(n_1994)
);

INVx4_ASAP7_75t_L g1995 ( 
.A(n_1657),
.Y(n_1995)
);

INVx2_ASAP7_75t_L g1996 ( 
.A(n_1663),
.Y(n_1996)
);

INVx1_ASAP7_75t_L g1997 ( 
.A(n_1669),
.Y(n_1997)
);

NAND2xp33_ASAP7_75t_L g1998 ( 
.A(n_1655),
.B(n_1077),
.Y(n_1998)
);

NAND2xp5_ASAP7_75t_L g1999 ( 
.A(n_1681),
.B(n_1032),
.Y(n_1999)
);

CKINVDCx5p33_ASAP7_75t_R g2000 ( 
.A(n_1681),
.Y(n_2000)
);

NAND2xp5_ASAP7_75t_L g2001 ( 
.A(n_1707),
.B(n_1034),
.Y(n_2001)
);

INVx1_ASAP7_75t_L g2002 ( 
.A(n_1707),
.Y(n_2002)
);

AOI22xp33_ASAP7_75t_L g2003 ( 
.A1(n_1697),
.A2(n_1047),
.B1(n_1048),
.B2(n_1038),
.Y(n_2003)
);

NAND2x1p5_ASAP7_75t_L g2004 ( 
.A(n_1576),
.B(n_1053),
.Y(n_2004)
);

AND2x6_ASAP7_75t_L g2005 ( 
.A(n_1487),
.B(n_912),
.Y(n_2005)
);

INVx5_ASAP7_75t_L g2006 ( 
.A(n_1576),
.Y(n_2006)
);

AND2x6_ASAP7_75t_SL g2007 ( 
.A(n_1627),
.B(n_1054),
.Y(n_2007)
);

INVx1_ASAP7_75t_L g2008 ( 
.A(n_1707),
.Y(n_2008)
);

NAND2xp5_ASAP7_75t_L g2009 ( 
.A(n_1707),
.B(n_1055),
.Y(n_2009)
);

NAND2xp5_ASAP7_75t_L g2010 ( 
.A(n_1707),
.B(n_1058),
.Y(n_2010)
);

AND2x4_ASAP7_75t_SL g2011 ( 
.A(n_1576),
.B(n_912),
.Y(n_2011)
);

AND2x2_ASAP7_75t_L g2012 ( 
.A(n_1551),
.B(n_1060),
.Y(n_2012)
);

BUFx6f_ASAP7_75t_L g2013 ( 
.A(n_1487),
.Y(n_2013)
);

AOI22xp33_ASAP7_75t_SL g2014 ( 
.A1(n_1516),
.A2(n_1157),
.B1(n_1160),
.B2(n_1150),
.Y(n_2014)
);

CKINVDCx5p33_ASAP7_75t_R g2015 ( 
.A(n_1709),
.Y(n_2015)
);

INVx1_ASAP7_75t_L g2016 ( 
.A(n_1707),
.Y(n_2016)
);

AND2x4_ASAP7_75t_L g2017 ( 
.A(n_1707),
.B(n_1064),
.Y(n_2017)
);

AND2x2_ASAP7_75t_L g2018 ( 
.A(n_1863),
.B(n_1176),
.Y(n_2018)
);

INVx2_ASAP7_75t_L g2019 ( 
.A(n_1877),
.Y(n_2019)
);

OAI21xp33_ASAP7_75t_L g2020 ( 
.A1(n_1938),
.A2(n_1082),
.B(n_1071),
.Y(n_2020)
);

O2A1O1Ixp33_ASAP7_75t_L g2021 ( 
.A1(n_1817),
.A2(n_1087),
.B(n_1091),
.C(n_1083),
.Y(n_2021)
);

OAI22xp5_ASAP7_75t_L g2022 ( 
.A1(n_1905),
.A2(n_1095),
.B1(n_1097),
.B2(n_1093),
.Y(n_2022)
);

OAI22xp5_ASAP7_75t_L g2023 ( 
.A1(n_1892),
.A2(n_1105),
.B1(n_1106),
.B2(n_1101),
.Y(n_2023)
);

BUFx2_ASAP7_75t_L g2024 ( 
.A(n_1843),
.Y(n_2024)
);

INVx1_ASAP7_75t_L g2025 ( 
.A(n_1753),
.Y(n_2025)
);

AND2x2_ASAP7_75t_L g2026 ( 
.A(n_1862),
.B(n_1143),
.Y(n_2026)
);

AOI21xp5_ASAP7_75t_L g2027 ( 
.A1(n_1770),
.A2(n_1127),
.B(n_1111),
.Y(n_2027)
);

AND2x2_ASAP7_75t_L g2028 ( 
.A(n_2012),
.B(n_1128),
.Y(n_2028)
);

NOR2xp33_ASAP7_75t_L g2029 ( 
.A(n_1752),
.B(n_1135),
.Y(n_2029)
);

NOR2xp33_ASAP7_75t_L g2030 ( 
.A(n_1745),
.B(n_1164),
.Y(n_2030)
);

CKINVDCx5p33_ASAP7_75t_R g2031 ( 
.A(n_1761),
.Y(n_2031)
);

NOR2xp33_ASAP7_75t_L g2032 ( 
.A(n_1797),
.B(n_1744),
.Y(n_2032)
);

BUFx6f_ASAP7_75t_SL g2033 ( 
.A(n_1740),
.Y(n_2033)
);

NAND2xp5_ASAP7_75t_L g2034 ( 
.A(n_1754),
.B(n_946),
.Y(n_2034)
);

NAND3xp33_ASAP7_75t_SL g2035 ( 
.A(n_1811),
.B(n_974),
.C(n_946),
.Y(n_2035)
);

NAND2xp5_ASAP7_75t_SL g2036 ( 
.A(n_1900),
.B(n_1878),
.Y(n_2036)
);

INVx1_ASAP7_75t_L g2037 ( 
.A(n_1742),
.Y(n_2037)
);

AND2x2_ASAP7_75t_L g2038 ( 
.A(n_2004),
.B(n_974),
.Y(n_2038)
);

INVx2_ASAP7_75t_L g2039 ( 
.A(n_1775),
.Y(n_2039)
);

O2A1O1Ixp33_ASAP7_75t_L g2040 ( 
.A1(n_1893),
.A2(n_1020),
.B(n_1040),
.C(n_1019),
.Y(n_2040)
);

AOI21xp5_ASAP7_75t_L g2041 ( 
.A1(n_1854),
.A2(n_1020),
.B(n_1019),
.Y(n_2041)
);

BUFx2_ASAP7_75t_L g2042 ( 
.A(n_1785),
.Y(n_2042)
);

BUFx6f_ASAP7_75t_L g2043 ( 
.A(n_1776),
.Y(n_2043)
);

AOI21xp5_ASAP7_75t_L g2044 ( 
.A1(n_1975),
.A2(n_1078),
.B(n_1146),
.Y(n_2044)
);

NAND2xp5_ASAP7_75t_L g2045 ( 
.A(n_1867),
.B(n_1146),
.Y(n_2045)
);

NAND2xp5_ASAP7_75t_L g2046 ( 
.A(n_1870),
.B(n_1146),
.Y(n_2046)
);

AO32x2_ASAP7_75t_L g2047 ( 
.A1(n_1886),
.A2(n_1146),
.A3(n_32),
.B1(n_28),
.B2(n_31),
.Y(n_2047)
);

INVx3_ASAP7_75t_L g2048 ( 
.A(n_1890),
.Y(n_2048)
);

A2O1A1Ixp33_ASAP7_75t_L g2049 ( 
.A1(n_1919),
.A2(n_33),
.B(n_31),
.C(n_32),
.Y(n_2049)
);

NAND2xp5_ASAP7_75t_L g2050 ( 
.A(n_1804),
.B(n_34),
.Y(n_2050)
);

BUFx12f_ASAP7_75t_L g2051 ( 
.A(n_1788),
.Y(n_2051)
);

OAI22xp5_ASAP7_75t_SL g2052 ( 
.A1(n_1921),
.A2(n_37),
.B1(n_35),
.B2(n_36),
.Y(n_2052)
);

OAI22xp5_ASAP7_75t_L g2053 ( 
.A1(n_1994),
.A2(n_38),
.B1(n_35),
.B2(n_36),
.Y(n_2053)
);

AOI22xp33_ASAP7_75t_L g2054 ( 
.A1(n_1923),
.A2(n_41),
.B1(n_39),
.B2(n_40),
.Y(n_2054)
);

INVx1_ASAP7_75t_L g2055 ( 
.A(n_1819),
.Y(n_2055)
);

NOR2xp33_ASAP7_75t_R g2056 ( 
.A(n_2015),
.B(n_39),
.Y(n_2056)
);

NOR2xp33_ASAP7_75t_L g2057 ( 
.A(n_1774),
.B(n_40),
.Y(n_2057)
);

NAND2xp5_ASAP7_75t_SL g2058 ( 
.A(n_1878),
.B(n_41),
.Y(n_2058)
);

AOI21xp5_ASAP7_75t_L g2059 ( 
.A1(n_1974),
.A2(n_677),
.B(n_676),
.Y(n_2059)
);

NOR2xp67_ASAP7_75t_L g2060 ( 
.A(n_1736),
.B(n_42),
.Y(n_2060)
);

BUFx2_ASAP7_75t_L g2061 ( 
.A(n_1749),
.Y(n_2061)
);

NAND2xp5_ASAP7_75t_SL g2062 ( 
.A(n_1878),
.B(n_43),
.Y(n_2062)
);

AND2x2_ASAP7_75t_SL g2063 ( 
.A(n_1807),
.B(n_1897),
.Y(n_2063)
);

O2A1O1Ixp33_ASAP7_75t_L g2064 ( 
.A1(n_1958),
.A2(n_46),
.B(n_44),
.C(n_45),
.Y(n_2064)
);

NAND3xp33_ASAP7_75t_SL g2065 ( 
.A(n_1738),
.B(n_44),
.C(n_45),
.Y(n_2065)
);

INVx1_ASAP7_75t_SL g2066 ( 
.A(n_2011),
.Y(n_2066)
);

CKINVDCx20_ASAP7_75t_R g2067 ( 
.A(n_1749),
.Y(n_2067)
);

OAI22xp5_ASAP7_75t_L g2068 ( 
.A1(n_1806),
.A2(n_54),
.B1(n_51),
.B2(n_52),
.Y(n_2068)
);

AOI22xp33_ASAP7_75t_L g2069 ( 
.A1(n_1829),
.A2(n_55),
.B1(n_51),
.B2(n_54),
.Y(n_2069)
);

A2O1A1Ixp33_ASAP7_75t_L g2070 ( 
.A1(n_1873),
.A2(n_58),
.B(n_56),
.C(n_57),
.Y(n_2070)
);

A2O1A1Ixp33_ASAP7_75t_L g2071 ( 
.A1(n_1907),
.A2(n_59),
.B(n_57),
.C(n_58),
.Y(n_2071)
);

OAI22x1_ASAP7_75t_L g2072 ( 
.A1(n_1828),
.A2(n_63),
.B1(n_61),
.B2(n_62),
.Y(n_2072)
);

NAND2xp5_ASAP7_75t_L g2073 ( 
.A(n_1813),
.B(n_62),
.Y(n_2073)
);

NAND2xp5_ASAP7_75t_L g2074 ( 
.A(n_1815),
.B(n_63),
.Y(n_2074)
);

BUFx6f_ASAP7_75t_L g2075 ( 
.A(n_1776),
.Y(n_2075)
);

INVx1_ASAP7_75t_L g2076 ( 
.A(n_1816),
.Y(n_2076)
);

O2A1O1Ixp33_ASAP7_75t_L g2077 ( 
.A1(n_1865),
.A2(n_66),
.B(n_64),
.C(n_65),
.Y(n_2077)
);

INVx3_ASAP7_75t_L g2078 ( 
.A(n_1890),
.Y(n_2078)
);

BUFx3_ASAP7_75t_L g2079 ( 
.A(n_1748),
.Y(n_2079)
);

A2O1A1Ixp33_ASAP7_75t_L g2080 ( 
.A1(n_1912),
.A2(n_67),
.B(n_65),
.C(n_66),
.Y(n_2080)
);

A2O1A1Ixp33_ASAP7_75t_L g2081 ( 
.A1(n_1932),
.A2(n_69),
.B(n_67),
.C(n_68),
.Y(n_2081)
);

NOR2x1_ASAP7_75t_SL g2082 ( 
.A(n_1757),
.B(n_69),
.Y(n_2082)
);

OAI22x1_ASAP7_75t_L g2083 ( 
.A1(n_1820),
.A2(n_1771),
.B1(n_1881),
.B2(n_1802),
.Y(n_2083)
);

BUFx12f_ASAP7_75t_L g2084 ( 
.A(n_1871),
.Y(n_2084)
);

NAND2xp5_ASAP7_75t_L g2085 ( 
.A(n_2017),
.B(n_68),
.Y(n_2085)
);

AND2x2_ASAP7_75t_L g2086 ( 
.A(n_1866),
.B(n_70),
.Y(n_2086)
);

CKINVDCx5p33_ASAP7_75t_R g2087 ( 
.A(n_1823),
.Y(n_2087)
);

AND2x4_ASAP7_75t_L g2088 ( 
.A(n_1735),
.B(n_71),
.Y(n_2088)
);

A2O1A1Ixp33_ASAP7_75t_L g2089 ( 
.A1(n_1940),
.A2(n_74),
.B(n_72),
.C(n_73),
.Y(n_2089)
);

INVxp67_ASAP7_75t_L g2090 ( 
.A(n_1737),
.Y(n_2090)
);

AND2x2_ASAP7_75t_L g2091 ( 
.A(n_2017),
.B(n_72),
.Y(n_2091)
);

BUFx3_ASAP7_75t_L g2092 ( 
.A(n_1772),
.Y(n_2092)
);

AOI21xp5_ASAP7_75t_L g2093 ( 
.A1(n_1891),
.A2(n_696),
.B(n_694),
.Y(n_2093)
);

INVxp33_ASAP7_75t_SL g2094 ( 
.A(n_1917),
.Y(n_2094)
);

INVxp67_ASAP7_75t_L g2095 ( 
.A(n_1739),
.Y(n_2095)
);

NAND2xp5_ASAP7_75t_L g2096 ( 
.A(n_1798),
.B(n_1809),
.Y(n_2096)
);

BUFx3_ASAP7_75t_L g2097 ( 
.A(n_1800),
.Y(n_2097)
);

INVx4_ASAP7_75t_L g2098 ( 
.A(n_1890),
.Y(n_2098)
);

NAND2xp5_ASAP7_75t_SL g2099 ( 
.A(n_1741),
.B(n_75),
.Y(n_2099)
);

CKINVDCx5p33_ASAP7_75t_R g2100 ( 
.A(n_1903),
.Y(n_2100)
);

OAI22xp5_ASAP7_75t_L g2101 ( 
.A1(n_1994),
.A2(n_79),
.B1(n_76),
.B2(n_78),
.Y(n_2101)
);

BUFx6f_ASAP7_75t_L g2102 ( 
.A(n_1776),
.Y(n_2102)
);

INVx2_ASAP7_75t_L g2103 ( 
.A(n_1904),
.Y(n_2103)
);

NAND2xp5_ASAP7_75t_SL g2104 ( 
.A(n_2002),
.B(n_76),
.Y(n_2104)
);

NOR2xp33_ASAP7_75t_L g2105 ( 
.A(n_1898),
.B(n_81),
.Y(n_2105)
);

INVx4_ASAP7_75t_L g2106 ( 
.A(n_1896),
.Y(n_2106)
);

INVx2_ASAP7_75t_SL g2107 ( 
.A(n_1839),
.Y(n_2107)
);

NAND2xp5_ASAP7_75t_SL g2108 ( 
.A(n_2008),
.B(n_81),
.Y(n_2108)
);

NOR2xp33_ASAP7_75t_L g2109 ( 
.A(n_1899),
.B(n_82),
.Y(n_2109)
);

CKINVDCx14_ASAP7_75t_R g2110 ( 
.A(n_1805),
.Y(n_2110)
);

INVxp67_ASAP7_75t_L g2111 ( 
.A(n_2016),
.Y(n_2111)
);

OAI22xp5_ASAP7_75t_L g2112 ( 
.A1(n_2001),
.A2(n_85),
.B1(n_83),
.B2(n_84),
.Y(n_2112)
);

AND2x4_ASAP7_75t_L g2113 ( 
.A(n_1855),
.B(n_83),
.Y(n_2113)
);

BUFx2_ASAP7_75t_L g2114 ( 
.A(n_1757),
.Y(n_2114)
);

BUFx2_ASAP7_75t_L g2115 ( 
.A(n_1765),
.Y(n_2115)
);

AND2x4_ASAP7_75t_L g2116 ( 
.A(n_1855),
.B(n_84),
.Y(n_2116)
);

NAND2xp5_ASAP7_75t_L g2117 ( 
.A(n_1798),
.B(n_86),
.Y(n_2117)
);

NAND2xp5_ASAP7_75t_L g2118 ( 
.A(n_1759),
.B(n_2003),
.Y(n_2118)
);

INVx1_ASAP7_75t_L g2119 ( 
.A(n_1784),
.Y(n_2119)
);

CKINVDCx5p33_ASAP7_75t_R g2120 ( 
.A(n_1934),
.Y(n_2120)
);

OR2x2_ASAP7_75t_L g2121 ( 
.A(n_1769),
.B(n_86),
.Y(n_2121)
);

INVx2_ASAP7_75t_L g2122 ( 
.A(n_1879),
.Y(n_2122)
);

INVx1_ASAP7_75t_L g2123 ( 
.A(n_1801),
.Y(n_2123)
);

OAI22xp5_ASAP7_75t_L g2124 ( 
.A1(n_2009),
.A2(n_89),
.B1(n_87),
.B2(n_88),
.Y(n_2124)
);

BUFx12f_ASAP7_75t_L g2125 ( 
.A(n_2007),
.Y(n_2125)
);

NOR2xp33_ASAP7_75t_L g2126 ( 
.A(n_1925),
.B(n_87),
.Y(n_2126)
);

AOI22xp5_ASAP7_75t_L g2127 ( 
.A1(n_1836),
.A2(n_92),
.B1(n_88),
.B2(n_91),
.Y(n_2127)
);

O2A1O1Ixp33_ASAP7_75t_L g2128 ( 
.A1(n_1908),
.A2(n_94),
.B(n_92),
.C(n_93),
.Y(n_2128)
);

OAI21xp5_ASAP7_75t_L g2129 ( 
.A1(n_1990),
.A2(n_1941),
.B(n_1962),
.Y(n_2129)
);

INVx2_ASAP7_75t_L g2130 ( 
.A(n_1880),
.Y(n_2130)
);

O2A1O1Ixp33_ASAP7_75t_L g2131 ( 
.A1(n_1976),
.A2(n_96),
.B(n_94),
.C(n_95),
.Y(n_2131)
);

NAND2xp5_ASAP7_75t_SL g2132 ( 
.A(n_1896),
.B(n_95),
.Y(n_2132)
);

INVx1_ASAP7_75t_L g2133 ( 
.A(n_1746),
.Y(n_2133)
);

NAND2xp5_ASAP7_75t_L g2134 ( 
.A(n_1780),
.B(n_96),
.Y(n_2134)
);

OAI21xp33_ASAP7_75t_SL g2135 ( 
.A1(n_1960),
.A2(n_97),
.B(n_98),
.Y(n_2135)
);

NAND2xp5_ASAP7_75t_L g2136 ( 
.A(n_1920),
.B(n_98),
.Y(n_2136)
);

BUFx2_ASAP7_75t_L g2137 ( 
.A(n_1765),
.Y(n_2137)
);

AO32x1_ASAP7_75t_L g2138 ( 
.A1(n_1986),
.A2(n_101),
.A3(n_99),
.B1(n_100),
.B2(n_103),
.Y(n_2138)
);

BUFx6f_ASAP7_75t_L g2139 ( 
.A(n_1792),
.Y(n_2139)
);

NOR2xp33_ASAP7_75t_L g2140 ( 
.A(n_1889),
.B(n_101),
.Y(n_2140)
);

NOR2xp33_ASAP7_75t_L g2141 ( 
.A(n_1778),
.B(n_104),
.Y(n_2141)
);

INVx4_ASAP7_75t_L g2142 ( 
.A(n_1896),
.Y(n_2142)
);

OR2x2_ASAP7_75t_L g2143 ( 
.A(n_1768),
.B(n_105),
.Y(n_2143)
);

NOR2xp33_ASAP7_75t_L g2144 ( 
.A(n_1796),
.B(n_106),
.Y(n_2144)
);

AOI22xp33_ASAP7_75t_L g2145 ( 
.A1(n_1845),
.A2(n_108),
.B1(n_106),
.B2(n_107),
.Y(n_2145)
);

NAND2xp5_ASAP7_75t_SL g2146 ( 
.A(n_1795),
.B(n_107),
.Y(n_2146)
);

NAND2xp5_ASAP7_75t_L g2147 ( 
.A(n_1920),
.B(n_109),
.Y(n_2147)
);

O2A1O1Ixp33_ASAP7_75t_L g2148 ( 
.A1(n_2010),
.A2(n_111),
.B(n_109),
.C(n_110),
.Y(n_2148)
);

AND2x2_ASAP7_75t_L g2149 ( 
.A(n_1758),
.B(n_110),
.Y(n_2149)
);

AND2x4_ASAP7_75t_SL g2150 ( 
.A(n_1762),
.B(n_111),
.Y(n_2150)
);

NOR2xp33_ASAP7_75t_R g2151 ( 
.A(n_1947),
.B(n_112),
.Y(n_2151)
);

CKINVDCx5p33_ASAP7_75t_R g2152 ( 
.A(n_1869),
.Y(n_2152)
);

AND2x2_ASAP7_75t_L g2153 ( 
.A(n_1874),
.B(n_115),
.Y(n_2153)
);

NAND2xp5_ASAP7_75t_SL g2154 ( 
.A(n_1789),
.B(n_115),
.Y(n_2154)
);

BUFx3_ASAP7_75t_L g2155 ( 
.A(n_1789),
.Y(n_2155)
);

NOR2xp33_ASAP7_75t_L g2156 ( 
.A(n_1972),
.B(n_116),
.Y(n_2156)
);

A2O1A1Ixp33_ASAP7_75t_L g2157 ( 
.A1(n_1838),
.A2(n_118),
.B(n_116),
.C(n_117),
.Y(n_2157)
);

NOR3xp33_ASAP7_75t_SL g2158 ( 
.A(n_1926),
.B(n_117),
.C(n_118),
.Y(n_2158)
);

AOI21xp5_ASAP7_75t_L g2159 ( 
.A1(n_1872),
.A2(n_710),
.B(n_709),
.Y(n_2159)
);

A2O1A1Ixp33_ASAP7_75t_L g2160 ( 
.A1(n_1946),
.A2(n_122),
.B(n_119),
.C(n_120),
.Y(n_2160)
);

BUFx6f_ASAP7_75t_L g2161 ( 
.A(n_1792),
.Y(n_2161)
);

A2O1A1Ixp33_ASAP7_75t_L g2162 ( 
.A1(n_1845),
.A2(n_123),
.B(n_120),
.C(n_122),
.Y(n_2162)
);

CKINVDCx5p33_ASAP7_75t_R g2163 ( 
.A(n_1924),
.Y(n_2163)
);

NAND2xp5_ASAP7_75t_L g2164 ( 
.A(n_1766),
.B(n_124),
.Y(n_2164)
);

OAI21xp33_ASAP7_75t_L g2165 ( 
.A1(n_1790),
.A2(n_125),
.B(n_128),
.Y(n_2165)
);

NAND2xp5_ASAP7_75t_L g2166 ( 
.A(n_1766),
.B(n_125),
.Y(n_2166)
);

OAI22x1_ASAP7_75t_L g2167 ( 
.A1(n_1895),
.A2(n_1985),
.B1(n_1763),
.B2(n_1789),
.Y(n_2167)
);

INVxp67_ASAP7_75t_L g2168 ( 
.A(n_1987),
.Y(n_2168)
);

HB1xp67_ASAP7_75t_L g2169 ( 
.A(n_1826),
.Y(n_2169)
);

INVx1_ASAP7_75t_L g2170 ( 
.A(n_1830),
.Y(n_2170)
);

INVx1_ASAP7_75t_L g2171 ( 
.A(n_1832),
.Y(n_2171)
);

INVx2_ASAP7_75t_SL g2172 ( 
.A(n_2006),
.Y(n_2172)
);

O2A1O1Ixp33_ASAP7_75t_L g2173 ( 
.A1(n_1773),
.A2(n_1787),
.B(n_1799),
.C(n_1786),
.Y(n_2173)
);

INVx1_ASAP7_75t_L g2174 ( 
.A(n_1844),
.Y(n_2174)
);

NAND2xp5_ASAP7_75t_L g2175 ( 
.A(n_1915),
.B(n_129),
.Y(n_2175)
);

NAND2xp5_ASAP7_75t_L g2176 ( 
.A(n_1915),
.B(n_130),
.Y(n_2176)
);

NOR2xp33_ASAP7_75t_L g2177 ( 
.A(n_1846),
.B(n_131),
.Y(n_2177)
);

NAND2xp5_ASAP7_75t_SL g2178 ( 
.A(n_2006),
.B(n_132),
.Y(n_2178)
);

BUFx3_ASAP7_75t_L g2179 ( 
.A(n_2006),
.Y(n_2179)
);

INVx1_ASAP7_75t_L g2180 ( 
.A(n_1851),
.Y(n_2180)
);

AOI22xp33_ASAP7_75t_L g2181 ( 
.A1(n_1831),
.A2(n_136),
.B1(n_133),
.B2(n_134),
.Y(n_2181)
);

HB1xp67_ASAP7_75t_L g2182 ( 
.A(n_1969),
.Y(n_2182)
);

BUFx2_ASAP7_75t_L g2183 ( 
.A(n_1779),
.Y(n_2183)
);

NAND2xp5_ASAP7_75t_L g2184 ( 
.A(n_1918),
.B(n_136),
.Y(n_2184)
);

NOR2xp33_ASAP7_75t_L g2185 ( 
.A(n_1782),
.B(n_137),
.Y(n_2185)
);

OR2x6_ASAP7_75t_L g2186 ( 
.A(n_1887),
.B(n_137),
.Y(n_2186)
);

INVx6_ASAP7_75t_L g2187 ( 
.A(n_1945),
.Y(n_2187)
);

INVx1_ASAP7_75t_L g2188 ( 
.A(n_1860),
.Y(n_2188)
);

AND2x2_ASAP7_75t_L g2189 ( 
.A(n_2014),
.B(n_139),
.Y(n_2189)
);

INVx1_ASAP7_75t_L g2190 ( 
.A(n_1991),
.Y(n_2190)
);

CKINVDCx5p33_ASAP7_75t_R g2191 ( 
.A(n_1936),
.Y(n_2191)
);

NAND2xp5_ASAP7_75t_L g2192 ( 
.A(n_1918),
.B(n_139),
.Y(n_2192)
);

NAND2xp5_ASAP7_75t_SL g2193 ( 
.A(n_1933),
.B(n_141),
.Y(n_2193)
);

INVx2_ASAP7_75t_L g2194 ( 
.A(n_1824),
.Y(n_2194)
);

BUFx2_ASAP7_75t_L g2195 ( 
.A(n_1779),
.Y(n_2195)
);

NAND2x1p5_ASAP7_75t_L g2196 ( 
.A(n_1948),
.B(n_1995),
.Y(n_2196)
);

AOI21xp33_ASAP7_75t_L g2197 ( 
.A1(n_1927),
.A2(n_141),
.B(n_144),
.Y(n_2197)
);

NAND2xp5_ASAP7_75t_SL g2198 ( 
.A(n_2000),
.B(n_144),
.Y(n_2198)
);

INVx3_ASAP7_75t_L g2199 ( 
.A(n_1948),
.Y(n_2199)
);

NOR3xp33_ASAP7_75t_SL g2200 ( 
.A(n_1837),
.B(n_146),
.C(n_147),
.Y(n_2200)
);

NAND2xp5_ASAP7_75t_L g2201 ( 
.A(n_1967),
.B(n_146),
.Y(n_2201)
);

NAND2xp5_ASAP7_75t_L g2202 ( 
.A(n_1968),
.B(n_148),
.Y(n_2202)
);

INVx3_ASAP7_75t_L g2203 ( 
.A(n_1948),
.Y(n_2203)
);

CKINVDCx5p33_ASAP7_75t_R g2204 ( 
.A(n_1942),
.Y(n_2204)
);

INVx3_ASAP7_75t_L g2205 ( 
.A(n_1894),
.Y(n_2205)
);

INVx2_ASAP7_75t_L g2206 ( 
.A(n_1840),
.Y(n_2206)
);

NOR2xp33_ASAP7_75t_L g2207 ( 
.A(n_1764),
.B(n_148),
.Y(n_2207)
);

NAND2xp5_ASAP7_75t_L g2208 ( 
.A(n_1956),
.B(n_149),
.Y(n_2208)
);

NAND2xp5_ASAP7_75t_L g2209 ( 
.A(n_1956),
.B(n_1822),
.Y(n_2209)
);

NOR2xp33_ASAP7_75t_L g2210 ( 
.A(n_1767),
.B(n_149),
.Y(n_2210)
);

INVx2_ASAP7_75t_L g2211 ( 
.A(n_1848),
.Y(n_2211)
);

INVx2_ASAP7_75t_L g2212 ( 
.A(n_1850),
.Y(n_2212)
);

NAND2xp5_ASAP7_75t_L g2213 ( 
.A(n_1827),
.B(n_150),
.Y(n_2213)
);

INVx1_ASAP7_75t_L g2214 ( 
.A(n_1906),
.Y(n_2214)
);

A2O1A1Ixp33_ASAP7_75t_L g2215 ( 
.A1(n_1831),
.A2(n_153),
.B(n_150),
.C(n_152),
.Y(n_2215)
);

CKINVDCx5p33_ASAP7_75t_R g2216 ( 
.A(n_1868),
.Y(n_2216)
);

NOR2xp33_ASAP7_75t_L g2217 ( 
.A(n_1833),
.B(n_154),
.Y(n_2217)
);

NOR2xp33_ASAP7_75t_L g2218 ( 
.A(n_1834),
.B(n_154),
.Y(n_2218)
);

INVx2_ASAP7_75t_L g2219 ( 
.A(n_1852),
.Y(n_2219)
);

OA22x2_ASAP7_75t_L g2220 ( 
.A1(n_1951),
.A2(n_157),
.B1(n_155),
.B2(n_156),
.Y(n_2220)
);

NAND2xp5_ASAP7_75t_SL g2221 ( 
.A(n_1803),
.B(n_157),
.Y(n_2221)
);

BUFx2_ASAP7_75t_L g2222 ( 
.A(n_1794),
.Y(n_2222)
);

BUFx12f_ASAP7_75t_L g2223 ( 
.A(n_1906),
.Y(n_2223)
);

CKINVDCx8_ASAP7_75t_R g2224 ( 
.A(n_1794),
.Y(n_2224)
);

O2A1O1Ixp33_ASAP7_75t_L g2225 ( 
.A1(n_1743),
.A2(n_160),
.B(n_158),
.C(n_159),
.Y(n_2225)
);

INVx2_ASAP7_75t_L g2226 ( 
.A(n_1858),
.Y(n_2226)
);

INVx1_ASAP7_75t_L g2227 ( 
.A(n_1861),
.Y(n_2227)
);

NOR2xp33_ASAP7_75t_L g2228 ( 
.A(n_1909),
.B(n_158),
.Y(n_2228)
);

NOR2xp33_ASAP7_75t_L g2229 ( 
.A(n_1952),
.B(n_159),
.Y(n_2229)
);

NOR2xp33_ASAP7_75t_R g2230 ( 
.A(n_1794),
.B(n_2005),
.Y(n_2230)
);

INVx1_ASAP7_75t_L g2231 ( 
.A(n_1750),
.Y(n_2231)
);

NAND2xp5_ASAP7_75t_L g2232 ( 
.A(n_1853),
.B(n_160),
.Y(n_2232)
);

NAND2xp5_ASAP7_75t_L g2233 ( 
.A(n_1781),
.B(n_161),
.Y(n_2233)
);

INVx1_ASAP7_75t_L g2234 ( 
.A(n_1756),
.Y(n_2234)
);

BUFx3_ASAP7_75t_L g2235 ( 
.A(n_1973),
.Y(n_2235)
);

AND2x2_ASAP7_75t_L g2236 ( 
.A(n_1814),
.B(n_161),
.Y(n_2236)
);

NOR2xp33_ASAP7_75t_L g2237 ( 
.A(n_1747),
.B(n_162),
.Y(n_2237)
);

OAI22x1_ASAP7_75t_L g2238 ( 
.A1(n_1955),
.A2(n_164),
.B1(n_162),
.B2(n_163),
.Y(n_2238)
);

BUFx4f_ASAP7_75t_L g2239 ( 
.A(n_1835),
.Y(n_2239)
);

NAND2xp5_ASAP7_75t_L g2240 ( 
.A(n_1963),
.B(n_163),
.Y(n_2240)
);

BUFx2_ASAP7_75t_L g2241 ( 
.A(n_1835),
.Y(n_2241)
);

HB1xp67_ASAP7_75t_L g2242 ( 
.A(n_1911),
.Y(n_2242)
);

AOI21xp5_ASAP7_75t_L g2243 ( 
.A1(n_1996),
.A2(n_720),
.B(n_718),
.Y(n_2243)
);

NOR2xp33_ASAP7_75t_R g2244 ( 
.A(n_1835),
.B(n_165),
.Y(n_2244)
);

NOR2xp33_ASAP7_75t_L g2245 ( 
.A(n_1964),
.B(n_166),
.Y(n_2245)
);

AOI21xp5_ASAP7_75t_L g2246 ( 
.A1(n_1901),
.A2(n_728),
.B(n_724),
.Y(n_2246)
);

INVx2_ASAP7_75t_L g2247 ( 
.A(n_1999),
.Y(n_2247)
);

INVx2_ASAP7_75t_L g2248 ( 
.A(n_1997),
.Y(n_2248)
);

INVx3_ASAP7_75t_L g2249 ( 
.A(n_2005),
.Y(n_2249)
);

INVx4_ASAP7_75t_L g2250 ( 
.A(n_2005),
.Y(n_2250)
);

CKINVDCx20_ASAP7_75t_R g2251 ( 
.A(n_1859),
.Y(n_2251)
);

INVx3_ASAP7_75t_L g2252 ( 
.A(n_1979),
.Y(n_2252)
);

AND2x2_ASAP7_75t_L g2253 ( 
.A(n_1875),
.B(n_170),
.Y(n_2253)
);

INVx1_ASAP7_75t_L g2254 ( 
.A(n_1760),
.Y(n_2254)
);

AOI22xp33_ASAP7_75t_L g2255 ( 
.A1(n_1755),
.A2(n_1929),
.B1(n_1939),
.B2(n_1930),
.Y(n_2255)
);

NOR2xp33_ASAP7_75t_L g2256 ( 
.A(n_1910),
.B(n_171),
.Y(n_2256)
);

O2A1O1Ixp33_ASAP7_75t_L g2257 ( 
.A1(n_1882),
.A2(n_174),
.B(n_172),
.C(n_173),
.Y(n_2257)
);

A2O1A1Ixp33_ASAP7_75t_L g2258 ( 
.A1(n_1864),
.A2(n_174),
.B(n_172),
.C(n_173),
.Y(n_2258)
);

NOR2xp33_ASAP7_75t_L g2259 ( 
.A(n_1902),
.B(n_177),
.Y(n_2259)
);

CKINVDCx20_ASAP7_75t_R g2260 ( 
.A(n_1884),
.Y(n_2260)
);

NAND2xp5_ASAP7_75t_L g2261 ( 
.A(n_1755),
.B(n_177),
.Y(n_2261)
);

AOI22xp33_ASAP7_75t_L g2262 ( 
.A1(n_1929),
.A2(n_1930),
.B1(n_1939),
.B2(n_1982),
.Y(n_2262)
);

INVx1_ASAP7_75t_L g2263 ( 
.A(n_1825),
.Y(n_2263)
);

BUFx6f_ASAP7_75t_SL g2264 ( 
.A(n_1982),
.Y(n_2264)
);

AND2x4_ASAP7_75t_SL g2265 ( 
.A(n_1810),
.B(n_178),
.Y(n_2265)
);

NAND2xp5_ASAP7_75t_L g2266 ( 
.A(n_1849),
.B(n_1953),
.Y(n_2266)
);

BUFx12f_ASAP7_75t_L g2267 ( 
.A(n_1949),
.Y(n_2267)
);

BUFx3_ASAP7_75t_L g2268 ( 
.A(n_1935),
.Y(n_2268)
);

INVx8_ASAP7_75t_L g2269 ( 
.A(n_1818),
.Y(n_2269)
);

NOR2xp33_ASAP7_75t_SL g2270 ( 
.A(n_1818),
.B(n_731),
.Y(n_2270)
);

BUFx2_ASAP7_75t_L g2271 ( 
.A(n_1856),
.Y(n_2271)
);

OAI22x1_ASAP7_75t_L g2272 ( 
.A1(n_1808),
.A2(n_180),
.B1(n_178),
.B2(n_179),
.Y(n_2272)
);

INVx4_ASAP7_75t_L g2273 ( 
.A(n_1841),
.Y(n_2273)
);

INVx2_ASAP7_75t_L g2274 ( 
.A(n_1957),
.Y(n_2274)
);

INVx5_ASAP7_75t_L g2275 ( 
.A(n_1841),
.Y(n_2275)
);

NAND2xp5_ASAP7_75t_L g2276 ( 
.A(n_1888),
.B(n_1970),
.Y(n_2276)
);

AND2x4_ASAP7_75t_L g2277 ( 
.A(n_1842),
.B(n_180),
.Y(n_2277)
);

NAND2xp5_ASAP7_75t_L g2278 ( 
.A(n_1959),
.B(n_182),
.Y(n_2278)
);

INVx1_ASAP7_75t_L g2279 ( 
.A(n_1876),
.Y(n_2279)
);

AND2x4_ASAP7_75t_L g2280 ( 
.A(n_1791),
.B(n_182),
.Y(n_2280)
);

OAI22xp5_ASAP7_75t_L g2281 ( 
.A1(n_1914),
.A2(n_185),
.B1(n_183),
.B2(n_184),
.Y(n_2281)
);

NAND2xp5_ASAP7_75t_L g2282 ( 
.A(n_1913),
.B(n_183),
.Y(n_2282)
);

NAND3xp33_ASAP7_75t_L g2283 ( 
.A(n_1931),
.B(n_184),
.C(n_185),
.Y(n_2283)
);

NOR2xp33_ASAP7_75t_L g2284 ( 
.A(n_1937),
.B(n_187),
.Y(n_2284)
);

NAND2xp5_ASAP7_75t_L g2285 ( 
.A(n_1916),
.B(n_188),
.Y(n_2285)
);

NAND2xp5_ASAP7_75t_L g2286 ( 
.A(n_1944),
.B(n_188),
.Y(n_2286)
);

NOR2xp33_ASAP7_75t_L g2287 ( 
.A(n_1965),
.B(n_189),
.Y(n_2287)
);

BUFx6f_ASAP7_75t_L g2288 ( 
.A(n_1883),
.Y(n_2288)
);

OAI221xp5_ASAP7_75t_L g2289 ( 
.A1(n_1943),
.A2(n_192),
.B1(n_190),
.B2(n_191),
.C(n_193),
.Y(n_2289)
);

OAI21xp5_ASAP7_75t_L g2290 ( 
.A1(n_1783),
.A2(n_193),
.B(n_194),
.Y(n_2290)
);

O2A1O1Ixp33_ASAP7_75t_L g2291 ( 
.A1(n_1821),
.A2(n_196),
.B(n_194),
.C(n_195),
.Y(n_2291)
);

BUFx12f_ASAP7_75t_L g2292 ( 
.A(n_1949),
.Y(n_2292)
);

NAND2xp5_ASAP7_75t_L g2293 ( 
.A(n_1950),
.B(n_195),
.Y(n_2293)
);

NOR2xp33_ASAP7_75t_L g2294 ( 
.A(n_1966),
.B(n_197),
.Y(n_2294)
);

INVx2_ASAP7_75t_SL g2295 ( 
.A(n_1885),
.Y(n_2295)
);

AOI22xp5_ASAP7_75t_L g2296 ( 
.A1(n_1977),
.A2(n_201),
.B1(n_199),
.B2(n_200),
.Y(n_2296)
);

NAND3xp33_ASAP7_75t_SL g2297 ( 
.A(n_1971),
.B(n_199),
.C(n_202),
.Y(n_2297)
);

NOR2xp67_ASAP7_75t_L g2298 ( 
.A(n_1961),
.B(n_202),
.Y(n_2298)
);

NOR2xp33_ASAP7_75t_L g2299 ( 
.A(n_1928),
.B(n_205),
.Y(n_2299)
);

AND2x2_ASAP7_75t_L g2300 ( 
.A(n_1980),
.B(n_206),
.Y(n_2300)
);

INVx2_ASAP7_75t_L g2301 ( 
.A(n_1978),
.Y(n_2301)
);

CKINVDCx5p33_ASAP7_75t_R g2302 ( 
.A(n_1954),
.Y(n_2302)
);

NAND2xp5_ASAP7_75t_L g2303 ( 
.A(n_1981),
.B(n_208),
.Y(n_2303)
);

NAND2xp5_ASAP7_75t_L g2304 ( 
.A(n_1847),
.B(n_208),
.Y(n_2304)
);

NOR2xp33_ASAP7_75t_L g2305 ( 
.A(n_1857),
.B(n_1983),
.Y(n_2305)
);

NAND2xp5_ASAP7_75t_L g2306 ( 
.A(n_1989),
.B(n_209),
.Y(n_2306)
);

INVx3_ASAP7_75t_SL g2307 ( 
.A(n_2013),
.Y(n_2307)
);

NOR2xp33_ASAP7_75t_L g2308 ( 
.A(n_1988),
.B(n_210),
.Y(n_2308)
);

AOI22xp5_ASAP7_75t_L g2309 ( 
.A1(n_1993),
.A2(n_1984),
.B1(n_1992),
.B2(n_1922),
.Y(n_2309)
);

BUFx12f_ASAP7_75t_L g2310 ( 
.A(n_2013),
.Y(n_2310)
);

INVx1_ASAP7_75t_L g2311 ( 
.A(n_1998),
.Y(n_2311)
);

O2A1O1Ixp33_ASAP7_75t_L g2312 ( 
.A1(n_1922),
.A2(n_213),
.B(n_211),
.C(n_212),
.Y(n_2312)
);

AOI21xp5_ASAP7_75t_L g2313 ( 
.A1(n_1770),
.A2(n_212),
.B(n_214),
.Y(n_2313)
);

BUFx6f_ASAP7_75t_L g2314 ( 
.A(n_1776),
.Y(n_2314)
);

NAND2xp5_ASAP7_75t_L g2315 ( 
.A(n_1751),
.B(n_215),
.Y(n_2315)
);

AOI21xp5_ASAP7_75t_L g2316 ( 
.A1(n_1770),
.A2(n_215),
.B(n_216),
.Y(n_2316)
);

NAND2xp5_ASAP7_75t_L g2317 ( 
.A(n_1751),
.B(n_217),
.Y(n_2317)
);

AOI21xp5_ASAP7_75t_L g2318 ( 
.A1(n_1770),
.A2(n_217),
.B(n_218),
.Y(n_2318)
);

INVx1_ASAP7_75t_L g2319 ( 
.A(n_1751),
.Y(n_2319)
);

O2A1O1Ixp33_ASAP7_75t_L g2320 ( 
.A1(n_1817),
.A2(n_222),
.B(n_218),
.C(n_219),
.Y(n_2320)
);

INVx3_ASAP7_75t_L g2321 ( 
.A(n_1890),
.Y(n_2321)
);

NOR2xp33_ASAP7_75t_L g2322 ( 
.A(n_1752),
.B(n_222),
.Y(n_2322)
);

NOR2xp33_ASAP7_75t_L g2323 ( 
.A(n_1752),
.B(n_223),
.Y(n_2323)
);

NOR2xp33_ASAP7_75t_L g2324 ( 
.A(n_1752),
.B(n_225),
.Y(n_2324)
);

INVx1_ASAP7_75t_L g2325 ( 
.A(n_1751),
.Y(n_2325)
);

NAND2xp5_ASAP7_75t_L g2326 ( 
.A(n_1751),
.B(n_228),
.Y(n_2326)
);

CKINVDCx8_ASAP7_75t_R g2327 ( 
.A(n_2007),
.Y(n_2327)
);

INVx3_ASAP7_75t_SL g2328 ( 
.A(n_1761),
.Y(n_2328)
);

BUFx2_ASAP7_75t_L g2329 ( 
.A(n_1843),
.Y(n_2329)
);

AOI21xp5_ASAP7_75t_L g2330 ( 
.A1(n_1770),
.A2(n_229),
.B(n_230),
.Y(n_2330)
);

OAI22xp5_ASAP7_75t_L g2331 ( 
.A1(n_1938),
.A2(n_234),
.B1(n_232),
.B2(n_233),
.Y(n_2331)
);

NAND2xp5_ASAP7_75t_L g2332 ( 
.A(n_1751),
.B(n_232),
.Y(n_2332)
);

NAND2xp5_ASAP7_75t_L g2333 ( 
.A(n_1751),
.B(n_235),
.Y(n_2333)
);

OAI21x1_ASAP7_75t_L g2334 ( 
.A1(n_1770),
.A2(n_235),
.B(n_236),
.Y(n_2334)
);

NOR2xp33_ASAP7_75t_L g2335 ( 
.A(n_1752),
.B(n_236),
.Y(n_2335)
);

INVx2_ASAP7_75t_L g2336 ( 
.A(n_1877),
.Y(n_2336)
);

AOI21xp5_ASAP7_75t_L g2337 ( 
.A1(n_1770),
.A2(n_237),
.B(n_238),
.Y(n_2337)
);

AOI21x1_ASAP7_75t_L g2338 ( 
.A1(n_1777),
.A2(n_237),
.B(n_239),
.Y(n_2338)
);

AOI22xp5_ASAP7_75t_L g2339 ( 
.A1(n_1892),
.A2(n_241),
.B1(n_239),
.B2(n_240),
.Y(n_2339)
);

INVx2_ASAP7_75t_L g2340 ( 
.A(n_1877),
.Y(n_2340)
);

AND2x2_ASAP7_75t_L g2341 ( 
.A(n_1793),
.B(n_240),
.Y(n_2341)
);

NAND2xp5_ASAP7_75t_L g2342 ( 
.A(n_1751),
.B(n_241),
.Y(n_2342)
);

INVx1_ASAP7_75t_L g2343 ( 
.A(n_1751),
.Y(n_2343)
);

INVx2_ASAP7_75t_L g2344 ( 
.A(n_1877),
.Y(n_2344)
);

AO21x1_ASAP7_75t_L g2345 ( 
.A1(n_1777),
.A2(n_243),
.B(n_244),
.Y(n_2345)
);

BUFx12f_ASAP7_75t_L g2346 ( 
.A(n_1788),
.Y(n_2346)
);

INVx4_ASAP7_75t_L g2347 ( 
.A(n_1740),
.Y(n_2347)
);

AO21x1_ASAP7_75t_L g2348 ( 
.A1(n_1777),
.A2(n_245),
.B(n_246),
.Y(n_2348)
);

AND2x2_ASAP7_75t_L g2349 ( 
.A(n_1793),
.B(n_247),
.Y(n_2349)
);

NAND2xp5_ASAP7_75t_L g2350 ( 
.A(n_1751),
.B(n_253),
.Y(n_2350)
);

INVx2_ASAP7_75t_L g2351 ( 
.A(n_1877),
.Y(n_2351)
);

AND2x2_ASAP7_75t_L g2352 ( 
.A(n_1793),
.B(n_255),
.Y(n_2352)
);

NOR2xp33_ASAP7_75t_L g2353 ( 
.A(n_1752),
.B(n_257),
.Y(n_2353)
);

AOI22xp5_ASAP7_75t_L g2354 ( 
.A1(n_1892),
.A2(n_260),
.B1(n_258),
.B2(n_259),
.Y(n_2354)
);

NOR3xp33_ASAP7_75t_SL g2355 ( 
.A(n_1820),
.B(n_259),
.C(n_261),
.Y(n_2355)
);

AOI21xp5_ASAP7_75t_L g2356 ( 
.A1(n_1770),
.A2(n_261),
.B(n_262),
.Y(n_2356)
);

INVx3_ASAP7_75t_L g2357 ( 
.A(n_1890),
.Y(n_2357)
);

BUFx6f_ASAP7_75t_L g2358 ( 
.A(n_1776),
.Y(n_2358)
);

NOR3xp33_ASAP7_75t_SL g2359 ( 
.A(n_1820),
.B(n_263),
.C(n_265),
.Y(n_2359)
);

AO21x1_ASAP7_75t_L g2360 ( 
.A1(n_1777),
.A2(n_265),
.B(n_266),
.Y(n_2360)
);

AOI21xp5_ASAP7_75t_L g2361 ( 
.A1(n_1770),
.A2(n_267),
.B(n_268),
.Y(n_2361)
);

INVx3_ASAP7_75t_L g2362 ( 
.A(n_1890),
.Y(n_2362)
);

INVx1_ASAP7_75t_SL g2363 ( 
.A(n_1807),
.Y(n_2363)
);

NAND2xp5_ASAP7_75t_SL g2364 ( 
.A(n_1793),
.B(n_267),
.Y(n_2364)
);

NAND2xp5_ASAP7_75t_L g2365 ( 
.A(n_1751),
.B(n_269),
.Y(n_2365)
);

AOI21xp5_ASAP7_75t_L g2366 ( 
.A1(n_1770),
.A2(n_269),
.B(n_270),
.Y(n_2366)
);

AOI22xp5_ASAP7_75t_L g2367 ( 
.A1(n_1892),
.A2(n_273),
.B1(n_270),
.B2(n_272),
.Y(n_2367)
);

NAND2xp5_ASAP7_75t_L g2368 ( 
.A(n_1751),
.B(n_273),
.Y(n_2368)
);

AND2x2_ASAP7_75t_SL g2369 ( 
.A(n_1843),
.B(n_274),
.Y(n_2369)
);

NOR2xp33_ASAP7_75t_L g2370 ( 
.A(n_1752),
.B(n_275),
.Y(n_2370)
);

AOI21xp5_ASAP7_75t_L g2371 ( 
.A1(n_1770),
.A2(n_276),
.B(n_277),
.Y(n_2371)
);

INVx2_ASAP7_75t_L g2372 ( 
.A(n_1877),
.Y(n_2372)
);

BUFx12f_ASAP7_75t_L g2373 ( 
.A(n_1788),
.Y(n_2373)
);

OAI22xp5_ASAP7_75t_L g2374 ( 
.A1(n_1938),
.A2(n_284),
.B1(n_281),
.B2(n_282),
.Y(n_2374)
);

BUFx6f_ASAP7_75t_L g2375 ( 
.A(n_1776),
.Y(n_2375)
);

INVx2_ASAP7_75t_L g2376 ( 
.A(n_1877),
.Y(n_2376)
);

NAND2xp5_ASAP7_75t_L g2377 ( 
.A(n_1751),
.B(n_281),
.Y(n_2377)
);

NAND2xp5_ASAP7_75t_SL g2378 ( 
.A(n_1793),
.B(n_282),
.Y(n_2378)
);

NAND2xp5_ASAP7_75t_L g2379 ( 
.A(n_1751),
.B(n_285),
.Y(n_2379)
);

BUFx2_ASAP7_75t_L g2380 ( 
.A(n_1843),
.Y(n_2380)
);

NAND2xp5_ASAP7_75t_L g2381 ( 
.A(n_1751),
.B(n_286),
.Y(n_2381)
);

NOR2xp33_ASAP7_75t_L g2382 ( 
.A(n_1752),
.B(n_287),
.Y(n_2382)
);

NAND2xp5_ASAP7_75t_L g2383 ( 
.A(n_1751),
.B(n_288),
.Y(n_2383)
);

BUFx4f_ASAP7_75t_L g2384 ( 
.A(n_1736),
.Y(n_2384)
);

OAI22xp5_ASAP7_75t_L g2385 ( 
.A1(n_1938),
.A2(n_292),
.B1(n_289),
.B2(n_290),
.Y(n_2385)
);

INVx1_ASAP7_75t_L g2386 ( 
.A(n_1751),
.Y(n_2386)
);

CKINVDCx6p67_ASAP7_75t_R g2387 ( 
.A(n_1785),
.Y(n_2387)
);

NAND2xp5_ASAP7_75t_SL g2388 ( 
.A(n_1793),
.B(n_298),
.Y(n_2388)
);

OAI22xp5_ASAP7_75t_L g2389 ( 
.A1(n_1938),
.A2(n_302),
.B1(n_299),
.B2(n_301),
.Y(n_2389)
);

AOI21xp5_ASAP7_75t_L g2390 ( 
.A1(n_1770),
.A2(n_303),
.B(n_304),
.Y(n_2390)
);

NAND2xp5_ASAP7_75t_SL g2391 ( 
.A(n_1793),
.B(n_303),
.Y(n_2391)
);

BUFx6f_ASAP7_75t_L g2392 ( 
.A(n_1776),
.Y(n_2392)
);

AND2x2_ASAP7_75t_L g2393 ( 
.A(n_1793),
.B(n_304),
.Y(n_2393)
);

INVx1_ASAP7_75t_L g2394 ( 
.A(n_1751),
.Y(n_2394)
);

BUFx2_ASAP7_75t_L g2395 ( 
.A(n_1843),
.Y(n_2395)
);

A2O1A1Ixp33_ASAP7_75t_L g2396 ( 
.A1(n_1817),
.A2(n_307),
.B(n_305),
.C(n_306),
.Y(n_2396)
);

AOI21x1_ASAP7_75t_L g2397 ( 
.A1(n_1777),
.A2(n_305),
.B(n_307),
.Y(n_2397)
);

OAI22xp5_ASAP7_75t_L g2398 ( 
.A1(n_1938),
.A2(n_310),
.B1(n_308),
.B2(n_309),
.Y(n_2398)
);

NAND3xp33_ASAP7_75t_L g2399 ( 
.A(n_1908),
.B(n_309),
.C(n_311),
.Y(n_2399)
);

INVx2_ASAP7_75t_L g2400 ( 
.A(n_1877),
.Y(n_2400)
);

AOI21xp5_ASAP7_75t_L g2401 ( 
.A1(n_1770),
.A2(n_312),
.B(n_313),
.Y(n_2401)
);

INVx4_ASAP7_75t_L g2402 ( 
.A(n_1740),
.Y(n_2402)
);

INVx1_ASAP7_75t_L g2403 ( 
.A(n_1751),
.Y(n_2403)
);

CKINVDCx5p33_ASAP7_75t_R g2404 ( 
.A(n_1761),
.Y(n_2404)
);

NOR2xp33_ASAP7_75t_R g2405 ( 
.A(n_1761),
.B(n_314),
.Y(n_2405)
);

NAND2xp5_ASAP7_75t_L g2406 ( 
.A(n_1751),
.B(n_314),
.Y(n_2406)
);

NAND2xp5_ASAP7_75t_L g2407 ( 
.A(n_1751),
.B(n_315),
.Y(n_2407)
);

INVx1_ASAP7_75t_L g2408 ( 
.A(n_1751),
.Y(n_2408)
);

INVx1_ASAP7_75t_L g2409 ( 
.A(n_1751),
.Y(n_2409)
);

NOR2xp33_ASAP7_75t_L g2410 ( 
.A(n_1752),
.B(n_316),
.Y(n_2410)
);

INVx1_ASAP7_75t_L g2411 ( 
.A(n_1751),
.Y(n_2411)
);

NAND2xp5_ASAP7_75t_SL g2412 ( 
.A(n_1793),
.B(n_317),
.Y(n_2412)
);

INVx5_ASAP7_75t_L g2413 ( 
.A(n_1779),
.Y(n_2413)
);

NAND2xp5_ASAP7_75t_SL g2414 ( 
.A(n_1793),
.B(n_317),
.Y(n_2414)
);

INVx1_ASAP7_75t_L g2415 ( 
.A(n_1751),
.Y(n_2415)
);

NAND2xp5_ASAP7_75t_L g2416 ( 
.A(n_1751),
.B(n_319),
.Y(n_2416)
);

NOR2xp33_ASAP7_75t_L g2417 ( 
.A(n_1752),
.B(n_321),
.Y(n_2417)
);

INVx1_ASAP7_75t_L g2418 ( 
.A(n_1751),
.Y(n_2418)
);

NAND3xp33_ASAP7_75t_L g2419 ( 
.A(n_1908),
.B(n_321),
.C(n_322),
.Y(n_2419)
);

AND2x2_ASAP7_75t_L g2420 ( 
.A(n_1793),
.B(n_323),
.Y(n_2420)
);

AOI221xp5_ASAP7_75t_L g2421 ( 
.A1(n_1809),
.A2(n_325),
.B1(n_323),
.B2(n_324),
.C(n_326),
.Y(n_2421)
);

NAND2xp5_ASAP7_75t_L g2422 ( 
.A(n_1751),
.B(n_327),
.Y(n_2422)
);

NAND2xp5_ASAP7_75t_L g2423 ( 
.A(n_1751),
.B(n_327),
.Y(n_2423)
);

AOI21xp5_ASAP7_75t_L g2424 ( 
.A1(n_1770),
.A2(n_328),
.B(n_329),
.Y(n_2424)
);

A2O1A1Ixp33_ASAP7_75t_SL g2425 ( 
.A1(n_1812),
.A2(n_332),
.B(n_330),
.C(n_331),
.Y(n_2425)
);

INVx1_ASAP7_75t_SL g2426 ( 
.A(n_1807),
.Y(n_2426)
);

BUFx3_ASAP7_75t_L g2427 ( 
.A(n_1740),
.Y(n_2427)
);

A2O1A1Ixp33_ASAP7_75t_L g2428 ( 
.A1(n_1817),
.A2(n_334),
.B(n_331),
.C(n_333),
.Y(n_2428)
);

A2O1A1Ixp33_ASAP7_75t_L g2429 ( 
.A1(n_1817),
.A2(n_336),
.B(n_334),
.C(n_335),
.Y(n_2429)
);

NOR2xp33_ASAP7_75t_L g2430 ( 
.A(n_1752),
.B(n_336),
.Y(n_2430)
);

A2O1A1Ixp33_ASAP7_75t_SL g2431 ( 
.A1(n_1812),
.A2(n_341),
.B(n_337),
.C(n_340),
.Y(n_2431)
);

AO21x2_ASAP7_75t_L g2432 ( 
.A1(n_1770),
.A2(n_342),
.B(n_343),
.Y(n_2432)
);

NAND2x1p5_ASAP7_75t_L g2433 ( 
.A(n_1878),
.B(n_342),
.Y(n_2433)
);

INVx1_ASAP7_75t_L g2434 ( 
.A(n_2025),
.Y(n_2434)
);

NAND2x1_ASAP7_75t_L g2435 ( 
.A(n_2199),
.B(n_347),
.Y(n_2435)
);

BUFx12f_ASAP7_75t_L g2436 ( 
.A(n_2051),
.Y(n_2436)
);

INVx1_ASAP7_75t_L g2437 ( 
.A(n_2319),
.Y(n_2437)
);

BUFx6f_ASAP7_75t_L g2438 ( 
.A(n_2310),
.Y(n_2438)
);

A2O1A1Ixp33_ASAP7_75t_L g2439 ( 
.A1(n_2173),
.A2(n_351),
.B(n_348),
.C(n_349),
.Y(n_2439)
);

BUFx2_ASAP7_75t_R g2440 ( 
.A(n_2031),
.Y(n_2440)
);

BUFx3_ASAP7_75t_L g2441 ( 
.A(n_2067),
.Y(n_2441)
);

HB1xp67_ASAP7_75t_L g2442 ( 
.A(n_2230),
.Y(n_2442)
);

NAND2xp5_ASAP7_75t_L g2443 ( 
.A(n_2055),
.B(n_352),
.Y(n_2443)
);

BUFx12f_ASAP7_75t_L g2444 ( 
.A(n_2346),
.Y(n_2444)
);

AOI22x1_ASAP7_75t_L g2445 ( 
.A1(n_2044),
.A2(n_354),
.B1(n_352),
.B2(n_353),
.Y(n_2445)
);

AND2x6_ASAP7_75t_L g2446 ( 
.A(n_2113),
.B(n_640),
.Y(n_2446)
);

INVx2_ASAP7_75t_L g2447 ( 
.A(n_2019),
.Y(n_2447)
);

HB1xp67_ASAP7_75t_L g2448 ( 
.A(n_2182),
.Y(n_2448)
);

BUFx8_ASAP7_75t_L g2449 ( 
.A(n_2033),
.Y(n_2449)
);

BUFx3_ASAP7_75t_L g2450 ( 
.A(n_2061),
.Y(n_2450)
);

INVx2_ASAP7_75t_L g2451 ( 
.A(n_2336),
.Y(n_2451)
);

BUFx6f_ASAP7_75t_L g2452 ( 
.A(n_2269),
.Y(n_2452)
);

INVx4_ASAP7_75t_L g2453 ( 
.A(n_2387),
.Y(n_2453)
);

INVx2_ASAP7_75t_L g2454 ( 
.A(n_2340),
.Y(n_2454)
);

AO21x2_ASAP7_75t_L g2455 ( 
.A1(n_2334),
.A2(n_353),
.B(n_354),
.Y(n_2455)
);

BUFx6f_ASAP7_75t_L g2456 ( 
.A(n_2269),
.Y(n_2456)
);

INVx1_ASAP7_75t_L g2457 ( 
.A(n_2325),
.Y(n_2457)
);

BUFx6f_ASAP7_75t_L g2458 ( 
.A(n_2269),
.Y(n_2458)
);

INVx1_ASAP7_75t_L g2459 ( 
.A(n_2343),
.Y(n_2459)
);

NAND2x1p5_ASAP7_75t_L g2460 ( 
.A(n_2413),
.B(n_2239),
.Y(n_2460)
);

INVx2_ASAP7_75t_L g2461 ( 
.A(n_2344),
.Y(n_2461)
);

INVx2_ASAP7_75t_L g2462 ( 
.A(n_2351),
.Y(n_2462)
);

INVx2_ASAP7_75t_L g2463 ( 
.A(n_2372),
.Y(n_2463)
);

INVx1_ASAP7_75t_L g2464 ( 
.A(n_2386),
.Y(n_2464)
);

INVx4_ASAP7_75t_SL g2465 ( 
.A(n_2307),
.Y(n_2465)
);

INVx1_ASAP7_75t_SL g2466 ( 
.A(n_2363),
.Y(n_2466)
);

BUFx6f_ASAP7_75t_SL g2467 ( 
.A(n_2079),
.Y(n_2467)
);

NOR2xp33_ASAP7_75t_L g2468 ( 
.A(n_2096),
.B(n_356),
.Y(n_2468)
);

BUFx3_ASAP7_75t_L g2469 ( 
.A(n_2427),
.Y(n_2469)
);

NAND2xp5_ASAP7_75t_L g2470 ( 
.A(n_2076),
.B(n_359),
.Y(n_2470)
);

INVx1_ASAP7_75t_L g2471 ( 
.A(n_2394),
.Y(n_2471)
);

BUFx8_ASAP7_75t_L g2472 ( 
.A(n_2033),
.Y(n_2472)
);

NAND2xp5_ASAP7_75t_L g2473 ( 
.A(n_2231),
.B(n_360),
.Y(n_2473)
);

AND2x4_ASAP7_75t_L g2474 ( 
.A(n_2234),
.B(n_362),
.Y(n_2474)
);

AO21x2_ASAP7_75t_L g2475 ( 
.A1(n_2432),
.A2(n_363),
.B(n_364),
.Y(n_2475)
);

CKINVDCx14_ASAP7_75t_R g2476 ( 
.A(n_2373),
.Y(n_2476)
);

OAI21xp5_ASAP7_75t_L g2477 ( 
.A1(n_2129),
.A2(n_365),
.B(n_366),
.Y(n_2477)
);

INVx3_ASAP7_75t_L g2478 ( 
.A(n_2196),
.Y(n_2478)
);

INVx2_ASAP7_75t_L g2479 ( 
.A(n_2376),
.Y(n_2479)
);

INVx1_ASAP7_75t_L g2480 ( 
.A(n_2403),
.Y(n_2480)
);

INVx2_ASAP7_75t_L g2481 ( 
.A(n_2400),
.Y(n_2481)
);

AO21x2_ASAP7_75t_L g2482 ( 
.A1(n_2432),
.A2(n_366),
.B(n_367),
.Y(n_2482)
);

CKINVDCx5p33_ASAP7_75t_R g2483 ( 
.A(n_2084),
.Y(n_2483)
);

INVx1_ASAP7_75t_L g2484 ( 
.A(n_2408),
.Y(n_2484)
);

BUFx3_ASAP7_75t_L g2485 ( 
.A(n_2042),
.Y(n_2485)
);

INVx2_ASAP7_75t_L g2486 ( 
.A(n_2039),
.Y(n_2486)
);

INVx3_ASAP7_75t_L g2487 ( 
.A(n_2196),
.Y(n_2487)
);

BUFx3_ASAP7_75t_L g2488 ( 
.A(n_2187),
.Y(n_2488)
);

NAND2xp5_ASAP7_75t_L g2489 ( 
.A(n_2254),
.B(n_368),
.Y(n_2489)
);

INVx1_ASAP7_75t_L g2490 ( 
.A(n_2409),
.Y(n_2490)
);

INVx1_ASAP7_75t_L g2491 ( 
.A(n_2411),
.Y(n_2491)
);

BUFx6f_ASAP7_75t_L g2492 ( 
.A(n_2043),
.Y(n_2492)
);

AO21x2_ASAP7_75t_L g2493 ( 
.A1(n_2338),
.A2(n_369),
.B(n_370),
.Y(n_2493)
);

CKINVDCx20_ASAP7_75t_R g2494 ( 
.A(n_2328),
.Y(n_2494)
);

BUFx12f_ASAP7_75t_L g2495 ( 
.A(n_2404),
.Y(n_2495)
);

INVx1_ASAP7_75t_L g2496 ( 
.A(n_2415),
.Y(n_2496)
);

INVx6_ASAP7_75t_L g2497 ( 
.A(n_2347),
.Y(n_2497)
);

INVx4_ASAP7_75t_L g2498 ( 
.A(n_2347),
.Y(n_2498)
);

BUFx3_ASAP7_75t_L g2499 ( 
.A(n_2187),
.Y(n_2499)
);

INVx2_ASAP7_75t_L g2500 ( 
.A(n_2248),
.Y(n_2500)
);

BUFx3_ASAP7_75t_L g2501 ( 
.A(n_2402),
.Y(n_2501)
);

INVx5_ASAP7_75t_L g2502 ( 
.A(n_2402),
.Y(n_2502)
);

INVx6_ASAP7_75t_L g2503 ( 
.A(n_2097),
.Y(n_2503)
);

AO21x2_ASAP7_75t_L g2504 ( 
.A1(n_2397),
.A2(n_372),
.B(n_373),
.Y(n_2504)
);

BUFx3_ASAP7_75t_L g2505 ( 
.A(n_2092),
.Y(n_2505)
);

NAND2x1p5_ASAP7_75t_L g2506 ( 
.A(n_2413),
.B(n_2239),
.Y(n_2506)
);

OAI21x1_ASAP7_75t_L g2507 ( 
.A1(n_2059),
.A2(n_373),
.B(n_376),
.Y(n_2507)
);

INVx1_ASAP7_75t_L g2508 ( 
.A(n_2418),
.Y(n_2508)
);

NAND2x1p5_ASAP7_75t_L g2509 ( 
.A(n_2413),
.B(n_376),
.Y(n_2509)
);

AND2x2_ASAP7_75t_L g2510 ( 
.A(n_2363),
.B(n_377),
.Y(n_2510)
);

AO21x2_ASAP7_75t_L g2511 ( 
.A1(n_2313),
.A2(n_377),
.B(n_378),
.Y(n_2511)
);

BUFx2_ASAP7_75t_R g2512 ( 
.A(n_2327),
.Y(n_2512)
);

OAI22x1_ASAP7_75t_L g2513 ( 
.A1(n_2433),
.A2(n_381),
.B1(n_379),
.B2(n_380),
.Y(n_2513)
);

NAND2xp5_ASAP7_75t_L g2514 ( 
.A(n_2119),
.B(n_379),
.Y(n_2514)
);

INVx2_ASAP7_75t_L g2515 ( 
.A(n_2123),
.Y(n_2515)
);

AND2x4_ASAP7_75t_L g2516 ( 
.A(n_2199),
.B(n_2203),
.Y(n_2516)
);

AOI22xp33_ASAP7_75t_SL g2517 ( 
.A1(n_2369),
.A2(n_384),
.B1(n_382),
.B2(n_383),
.Y(n_2517)
);

INVx1_ASAP7_75t_SL g2518 ( 
.A(n_2426),
.Y(n_2518)
);

NAND2x1p5_ASAP7_75t_L g2519 ( 
.A(n_2098),
.B(n_385),
.Y(n_2519)
);

AO21x2_ASAP7_75t_L g2520 ( 
.A1(n_2316),
.A2(n_385),
.B(n_386),
.Y(n_2520)
);

AO21x2_ASAP7_75t_L g2521 ( 
.A1(n_2318),
.A2(n_387),
.B(n_388),
.Y(n_2521)
);

AND2x2_ASAP7_75t_L g2522 ( 
.A(n_2426),
.B(n_387),
.Y(n_2522)
);

INVx5_ASAP7_75t_L g2523 ( 
.A(n_2098),
.Y(n_2523)
);

BUFx3_ASAP7_75t_L g2524 ( 
.A(n_2024),
.Y(n_2524)
);

OAI21x1_ASAP7_75t_L g2525 ( 
.A1(n_2243),
.A2(n_388),
.B(n_389),
.Y(n_2525)
);

INVx1_ASAP7_75t_L g2526 ( 
.A(n_2037),
.Y(n_2526)
);

AOI22x1_ASAP7_75t_L g2527 ( 
.A1(n_2246),
.A2(n_392),
.B1(n_390),
.B2(n_391),
.Y(n_2527)
);

OAI21xp5_ASAP7_75t_L g2528 ( 
.A1(n_2135),
.A2(n_392),
.B(n_393),
.Y(n_2528)
);

AO21x2_ASAP7_75t_L g2529 ( 
.A1(n_2330),
.A2(n_393),
.B(n_394),
.Y(n_2529)
);

AO21x2_ASAP7_75t_L g2530 ( 
.A1(n_2337),
.A2(n_394),
.B(n_395),
.Y(n_2530)
);

INVx2_ASAP7_75t_L g2531 ( 
.A(n_2170),
.Y(n_2531)
);

NOR2xp33_ASAP7_75t_L g2532 ( 
.A(n_2032),
.B(n_2260),
.Y(n_2532)
);

BUFx3_ASAP7_75t_L g2533 ( 
.A(n_2329),
.Y(n_2533)
);

NOR2xp33_ASAP7_75t_L g2534 ( 
.A(n_2090),
.B(n_395),
.Y(n_2534)
);

AOI21xp5_ASAP7_75t_L g2535 ( 
.A1(n_2045),
.A2(n_397),
.B(n_398),
.Y(n_2535)
);

OAI21x1_ASAP7_75t_SL g2536 ( 
.A1(n_2290),
.A2(n_397),
.B(n_399),
.Y(n_2536)
);

INVxp67_ASAP7_75t_L g2537 ( 
.A(n_2380),
.Y(n_2537)
);

INVx3_ASAP7_75t_L g2538 ( 
.A(n_2203),
.Y(n_2538)
);

BUFx2_ASAP7_75t_L g2539 ( 
.A(n_2395),
.Y(n_2539)
);

NAND2xp5_ASAP7_75t_L g2540 ( 
.A(n_2118),
.B(n_400),
.Y(n_2540)
);

BUFx2_ASAP7_75t_L g2541 ( 
.A(n_2223),
.Y(n_2541)
);

NAND2xp5_ASAP7_75t_SL g2542 ( 
.A(n_2063),
.B(n_2244),
.Y(n_2542)
);

AND2x4_ASAP7_75t_L g2543 ( 
.A(n_2106),
.B(n_400),
.Y(n_2543)
);

AOI22x1_ASAP7_75t_L g2544 ( 
.A1(n_2093),
.A2(n_403),
.B1(n_401),
.B2(n_402),
.Y(n_2544)
);

BUFx2_ASAP7_75t_L g2545 ( 
.A(n_2267),
.Y(n_2545)
);

AND2x2_ASAP7_75t_L g2546 ( 
.A(n_2038),
.B(n_401),
.Y(n_2546)
);

INVx1_ASAP7_75t_SL g2547 ( 
.A(n_2066),
.Y(n_2547)
);

HB1xp67_ASAP7_75t_L g2548 ( 
.A(n_2275),
.Y(n_2548)
);

NOR2xp33_ASAP7_75t_L g2549 ( 
.A(n_2251),
.B(n_405),
.Y(n_2549)
);

INVx2_ASAP7_75t_L g2550 ( 
.A(n_2171),
.Y(n_2550)
);

AND2x4_ASAP7_75t_L g2551 ( 
.A(n_2106),
.B(n_407),
.Y(n_2551)
);

AO21x2_ASAP7_75t_L g2552 ( 
.A1(n_2356),
.A2(n_407),
.B(n_409),
.Y(n_2552)
);

NAND2xp5_ASAP7_75t_L g2553 ( 
.A(n_2133),
.B(n_409),
.Y(n_2553)
);

AND2x2_ASAP7_75t_L g2554 ( 
.A(n_2255),
.B(n_2018),
.Y(n_2554)
);

AND2x2_ASAP7_75t_L g2555 ( 
.A(n_2086),
.B(n_410),
.Y(n_2555)
);

CKINVDCx16_ASAP7_75t_R g2556 ( 
.A(n_2405),
.Y(n_2556)
);

INVx3_ASAP7_75t_L g2557 ( 
.A(n_2142),
.Y(n_2557)
);

BUFx2_ASAP7_75t_R g2558 ( 
.A(n_2087),
.Y(n_2558)
);

HB1xp67_ASAP7_75t_L g2559 ( 
.A(n_2275),
.Y(n_2559)
);

INVx1_ASAP7_75t_L g2560 ( 
.A(n_2174),
.Y(n_2560)
);

BUFx12f_ASAP7_75t_L g2561 ( 
.A(n_2100),
.Y(n_2561)
);

INVx1_ASAP7_75t_L g2562 ( 
.A(n_2180),
.Y(n_2562)
);

NAND2x1p5_ASAP7_75t_L g2563 ( 
.A(n_2142),
.B(n_412),
.Y(n_2563)
);

INVxp67_ASAP7_75t_SL g2564 ( 
.A(n_2043),
.Y(n_2564)
);

AND2x4_ASAP7_75t_L g2565 ( 
.A(n_2155),
.B(n_412),
.Y(n_2565)
);

BUFx3_ASAP7_75t_L g2566 ( 
.A(n_2384),
.Y(n_2566)
);

OAI22xp33_ASAP7_75t_SL g2567 ( 
.A1(n_2339),
.A2(n_416),
.B1(n_414),
.B2(n_415),
.Y(n_2567)
);

AO21x2_ASAP7_75t_L g2568 ( 
.A1(n_2361),
.A2(n_414),
.B(n_415),
.Y(n_2568)
);

BUFx3_ASAP7_75t_L g2569 ( 
.A(n_2384),
.Y(n_2569)
);

INVx2_ASAP7_75t_L g2570 ( 
.A(n_2188),
.Y(n_2570)
);

INVx3_ASAP7_75t_L g2571 ( 
.A(n_2250),
.Y(n_2571)
);

BUFx2_ASAP7_75t_SL g2572 ( 
.A(n_2224),
.Y(n_2572)
);

INVx1_ASAP7_75t_L g2573 ( 
.A(n_2315),
.Y(n_2573)
);

INVx1_ASAP7_75t_L g2574 ( 
.A(n_2317),
.Y(n_2574)
);

INVx1_ASAP7_75t_L g2575 ( 
.A(n_2326),
.Y(n_2575)
);

OAI21xp5_ASAP7_75t_L g2576 ( 
.A1(n_2135),
.A2(n_417),
.B(n_418),
.Y(n_2576)
);

INVx1_ASAP7_75t_L g2577 ( 
.A(n_2332),
.Y(n_2577)
);

OAI21x1_ASAP7_75t_L g2578 ( 
.A1(n_2159),
.A2(n_417),
.B(n_418),
.Y(n_2578)
);

AO21x2_ASAP7_75t_L g2579 ( 
.A1(n_2366),
.A2(n_419),
.B(n_420),
.Y(n_2579)
);

BUFx3_ASAP7_75t_L g2580 ( 
.A(n_2268),
.Y(n_2580)
);

BUFx2_ASAP7_75t_L g2581 ( 
.A(n_2292),
.Y(n_2581)
);

OR2x2_ASAP7_75t_L g2582 ( 
.A(n_2204),
.B(n_421),
.Y(n_2582)
);

AO22x1_ASAP7_75t_L g2583 ( 
.A1(n_2094),
.A2(n_424),
.B1(n_422),
.B2(n_423),
.Y(n_2583)
);

BUFx2_ASAP7_75t_SL g2584 ( 
.A(n_2264),
.Y(n_2584)
);

INVx8_ASAP7_75t_L g2585 ( 
.A(n_2186),
.Y(n_2585)
);

NAND2x1p5_ASAP7_75t_L g2586 ( 
.A(n_2250),
.B(n_422),
.Y(n_2586)
);

INVx3_ASAP7_75t_L g2587 ( 
.A(n_2048),
.Y(n_2587)
);

BUFx2_ASAP7_75t_R g2588 ( 
.A(n_2216),
.Y(n_2588)
);

AND2x4_ASAP7_75t_L g2589 ( 
.A(n_2179),
.B(n_424),
.Y(n_2589)
);

INVx1_ASAP7_75t_SL g2590 ( 
.A(n_2066),
.Y(n_2590)
);

OAI21x1_ASAP7_75t_L g2591 ( 
.A1(n_2311),
.A2(n_425),
.B(n_426),
.Y(n_2591)
);

BUFx3_ASAP7_75t_L g2592 ( 
.A(n_2235),
.Y(n_2592)
);

BUFx3_ASAP7_75t_L g2593 ( 
.A(n_2114),
.Y(n_2593)
);

BUFx10_ASAP7_75t_L g2594 ( 
.A(n_2264),
.Y(n_2594)
);

AOI21xp5_ASAP7_75t_L g2595 ( 
.A1(n_2046),
.A2(n_426),
.B(n_427),
.Y(n_2595)
);

INVx3_ASAP7_75t_L g2596 ( 
.A(n_2048),
.Y(n_2596)
);

INVx8_ASAP7_75t_L g2597 ( 
.A(n_2186),
.Y(n_2597)
);

NAND2xp5_ASAP7_75t_SL g2598 ( 
.A(n_2115),
.B(n_427),
.Y(n_2598)
);

NOR2xp33_ASAP7_75t_L g2599 ( 
.A(n_2168),
.B(n_428),
.Y(n_2599)
);

NAND2x1p5_ASAP7_75t_L g2600 ( 
.A(n_2275),
.B(n_429),
.Y(n_2600)
);

INVx4_ASAP7_75t_L g2601 ( 
.A(n_2186),
.Y(n_2601)
);

AO21x2_ASAP7_75t_L g2602 ( 
.A1(n_2371),
.A2(n_429),
.B(n_430),
.Y(n_2602)
);

INVx6_ASAP7_75t_SL g2603 ( 
.A(n_2088),
.Y(n_2603)
);

NOR2xp33_ASAP7_75t_L g2604 ( 
.A(n_2209),
.B(n_432),
.Y(n_2604)
);

NAND2xp5_ASAP7_75t_L g2605 ( 
.A(n_2020),
.B(n_433),
.Y(n_2605)
);

INVx2_ASAP7_75t_SL g2606 ( 
.A(n_2150),
.Y(n_2606)
);

INVx5_ASAP7_75t_L g2607 ( 
.A(n_2075),
.Y(n_2607)
);

AOI21xp5_ASAP7_75t_L g2608 ( 
.A1(n_2020),
.A2(n_437),
.B(n_438),
.Y(n_2608)
);

INVx8_ASAP7_75t_L g2609 ( 
.A(n_2088),
.Y(n_2609)
);

INVxp67_ASAP7_75t_SL g2610 ( 
.A(n_2075),
.Y(n_2610)
);

CKINVDCx5p33_ASAP7_75t_R g2611 ( 
.A(n_2120),
.Y(n_2611)
);

INVxp67_ASAP7_75t_SL g2612 ( 
.A(n_2102),
.Y(n_2612)
);

AOI22xp5_ASAP7_75t_L g2613 ( 
.A1(n_2030),
.A2(n_443),
.B1(n_439),
.B2(n_442),
.Y(n_2613)
);

BUFx2_ASAP7_75t_L g2614 ( 
.A(n_2137),
.Y(n_2614)
);

INVx1_ASAP7_75t_SL g2615 ( 
.A(n_2242),
.Y(n_2615)
);

NAND2xp5_ASAP7_75t_L g2616 ( 
.A(n_2227),
.B(n_442),
.Y(n_2616)
);

NAND2xp5_ASAP7_75t_L g2617 ( 
.A(n_2263),
.B(n_443),
.Y(n_2617)
);

CKINVDCx20_ASAP7_75t_R g2618 ( 
.A(n_2302),
.Y(n_2618)
);

INVx3_ASAP7_75t_L g2619 ( 
.A(n_2078),
.Y(n_2619)
);

INVx1_ASAP7_75t_L g2620 ( 
.A(n_2333),
.Y(n_2620)
);

BUFx3_ASAP7_75t_L g2621 ( 
.A(n_2078),
.Y(n_2621)
);

AND2x4_ASAP7_75t_L g2622 ( 
.A(n_2321),
.B(n_446),
.Y(n_2622)
);

BUFx2_ASAP7_75t_L g2623 ( 
.A(n_2183),
.Y(n_2623)
);

INVx1_ASAP7_75t_L g2624 ( 
.A(n_2342),
.Y(n_2624)
);

INVx1_ASAP7_75t_L g2625 ( 
.A(n_2350),
.Y(n_2625)
);

BUFx12f_ASAP7_75t_L g2626 ( 
.A(n_2125),
.Y(n_2626)
);

AO21x2_ASAP7_75t_L g2627 ( 
.A1(n_2390),
.A2(n_447),
.B(n_449),
.Y(n_2627)
);

BUFx3_ASAP7_75t_L g2628 ( 
.A(n_2321),
.Y(n_2628)
);

BUFx3_ASAP7_75t_L g2629 ( 
.A(n_2357),
.Y(n_2629)
);

OAI21xp5_ASAP7_75t_L g2630 ( 
.A1(n_2027),
.A2(n_450),
.B(n_451),
.Y(n_2630)
);

AOI22xp33_ASAP7_75t_L g2631 ( 
.A1(n_2052),
.A2(n_452),
.B1(n_450),
.B2(n_451),
.Y(n_2631)
);

BUFx2_ASAP7_75t_L g2632 ( 
.A(n_2195),
.Y(n_2632)
);

AND2x2_ASAP7_75t_L g2633 ( 
.A(n_2091),
.B(n_453),
.Y(n_2633)
);

BUFx3_ASAP7_75t_L g2634 ( 
.A(n_2357),
.Y(n_2634)
);

INVx2_ASAP7_75t_SL g2635 ( 
.A(n_2362),
.Y(n_2635)
);

INVx1_ASAP7_75t_L g2636 ( 
.A(n_2365),
.Y(n_2636)
);

AO21x2_ASAP7_75t_L g2637 ( 
.A1(n_2401),
.A2(n_453),
.B(n_454),
.Y(n_2637)
);

INVx1_ASAP7_75t_SL g2638 ( 
.A(n_2222),
.Y(n_2638)
);

BUFx3_ASAP7_75t_L g2639 ( 
.A(n_2362),
.Y(n_2639)
);

INVx2_ASAP7_75t_SL g2640 ( 
.A(n_2277),
.Y(n_2640)
);

INVx1_ASAP7_75t_SL g2641 ( 
.A(n_2241),
.Y(n_2641)
);

INVx4_ASAP7_75t_SL g2642 ( 
.A(n_2139),
.Y(n_2642)
);

INVx1_ASAP7_75t_L g2643 ( 
.A(n_2368),
.Y(n_2643)
);

INVx2_ASAP7_75t_L g2644 ( 
.A(n_2103),
.Y(n_2644)
);

INVx4_ASAP7_75t_L g2645 ( 
.A(n_2433),
.Y(n_2645)
);

INVx1_ASAP7_75t_L g2646 ( 
.A(n_2377),
.Y(n_2646)
);

INVx1_ASAP7_75t_L g2647 ( 
.A(n_2379),
.Y(n_2647)
);

AOI22xp33_ASAP7_75t_L g2648 ( 
.A1(n_2052),
.A2(n_2165),
.B1(n_2121),
.B2(n_2140),
.Y(n_2648)
);

BUFx2_ASAP7_75t_SL g2649 ( 
.A(n_2277),
.Y(n_2649)
);

INVx2_ASAP7_75t_SL g2650 ( 
.A(n_2265),
.Y(n_2650)
);

BUFx3_ASAP7_75t_L g2651 ( 
.A(n_2271),
.Y(n_2651)
);

BUFx3_ASAP7_75t_L g2652 ( 
.A(n_2252),
.Y(n_2652)
);

INVx3_ASAP7_75t_SL g2653 ( 
.A(n_2152),
.Y(n_2653)
);

CKINVDCx20_ASAP7_75t_R g2654 ( 
.A(n_2056),
.Y(n_2654)
);

OAI21xp5_ASAP7_75t_L g2655 ( 
.A1(n_2424),
.A2(n_455),
.B(n_458),
.Y(n_2655)
);

AO21x1_ASAP7_75t_L g2656 ( 
.A1(n_2290),
.A2(n_460),
.B(n_461),
.Y(n_2656)
);

OR2x4_ASAP7_75t_L g2657 ( 
.A(n_2035),
.B(n_460),
.Y(n_2657)
);

INVx1_ASAP7_75t_L g2658 ( 
.A(n_2381),
.Y(n_2658)
);

BUFx4_ASAP7_75t_SL g2659 ( 
.A(n_2163),
.Y(n_2659)
);

BUFx3_ASAP7_75t_L g2660 ( 
.A(n_2252),
.Y(n_2660)
);

AO21x1_ASAP7_75t_L g2661 ( 
.A1(n_2068),
.A2(n_461),
.B(n_462),
.Y(n_2661)
);

NAND2x1p5_ASAP7_75t_L g2662 ( 
.A(n_2249),
.B(n_462),
.Y(n_2662)
);

HB1xp67_ASAP7_75t_L g2663 ( 
.A(n_2169),
.Y(n_2663)
);

INVx1_ASAP7_75t_L g2664 ( 
.A(n_2383),
.Y(n_2664)
);

INVx2_ASAP7_75t_SL g2665 ( 
.A(n_2172),
.Y(n_2665)
);

CKINVDCx16_ASAP7_75t_R g2666 ( 
.A(n_2151),
.Y(n_2666)
);

INVx4_ASAP7_75t_L g2667 ( 
.A(n_2139),
.Y(n_2667)
);

OA21x2_ASAP7_75t_L g2668 ( 
.A1(n_2345),
.A2(n_464),
.B(n_465),
.Y(n_2668)
);

BUFx2_ASAP7_75t_L g2669 ( 
.A(n_2205),
.Y(n_2669)
);

OA21x2_ASAP7_75t_L g2670 ( 
.A1(n_2348),
.A2(n_466),
.B(n_467),
.Y(n_2670)
);

OR2x6_ASAP7_75t_L g2671 ( 
.A(n_2113),
.B(n_466),
.Y(n_2671)
);

INVx2_ASAP7_75t_L g2672 ( 
.A(n_2122),
.Y(n_2672)
);

OAI21x1_ASAP7_75t_SL g2673 ( 
.A1(n_2082),
.A2(n_469),
.B(n_470),
.Y(n_2673)
);

INVx1_ASAP7_75t_L g2674 ( 
.A(n_2406),
.Y(n_2674)
);

BUFx4_ASAP7_75t_SL g2675 ( 
.A(n_2191),
.Y(n_2675)
);

BUFx3_ASAP7_75t_L g2676 ( 
.A(n_2107),
.Y(n_2676)
);

BUFx5_ASAP7_75t_L g2677 ( 
.A(n_2279),
.Y(n_2677)
);

OAI21x1_ASAP7_75t_SL g2678 ( 
.A1(n_2339),
.A2(n_2367),
.B(n_2354),
.Y(n_2678)
);

INVx1_ASAP7_75t_L g2679 ( 
.A(n_2407),
.Y(n_2679)
);

AND2x2_ASAP7_75t_L g2680 ( 
.A(n_2189),
.B(n_471),
.Y(n_2680)
);

INVx2_ASAP7_75t_L g2681 ( 
.A(n_2130),
.Y(n_2681)
);

INVx2_ASAP7_75t_L g2682 ( 
.A(n_2194),
.Y(n_2682)
);

BUFx3_ASAP7_75t_L g2683 ( 
.A(n_2205),
.Y(n_2683)
);

BUFx2_ASAP7_75t_L g2684 ( 
.A(n_2116),
.Y(n_2684)
);

INVx1_ASAP7_75t_L g2685 ( 
.A(n_2416),
.Y(n_2685)
);

OAI21xp5_ASAP7_75t_L g2686 ( 
.A1(n_2040),
.A2(n_2021),
.B(n_2041),
.Y(n_2686)
);

INVx2_ASAP7_75t_SL g2687 ( 
.A(n_2116),
.Y(n_2687)
);

INVx1_ASAP7_75t_L g2688 ( 
.A(n_2422),
.Y(n_2688)
);

AND2x2_ASAP7_75t_L g2689 ( 
.A(n_2262),
.B(n_473),
.Y(n_2689)
);

INVx6_ASAP7_75t_L g2690 ( 
.A(n_2280),
.Y(n_2690)
);

AND2x2_ASAP7_75t_L g2691 ( 
.A(n_2028),
.B(n_474),
.Y(n_2691)
);

INVx1_ASAP7_75t_L g2692 ( 
.A(n_2423),
.Y(n_2692)
);

AND2x2_ASAP7_75t_L g2693 ( 
.A(n_2341),
.B(n_474),
.Y(n_2693)
);

BUFx3_ASAP7_75t_L g2694 ( 
.A(n_2083),
.Y(n_2694)
);

AO21x2_ASAP7_75t_L g2695 ( 
.A1(n_2360),
.A2(n_475),
.B(n_476),
.Y(n_2695)
);

INVx1_ASAP7_75t_SL g2696 ( 
.A(n_2161),
.Y(n_2696)
);

NAND2xp5_ASAP7_75t_L g2697 ( 
.A(n_2190),
.B(n_476),
.Y(n_2697)
);

CKINVDCx20_ASAP7_75t_R g2698 ( 
.A(n_2110),
.Y(n_2698)
);

OAI21xp5_ASAP7_75t_L g2699 ( 
.A1(n_2050),
.A2(n_477),
.B(n_478),
.Y(n_2699)
);

BUFx3_ASAP7_75t_L g2700 ( 
.A(n_2295),
.Y(n_2700)
);

AOI22x1_ASAP7_75t_L g2701 ( 
.A1(n_2167),
.A2(n_477),
.B1(n_479),
.B2(n_480),
.Y(n_2701)
);

INVx5_ASAP7_75t_L g2702 ( 
.A(n_2161),
.Y(n_2702)
);

INVx8_ASAP7_75t_L g2703 ( 
.A(n_2161),
.Y(n_2703)
);

INVx5_ASAP7_75t_L g2704 ( 
.A(n_2288),
.Y(n_2704)
);

OAI21x1_ASAP7_75t_L g2705 ( 
.A1(n_2309),
.A2(n_480),
.B(n_481),
.Y(n_2705)
);

INVx1_ASAP7_75t_SL g2706 ( 
.A(n_2288),
.Y(n_2706)
);

INVx2_ASAP7_75t_L g2707 ( 
.A(n_2206),
.Y(n_2707)
);

AOI31xp33_ASAP7_75t_L g2708 ( 
.A1(n_2068),
.A2(n_481),
.A3(n_482),
.B(n_483),
.Y(n_2708)
);

NAND2xp5_ASAP7_75t_L g2709 ( 
.A(n_2211),
.B(n_483),
.Y(n_2709)
);

AND2x2_ASAP7_75t_L g2710 ( 
.A(n_2349),
.B(n_484),
.Y(n_2710)
);

INVxp67_ASAP7_75t_SL g2711 ( 
.A(n_2314),
.Y(n_2711)
);

NAND2x1p5_ASAP7_75t_L g2712 ( 
.A(n_2249),
.B(n_484),
.Y(n_2712)
);

INVx2_ASAP7_75t_L g2713 ( 
.A(n_2212),
.Y(n_2713)
);

OAI21xp5_ASAP7_75t_L g2714 ( 
.A1(n_2073),
.A2(n_485),
.B(n_486),
.Y(n_2714)
);

INVx3_ASAP7_75t_SL g2715 ( 
.A(n_2280),
.Y(n_2715)
);

OAI21x1_ASAP7_75t_L g2716 ( 
.A1(n_2309),
.A2(n_485),
.B(n_487),
.Y(n_2716)
);

INVx1_ASAP7_75t_L g2717 ( 
.A(n_2074),
.Y(n_2717)
);

OAI21x1_ASAP7_75t_L g2718 ( 
.A1(n_2221),
.A2(n_488),
.B(n_489),
.Y(n_2718)
);

NAND2x1p5_ASAP7_75t_L g2719 ( 
.A(n_2273),
.B(n_488),
.Y(n_2719)
);

AO21x2_ASAP7_75t_L g2720 ( 
.A1(n_2425),
.A2(n_490),
.B(n_492),
.Y(n_2720)
);

OAI21xp5_ASAP7_75t_L g2721 ( 
.A1(n_2278),
.A2(n_490),
.B(n_492),
.Y(n_2721)
);

NAND2x1p5_ASAP7_75t_L g2722 ( 
.A(n_2273),
.B(n_493),
.Y(n_2722)
);

BUFx3_ASAP7_75t_L g2723 ( 
.A(n_2352),
.Y(n_2723)
);

INVx1_ASAP7_75t_L g2724 ( 
.A(n_2214),
.Y(n_2724)
);

BUFx12f_ASAP7_75t_L g2725 ( 
.A(n_2026),
.Y(n_2725)
);

BUFx10_ASAP7_75t_L g2726 ( 
.A(n_2229),
.Y(n_2726)
);

BUFx10_ASAP7_75t_L g2727 ( 
.A(n_2126),
.Y(n_2727)
);

CKINVDCx20_ASAP7_75t_R g2728 ( 
.A(n_2036),
.Y(n_2728)
);

BUFx3_ASAP7_75t_L g2729 ( 
.A(n_2393),
.Y(n_2729)
);

AOI22x1_ASAP7_75t_L g2730 ( 
.A1(n_2272),
.A2(n_496),
.B1(n_497),
.B2(n_498),
.Y(n_2730)
);

BUFx8_ASAP7_75t_L g2731 ( 
.A(n_2047),
.Y(n_2731)
);

BUFx2_ASAP7_75t_L g2732 ( 
.A(n_2095),
.Y(n_2732)
);

INVx6_ASAP7_75t_L g2733 ( 
.A(n_2420),
.Y(n_2733)
);

HB1xp67_ASAP7_75t_L g2734 ( 
.A(n_2358),
.Y(n_2734)
);

NOR2xp33_ASAP7_75t_L g2735 ( 
.A(n_2266),
.B(n_2029),
.Y(n_2735)
);

BUFx3_ASAP7_75t_L g2736 ( 
.A(n_2219),
.Y(n_2736)
);

NOR2xp33_ASAP7_75t_L g2737 ( 
.A(n_2276),
.B(n_2105),
.Y(n_2737)
);

BUFx2_ASAP7_75t_L g2738 ( 
.A(n_2111),
.Y(n_2738)
);

INVx6_ASAP7_75t_L g2739 ( 
.A(n_2358),
.Y(n_2739)
);

NAND3xp33_ASAP7_75t_L g2740 ( 
.A(n_2200),
.B(n_499),
.C(n_500),
.Y(n_2740)
);

INVx3_ASAP7_75t_L g2741 ( 
.A(n_2375),
.Y(n_2741)
);

OR3x4_ASAP7_75t_SL g2742 ( 
.A(n_2355),
.B(n_2359),
.C(n_2220),
.Y(n_2742)
);

BUFx2_ASAP7_75t_L g2743 ( 
.A(n_2226),
.Y(n_2743)
);

INVx1_ASAP7_75t_L g2744 ( 
.A(n_2201),
.Y(n_2744)
);

NOR2xp33_ASAP7_75t_R g2745 ( 
.A(n_2297),
.B(n_502),
.Y(n_2745)
);

AO21x2_ASAP7_75t_L g2746 ( 
.A1(n_2431),
.A2(n_503),
.B(n_504),
.Y(n_2746)
);

NAND2x1p5_ASAP7_75t_L g2747 ( 
.A(n_2392),
.B(n_505),
.Y(n_2747)
);

OAI21xp5_ASAP7_75t_L g2748 ( 
.A1(n_2213),
.A2(n_506),
.B(n_507),
.Y(n_2748)
);

NAND2xp5_ASAP7_75t_L g2749 ( 
.A(n_2247),
.B(n_507),
.Y(n_2749)
);

NAND2x1p5_ASAP7_75t_L g2750 ( 
.A(n_2392),
.B(n_508),
.Y(n_2750)
);

AND2x2_ASAP7_75t_L g2751 ( 
.A(n_2253),
.B(n_508),
.Y(n_2751)
);

BUFx4f_ASAP7_75t_SL g2752 ( 
.A(n_2132),
.Y(n_2752)
);

INVx1_ASAP7_75t_L g2753 ( 
.A(n_2202),
.Y(n_2753)
);

INVx2_ASAP7_75t_L g2754 ( 
.A(n_2301),
.Y(n_2754)
);

BUFx10_ASAP7_75t_L g2755 ( 
.A(n_2299),
.Y(n_2755)
);

HB1xp67_ASAP7_75t_L g2756 ( 
.A(n_2300),
.Y(n_2756)
);

AO21x2_ASAP7_75t_L g2757 ( 
.A1(n_2283),
.A2(n_509),
.B(n_510),
.Y(n_2757)
);

CKINVDCx8_ASAP7_75t_R g2758 ( 
.A(n_2057),
.Y(n_2758)
);

BUFx3_ASAP7_75t_L g2759 ( 
.A(n_2274),
.Y(n_2759)
);

NAND3xp33_ASAP7_75t_L g2760 ( 
.A(n_2127),
.B(n_510),
.C(n_511),
.Y(n_2760)
);

INVx2_ASAP7_75t_SL g2761 ( 
.A(n_2149),
.Y(n_2761)
);

INVx3_ASAP7_75t_L g2762 ( 
.A(n_2143),
.Y(n_2762)
);

INVx1_ASAP7_75t_L g2763 ( 
.A(n_2034),
.Y(n_2763)
);

INVx3_ASAP7_75t_L g2764 ( 
.A(n_2153),
.Y(n_2764)
);

BUFx2_ASAP7_75t_R g2765 ( 
.A(n_2146),
.Y(n_2765)
);

BUFx2_ASAP7_75t_L g2766 ( 
.A(n_2085),
.Y(n_2766)
);

BUFx12f_ASAP7_75t_L g2767 ( 
.A(n_2236),
.Y(n_2767)
);

BUFx3_ASAP7_75t_L g2768 ( 
.A(n_2240),
.Y(n_2768)
);

INVx1_ASAP7_75t_SL g2769 ( 
.A(n_2136),
.Y(n_2769)
);

AND2x4_ASAP7_75t_L g2770 ( 
.A(n_2305),
.B(n_511),
.Y(n_2770)
);

OA21x2_ASAP7_75t_L g2771 ( 
.A1(n_2283),
.A2(n_512),
.B(n_513),
.Y(n_2771)
);

CKINVDCx11_ASAP7_75t_R g2772 ( 
.A(n_2053),
.Y(n_2772)
);

AOI22xp33_ASAP7_75t_L g2773 ( 
.A1(n_2165),
.A2(n_2144),
.B1(n_2323),
.B2(n_2322),
.Y(n_2773)
);

AND2x2_ASAP7_75t_L g2774 ( 
.A(n_2245),
.B(n_514),
.Y(n_2774)
);

AOI21xp5_ASAP7_75t_L g2775 ( 
.A1(n_2134),
.A2(n_515),
.B(n_517),
.Y(n_2775)
);

INVx1_ASAP7_75t_L g2776 ( 
.A(n_2147),
.Y(n_2776)
);

INVx2_ASAP7_75t_L g2777 ( 
.A(n_2293),
.Y(n_2777)
);

AOI22x1_ASAP7_75t_L g2778 ( 
.A1(n_2238),
.A2(n_515),
.B1(n_518),
.B2(n_520),
.Y(n_2778)
);

AO21x2_ASAP7_75t_L g2779 ( 
.A1(n_2303),
.A2(n_518),
.B(n_521),
.Y(n_2779)
);

INVx1_ASAP7_75t_L g2780 ( 
.A(n_2164),
.Y(n_2780)
);

OA21x2_ASAP7_75t_L g2781 ( 
.A1(n_2258),
.A2(n_521),
.B(n_524),
.Y(n_2781)
);

CKINVDCx6p67_ASAP7_75t_R g2782 ( 
.A(n_2072),
.Y(n_2782)
);

OAI21x1_ASAP7_75t_L g2783 ( 
.A1(n_2312),
.A2(n_524),
.B(n_525),
.Y(n_2783)
);

AND2x4_ASAP7_75t_L g2784 ( 
.A(n_2060),
.B(n_525),
.Y(n_2784)
);

AND2x2_ASAP7_75t_L g2785 ( 
.A(n_2109),
.B(n_526),
.Y(n_2785)
);

BUFx10_ASAP7_75t_L g2786 ( 
.A(n_2259),
.Y(n_2786)
);

AND2x4_ASAP7_75t_L g2787 ( 
.A(n_2166),
.B(n_526),
.Y(n_2787)
);

BUFx6f_ASAP7_75t_L g2788 ( 
.A(n_2154),
.Y(n_2788)
);

AO21x2_ASAP7_75t_L g2789 ( 
.A1(n_2399),
.A2(n_527),
.B(n_529),
.Y(n_2789)
);

HB1xp67_ASAP7_75t_L g2790 ( 
.A(n_2175),
.Y(n_2790)
);

INVxp67_ASAP7_75t_SL g2791 ( 
.A(n_2354),
.Y(n_2791)
);

OAI21x1_ASAP7_75t_L g2792 ( 
.A1(n_2178),
.A2(n_531),
.B(n_532),
.Y(n_2792)
);

NAND2xp5_ASAP7_75t_L g2793 ( 
.A(n_2207),
.B(n_533),
.Y(n_2793)
);

BUFx2_ASAP7_75t_SL g2794 ( 
.A(n_2298),
.Y(n_2794)
);

NAND2x1p5_ASAP7_75t_L g2795 ( 
.A(n_2058),
.B(n_534),
.Y(n_2795)
);

INVx3_ASAP7_75t_L g2796 ( 
.A(n_2304),
.Y(n_2796)
);

OR3x4_ASAP7_75t_SL g2797 ( 
.A(n_2158),
.B(n_2069),
.C(n_2197),
.Y(n_2797)
);

BUFx2_ASAP7_75t_L g2798 ( 
.A(n_2117),
.Y(n_2798)
);

INVx1_ASAP7_75t_L g2799 ( 
.A(n_2367),
.Y(n_2799)
);

NAND2x1p5_ASAP7_75t_L g2800 ( 
.A(n_2062),
.B(n_536),
.Y(n_2800)
);

OAI21x1_ASAP7_75t_L g2801 ( 
.A1(n_2320),
.A2(n_537),
.B(n_538),
.Y(n_2801)
);

INVx2_ASAP7_75t_L g2802 ( 
.A(n_2486),
.Y(n_2802)
);

INVx1_ASAP7_75t_L g2803 ( 
.A(n_2434),
.Y(n_2803)
);

INVx1_ASAP7_75t_L g2804 ( 
.A(n_2437),
.Y(n_2804)
);

INVx1_ASAP7_75t_L g2805 ( 
.A(n_2457),
.Y(n_2805)
);

AO21x1_ASAP7_75t_L g2806 ( 
.A1(n_2708),
.A2(n_2101),
.B(n_2127),
.Y(n_2806)
);

INVx2_ASAP7_75t_L g2807 ( 
.A(n_2500),
.Y(n_2807)
);

INVx1_ASAP7_75t_L g2808 ( 
.A(n_2459),
.Y(n_2808)
);

INVx1_ASAP7_75t_L g2809 ( 
.A(n_2464),
.Y(n_2809)
);

INVx1_ASAP7_75t_L g2810 ( 
.A(n_2471),
.Y(n_2810)
);

INVx1_ASAP7_75t_L g2811 ( 
.A(n_2480),
.Y(n_2811)
);

INVx1_ASAP7_75t_L g2812 ( 
.A(n_2484),
.Y(n_2812)
);

INVx2_ASAP7_75t_L g2813 ( 
.A(n_2515),
.Y(n_2813)
);

INVx2_ASAP7_75t_L g2814 ( 
.A(n_2531),
.Y(n_2814)
);

AO21x1_ASAP7_75t_SL g2815 ( 
.A1(n_2548),
.A2(n_2559),
.B(n_2442),
.Y(n_2815)
);

AND2x2_ASAP7_75t_L g2816 ( 
.A(n_2554),
.B(n_2691),
.Y(n_2816)
);

BUFx12f_ASAP7_75t_L g2817 ( 
.A(n_2449),
.Y(n_2817)
);

INVx1_ASAP7_75t_L g2818 ( 
.A(n_2490),
.Y(n_2818)
);

AO21x1_ASAP7_75t_SL g2819 ( 
.A1(n_2548),
.A2(n_2296),
.B(n_2184),
.Y(n_2819)
);

OAI22xp5_ASAP7_75t_SL g2820 ( 
.A1(n_2654),
.A2(n_2335),
.B1(n_2353),
.B2(n_2324),
.Y(n_2820)
);

INVx1_ASAP7_75t_L g2821 ( 
.A(n_2491),
.Y(n_2821)
);

INVx8_ASAP7_75t_L g2822 ( 
.A(n_2502),
.Y(n_2822)
);

HB1xp67_ASAP7_75t_L g2823 ( 
.A(n_2448),
.Y(n_2823)
);

INVx2_ASAP7_75t_L g2824 ( 
.A(n_2550),
.Y(n_2824)
);

INVx1_ASAP7_75t_L g2825 ( 
.A(n_2496),
.Y(n_2825)
);

NAND2x1p5_ASAP7_75t_L g2826 ( 
.A(n_2502),
.B(n_2198),
.Y(n_2826)
);

INVx1_ASAP7_75t_L g2827 ( 
.A(n_2508),
.Y(n_2827)
);

INVx1_ASAP7_75t_L g2828 ( 
.A(n_2526),
.Y(n_2828)
);

INVx1_ASAP7_75t_L g2829 ( 
.A(n_2560),
.Y(n_2829)
);

INVx2_ASAP7_75t_L g2830 ( 
.A(n_2570),
.Y(n_2830)
);

OAI22xp5_ASAP7_75t_L g2831 ( 
.A1(n_2671),
.A2(n_2296),
.B1(n_2419),
.B2(n_2399),
.Y(n_2831)
);

INVx2_ASAP7_75t_L g2832 ( 
.A(n_2447),
.Y(n_2832)
);

NAND2x1p5_ASAP7_75t_L g2833 ( 
.A(n_2502),
.B(n_2193),
.Y(n_2833)
);

OAI22xp33_ASAP7_75t_L g2834 ( 
.A1(n_2671),
.A2(n_2065),
.B1(n_2289),
.B2(n_2192),
.Y(n_2834)
);

CKINVDCx20_ASAP7_75t_R g2835 ( 
.A(n_2494),
.Y(n_2835)
);

AND2x2_ASAP7_75t_L g2836 ( 
.A(n_2756),
.B(n_2156),
.Y(n_2836)
);

AOI22xp5_ASAP7_75t_L g2837 ( 
.A1(n_2735),
.A2(n_2370),
.B1(n_2410),
.B2(n_2382),
.Y(n_2837)
);

HB1xp67_ASAP7_75t_L g2838 ( 
.A(n_2448),
.Y(n_2838)
);

INVx6_ASAP7_75t_L g2839 ( 
.A(n_2438),
.Y(n_2839)
);

INVx1_ASAP7_75t_L g2840 ( 
.A(n_2562),
.Y(n_2840)
);

AOI22xp33_ASAP7_75t_L g2841 ( 
.A1(n_2678),
.A2(n_2417),
.B1(n_2430),
.B2(n_2228),
.Y(n_2841)
);

OAI22xp5_ASAP7_75t_L g2842 ( 
.A1(n_2671),
.A2(n_2054),
.B1(n_2208),
.B2(n_2176),
.Y(n_2842)
);

INVx3_ASAP7_75t_L g2843 ( 
.A(n_2645),
.Y(n_2843)
);

INVx2_ASAP7_75t_L g2844 ( 
.A(n_2451),
.Y(n_2844)
);

INVx3_ASAP7_75t_L g2845 ( 
.A(n_2645),
.Y(n_2845)
);

CKINVDCx5p33_ASAP7_75t_R g2846 ( 
.A(n_2483),
.Y(n_2846)
);

INVx2_ASAP7_75t_L g2847 ( 
.A(n_2454),
.Y(n_2847)
);

INVx2_ASAP7_75t_L g2848 ( 
.A(n_2461),
.Y(n_2848)
);

OAI22xp5_ASAP7_75t_L g2849 ( 
.A1(n_2648),
.A2(n_2181),
.B1(n_2145),
.B2(n_2294),
.Y(n_2849)
);

AOI22xp33_ASAP7_75t_L g2850 ( 
.A1(n_2648),
.A2(n_2217),
.B1(n_2218),
.B2(n_2210),
.Y(n_2850)
);

INVx2_ASAP7_75t_L g2851 ( 
.A(n_2462),
.Y(n_2851)
);

INVx1_ASAP7_75t_SL g2852 ( 
.A(n_2501),
.Y(n_2852)
);

INVx2_ASAP7_75t_L g2853 ( 
.A(n_2463),
.Y(n_2853)
);

INVx1_ASAP7_75t_L g2854 ( 
.A(n_2443),
.Y(n_2854)
);

INVx1_ASAP7_75t_L g2855 ( 
.A(n_2470),
.Y(n_2855)
);

INVx2_ASAP7_75t_L g2856 ( 
.A(n_2479),
.Y(n_2856)
);

INVx1_ASAP7_75t_L g2857 ( 
.A(n_2470),
.Y(n_2857)
);

CKINVDCx5p33_ASAP7_75t_R g2858 ( 
.A(n_2449),
.Y(n_2858)
);

INVx2_ASAP7_75t_L g2859 ( 
.A(n_2481),
.Y(n_2859)
);

AOI22xp33_ASAP7_75t_L g2860 ( 
.A1(n_2791),
.A2(n_2256),
.B1(n_2185),
.B2(n_2141),
.Y(n_2860)
);

BUFx6f_ASAP7_75t_L g2861 ( 
.A(n_2452),
.Y(n_2861)
);

AO21x1_ASAP7_75t_L g2862 ( 
.A1(n_2708),
.A2(n_2281),
.B(n_2331),
.Y(n_2862)
);

HB1xp67_ASAP7_75t_L g2863 ( 
.A(n_2466),
.Y(n_2863)
);

BUFx3_ASAP7_75t_L g2864 ( 
.A(n_2438),
.Y(n_2864)
);

CKINVDCx5p33_ASAP7_75t_R g2865 ( 
.A(n_2472),
.Y(n_2865)
);

AOI22xp5_ASAP7_75t_L g2866 ( 
.A1(n_2532),
.A2(n_2284),
.B1(n_2177),
.B2(n_2287),
.Y(n_2866)
);

AOI22xp33_ASAP7_75t_L g2867 ( 
.A1(n_2791),
.A2(n_2799),
.B1(n_2772),
.B2(n_2446),
.Y(n_2867)
);

CKINVDCx20_ASAP7_75t_R g2868 ( 
.A(n_2472),
.Y(n_2868)
);

NAND2xp5_ASAP7_75t_L g2869 ( 
.A(n_2468),
.B(n_2737),
.Y(n_2869)
);

AOI22xp33_ASAP7_75t_SL g2870 ( 
.A1(n_2585),
.A2(n_2385),
.B1(n_2374),
.B2(n_2389),
.Y(n_2870)
);

AND2x4_ASAP7_75t_L g2871 ( 
.A(n_2478),
.B(n_2099),
.Y(n_2871)
);

BUFx2_ASAP7_75t_SL g2872 ( 
.A(n_2453),
.Y(n_2872)
);

AOI22xp5_ASAP7_75t_L g2873 ( 
.A1(n_2446),
.A2(n_2767),
.B1(n_2725),
.B2(n_2474),
.Y(n_2873)
);

BUFx3_ASAP7_75t_L g2874 ( 
.A(n_2438),
.Y(n_2874)
);

INVx4_ASAP7_75t_L g2875 ( 
.A(n_2453),
.Y(n_2875)
);

INVx1_ASAP7_75t_L g2876 ( 
.A(n_2514),
.Y(n_2876)
);

OAI21xp5_ASAP7_75t_L g2877 ( 
.A1(n_2773),
.A2(n_2237),
.B(n_2023),
.Y(n_2877)
);

AOI22xp33_ASAP7_75t_L g2878 ( 
.A1(n_2446),
.A2(n_2364),
.B1(n_2378),
.B2(n_2414),
.Y(n_2878)
);

CKINVDCx5p33_ASAP7_75t_R g2879 ( 
.A(n_2436),
.Y(n_2879)
);

CKINVDCx11_ASAP7_75t_R g2880 ( 
.A(n_2444),
.Y(n_2880)
);

INVx1_ASAP7_75t_L g2881 ( 
.A(n_2553),
.Y(n_2881)
);

OAI22xp5_ASAP7_75t_L g2882 ( 
.A1(n_2649),
.A2(n_2631),
.B1(n_2715),
.B2(n_2609),
.Y(n_2882)
);

AND2x4_ASAP7_75t_L g2883 ( 
.A(n_2478),
.B(n_2104),
.Y(n_2883)
);

AOI22xp5_ASAP7_75t_L g2884 ( 
.A1(n_2446),
.A2(n_2233),
.B1(n_2388),
.B2(n_2412),
.Y(n_2884)
);

NAND2x1p5_ASAP7_75t_L g2885 ( 
.A(n_2498),
.B(n_2391),
.Y(n_2885)
);

BUFx2_ASAP7_75t_L g2886 ( 
.A(n_2603),
.Y(n_2886)
);

OAI22xp5_ASAP7_75t_L g2887 ( 
.A1(n_2631),
.A2(n_2215),
.B1(n_2162),
.B2(n_2428),
.Y(n_2887)
);

BUFx3_ASAP7_75t_L g2888 ( 
.A(n_2469),
.Y(n_2888)
);

NOR2xp33_ASAP7_75t_L g2889 ( 
.A(n_2601),
.B(n_2261),
.Y(n_2889)
);

AND2x4_ASAP7_75t_L g2890 ( 
.A(n_2487),
.B(n_2108),
.Y(n_2890)
);

AOI22xp33_ASAP7_75t_L g2891 ( 
.A1(n_2756),
.A2(n_2308),
.B1(n_2421),
.B2(n_2232),
.Y(n_2891)
);

INVx1_ASAP7_75t_L g2892 ( 
.A(n_2475),
.Y(n_2892)
);

NAND2xp5_ASAP7_75t_L g2893 ( 
.A(n_2689),
.B(n_2022),
.Y(n_2893)
);

AOI22xp33_ASAP7_75t_SL g2894 ( 
.A1(n_2585),
.A2(n_2398),
.B1(n_2124),
.B2(n_2112),
.Y(n_2894)
);

INVx1_ASAP7_75t_L g2895 ( 
.A(n_2475),
.Y(n_2895)
);

INVx1_ASAP7_75t_L g2896 ( 
.A(n_2482),
.Y(n_2896)
);

INVx2_ASAP7_75t_L g2897 ( 
.A(n_2644),
.Y(n_2897)
);

AND2x2_ASAP7_75t_L g2898 ( 
.A(n_2546),
.B(n_2047),
.Y(n_2898)
);

INVx3_ASAP7_75t_L g2899 ( 
.A(n_2487),
.Y(n_2899)
);

AOI22xp5_ASAP7_75t_L g2900 ( 
.A1(n_2474),
.A2(n_2770),
.B1(n_2690),
.B2(n_2751),
.Y(n_2900)
);

INVx1_ASAP7_75t_L g2901 ( 
.A(n_2553),
.Y(n_2901)
);

AOI22xp33_ASAP7_75t_L g2902 ( 
.A1(n_2585),
.A2(n_2282),
.B1(n_2285),
.B2(n_2286),
.Y(n_2902)
);

CKINVDCx11_ASAP7_75t_R g2903 ( 
.A(n_2495),
.Y(n_2903)
);

INVx2_ASAP7_75t_L g2904 ( 
.A(n_2672),
.Y(n_2904)
);

INVx2_ASAP7_75t_L g2905 ( 
.A(n_2681),
.Y(n_2905)
);

INVx2_ASAP7_75t_L g2906 ( 
.A(n_2682),
.Y(n_2906)
);

INVx4_ASAP7_75t_L g2907 ( 
.A(n_2465),
.Y(n_2907)
);

INVx1_ASAP7_75t_SL g2908 ( 
.A(n_2497),
.Y(n_2908)
);

BUFx8_ASAP7_75t_L g2909 ( 
.A(n_2467),
.Y(n_2909)
);

CKINVDCx20_ASAP7_75t_R g2910 ( 
.A(n_2476),
.Y(n_2910)
);

AND2x4_ASAP7_75t_L g2911 ( 
.A(n_2601),
.B(n_2396),
.Y(n_2911)
);

OAI21x1_ASAP7_75t_SL g2912 ( 
.A1(n_2528),
.A2(n_2131),
.B(n_2148),
.Y(n_2912)
);

NOR2xp33_ASAP7_75t_L g2913 ( 
.A(n_2758),
.B(n_2306),
.Y(n_2913)
);

OAI21xp5_ASAP7_75t_L g2914 ( 
.A1(n_2773),
.A2(n_2429),
.B(n_2157),
.Y(n_2914)
);

INVx1_ASAP7_75t_L g2915 ( 
.A(n_2617),
.Y(n_2915)
);

AOI22xp33_ASAP7_75t_L g2916 ( 
.A1(n_2597),
.A2(n_2782),
.B1(n_2690),
.B2(n_2770),
.Y(n_2916)
);

INVx2_ASAP7_75t_L g2917 ( 
.A(n_2707),
.Y(n_2917)
);

NAND2xp5_ASAP7_75t_L g2918 ( 
.A(n_2604),
.B(n_2762),
.Y(n_2918)
);

BUFx2_ASAP7_75t_L g2919 ( 
.A(n_2603),
.Y(n_2919)
);

INVx1_ASAP7_75t_L g2920 ( 
.A(n_2754),
.Y(n_2920)
);

CKINVDCx20_ASAP7_75t_R g2921 ( 
.A(n_2441),
.Y(n_2921)
);

CKINVDCx20_ASAP7_75t_R g2922 ( 
.A(n_2618),
.Y(n_2922)
);

INVx2_ASAP7_75t_L g2923 ( 
.A(n_2713),
.Y(n_2923)
);

BUFx2_ASAP7_75t_L g2924 ( 
.A(n_2498),
.Y(n_2924)
);

AND2x2_ASAP7_75t_L g2925 ( 
.A(n_2466),
.B(n_2047),
.Y(n_2925)
);

AO21x1_ASAP7_75t_L g2926 ( 
.A1(n_2567),
.A2(n_2257),
.B(n_2225),
.Y(n_2926)
);

NAND2xp5_ASAP7_75t_L g2927 ( 
.A(n_2762),
.B(n_2160),
.Y(n_2927)
);

HB1xp67_ASAP7_75t_L g2928 ( 
.A(n_2518),
.Y(n_2928)
);

NAND2x1p5_ASAP7_75t_L g2929 ( 
.A(n_2566),
.B(n_2569),
.Y(n_2929)
);

INVx2_ASAP7_75t_L g2930 ( 
.A(n_2724),
.Y(n_2930)
);

INVx1_ASAP7_75t_L g2931 ( 
.A(n_2473),
.Y(n_2931)
);

BUFx2_ASAP7_75t_R g2932 ( 
.A(n_2611),
.Y(n_2932)
);

INVx1_ASAP7_75t_L g2933 ( 
.A(n_2473),
.Y(n_2933)
);

OAI22xp5_ASAP7_75t_L g2934 ( 
.A1(n_2609),
.A2(n_2049),
.B1(n_2080),
.B2(n_2071),
.Y(n_2934)
);

INVx3_ASAP7_75t_L g2935 ( 
.A(n_2523),
.Y(n_2935)
);

INVx1_ASAP7_75t_L g2936 ( 
.A(n_2489),
.Y(n_2936)
);

AOI22xp5_ASAP7_75t_L g2937 ( 
.A1(n_2761),
.A2(n_2070),
.B1(n_2089),
.B2(n_2081),
.Y(n_2937)
);

INVx1_ASAP7_75t_L g2938 ( 
.A(n_2489),
.Y(n_2938)
);

INVx1_ASAP7_75t_L g2939 ( 
.A(n_2697),
.Y(n_2939)
);

BUFx3_ASAP7_75t_L g2940 ( 
.A(n_2497),
.Y(n_2940)
);

HB1xp67_ASAP7_75t_L g2941 ( 
.A(n_2518),
.Y(n_2941)
);

NAND2x1p5_ASAP7_75t_L g2942 ( 
.A(n_2523),
.B(n_2270),
.Y(n_2942)
);

NAND2x1p5_ASAP7_75t_L g2943 ( 
.A(n_2523),
.B(n_2270),
.Y(n_2943)
);

BUFx12f_ASAP7_75t_L g2944 ( 
.A(n_2626),
.Y(n_2944)
);

NAND2xp5_ASAP7_75t_L g2945 ( 
.A(n_2684),
.B(n_2077),
.Y(n_2945)
);

INVx3_ASAP7_75t_L g2946 ( 
.A(n_2460),
.Y(n_2946)
);

OAI22xp5_ASAP7_75t_L g2947 ( 
.A1(n_2609),
.A2(n_2064),
.B1(n_2128),
.B2(n_2291),
.Y(n_2947)
);

INVx1_ASAP7_75t_L g2948 ( 
.A(n_2616),
.Y(n_2948)
);

INVx2_ASAP7_75t_L g2949 ( 
.A(n_2743),
.Y(n_2949)
);

BUFx6f_ASAP7_75t_SL g2950 ( 
.A(n_2594),
.Y(n_2950)
);

INVx1_ASAP7_75t_L g2951 ( 
.A(n_2482),
.Y(n_2951)
);

NAND2xp5_ASAP7_75t_L g2952 ( 
.A(n_2776),
.B(n_2687),
.Y(n_2952)
);

AOI22xp33_ASAP7_75t_L g2953 ( 
.A1(n_2597),
.A2(n_2138),
.B1(n_540),
.B2(n_541),
.Y(n_2953)
);

INVx1_ASAP7_75t_L g2954 ( 
.A(n_2455),
.Y(n_2954)
);

INVx1_ASAP7_75t_L g2955 ( 
.A(n_2455),
.Y(n_2955)
);

BUFx2_ASAP7_75t_L g2956 ( 
.A(n_2465),
.Y(n_2956)
);

BUFx3_ASAP7_75t_L g2957 ( 
.A(n_2505),
.Y(n_2957)
);

OAI22xp5_ASAP7_75t_L g2958 ( 
.A1(n_2597),
.A2(n_537),
.B1(n_541),
.B2(n_542),
.Y(n_2958)
);

BUFx3_ASAP7_75t_L g2959 ( 
.A(n_2450),
.Y(n_2959)
);

INVx2_ASAP7_75t_L g2960 ( 
.A(n_2736),
.Y(n_2960)
);

INVx11_ASAP7_75t_L g2961 ( 
.A(n_2561),
.Y(n_2961)
);

OAI22xp5_ASAP7_75t_L g2962 ( 
.A1(n_2517),
.A2(n_545),
.B1(n_546),
.B2(n_547),
.Y(n_2962)
);

OAI21x1_ASAP7_75t_SL g2963 ( 
.A1(n_2576),
.A2(n_545),
.B(n_546),
.Y(n_2963)
);

AND2x2_ASAP7_75t_L g2964 ( 
.A(n_2510),
.B(n_547),
.Y(n_2964)
);

INVx1_ASAP7_75t_L g2965 ( 
.A(n_2591),
.Y(n_2965)
);

OAI22xp5_ASAP7_75t_L g2966 ( 
.A1(n_2517),
.A2(n_548),
.B1(n_549),
.B2(n_550),
.Y(n_2966)
);

AOI22xp33_ASAP7_75t_L g2967 ( 
.A1(n_2768),
.A2(n_549),
.B1(n_550),
.B2(n_551),
.Y(n_2967)
);

OA21x2_ASAP7_75t_L g2968 ( 
.A1(n_2477),
.A2(n_551),
.B(n_552),
.Y(n_2968)
);

INVx3_ASAP7_75t_L g2969 ( 
.A(n_2460),
.Y(n_2969)
);

AOI22xp33_ASAP7_75t_L g2970 ( 
.A1(n_2764),
.A2(n_552),
.B1(n_553),
.B2(n_554),
.Y(n_2970)
);

AOI22xp33_ASAP7_75t_L g2971 ( 
.A1(n_2764),
.A2(n_554),
.B1(n_555),
.B2(n_556),
.Y(n_2971)
);

INVx1_ASAP7_75t_L g2972 ( 
.A(n_2668),
.Y(n_2972)
);

BUFx3_ASAP7_75t_L g2973 ( 
.A(n_2485),
.Y(n_2973)
);

INVx1_ASAP7_75t_L g2974 ( 
.A(n_2668),
.Y(n_2974)
);

NAND2xp5_ASAP7_75t_L g2975 ( 
.A(n_2763),
.B(n_640),
.Y(n_2975)
);

INVx1_ASAP7_75t_L g2976 ( 
.A(n_2670),
.Y(n_2976)
);

INVx1_ASAP7_75t_L g2977 ( 
.A(n_2670),
.Y(n_2977)
);

CKINVDCx6p67_ASAP7_75t_R g2978 ( 
.A(n_2467),
.Y(n_2978)
);

AND2x4_ASAP7_75t_L g2979 ( 
.A(n_2557),
.B(n_556),
.Y(n_2979)
);

AOI22xp33_ASAP7_75t_L g2980 ( 
.A1(n_2740),
.A2(n_557),
.B1(n_558),
.B2(n_559),
.Y(n_2980)
);

BUFx10_ASAP7_75t_L g2981 ( 
.A(n_2503),
.Y(n_2981)
);

INVx2_ASAP7_75t_L g2982 ( 
.A(n_2749),
.Y(n_2982)
);

OAI21xp5_ASAP7_75t_L g2983 ( 
.A1(n_2760),
.A2(n_558),
.B(n_560),
.Y(n_2983)
);

INVx1_ASAP7_75t_L g2984 ( 
.A(n_2616),
.Y(n_2984)
);

BUFx6f_ASAP7_75t_L g2985 ( 
.A(n_2452),
.Y(n_2985)
);

INVx2_ASAP7_75t_SL g2986 ( 
.A(n_2594),
.Y(n_2986)
);

INVx3_ASAP7_75t_L g2987 ( 
.A(n_2506),
.Y(n_2987)
);

INVx3_ASAP7_75t_L g2988 ( 
.A(n_2506),
.Y(n_2988)
);

BUFx3_ASAP7_75t_L g2989 ( 
.A(n_2592),
.Y(n_2989)
);

INVx1_ASAP7_75t_L g2990 ( 
.A(n_2709),
.Y(n_2990)
);

AO21x1_ASAP7_75t_L g2991 ( 
.A1(n_2567),
.A2(n_560),
.B(n_561),
.Y(n_2991)
);

INVx1_ASAP7_75t_L g2992 ( 
.A(n_2709),
.Y(n_2992)
);

INVx3_ASAP7_75t_SL g2993 ( 
.A(n_2653),
.Y(n_2993)
);

BUFx10_ASAP7_75t_L g2994 ( 
.A(n_2503),
.Y(n_2994)
);

INVx1_ASAP7_75t_L g2995 ( 
.A(n_2622),
.Y(n_2995)
);

INVx1_ASAP7_75t_L g2996 ( 
.A(n_2622),
.Y(n_2996)
);

BUFx2_ASAP7_75t_L g2997 ( 
.A(n_2465),
.Y(n_2997)
);

AO21x1_ASAP7_75t_SL g2998 ( 
.A1(n_2559),
.A2(n_561),
.B(n_562),
.Y(n_2998)
);

CKINVDCx6p67_ASAP7_75t_R g2999 ( 
.A(n_2556),
.Y(n_2999)
);

INVx1_ASAP7_75t_L g3000 ( 
.A(n_2522),
.Y(n_3000)
);

BUFx6f_ASAP7_75t_SL g3001 ( 
.A(n_2694),
.Y(n_3001)
);

INVx1_ASAP7_75t_L g3002 ( 
.A(n_2519),
.Y(n_3002)
);

BUFx2_ASAP7_75t_R g3003 ( 
.A(n_2542),
.Y(n_3003)
);

OA21x2_ASAP7_75t_L g3004 ( 
.A1(n_2477),
.A2(n_562),
.B(n_563),
.Y(n_3004)
);

HB1xp67_ASAP7_75t_L g3005 ( 
.A(n_2663),
.Y(n_3005)
);

OA21x2_ASAP7_75t_L g3006 ( 
.A1(n_2705),
.A2(n_563),
.B(n_564),
.Y(n_3006)
);

INVx1_ASAP7_75t_L g3007 ( 
.A(n_2519),
.Y(n_3007)
);

HB1xp67_ASAP7_75t_L g3008 ( 
.A(n_2663),
.Y(n_3008)
);

OAI21x1_ASAP7_75t_L g3009 ( 
.A1(n_2741),
.A2(n_564),
.B(n_565),
.Y(n_3009)
);

BUFx6f_ASAP7_75t_L g3010 ( 
.A(n_2452),
.Y(n_3010)
);

INVx3_ASAP7_75t_L g3011 ( 
.A(n_2456),
.Y(n_3011)
);

INVx1_ASAP7_75t_L g3012 ( 
.A(n_2563),
.Y(n_3012)
);

BUFx2_ASAP7_75t_L g3013 ( 
.A(n_2524),
.Y(n_3013)
);

INVx1_ASAP7_75t_L g3014 ( 
.A(n_2695),
.Y(n_3014)
);

AND2x4_ASAP7_75t_L g3015 ( 
.A(n_2557),
.B(n_2516),
.Y(n_3015)
);

NAND2x1p5_ASAP7_75t_L g3016 ( 
.A(n_2456),
.B(n_639),
.Y(n_3016)
);

BUFx2_ASAP7_75t_L g3017 ( 
.A(n_2533),
.Y(n_3017)
);

INVx1_ASAP7_75t_L g3018 ( 
.A(n_2695),
.Y(n_3018)
);

BUFx4f_ASAP7_75t_SL g3019 ( 
.A(n_2698),
.Y(n_3019)
);

INVx1_ASAP7_75t_L g3020 ( 
.A(n_2656),
.Y(n_3020)
);

AOI22xp33_ASAP7_75t_L g3021 ( 
.A1(n_2740),
.A2(n_565),
.B1(n_566),
.B2(n_567),
.Y(n_3021)
);

BUFx6f_ASAP7_75t_L g3022 ( 
.A(n_2456),
.Y(n_3022)
);

AO21x2_ASAP7_75t_L g3023 ( 
.A1(n_2536),
.A2(n_638),
.B(n_567),
.Y(n_3023)
);

BUFx6f_ASAP7_75t_L g3024 ( 
.A(n_2458),
.Y(n_3024)
);

AOI22xp33_ASAP7_75t_L g3025 ( 
.A1(n_2766),
.A2(n_566),
.B1(n_569),
.B2(n_571),
.Y(n_3025)
);

OAI21xp5_ASAP7_75t_L g3026 ( 
.A1(n_2760),
.A2(n_569),
.B(n_571),
.Y(n_3026)
);

INVx1_ASAP7_75t_L g3027 ( 
.A(n_2563),
.Y(n_3027)
);

INVx1_ASAP7_75t_L g3028 ( 
.A(n_2719),
.Y(n_3028)
);

INVx1_ASAP7_75t_L g3029 ( 
.A(n_2719),
.Y(n_3029)
);

INVxp67_ASAP7_75t_L g3030 ( 
.A(n_2539),
.Y(n_3030)
);

INVxp67_ASAP7_75t_SL g3031 ( 
.A(n_2537),
.Y(n_3031)
);

INVx2_ASAP7_75t_L g3032 ( 
.A(n_2445),
.Y(n_3032)
);

CKINVDCx11_ASAP7_75t_R g3033 ( 
.A(n_2541),
.Y(n_3033)
);

INVx1_ASAP7_75t_L g3034 ( 
.A(n_2722),
.Y(n_3034)
);

INVx1_ASAP7_75t_L g3035 ( 
.A(n_2722),
.Y(n_3035)
);

BUFx3_ASAP7_75t_L g3036 ( 
.A(n_2580),
.Y(n_3036)
);

AO21x1_ASAP7_75t_L g3037 ( 
.A1(n_2576),
.A2(n_572),
.B(n_573),
.Y(n_3037)
);

BUFx4_ASAP7_75t_R g3038 ( 
.A(n_2651),
.Y(n_3038)
);

INVx1_ASAP7_75t_L g3039 ( 
.A(n_2493),
.Y(n_3039)
);

INVx2_ASAP7_75t_L g3040 ( 
.A(n_2747),
.Y(n_3040)
);

INVx1_ASAP7_75t_L g3041 ( 
.A(n_2493),
.Y(n_3041)
);

AO21x1_ASAP7_75t_L g3042 ( 
.A1(n_2608),
.A2(n_572),
.B(n_573),
.Y(n_3042)
);

AOI22xp33_ASAP7_75t_SL g3043 ( 
.A1(n_2778),
.A2(n_574),
.B1(n_575),
.B2(n_576),
.Y(n_3043)
);

INVx1_ASAP7_75t_L g3044 ( 
.A(n_2504),
.Y(n_3044)
);

INVxp67_ASAP7_75t_SL g3045 ( 
.A(n_2537),
.Y(n_3045)
);

INVx2_ASAP7_75t_L g3046 ( 
.A(n_2747),
.Y(n_3046)
);

INVx1_ASAP7_75t_L g3047 ( 
.A(n_2732),
.Y(n_3047)
);

HB1xp67_ASAP7_75t_L g3048 ( 
.A(n_2738),
.Y(n_3048)
);

INVx3_ASAP7_75t_L g3049 ( 
.A(n_2458),
.Y(n_3049)
);

BUFx3_ASAP7_75t_L g3050 ( 
.A(n_2488),
.Y(n_3050)
);

INVx1_ASAP7_75t_L g3051 ( 
.A(n_2543),
.Y(n_3051)
);

INVx2_ASAP7_75t_L g3052 ( 
.A(n_2750),
.Y(n_3052)
);

BUFx2_ASAP7_75t_L g3053 ( 
.A(n_2458),
.Y(n_3053)
);

INVx1_ASAP7_75t_L g3054 ( 
.A(n_2543),
.Y(n_3054)
);

INVx1_ASAP7_75t_L g3055 ( 
.A(n_2551),
.Y(n_3055)
);

BUFx2_ASAP7_75t_L g3056 ( 
.A(n_2442),
.Y(n_3056)
);

BUFx6f_ASAP7_75t_L g3057 ( 
.A(n_2703),
.Y(n_3057)
);

OR2x2_ASAP7_75t_L g3058 ( 
.A(n_2615),
.B(n_574),
.Y(n_3058)
);

AOI21x1_ASAP7_75t_L g3059 ( 
.A1(n_2734),
.A2(n_576),
.B(n_578),
.Y(n_3059)
);

CKINVDCx11_ASAP7_75t_R g3060 ( 
.A(n_2545),
.Y(n_3060)
);

HB1xp67_ASAP7_75t_L g3061 ( 
.A(n_2615),
.Y(n_3061)
);

INVx2_ASAP7_75t_SL g3062 ( 
.A(n_2659),
.Y(n_3062)
);

INVx2_ASAP7_75t_L g3063 ( 
.A(n_2750),
.Y(n_3063)
);

INVx3_ASAP7_75t_L g3064 ( 
.A(n_2703),
.Y(n_3064)
);

INVx1_ASAP7_75t_L g3065 ( 
.A(n_2551),
.Y(n_3065)
);

CKINVDCx20_ASAP7_75t_R g3066 ( 
.A(n_2666),
.Y(n_3066)
);

INVx3_ASAP7_75t_L g3067 ( 
.A(n_2703),
.Y(n_3067)
);

INVx3_ASAP7_75t_L g3068 ( 
.A(n_2571),
.Y(n_3068)
);

INVx1_ASAP7_75t_L g3069 ( 
.A(n_2586),
.Y(n_3069)
);

AND2x2_ASAP7_75t_L g3070 ( 
.A(n_2680),
.B(n_579),
.Y(n_3070)
);

INVx1_ASAP7_75t_L g3071 ( 
.A(n_2586),
.Y(n_3071)
);

BUFx4_ASAP7_75t_R g3072 ( 
.A(n_2755),
.Y(n_3072)
);

AND2x2_ASAP7_75t_L g3073 ( 
.A(n_2633),
.B(n_579),
.Y(n_3073)
);

INVx1_ASAP7_75t_L g3074 ( 
.A(n_2600),
.Y(n_3074)
);

INVx1_ASAP7_75t_L g3075 ( 
.A(n_2600),
.Y(n_3075)
);

AOI22xp33_ASAP7_75t_L g3076 ( 
.A1(n_2798),
.A2(n_2790),
.B1(n_2731),
.B2(n_2774),
.Y(n_3076)
);

AOI22xp33_ASAP7_75t_L g3077 ( 
.A1(n_2790),
.A2(n_580),
.B1(n_581),
.B2(n_582),
.Y(n_3077)
);

AND2x2_ASAP7_75t_L g3078 ( 
.A(n_2555),
.B(n_580),
.Y(n_3078)
);

INVx1_ASAP7_75t_L g3079 ( 
.A(n_2504),
.Y(n_3079)
);

AO21x1_ASAP7_75t_L g3080 ( 
.A1(n_2608),
.A2(n_581),
.B(n_583),
.Y(n_3080)
);

BUFx10_ASAP7_75t_L g3081 ( 
.A(n_2565),
.Y(n_3081)
);

AND2x2_ASAP7_75t_L g3082 ( 
.A(n_2693),
.B(n_583),
.Y(n_3082)
);

INVx1_ASAP7_75t_L g3083 ( 
.A(n_2771),
.Y(n_3083)
);

INVx1_ASAP7_75t_L g3084 ( 
.A(n_2771),
.Y(n_3084)
);

AND2x2_ASAP7_75t_L g3085 ( 
.A(n_2710),
.B(n_584),
.Y(n_3085)
);

INVx3_ASAP7_75t_L g3086 ( 
.A(n_2571),
.Y(n_3086)
);

AOI22xp33_ASAP7_75t_L g3087 ( 
.A1(n_2731),
.A2(n_584),
.B1(n_585),
.B2(n_586),
.Y(n_3087)
);

INVx1_ASAP7_75t_L g3088 ( 
.A(n_2716),
.Y(n_3088)
);

BUFx3_ASAP7_75t_L g3089 ( 
.A(n_2499),
.Y(n_3089)
);

INVx3_ASAP7_75t_L g3090 ( 
.A(n_2607),
.Y(n_3090)
);

AND2x2_ASAP7_75t_L g3091 ( 
.A(n_2549),
.B(n_2565),
.Y(n_3091)
);

AND2x2_ASAP7_75t_L g3092 ( 
.A(n_2589),
.B(n_586),
.Y(n_3092)
);

INVx1_ASAP7_75t_L g3093 ( 
.A(n_2662),
.Y(n_3093)
);

INVx1_ASAP7_75t_L g3094 ( 
.A(n_2662),
.Y(n_3094)
);

INVx3_ASAP7_75t_L g3095 ( 
.A(n_2607),
.Y(n_3095)
);

HB1xp67_ASAP7_75t_L g3096 ( 
.A(n_2759),
.Y(n_3096)
);

INVx1_ASAP7_75t_L g3097 ( 
.A(n_2712),
.Y(n_3097)
);

OA21x2_ASAP7_75t_L g3098 ( 
.A1(n_2655),
.A2(n_587),
.B(n_588),
.Y(n_3098)
);

INVx1_ASAP7_75t_L g3099 ( 
.A(n_2789),
.Y(n_3099)
);

BUFx2_ASAP7_75t_L g3100 ( 
.A(n_2650),
.Y(n_3100)
);

CKINVDCx20_ASAP7_75t_R g3101 ( 
.A(n_2581),
.Y(n_3101)
);

AOI22xp5_ASAP7_75t_L g3102 ( 
.A1(n_2534),
.A2(n_2599),
.B1(n_2769),
.B2(n_2785),
.Y(n_3102)
);

INVx1_ASAP7_75t_L g3103 ( 
.A(n_2789),
.Y(n_3103)
);

CKINVDCx5p33_ASAP7_75t_R g3104 ( 
.A(n_2675),
.Y(n_3104)
);

OAI22xp5_ASAP7_75t_L g3105 ( 
.A1(n_2613),
.A2(n_587),
.B1(n_588),
.B2(n_589),
.Y(n_3105)
);

INVx2_ASAP7_75t_L g3106 ( 
.A(n_2511),
.Y(n_3106)
);

AOI22xp33_ASAP7_75t_SL g3107 ( 
.A1(n_2730),
.A2(n_589),
.B1(n_590),
.B2(n_591),
.Y(n_3107)
);

BUFx3_ASAP7_75t_L g3108 ( 
.A(n_2676),
.Y(n_3108)
);

CKINVDCx11_ASAP7_75t_R g3109 ( 
.A(n_2755),
.Y(n_3109)
);

AOI22xp33_ASAP7_75t_SL g3110 ( 
.A1(n_2701),
.A2(n_590),
.B1(n_592),
.B2(n_593),
.Y(n_3110)
);

AOI22xp33_ASAP7_75t_L g3111 ( 
.A1(n_2752),
.A2(n_592),
.B1(n_594),
.B2(n_595),
.Y(n_3111)
);

INVx2_ASAP7_75t_L g3112 ( 
.A(n_2520),
.Y(n_3112)
);

BUFx2_ASAP7_75t_L g3113 ( 
.A(n_2593),
.Y(n_3113)
);

INVx2_ASAP7_75t_SL g3114 ( 
.A(n_2659),
.Y(n_3114)
);

OAI21x1_ASAP7_75t_SL g3115 ( 
.A1(n_2661),
.A2(n_2673),
.B(n_2630),
.Y(n_3115)
);

INVx1_ASAP7_75t_L g3116 ( 
.A(n_2677),
.Y(n_3116)
);

NAND2xp5_ASAP7_75t_SL g3117 ( 
.A(n_2607),
.B(n_594),
.Y(n_3117)
);

INVx1_ASAP7_75t_L g3118 ( 
.A(n_2677),
.Y(n_3118)
);

CKINVDCx20_ASAP7_75t_R g3119 ( 
.A(n_2584),
.Y(n_3119)
);

BUFx2_ASAP7_75t_L g3120 ( 
.A(n_2606),
.Y(n_3120)
);

NAND2xp5_ASAP7_75t_SL g3121 ( 
.A(n_2924),
.B(n_2589),
.Y(n_3121)
);

INVx1_ASAP7_75t_L g3122 ( 
.A(n_2803),
.Y(n_3122)
);

INVx1_ASAP7_75t_L g3123 ( 
.A(n_2803),
.Y(n_3123)
);

CKINVDCx5p33_ASAP7_75t_R g3124 ( 
.A(n_2880),
.Y(n_3124)
);

AND2x4_ASAP7_75t_SL g3125 ( 
.A(n_2875),
.B(n_2516),
.Y(n_3125)
);

NOR2xp33_ASAP7_75t_L g3126 ( 
.A(n_2869),
.B(n_2582),
.Y(n_3126)
);

INVx1_ASAP7_75t_L g3127 ( 
.A(n_2804),
.Y(n_3127)
);

INVx1_ASAP7_75t_L g3128 ( 
.A(n_2804),
.Y(n_3128)
);

AND2x2_ASAP7_75t_L g3129 ( 
.A(n_2816),
.B(n_2669),
.Y(n_3129)
);

INVx1_ASAP7_75t_L g3130 ( 
.A(n_2805),
.Y(n_3130)
);

BUFx2_ASAP7_75t_L g3131 ( 
.A(n_2822),
.Y(n_3131)
);

NAND3xp33_ASAP7_75t_SL g3132 ( 
.A(n_2873),
.B(n_2745),
.C(n_2613),
.Y(n_3132)
);

INVx2_ASAP7_75t_L g3133 ( 
.A(n_2802),
.Y(n_3133)
);

NAND2xp5_ASAP7_75t_L g3134 ( 
.A(n_2840),
.B(n_2769),
.Y(n_3134)
);

NOR2xp33_ASAP7_75t_R g3135 ( 
.A(n_2868),
.B(n_2728),
.Y(n_3135)
);

BUFx3_ASAP7_75t_L g3136 ( 
.A(n_2864),
.Y(n_3136)
);

OAI22xp5_ASAP7_75t_L g3137 ( 
.A1(n_2867),
.A2(n_2657),
.B1(n_2509),
.B2(n_2765),
.Y(n_3137)
);

INVx1_ASAP7_75t_L g3138 ( 
.A(n_2808),
.Y(n_3138)
);

HB1xp67_ASAP7_75t_L g3139 ( 
.A(n_3061),
.Y(n_3139)
);

OR2x2_ASAP7_75t_L g3140 ( 
.A(n_2823),
.B(n_2547),
.Y(n_3140)
);

INVx1_ASAP7_75t_L g3141 ( 
.A(n_2808),
.Y(n_3141)
);

AND2x4_ASAP7_75t_SL g3142 ( 
.A(n_2875),
.B(n_2538),
.Y(n_3142)
);

AND2x2_ASAP7_75t_L g3143 ( 
.A(n_3078),
.B(n_2547),
.Y(n_3143)
);

INVx3_ASAP7_75t_L g3144 ( 
.A(n_2822),
.Y(n_3144)
);

INVx1_ASAP7_75t_L g3145 ( 
.A(n_2809),
.Y(n_3145)
);

AND2x2_ASAP7_75t_SL g3146 ( 
.A(n_2907),
.B(n_2784),
.Y(n_3146)
);

AND2x2_ASAP7_75t_L g3147 ( 
.A(n_3070),
.B(n_2590),
.Y(n_3147)
);

OR2x2_ASAP7_75t_L g3148 ( 
.A(n_2838),
.B(n_2590),
.Y(n_3148)
);

INVx1_ASAP7_75t_L g3149 ( 
.A(n_2809),
.Y(n_3149)
);

NAND2xp33_ASAP7_75t_R g3150 ( 
.A(n_2956),
.B(n_2784),
.Y(n_3150)
);

CKINVDCx16_ASAP7_75t_R g3151 ( 
.A(n_2817),
.Y(n_3151)
);

OR2x6_ASAP7_75t_L g3152 ( 
.A(n_2872),
.B(n_2572),
.Y(n_3152)
);

AND2x2_ASAP7_75t_L g3153 ( 
.A(n_3073),
.B(n_2665),
.Y(n_3153)
);

NAND2xp33_ASAP7_75t_R g3154 ( 
.A(n_2997),
.B(n_2614),
.Y(n_3154)
);

CKINVDCx5p33_ASAP7_75t_R g3155 ( 
.A(n_2944),
.Y(n_3155)
);

OR2x6_ASAP7_75t_L g3156 ( 
.A(n_2907),
.B(n_2583),
.Y(n_3156)
);

INVx2_ASAP7_75t_L g3157 ( 
.A(n_2807),
.Y(n_3157)
);

INVx2_ASAP7_75t_L g3158 ( 
.A(n_2832),
.Y(n_3158)
);

CKINVDCx20_ASAP7_75t_R g3159 ( 
.A(n_2910),
.Y(n_3159)
);

INVx1_ASAP7_75t_L g3160 ( 
.A(n_2810),
.Y(n_3160)
);

NOR2xp33_ASAP7_75t_R g3161 ( 
.A(n_2858),
.B(n_2752),
.Y(n_3161)
);

HB1xp67_ASAP7_75t_L g3162 ( 
.A(n_3005),
.Y(n_3162)
);

OR2x6_ASAP7_75t_L g3163 ( 
.A(n_3062),
.B(n_2509),
.Y(n_3163)
);

INVx2_ASAP7_75t_L g3164 ( 
.A(n_2844),
.Y(n_3164)
);

INVx1_ASAP7_75t_L g3165 ( 
.A(n_2811),
.Y(n_3165)
);

NOR2xp33_ASAP7_75t_R g3166 ( 
.A(n_2865),
.B(n_2640),
.Y(n_3166)
);

BUFx10_ASAP7_75t_L g3167 ( 
.A(n_2950),
.Y(n_3167)
);

AND2x2_ASAP7_75t_SL g3168 ( 
.A(n_2916),
.B(n_2605),
.Y(n_3168)
);

NOR2x1_ASAP7_75t_SL g3169 ( 
.A(n_2815),
.B(n_2702),
.Y(n_3169)
);

NOR3xp33_ASAP7_75t_SL g3170 ( 
.A(n_3104),
.B(n_2598),
.C(n_2793),
.Y(n_3170)
);

INVx3_ASAP7_75t_L g3171 ( 
.A(n_2935),
.Y(n_3171)
);

NAND2xp5_ASAP7_75t_L g3172 ( 
.A(n_2812),
.B(n_2780),
.Y(n_3172)
);

INVx1_ASAP7_75t_L g3173 ( 
.A(n_2812),
.Y(n_3173)
);

INVxp67_ASAP7_75t_L g3174 ( 
.A(n_3013),
.Y(n_3174)
);

AND2x4_ASAP7_75t_L g3175 ( 
.A(n_2843),
.B(n_2642),
.Y(n_3175)
);

HB1xp67_ASAP7_75t_L g3176 ( 
.A(n_3008),
.Y(n_3176)
);

AOI22xp33_ASAP7_75t_L g3177 ( 
.A1(n_2806),
.A2(n_2686),
.B1(n_2513),
.B2(n_2796),
.Y(n_3177)
);

INVx3_ASAP7_75t_L g3178 ( 
.A(n_2935),
.Y(n_3178)
);

INVx2_ASAP7_75t_L g3179 ( 
.A(n_2847),
.Y(n_3179)
);

AND2x2_ASAP7_75t_L g3180 ( 
.A(n_3082),
.B(n_2621),
.Y(n_3180)
);

NAND2xp5_ASAP7_75t_L g3181 ( 
.A(n_2818),
.B(n_2540),
.Y(n_3181)
);

INVx2_ASAP7_75t_L g3182 ( 
.A(n_2848),
.Y(n_3182)
);

INVx2_ASAP7_75t_L g3183 ( 
.A(n_2851),
.Y(n_3183)
);

INVx1_ASAP7_75t_L g3184 ( 
.A(n_2818),
.Y(n_3184)
);

INVx2_ASAP7_75t_L g3185 ( 
.A(n_2853),
.Y(n_3185)
);

INVx1_ASAP7_75t_L g3186 ( 
.A(n_2821),
.Y(n_3186)
);

CKINVDCx16_ASAP7_75t_R g3187 ( 
.A(n_2835),
.Y(n_3187)
);

AOI22xp33_ASAP7_75t_L g3188 ( 
.A1(n_2862),
.A2(n_2686),
.B1(n_2796),
.B2(n_2787),
.Y(n_3188)
);

NOR3xp33_ASAP7_75t_SL g3189 ( 
.A(n_2879),
.B(n_2793),
.C(n_2748),
.Y(n_3189)
);

OAI222xp33_ASAP7_75t_L g3190 ( 
.A1(n_2900),
.A2(n_2712),
.B1(n_2800),
.B2(n_2795),
.C1(n_2605),
.C2(n_2435),
.Y(n_3190)
);

BUFx3_ASAP7_75t_L g3191 ( 
.A(n_2874),
.Y(n_3191)
);

NAND2xp5_ASAP7_75t_L g3192 ( 
.A(n_2821),
.B(n_2540),
.Y(n_3192)
);

INVx3_ASAP7_75t_L g3193 ( 
.A(n_2843),
.Y(n_3193)
);

AOI22xp5_ASAP7_75t_L g3194 ( 
.A1(n_2820),
.A2(n_2657),
.B1(n_2787),
.B2(n_2573),
.Y(n_3194)
);

HB1xp67_ASAP7_75t_L g3195 ( 
.A(n_3048),
.Y(n_3195)
);

OR2x2_ASAP7_75t_L g3196 ( 
.A(n_2949),
.B(n_2638),
.Y(n_3196)
);

XNOR2xp5_ASAP7_75t_L g3197 ( 
.A(n_2846),
.B(n_2512),
.Y(n_3197)
);

INVx1_ASAP7_75t_L g3198 ( 
.A(n_2825),
.Y(n_3198)
);

AND2x4_ASAP7_75t_L g3199 ( 
.A(n_2845),
.B(n_2642),
.Y(n_3199)
);

AND2x4_ASAP7_75t_L g3200 ( 
.A(n_2845),
.B(n_2642),
.Y(n_3200)
);

AND2x2_ASAP7_75t_L g3201 ( 
.A(n_3085),
.B(n_2628),
.Y(n_3201)
);

NOR2xp33_ASAP7_75t_R g3202 ( 
.A(n_2922),
.B(n_2440),
.Y(n_3202)
);

AND2x2_ASAP7_75t_L g3203 ( 
.A(n_3092),
.B(n_2629),
.Y(n_3203)
);

AO31x2_ASAP7_75t_L g3204 ( 
.A1(n_3106),
.A2(n_2439),
.A3(n_2777),
.B(n_2595),
.Y(n_3204)
);

NOR2xp33_ASAP7_75t_R g3205 ( 
.A(n_3119),
.B(n_2440),
.Y(n_3205)
);

HB1xp67_ASAP7_75t_L g3206 ( 
.A(n_2863),
.Y(n_3206)
);

BUFx6f_ASAP7_75t_L g3207 ( 
.A(n_3057),
.Y(n_3207)
);

INVx2_ASAP7_75t_L g3208 ( 
.A(n_2856),
.Y(n_3208)
);

AND2x2_ASAP7_75t_L g3209 ( 
.A(n_2964),
.B(n_2634),
.Y(n_3209)
);

AND2x2_ASAP7_75t_L g3210 ( 
.A(n_3096),
.B(n_2639),
.Y(n_3210)
);

HB1xp67_ASAP7_75t_L g3211 ( 
.A(n_2928),
.Y(n_3211)
);

CKINVDCx5p33_ASAP7_75t_R g3212 ( 
.A(n_2903),
.Y(n_3212)
);

AOI22xp33_ASAP7_75t_L g3213 ( 
.A1(n_2870),
.A2(n_2729),
.B1(n_2723),
.B2(n_2574),
.Y(n_3213)
);

NOR3xp33_ASAP7_75t_SL g3214 ( 
.A(n_2882),
.B(n_2748),
.C(n_2721),
.Y(n_3214)
);

NOR3xp33_ASAP7_75t_SL g3215 ( 
.A(n_2913),
.B(n_2721),
.C(n_2775),
.Y(n_3215)
);

BUFx6f_ASAP7_75t_L g3216 ( 
.A(n_3057),
.Y(n_3216)
);

OAI22xp5_ASAP7_75t_L g3217 ( 
.A1(n_2841),
.A2(n_2765),
.B1(n_2800),
.B2(n_2795),
.Y(n_3217)
);

OR2x6_ASAP7_75t_L g3218 ( 
.A(n_3114),
.B(n_2794),
.Y(n_3218)
);

AND2x4_ASAP7_75t_L g3219 ( 
.A(n_3116),
.B(n_2702),
.Y(n_3219)
);

AND2x4_ASAP7_75t_L g3220 ( 
.A(n_3116),
.B(n_2702),
.Y(n_3220)
);

NAND2xp33_ASAP7_75t_L g3221 ( 
.A(n_3057),
.B(n_2677),
.Y(n_3221)
);

AND2x2_ASAP7_75t_L g3222 ( 
.A(n_3091),
.B(n_2652),
.Y(n_3222)
);

NAND2xp33_ASAP7_75t_SL g3223 ( 
.A(n_2993),
.B(n_2623),
.Y(n_3223)
);

NOR2xp33_ASAP7_75t_R g3224 ( 
.A(n_2909),
.B(n_2538),
.Y(n_3224)
);

CKINVDCx11_ASAP7_75t_R g3225 ( 
.A(n_3060),
.Y(n_3225)
);

NOR2x1_ASAP7_75t_SL g3226 ( 
.A(n_2819),
.B(n_2704),
.Y(n_3226)
);

BUFx3_ASAP7_75t_L g3227 ( 
.A(n_2888),
.Y(n_3227)
);

NAND3xp33_ASAP7_75t_SL g3228 ( 
.A(n_2852),
.B(n_2630),
.C(n_2699),
.Y(n_3228)
);

NAND2xp33_ASAP7_75t_R g3229 ( 
.A(n_2979),
.B(n_2632),
.Y(n_3229)
);

CKINVDCx5p33_ASAP7_75t_R g3230 ( 
.A(n_2909),
.Y(n_3230)
);

AND2x2_ASAP7_75t_L g3231 ( 
.A(n_3000),
.B(n_2660),
.Y(n_3231)
);

AOI222xp33_ASAP7_75t_L g3232 ( 
.A1(n_2962),
.A2(n_2966),
.B1(n_2836),
.B2(n_3105),
.C1(n_2849),
.C2(n_2893),
.Y(n_3232)
);

AND2x2_ASAP7_75t_L g3233 ( 
.A(n_2960),
.B(n_2635),
.Y(n_3233)
);

OR2x2_ASAP7_75t_L g3234 ( 
.A(n_2941),
.B(n_2638),
.Y(n_3234)
);

HB1xp67_ASAP7_75t_L g3235 ( 
.A(n_3031),
.Y(n_3235)
);

HB1xp67_ASAP7_75t_L g3236 ( 
.A(n_3045),
.Y(n_3236)
);

AND2x2_ASAP7_75t_L g3237 ( 
.A(n_3053),
.B(n_2683),
.Y(n_3237)
);

INVx3_ASAP7_75t_L g3238 ( 
.A(n_2861),
.Y(n_3238)
);

AND2x2_ASAP7_75t_L g3239 ( 
.A(n_3017),
.B(n_2587),
.Y(n_3239)
);

CKINVDCx5p33_ASAP7_75t_R g3240 ( 
.A(n_3033),
.Y(n_3240)
);

NAND2xp33_ASAP7_75t_SL g3241 ( 
.A(n_2950),
.B(n_2788),
.Y(n_3241)
);

AND2x2_ASAP7_75t_L g3242 ( 
.A(n_2973),
.B(n_2587),
.Y(n_3242)
);

NAND2xp5_ASAP7_75t_L g3243 ( 
.A(n_2827),
.B(n_2575),
.Y(n_3243)
);

INVx3_ASAP7_75t_L g3244 ( 
.A(n_2861),
.Y(n_3244)
);

INVx2_ASAP7_75t_L g3245 ( 
.A(n_2859),
.Y(n_3245)
);

NAND3xp33_ASAP7_75t_SL g3246 ( 
.A(n_3101),
.B(n_2714),
.C(n_2699),
.Y(n_3246)
);

NAND3xp33_ASAP7_75t_SL g3247 ( 
.A(n_2921),
.B(n_2714),
.C(n_2775),
.Y(n_3247)
);

BUFx2_ASAP7_75t_L g3248 ( 
.A(n_3113),
.Y(n_3248)
);

NAND2xp5_ASAP7_75t_L g3249 ( 
.A(n_2828),
.B(n_2577),
.Y(n_3249)
);

HB1xp67_ASAP7_75t_L g3250 ( 
.A(n_3038),
.Y(n_3250)
);

AND2x2_ASAP7_75t_L g3251 ( 
.A(n_2813),
.B(n_2596),
.Y(n_3251)
);

AND2x2_ASAP7_75t_L g3252 ( 
.A(n_2814),
.B(n_2596),
.Y(n_3252)
);

NAND2xp5_ASAP7_75t_L g3253 ( 
.A(n_2829),
.B(n_2620),
.Y(n_3253)
);

HB1xp67_ASAP7_75t_L g3254 ( 
.A(n_3056),
.Y(n_3254)
);

INVx1_ASAP7_75t_SL g3255 ( 
.A(n_2839),
.Y(n_3255)
);

OR2x2_ASAP7_75t_L g3256 ( 
.A(n_2824),
.B(n_2830),
.Y(n_3256)
);

NOR2xp33_ASAP7_75t_R g3257 ( 
.A(n_2978),
.B(n_3066),
.Y(n_3257)
);

AND2x2_ASAP7_75t_L g3258 ( 
.A(n_3047),
.B(n_2619),
.Y(n_3258)
);

INVx1_ASAP7_75t_L g3259 ( 
.A(n_2829),
.Y(n_3259)
);

INVx5_ASAP7_75t_SL g3260 ( 
.A(n_2961),
.Y(n_3260)
);

AND2x4_ASAP7_75t_L g3261 ( 
.A(n_3118),
.B(n_2704),
.Y(n_3261)
);

NOR3xp33_ASAP7_75t_L g3262 ( 
.A(n_2834),
.B(n_2655),
.C(n_2625),
.Y(n_3262)
);

OR2x2_ASAP7_75t_L g3263 ( 
.A(n_3058),
.B(n_2920),
.Y(n_3263)
);

AND2x4_ASAP7_75t_L g3264 ( 
.A(n_3118),
.B(n_2704),
.Y(n_3264)
);

INVx1_ASAP7_75t_L g3265 ( 
.A(n_2930),
.Y(n_3265)
);

NAND2x1_ASAP7_75t_L g3266 ( 
.A(n_3002),
.B(n_2667),
.Y(n_3266)
);

INVx1_ASAP7_75t_SL g3267 ( 
.A(n_2839),
.Y(n_3267)
);

AOI22xp33_ASAP7_75t_L g3268 ( 
.A1(n_2894),
.A2(n_2664),
.B1(n_2624),
.B2(n_2636),
.Y(n_3268)
);

INVx4_ASAP7_75t_L g3269 ( 
.A(n_3072),
.Y(n_3269)
);

AND2x2_ASAP7_75t_L g3270 ( 
.A(n_2908),
.B(n_2619),
.Y(n_3270)
);

OR2x2_ASAP7_75t_L g3271 ( 
.A(n_3030),
.B(n_2641),
.Y(n_3271)
);

AOI22xp33_ASAP7_75t_L g3272 ( 
.A1(n_2911),
.A2(n_2647),
.B1(n_2658),
.B2(n_2674),
.Y(n_3272)
);

AOI22xp5_ASAP7_75t_L g3273 ( 
.A1(n_2837),
.A2(n_2692),
.B1(n_2643),
.B2(n_2646),
.Y(n_3273)
);

OAI21xp33_ASAP7_75t_L g3274 ( 
.A1(n_2850),
.A2(n_2512),
.B(n_2700),
.Y(n_3274)
);

AND2x2_ASAP7_75t_L g3275 ( 
.A(n_2959),
.B(n_2641),
.Y(n_3275)
);

OR2x2_ASAP7_75t_L g3276 ( 
.A(n_2897),
.B(n_2679),
.Y(n_3276)
);

INVx3_ASAP7_75t_L g3277 ( 
.A(n_2861),
.Y(n_3277)
);

NAND3xp33_ASAP7_75t_SL g3278 ( 
.A(n_3037),
.B(n_2595),
.C(n_2535),
.Y(n_3278)
);

CKINVDCx5p33_ASAP7_75t_R g3279 ( 
.A(n_2999),
.Y(n_3279)
);

HB1xp67_ASAP7_75t_L g3280 ( 
.A(n_2904),
.Y(n_3280)
);

BUFx10_ASAP7_75t_L g3281 ( 
.A(n_2986),
.Y(n_3281)
);

AND2x2_ASAP7_75t_L g3282 ( 
.A(n_2979),
.B(n_596),
.Y(n_3282)
);

HB1xp67_ASAP7_75t_L g3283 ( 
.A(n_2905),
.Y(n_3283)
);

INVx1_ASAP7_75t_L g3284 ( 
.A(n_2906),
.Y(n_3284)
);

INVx1_ASAP7_75t_L g3285 ( 
.A(n_2917),
.Y(n_3285)
);

INVx1_ASAP7_75t_L g3286 ( 
.A(n_2923),
.Y(n_3286)
);

AOI22xp33_ASAP7_75t_L g3287 ( 
.A1(n_2911),
.A2(n_2860),
.B1(n_2831),
.B2(n_2842),
.Y(n_3287)
);

INVx1_ASAP7_75t_L g3288 ( 
.A(n_2952),
.Y(n_3288)
);

BUFx2_ASAP7_75t_L g3289 ( 
.A(n_2985),
.Y(n_3289)
);

INVx1_ASAP7_75t_L g3290 ( 
.A(n_2995),
.Y(n_3290)
);

NAND2xp5_ASAP7_75t_L g3291 ( 
.A(n_2939),
.B(n_2685),
.Y(n_3291)
);

CKINVDCx5p33_ASAP7_75t_R g3292 ( 
.A(n_3019),
.Y(n_3292)
);

CKINVDCx16_ASAP7_75t_R g3293 ( 
.A(n_2957),
.Y(n_3293)
);

INVx3_ASAP7_75t_L g3294 ( 
.A(n_2985),
.Y(n_3294)
);

OR2x2_ASAP7_75t_L g3295 ( 
.A(n_3108),
.B(n_2688),
.Y(n_3295)
);

INVx1_ASAP7_75t_L g3296 ( 
.A(n_2996),
.Y(n_3296)
);

OAI21xp5_ASAP7_75t_L g3297 ( 
.A1(n_2877),
.A2(n_2783),
.B(n_2535),
.Y(n_3297)
);

AND2x2_ASAP7_75t_L g3298 ( 
.A(n_2998),
.B(n_3011),
.Y(n_3298)
);

AND2x2_ASAP7_75t_L g3299 ( 
.A(n_3011),
.B(n_597),
.Y(n_3299)
);

BUFx3_ASAP7_75t_L g3300 ( 
.A(n_3036),
.Y(n_3300)
);

INVx1_ASAP7_75t_L g3301 ( 
.A(n_3051),
.Y(n_3301)
);

HB1xp67_ASAP7_75t_L g3302 ( 
.A(n_3015),
.Y(n_3302)
);

INVx1_ASAP7_75t_L g3303 ( 
.A(n_3054),
.Y(n_3303)
);

AOI22xp33_ASAP7_75t_L g3304 ( 
.A1(n_2887),
.A2(n_2717),
.B1(n_2733),
.B2(n_2753),
.Y(n_3304)
);

O2A1O1Ixp33_ASAP7_75t_L g3305 ( 
.A1(n_2918),
.A2(n_2744),
.B(n_2742),
.C(n_2720),
.Y(n_3305)
);

BUFx3_ASAP7_75t_L g3306 ( 
.A(n_2989),
.Y(n_3306)
);

XOR2xp5_ASAP7_75t_L g3307 ( 
.A(n_2932),
.B(n_2588),
.Y(n_3307)
);

NAND2xp33_ASAP7_75t_R g3308 ( 
.A(n_3090),
.B(n_2781),
.Y(n_3308)
);

OAI21xp5_ASAP7_75t_SL g3309 ( 
.A1(n_3076),
.A2(n_2797),
.B(n_2788),
.Y(n_3309)
);

BUFx3_ASAP7_75t_L g3310 ( 
.A(n_2981),
.Y(n_3310)
);

AND2x2_ASAP7_75t_L g3311 ( 
.A(n_3049),
.B(n_598),
.Y(n_3311)
);

BUFx12f_ASAP7_75t_L g3312 ( 
.A(n_3109),
.Y(n_3312)
);

INVx1_ASAP7_75t_L g3313 ( 
.A(n_3055),
.Y(n_3313)
);

BUFx2_ASAP7_75t_L g3314 ( 
.A(n_2985),
.Y(n_3314)
);

AND2x2_ASAP7_75t_L g3315 ( 
.A(n_3049),
.B(n_599),
.Y(n_3315)
);

INVxp67_ASAP7_75t_L g3316 ( 
.A(n_2940),
.Y(n_3316)
);

OAI21xp5_ASAP7_75t_SL g3317 ( 
.A1(n_3087),
.A2(n_2788),
.B(n_2558),
.Y(n_3317)
);

INVx2_ASAP7_75t_L g3318 ( 
.A(n_3009),
.Y(n_3318)
);

OAI22xp33_ASAP7_75t_L g3319 ( 
.A1(n_3102),
.A2(n_2733),
.B1(n_2781),
.B2(n_2544),
.Y(n_3319)
);

CKINVDCx16_ASAP7_75t_R g3320 ( 
.A(n_2981),
.Y(n_3320)
);

CKINVDCx5p33_ASAP7_75t_R g3321 ( 
.A(n_3001),
.Y(n_3321)
);

INVx1_ASAP7_75t_L g3322 ( 
.A(n_3065),
.Y(n_3322)
);

AND2x2_ASAP7_75t_L g3323 ( 
.A(n_3015),
.B(n_599),
.Y(n_3323)
);

AND2x2_ASAP7_75t_L g3324 ( 
.A(n_3081),
.B(n_600),
.Y(n_3324)
);

CKINVDCx16_ASAP7_75t_R g3325 ( 
.A(n_2994),
.Y(n_3325)
);

NAND2xp5_ASAP7_75t_L g3326 ( 
.A(n_2854),
.B(n_2779),
.Y(n_3326)
);

AND2x2_ASAP7_75t_L g3327 ( 
.A(n_3081),
.B(n_601),
.Y(n_3327)
);

OA21x2_ASAP7_75t_L g3328 ( 
.A1(n_3083),
.A2(n_2801),
.B(n_2525),
.Y(n_3328)
);

AOI221xp5_ASAP7_75t_L g3329 ( 
.A1(n_2958),
.A2(n_2568),
.B1(n_2579),
.B2(n_2602),
.C(n_2552),
.Y(n_3329)
);

NAND4xp25_ASAP7_75t_L g3330 ( 
.A(n_2866),
.B(n_2588),
.C(n_2727),
.D(n_2558),
.Y(n_3330)
);

OR2x6_ASAP7_75t_L g3331 ( 
.A(n_2929),
.B(n_2792),
.Y(n_3331)
);

HB1xp67_ASAP7_75t_L g3332 ( 
.A(n_3007),
.Y(n_3332)
);

NAND2xp33_ASAP7_75t_R g3333 ( 
.A(n_3090),
.B(n_602),
.Y(n_3333)
);

XNOR2xp5_ASAP7_75t_L g3334 ( 
.A(n_3120),
.B(n_2675),
.Y(n_3334)
);

CKINVDCx5p33_ASAP7_75t_R g3335 ( 
.A(n_3001),
.Y(n_3335)
);

NAND2xp5_ASAP7_75t_L g3336 ( 
.A(n_2855),
.B(n_2857),
.Y(n_3336)
);

INVx1_ASAP7_75t_L g3337 ( 
.A(n_2975),
.Y(n_3337)
);

AND2x2_ASAP7_75t_L g3338 ( 
.A(n_3100),
.B(n_603),
.Y(n_3338)
);

NAND2xp33_ASAP7_75t_SL g3339 ( 
.A(n_3012),
.B(n_3027),
.Y(n_3339)
);

HB1xp67_ASAP7_75t_L g3340 ( 
.A(n_3069),
.Y(n_3340)
);

INVx1_ASAP7_75t_SL g3341 ( 
.A(n_2994),
.Y(n_3341)
);

CKINVDCx8_ASAP7_75t_R g3342 ( 
.A(n_3010),
.Y(n_3342)
);

NAND2xp33_ASAP7_75t_R g3343 ( 
.A(n_3095),
.B(n_603),
.Y(n_3343)
);

OAI22xp33_ASAP7_75t_SL g3344 ( 
.A1(n_3071),
.A2(n_2527),
.B1(n_2739),
.B2(n_2667),
.Y(n_3344)
);

INVx1_ASAP7_75t_L g3345 ( 
.A(n_3059),
.Y(n_3345)
);

AOI22xp33_ASAP7_75t_L g3346 ( 
.A1(n_2912),
.A2(n_2727),
.B1(n_2786),
.B2(n_2726),
.Y(n_3346)
);

HB1xp67_ASAP7_75t_L g3347 ( 
.A(n_3028),
.Y(n_3347)
);

INVx2_ASAP7_75t_L g3348 ( 
.A(n_3010),
.Y(n_3348)
);

AND2x4_ASAP7_75t_L g3349 ( 
.A(n_3029),
.B(n_3034),
.Y(n_3349)
);

AND2x2_ASAP7_75t_L g3350 ( 
.A(n_3010),
.B(n_604),
.Y(n_3350)
);

AOI22xp33_ASAP7_75t_L g3351 ( 
.A1(n_2963),
.A2(n_2786),
.B1(n_2726),
.B2(n_2529),
.Y(n_3351)
);

INVx3_ASAP7_75t_L g3352 ( 
.A(n_3022),
.Y(n_3352)
);

BUFx2_ASAP7_75t_L g3353 ( 
.A(n_3022),
.Y(n_3353)
);

OR2x2_ASAP7_75t_L g3354 ( 
.A(n_2982),
.B(n_2564),
.Y(n_3354)
);

BUFx6f_ASAP7_75t_L g3355 ( 
.A(n_3022),
.Y(n_3355)
);

CKINVDCx20_ASAP7_75t_R g3356 ( 
.A(n_3050),
.Y(n_3356)
);

NOR2xp33_ASAP7_75t_R g3357 ( 
.A(n_2946),
.B(n_2741),
.Y(n_3357)
);

OAI21xp33_ASAP7_75t_L g3358 ( 
.A1(n_2953),
.A2(n_2507),
.B(n_2578),
.Y(n_3358)
);

NAND3xp33_ASAP7_75t_L g3359 ( 
.A(n_3020),
.B(n_2711),
.C(n_2564),
.Y(n_3359)
);

BUFx3_ASAP7_75t_L g3360 ( 
.A(n_3089),
.Y(n_3360)
);

CKINVDCx5p33_ASAP7_75t_R g3361 ( 
.A(n_3003),
.Y(n_3361)
);

AND2x4_ASAP7_75t_L g3362 ( 
.A(n_3035),
.B(n_3095),
.Y(n_3362)
);

CKINVDCx16_ASAP7_75t_R g3363 ( 
.A(n_3024),
.Y(n_3363)
);

INVx2_ASAP7_75t_L g3364 ( 
.A(n_3024),
.Y(n_3364)
);

NAND3xp33_ASAP7_75t_SL g3365 ( 
.A(n_2991),
.B(n_2696),
.C(n_2706),
.Y(n_3365)
);

NAND2xp5_ASAP7_75t_L g3366 ( 
.A(n_2876),
.B(n_2881),
.Y(n_3366)
);

NOR2xp33_ASAP7_75t_R g3367 ( 
.A(n_2946),
.B(n_2739),
.Y(n_3367)
);

INVx1_ASAP7_75t_L g3368 ( 
.A(n_2901),
.Y(n_3368)
);

NOR2xp33_ASAP7_75t_R g3369 ( 
.A(n_2969),
.B(n_2492),
.Y(n_3369)
);

NAND2xp33_ASAP7_75t_R g3370 ( 
.A(n_2886),
.B(n_605),
.Y(n_3370)
);

HB1xp67_ASAP7_75t_L g3371 ( 
.A(n_3024),
.Y(n_3371)
);

AND2x4_ASAP7_75t_L g3372 ( 
.A(n_3093),
.B(n_2610),
.Y(n_3372)
);

INVx1_ASAP7_75t_L g3373 ( 
.A(n_2915),
.Y(n_3373)
);

CKINVDCx5p33_ASAP7_75t_R g3374 ( 
.A(n_2919),
.Y(n_3374)
);

INVxp67_ASAP7_75t_SL g3375 ( 
.A(n_3094),
.Y(n_3375)
);

NAND2xp33_ASAP7_75t_R g3376 ( 
.A(n_2987),
.B(n_2988),
.Y(n_3376)
);

AO21x1_ASAP7_75t_L g3377 ( 
.A1(n_3020),
.A2(n_2612),
.B(n_2711),
.Y(n_3377)
);

AND2x4_ASAP7_75t_L g3378 ( 
.A(n_3097),
.B(n_2610),
.Y(n_3378)
);

AND2x2_ASAP7_75t_L g3379 ( 
.A(n_3064),
.B(n_607),
.Y(n_3379)
);

AND2x2_ASAP7_75t_L g3380 ( 
.A(n_3064),
.B(n_3067),
.Y(n_3380)
);

HB1xp67_ASAP7_75t_L g3381 ( 
.A(n_3074),
.Y(n_3381)
);

OR2x6_ASAP7_75t_L g3382 ( 
.A(n_2987),
.B(n_2718),
.Y(n_3382)
);

HB1xp67_ASAP7_75t_L g3383 ( 
.A(n_3075),
.Y(n_3383)
);

CKINVDCx16_ASAP7_75t_R g3384 ( 
.A(n_2889),
.Y(n_3384)
);

CKINVDCx20_ASAP7_75t_R g3385 ( 
.A(n_3067),
.Y(n_3385)
);

INVx1_ASAP7_75t_L g3386 ( 
.A(n_2931),
.Y(n_3386)
);

NAND2xp5_ASAP7_75t_L g3387 ( 
.A(n_2933),
.B(n_2521),
.Y(n_3387)
);

BUFx3_ASAP7_75t_L g3388 ( 
.A(n_2988),
.Y(n_3388)
);

NAND2xp33_ASAP7_75t_R g3389 ( 
.A(n_3098),
.B(n_607),
.Y(n_3389)
);

AOI22xp33_ASAP7_75t_L g3390 ( 
.A1(n_2891),
.A2(n_2579),
.B1(n_2637),
.B2(n_2627),
.Y(n_3390)
);

AND2x2_ASAP7_75t_L g3391 ( 
.A(n_3129),
.B(n_2898),
.Y(n_3391)
);

INVx1_ASAP7_75t_L g3392 ( 
.A(n_3122),
.Y(n_3392)
);

HB1xp67_ASAP7_75t_L g3393 ( 
.A(n_3235),
.Y(n_3393)
);

AND2x2_ASAP7_75t_L g3394 ( 
.A(n_3143),
.B(n_2925),
.Y(n_3394)
);

OAI22xp33_ASAP7_75t_L g3395 ( 
.A1(n_3229),
.A2(n_2983),
.B1(n_3026),
.B2(n_2884),
.Y(n_3395)
);

INVx2_ASAP7_75t_L g3396 ( 
.A(n_3280),
.Y(n_3396)
);

NAND2xp5_ASAP7_75t_L g3397 ( 
.A(n_3123),
.B(n_3127),
.Y(n_3397)
);

INVx4_ASAP7_75t_SL g3398 ( 
.A(n_3156),
.Y(n_3398)
);

BUFx3_ASAP7_75t_L g3399 ( 
.A(n_3356),
.Y(n_3399)
);

OR2x2_ASAP7_75t_L g3400 ( 
.A(n_3162),
.B(n_2936),
.Y(n_3400)
);

OR2x2_ASAP7_75t_L g3401 ( 
.A(n_3176),
.B(n_2938),
.Y(n_3401)
);

INVx3_ASAP7_75t_L g3402 ( 
.A(n_3193),
.Y(n_3402)
);

INVx2_ASAP7_75t_L g3403 ( 
.A(n_3283),
.Y(n_3403)
);

INVx3_ASAP7_75t_L g3404 ( 
.A(n_3193),
.Y(n_3404)
);

INVx1_ASAP7_75t_L g3405 ( 
.A(n_3128),
.Y(n_3405)
);

INVx1_ASAP7_75t_L g3406 ( 
.A(n_3130),
.Y(n_3406)
);

BUFx3_ASAP7_75t_L g3407 ( 
.A(n_3227),
.Y(n_3407)
);

INVx1_ASAP7_75t_L g3408 ( 
.A(n_3138),
.Y(n_3408)
);

INVx2_ASAP7_75t_L g3409 ( 
.A(n_3256),
.Y(n_3409)
);

AND2x2_ASAP7_75t_L g3410 ( 
.A(n_3147),
.B(n_2948),
.Y(n_3410)
);

BUFx3_ASAP7_75t_L g3411 ( 
.A(n_3300),
.Y(n_3411)
);

INVx1_ASAP7_75t_L g3412 ( 
.A(n_3141),
.Y(n_3412)
);

BUFx3_ASAP7_75t_L g3413 ( 
.A(n_3306),
.Y(n_3413)
);

AOI221xp5_ASAP7_75t_L g3414 ( 
.A1(n_3268),
.A2(n_2984),
.B1(n_2914),
.B2(n_3025),
.C(n_3077),
.Y(n_3414)
);

INVx2_ASAP7_75t_L g3415 ( 
.A(n_3133),
.Y(n_3415)
);

AND2x4_ASAP7_75t_SL g3416 ( 
.A(n_3152),
.B(n_2899),
.Y(n_3416)
);

INVx1_ASAP7_75t_L g3417 ( 
.A(n_3145),
.Y(n_3417)
);

AOI22xp33_ASAP7_75t_SL g3418 ( 
.A1(n_3146),
.A2(n_3115),
.B1(n_3098),
.B2(n_3023),
.Y(n_3418)
);

AND2x2_ASAP7_75t_L g3419 ( 
.A(n_3222),
.B(n_3023),
.Y(n_3419)
);

HB1xp67_ASAP7_75t_L g3420 ( 
.A(n_3236),
.Y(n_3420)
);

INVx2_ASAP7_75t_L g3421 ( 
.A(n_3157),
.Y(n_3421)
);

INVx1_ASAP7_75t_L g3422 ( 
.A(n_3149),
.Y(n_3422)
);

INVx2_ASAP7_75t_L g3423 ( 
.A(n_3158),
.Y(n_3423)
);

AND2x2_ASAP7_75t_L g3424 ( 
.A(n_3248),
.B(n_2899),
.Y(n_3424)
);

AND2x2_ASAP7_75t_L g3425 ( 
.A(n_3275),
.B(n_2990),
.Y(n_3425)
);

BUFx2_ASAP7_75t_L g3426 ( 
.A(n_3250),
.Y(n_3426)
);

INVxp67_ASAP7_75t_SL g3427 ( 
.A(n_3377),
.Y(n_3427)
);

INVx2_ASAP7_75t_L g3428 ( 
.A(n_3164),
.Y(n_3428)
);

AOI33xp33_ASAP7_75t_L g3429 ( 
.A1(n_3213),
.A2(n_3111),
.A3(n_2967),
.B1(n_2970),
.B2(n_2971),
.B3(n_3021),
.Y(n_3429)
);

BUFx2_ASAP7_75t_L g3430 ( 
.A(n_3223),
.Y(n_3430)
);

INVx2_ASAP7_75t_L g3431 ( 
.A(n_3179),
.Y(n_3431)
);

INVx1_ASAP7_75t_L g3432 ( 
.A(n_3160),
.Y(n_3432)
);

INVx2_ASAP7_75t_SL g3433 ( 
.A(n_3131),
.Y(n_3433)
);

INVx2_ASAP7_75t_L g3434 ( 
.A(n_3182),
.Y(n_3434)
);

INVx1_ASAP7_75t_L g3435 ( 
.A(n_3165),
.Y(n_3435)
);

OR2x2_ASAP7_75t_SL g3436 ( 
.A(n_3293),
.B(n_2968),
.Y(n_3436)
);

INVx2_ASAP7_75t_L g3437 ( 
.A(n_3183),
.Y(n_3437)
);

INVx1_ASAP7_75t_L g3438 ( 
.A(n_3173),
.Y(n_3438)
);

OR2x2_ASAP7_75t_L g3439 ( 
.A(n_3139),
.B(n_2892),
.Y(n_3439)
);

INVx2_ASAP7_75t_L g3440 ( 
.A(n_3185),
.Y(n_3440)
);

INVx2_ASAP7_75t_L g3441 ( 
.A(n_3208),
.Y(n_3441)
);

OAI211xp5_ASAP7_75t_SL g3442 ( 
.A1(n_3189),
.A2(n_2902),
.B(n_2878),
.C(n_2980),
.Y(n_3442)
);

INVx2_ASAP7_75t_L g3443 ( 
.A(n_3245),
.Y(n_3443)
);

INVx1_ASAP7_75t_L g3444 ( 
.A(n_3184),
.Y(n_3444)
);

INVx2_ASAP7_75t_SL g3445 ( 
.A(n_3281),
.Y(n_3445)
);

NAND3xp33_ASAP7_75t_L g3446 ( 
.A(n_3177),
.B(n_3043),
.C(n_3107),
.Y(n_3446)
);

AOI21xp5_ASAP7_75t_L g3447 ( 
.A1(n_3319),
.A2(n_3339),
.B(n_3344),
.Y(n_3447)
);

AND2x2_ASAP7_75t_L g3448 ( 
.A(n_3258),
.B(n_2992),
.Y(n_3448)
);

INVx1_ASAP7_75t_L g3449 ( 
.A(n_3186),
.Y(n_3449)
);

AND2x4_ASAP7_75t_L g3450 ( 
.A(n_3169),
.B(n_2954),
.Y(n_3450)
);

INVx1_ASAP7_75t_L g3451 ( 
.A(n_3198),
.Y(n_3451)
);

AND2x2_ASAP7_75t_L g3452 ( 
.A(n_3231),
.B(n_2895),
.Y(n_3452)
);

BUFx3_ASAP7_75t_L g3453 ( 
.A(n_3360),
.Y(n_3453)
);

AND2x2_ASAP7_75t_L g3454 ( 
.A(n_3254),
.B(n_2896),
.Y(n_3454)
);

NOR2x1p5_ASAP7_75t_L g3455 ( 
.A(n_3269),
.B(n_3068),
.Y(n_3455)
);

AND2x4_ASAP7_75t_SL g3456 ( 
.A(n_3152),
.B(n_3068),
.Y(n_3456)
);

AND2x4_ASAP7_75t_L g3457 ( 
.A(n_3169),
.B(n_2954),
.Y(n_3457)
);

AND2x2_ASAP7_75t_L g3458 ( 
.A(n_3233),
.B(n_3239),
.Y(n_3458)
);

INVx1_ASAP7_75t_L g3459 ( 
.A(n_3259),
.Y(n_3459)
);

AND2x2_ASAP7_75t_L g3460 ( 
.A(n_3153),
.B(n_2951),
.Y(n_3460)
);

INVx1_ASAP7_75t_L g3461 ( 
.A(n_3265),
.Y(n_3461)
);

NAND2xp5_ASAP7_75t_L g3462 ( 
.A(n_3368),
.B(n_2955),
.Y(n_3462)
);

NAND2xp5_ASAP7_75t_L g3463 ( 
.A(n_3373),
.B(n_3014),
.Y(n_3463)
);

OR2x2_ASAP7_75t_L g3464 ( 
.A(n_3206),
.B(n_3211),
.Y(n_3464)
);

AND2x2_ASAP7_75t_L g3465 ( 
.A(n_3384),
.B(n_3196),
.Y(n_3465)
);

AND2x2_ASAP7_75t_L g3466 ( 
.A(n_3180),
.B(n_3040),
.Y(n_3466)
);

AOI22xp33_ASAP7_75t_L g3467 ( 
.A1(n_3132),
.A2(n_3262),
.B1(n_3246),
.B2(n_3287),
.Y(n_3467)
);

OAI211xp5_ASAP7_75t_L g3468 ( 
.A1(n_3274),
.A2(n_3110),
.B(n_3117),
.C(n_2937),
.Y(n_3468)
);

INVx2_ASAP7_75t_SL g3469 ( 
.A(n_3281),
.Y(n_3469)
);

INVx1_ASAP7_75t_L g3470 ( 
.A(n_3386),
.Y(n_3470)
);

AND2x2_ASAP7_75t_L g3471 ( 
.A(n_3201),
.B(n_3288),
.Y(n_3471)
);

INVx1_ASAP7_75t_L g3472 ( 
.A(n_3134),
.Y(n_3472)
);

HB1xp67_ASAP7_75t_L g3473 ( 
.A(n_3354),
.Y(n_3473)
);

AND2x2_ASAP7_75t_L g3474 ( 
.A(n_3209),
.B(n_3046),
.Y(n_3474)
);

AND2x2_ASAP7_75t_L g3475 ( 
.A(n_3195),
.B(n_3052),
.Y(n_3475)
);

INVx1_ASAP7_75t_L g3476 ( 
.A(n_3140),
.Y(n_3476)
);

INVx1_ASAP7_75t_L g3477 ( 
.A(n_3148),
.Y(n_3477)
);

INVx3_ASAP7_75t_L g3478 ( 
.A(n_3175),
.Y(n_3478)
);

HB1xp67_ASAP7_75t_L g3479 ( 
.A(n_3375),
.Y(n_3479)
);

OR2x2_ASAP7_75t_L g3480 ( 
.A(n_3234),
.B(n_3018),
.Y(n_3480)
);

OR2x2_ASAP7_75t_L g3481 ( 
.A(n_3263),
.B(n_3039),
.Y(n_3481)
);

AND2x2_ASAP7_75t_L g3482 ( 
.A(n_3210),
.B(n_3063),
.Y(n_3482)
);

AND2x2_ASAP7_75t_L g3483 ( 
.A(n_3332),
.B(n_3039),
.Y(n_3483)
);

NAND2xp5_ASAP7_75t_SL g3484 ( 
.A(n_3217),
.B(n_3086),
.Y(n_3484)
);

AND2x2_ASAP7_75t_L g3485 ( 
.A(n_3340),
.B(n_3041),
.Y(n_3485)
);

INVx2_ASAP7_75t_SL g3486 ( 
.A(n_3167),
.Y(n_3486)
);

INVx3_ASAP7_75t_L g3487 ( 
.A(n_3175),
.Y(n_3487)
);

INVx1_ASAP7_75t_L g3488 ( 
.A(n_3301),
.Y(n_3488)
);

BUFx3_ASAP7_75t_L g3489 ( 
.A(n_3385),
.Y(n_3489)
);

INVx2_ASAP7_75t_L g3490 ( 
.A(n_3284),
.Y(n_3490)
);

INVx3_ASAP7_75t_L g3491 ( 
.A(n_3199),
.Y(n_3491)
);

INVx2_ASAP7_75t_L g3492 ( 
.A(n_3285),
.Y(n_3492)
);

INVx3_ASAP7_75t_SL g3493 ( 
.A(n_3320),
.Y(n_3493)
);

AND2x2_ASAP7_75t_L g3494 ( 
.A(n_3347),
.B(n_3041),
.Y(n_3494)
);

AOI22xp33_ASAP7_75t_SL g3495 ( 
.A1(n_3269),
.A2(n_3004),
.B1(n_2968),
.B2(n_3016),
.Y(n_3495)
);

INVx2_ASAP7_75t_L g3496 ( 
.A(n_3286),
.Y(n_3496)
);

INVx1_ASAP7_75t_L g3497 ( 
.A(n_3303),
.Y(n_3497)
);

AND2x2_ASAP7_75t_L g3498 ( 
.A(n_3381),
.B(n_3044),
.Y(n_3498)
);

NAND2xp5_ASAP7_75t_L g3499 ( 
.A(n_3387),
.B(n_3044),
.Y(n_3499)
);

INVx1_ASAP7_75t_L g3500 ( 
.A(n_3313),
.Y(n_3500)
);

INVxp67_ASAP7_75t_SL g3501 ( 
.A(n_3359),
.Y(n_3501)
);

AND2x2_ASAP7_75t_L g3502 ( 
.A(n_3383),
.B(n_3079),
.Y(n_3502)
);

AND2x2_ASAP7_75t_L g3503 ( 
.A(n_3251),
.B(n_3079),
.Y(n_3503)
);

INVx3_ASAP7_75t_L g3504 ( 
.A(n_3199),
.Y(n_3504)
);

AOI22xp5_ASAP7_75t_L g3505 ( 
.A1(n_3232),
.A2(n_2945),
.B1(n_2927),
.B2(n_2934),
.Y(n_3505)
);

AND2x2_ASAP7_75t_L g3506 ( 
.A(n_3252),
.B(n_3086),
.Y(n_3506)
);

INVx1_ASAP7_75t_L g3507 ( 
.A(n_3322),
.Y(n_3507)
);

AND2x2_ASAP7_75t_L g3508 ( 
.A(n_3242),
.B(n_3088),
.Y(n_3508)
);

AND2x2_ASAP7_75t_L g3509 ( 
.A(n_3302),
.B(n_3088),
.Y(n_3509)
);

INVx1_ASAP7_75t_L g3510 ( 
.A(n_3336),
.Y(n_3510)
);

AND2x4_ASAP7_75t_L g3511 ( 
.A(n_3226),
.B(n_3112),
.Y(n_3511)
);

INVx1_ASAP7_75t_L g3512 ( 
.A(n_3366),
.Y(n_3512)
);

INVx2_ASAP7_75t_L g3513 ( 
.A(n_3290),
.Y(n_3513)
);

BUFx2_ASAP7_75t_L g3514 ( 
.A(n_3357),
.Y(n_3514)
);

AND2x4_ASAP7_75t_L g3515 ( 
.A(n_3226),
.B(n_3083),
.Y(n_3515)
);

INVxp67_ASAP7_75t_L g3516 ( 
.A(n_3308),
.Y(n_3516)
);

OR2x2_ASAP7_75t_L g3517 ( 
.A(n_3174),
.B(n_2972),
.Y(n_3517)
);

INVx2_ASAP7_75t_L g3518 ( 
.A(n_3296),
.Y(n_3518)
);

AND2x2_ASAP7_75t_L g3519 ( 
.A(n_3270),
.B(n_2972),
.Y(n_3519)
);

OAI22xp5_ASAP7_75t_L g3520 ( 
.A1(n_3188),
.A2(n_3004),
.B1(n_2942),
.B2(n_2943),
.Y(n_3520)
);

INVx1_ASAP7_75t_L g3521 ( 
.A(n_3243),
.Y(n_3521)
);

BUFx3_ASAP7_75t_L g3522 ( 
.A(n_3310),
.Y(n_3522)
);

BUFx3_ASAP7_75t_L g3523 ( 
.A(n_3136),
.Y(n_3523)
);

HB1xp67_ASAP7_75t_L g3524 ( 
.A(n_3326),
.Y(n_3524)
);

AND2x2_ASAP7_75t_L g3525 ( 
.A(n_3203),
.B(n_2974),
.Y(n_3525)
);

OAI22xp5_ASAP7_75t_L g3526 ( 
.A1(n_3214),
.A2(n_2885),
.B1(n_2826),
.B2(n_3006),
.Y(n_3526)
);

AND2x2_ASAP7_75t_L g3527 ( 
.A(n_3271),
.B(n_2976),
.Y(n_3527)
);

AND2x2_ASAP7_75t_L g3528 ( 
.A(n_3349),
.B(n_2976),
.Y(n_3528)
);

AND2x2_ASAP7_75t_L g3529 ( 
.A(n_3349),
.B(n_2977),
.Y(n_3529)
);

AND2x2_ASAP7_75t_L g3530 ( 
.A(n_3295),
.B(n_3282),
.Y(n_3530)
);

INVx2_ASAP7_75t_L g3531 ( 
.A(n_3276),
.Y(n_3531)
);

CKINVDCx20_ASAP7_75t_R g3532 ( 
.A(n_3159),
.Y(n_3532)
);

BUFx2_ASAP7_75t_L g3533 ( 
.A(n_3369),
.Y(n_3533)
);

OR2x2_ASAP7_75t_L g3534 ( 
.A(n_3249),
.B(n_3253),
.Y(n_3534)
);

AND2x2_ASAP7_75t_L g3535 ( 
.A(n_3237),
.B(n_2977),
.Y(n_3535)
);

OR2x2_ASAP7_75t_L g3536 ( 
.A(n_3172),
.B(n_3103),
.Y(n_3536)
);

NAND2x1_ASAP7_75t_L g3537 ( 
.A(n_3156),
.B(n_2965),
.Y(n_3537)
);

AND2x2_ASAP7_75t_L g3538 ( 
.A(n_3362),
.B(n_2871),
.Y(n_3538)
);

AND2x2_ASAP7_75t_L g3539 ( 
.A(n_3362),
.B(n_2871),
.Y(n_3539)
);

INVx2_ASAP7_75t_L g3540 ( 
.A(n_3372),
.Y(n_3540)
);

INVxp67_ASAP7_75t_SL g3541 ( 
.A(n_3328),
.Y(n_3541)
);

OAI31xp33_ASAP7_75t_SL g3542 ( 
.A1(n_3137),
.A2(n_3228),
.A3(n_3247),
.B(n_3121),
.Y(n_3542)
);

BUFx3_ASAP7_75t_L g3543 ( 
.A(n_3191),
.Y(n_3543)
);

INVx3_ASAP7_75t_L g3544 ( 
.A(n_3200),
.Y(n_3544)
);

AO21x2_ASAP7_75t_L g3545 ( 
.A1(n_3345),
.A2(n_3365),
.B(n_3297),
.Y(n_3545)
);

NAND2xp5_ASAP7_75t_L g3546 ( 
.A(n_3181),
.B(n_3099),
.Y(n_3546)
);

AOI21xp33_ASAP7_75t_L g3547 ( 
.A1(n_3389),
.A2(n_2746),
.B(n_2530),
.Y(n_3547)
);

BUFx3_ASAP7_75t_L g3548 ( 
.A(n_3144),
.Y(n_3548)
);

INVx2_ASAP7_75t_L g3549 ( 
.A(n_3372),
.Y(n_3549)
);

AND2x2_ASAP7_75t_L g3550 ( 
.A(n_3378),
.B(n_2883),
.Y(n_3550)
);

INVx2_ASAP7_75t_L g3551 ( 
.A(n_3378),
.Y(n_3551)
);

INVx2_ASAP7_75t_L g3552 ( 
.A(n_3171),
.Y(n_3552)
);

INVx2_ASAP7_75t_L g3553 ( 
.A(n_3171),
.Y(n_3553)
);

INVx2_ASAP7_75t_L g3554 ( 
.A(n_3178),
.Y(n_3554)
);

HB1xp67_ASAP7_75t_L g3555 ( 
.A(n_3371),
.Y(n_3555)
);

AND2x2_ASAP7_75t_L g3556 ( 
.A(n_3323),
.B(n_3363),
.Y(n_3556)
);

AND2x2_ASAP7_75t_L g3557 ( 
.A(n_3338),
.B(n_2883),
.Y(n_3557)
);

NAND2xp5_ASAP7_75t_L g3558 ( 
.A(n_3192),
.B(n_3099),
.Y(n_3558)
);

AND2x2_ASAP7_75t_L g3559 ( 
.A(n_3219),
.B(n_2890),
.Y(n_3559)
);

INVx4_ASAP7_75t_L g3560 ( 
.A(n_3200),
.Y(n_3560)
);

OR2x2_ASAP7_75t_L g3561 ( 
.A(n_3291),
.B(n_3103),
.Y(n_3561)
);

NAND2xp5_ASAP7_75t_L g3562 ( 
.A(n_3524),
.B(n_3390),
.Y(n_3562)
);

AND2x4_ASAP7_75t_L g3563 ( 
.A(n_3398),
.B(n_3298),
.Y(n_3563)
);

NAND2xp5_ASAP7_75t_SL g3564 ( 
.A(n_3430),
.B(n_3178),
.Y(n_3564)
);

AND2x4_ASAP7_75t_L g3565 ( 
.A(n_3398),
.B(n_3219),
.Y(n_3565)
);

INVx2_ASAP7_75t_L g3566 ( 
.A(n_3479),
.Y(n_3566)
);

NAND2xp5_ASAP7_75t_L g3567 ( 
.A(n_3524),
.B(n_3329),
.Y(n_3567)
);

AND2x2_ASAP7_75t_L g3568 ( 
.A(n_3458),
.B(n_3391),
.Y(n_3568)
);

NAND2xp5_ASAP7_75t_SL g3569 ( 
.A(n_3447),
.B(n_3220),
.Y(n_3569)
);

AND2x2_ASAP7_75t_L g3570 ( 
.A(n_3394),
.B(n_3289),
.Y(n_3570)
);

INVx1_ASAP7_75t_L g3571 ( 
.A(n_3393),
.Y(n_3571)
);

OR2x2_ASAP7_75t_L g3572 ( 
.A(n_3473),
.B(n_3325),
.Y(n_3572)
);

INVx2_ASAP7_75t_L g3573 ( 
.A(n_3415),
.Y(n_3573)
);

INVx1_ASAP7_75t_L g3574 ( 
.A(n_3393),
.Y(n_3574)
);

INVxp67_ASAP7_75t_SL g3575 ( 
.A(n_3479),
.Y(n_3575)
);

AND2x4_ASAP7_75t_SL g3576 ( 
.A(n_3560),
.B(n_3167),
.Y(n_3576)
);

AND2x2_ASAP7_75t_L g3577 ( 
.A(n_3530),
.B(n_3314),
.Y(n_3577)
);

HB1xp67_ASAP7_75t_L g3578 ( 
.A(n_3420),
.Y(n_3578)
);

AND2x2_ASAP7_75t_L g3579 ( 
.A(n_3460),
.B(n_3353),
.Y(n_3579)
);

AND2x2_ASAP7_75t_L g3580 ( 
.A(n_3465),
.B(n_3525),
.Y(n_3580)
);

NAND2x1_ASAP7_75t_L g3581 ( 
.A(n_3560),
.B(n_3218),
.Y(n_3581)
);

NAND2xp5_ASAP7_75t_L g3582 ( 
.A(n_3420),
.B(n_3084),
.Y(n_3582)
);

INVx2_ASAP7_75t_L g3583 ( 
.A(n_3396),
.Y(n_3583)
);

NAND2xp5_ASAP7_75t_L g3584 ( 
.A(n_3521),
.B(n_3168),
.Y(n_3584)
);

INVx1_ASAP7_75t_L g3585 ( 
.A(n_3470),
.Y(n_3585)
);

AND2x4_ASAP7_75t_L g3586 ( 
.A(n_3398),
.B(n_3220),
.Y(n_3586)
);

AND2x4_ASAP7_75t_L g3587 ( 
.A(n_3450),
.B(n_3261),
.Y(n_3587)
);

AND2x2_ASAP7_75t_L g3588 ( 
.A(n_3471),
.B(n_3261),
.Y(n_3588)
);

NAND2xp5_ASAP7_75t_L g3589 ( 
.A(n_3510),
.B(n_3337),
.Y(n_3589)
);

AOI22xp33_ASAP7_75t_SL g3590 ( 
.A1(n_3426),
.A2(n_3205),
.B1(n_3202),
.B2(n_3224),
.Y(n_3590)
);

AND2x2_ASAP7_75t_L g3591 ( 
.A(n_3476),
.B(n_3264),
.Y(n_3591)
);

AND2x2_ASAP7_75t_L g3592 ( 
.A(n_3477),
.B(n_3264),
.Y(n_3592)
);

INVx1_ASAP7_75t_L g3593 ( 
.A(n_3400),
.Y(n_3593)
);

INVx2_ASAP7_75t_L g3594 ( 
.A(n_3403),
.Y(n_3594)
);

AND2x2_ASAP7_75t_L g3595 ( 
.A(n_3473),
.B(n_3348),
.Y(n_3595)
);

NAND2xp5_ASAP7_75t_L g3596 ( 
.A(n_3512),
.B(n_3272),
.Y(n_3596)
);

INVx2_ASAP7_75t_L g3597 ( 
.A(n_3555),
.Y(n_3597)
);

NAND2xp5_ASAP7_75t_L g3598 ( 
.A(n_3546),
.B(n_3305),
.Y(n_3598)
);

NOR2xp33_ASAP7_75t_SL g3599 ( 
.A(n_3493),
.B(n_3312),
.Y(n_3599)
);

AND2x2_ASAP7_75t_L g3600 ( 
.A(n_3452),
.B(n_3364),
.Y(n_3600)
);

INVx1_ASAP7_75t_L g3601 ( 
.A(n_3401),
.Y(n_3601)
);

INVx2_ASAP7_75t_L g3602 ( 
.A(n_3421),
.Y(n_3602)
);

AND2x2_ASAP7_75t_L g3603 ( 
.A(n_3482),
.B(n_3316),
.Y(n_3603)
);

AND2x2_ASAP7_75t_L g3604 ( 
.A(n_3425),
.B(n_3475),
.Y(n_3604)
);

AND2x2_ASAP7_75t_L g3605 ( 
.A(n_3466),
.B(n_3474),
.Y(n_3605)
);

NAND2xp5_ASAP7_75t_L g3606 ( 
.A(n_3546),
.B(n_3273),
.Y(n_3606)
);

NAND2xp5_ASAP7_75t_L g3607 ( 
.A(n_3558),
.B(n_3351),
.Y(n_3607)
);

INVx1_ASAP7_75t_L g3608 ( 
.A(n_3461),
.Y(n_3608)
);

AND2x2_ASAP7_75t_L g3609 ( 
.A(n_3410),
.B(n_3324),
.Y(n_3609)
);

AND2x4_ASAP7_75t_L g3610 ( 
.A(n_3450),
.B(n_3144),
.Y(n_3610)
);

NAND2xp5_ASAP7_75t_L g3611 ( 
.A(n_3558),
.B(n_3215),
.Y(n_3611)
);

AND2x2_ASAP7_75t_L g3612 ( 
.A(n_3535),
.B(n_3327),
.Y(n_3612)
);

OR2x2_ASAP7_75t_L g3613 ( 
.A(n_3409),
.B(n_3341),
.Y(n_3613)
);

INVx1_ASAP7_75t_L g3614 ( 
.A(n_3397),
.Y(n_3614)
);

HB1xp67_ASAP7_75t_L g3615 ( 
.A(n_3555),
.Y(n_3615)
);

AND2x2_ASAP7_75t_L g3616 ( 
.A(n_3508),
.B(n_3350),
.Y(n_3616)
);

AND2x2_ASAP7_75t_L g3617 ( 
.A(n_3519),
.B(n_3550),
.Y(n_3617)
);

AND2x2_ASAP7_75t_L g3618 ( 
.A(n_3540),
.B(n_3255),
.Y(n_3618)
);

INVx2_ASAP7_75t_L g3619 ( 
.A(n_3423),
.Y(n_3619)
);

AND2x2_ASAP7_75t_L g3620 ( 
.A(n_3549),
.B(n_3267),
.Y(n_3620)
);

INVx2_ASAP7_75t_L g3621 ( 
.A(n_3428),
.Y(n_3621)
);

AND2x2_ASAP7_75t_L g3622 ( 
.A(n_3551),
.B(n_3557),
.Y(n_3622)
);

OR2x6_ASAP7_75t_L g3623 ( 
.A(n_3537),
.B(n_3163),
.Y(n_3623)
);

AND2x2_ASAP7_75t_L g3624 ( 
.A(n_3424),
.B(n_3346),
.Y(n_3624)
);

AND2x4_ASAP7_75t_L g3625 ( 
.A(n_3457),
.B(n_3125),
.Y(n_3625)
);

NOR2xp67_ASAP7_75t_L g3626 ( 
.A(n_3516),
.B(n_3330),
.Y(n_3626)
);

NAND2xp5_ASAP7_75t_L g3627 ( 
.A(n_3472),
.B(n_3204),
.Y(n_3627)
);

OAI22xp5_ASAP7_75t_L g3628 ( 
.A1(n_3467),
.A2(n_3304),
.B1(n_3163),
.B2(n_3194),
.Y(n_3628)
);

INVx2_ASAP7_75t_L g3629 ( 
.A(n_3431),
.Y(n_3629)
);

INVx1_ASAP7_75t_L g3630 ( 
.A(n_3397),
.Y(n_3630)
);

HB1xp67_ASAP7_75t_L g3631 ( 
.A(n_3434),
.Y(n_3631)
);

INVx1_ASAP7_75t_L g3632 ( 
.A(n_3488),
.Y(n_3632)
);

INVx2_ASAP7_75t_L g3633 ( 
.A(n_3437),
.Y(n_3633)
);

AND2x2_ASAP7_75t_L g3634 ( 
.A(n_3531),
.B(n_3238),
.Y(n_3634)
);

INVx1_ASAP7_75t_L g3635 ( 
.A(n_3497),
.Y(n_3635)
);

AND2x4_ASAP7_75t_L g3636 ( 
.A(n_3457),
.B(n_3142),
.Y(n_3636)
);

INVx1_ASAP7_75t_L g3637 ( 
.A(n_3500),
.Y(n_3637)
);

AND2x2_ASAP7_75t_L g3638 ( 
.A(n_3506),
.B(n_3238),
.Y(n_3638)
);

INVx1_ASAP7_75t_L g3639 ( 
.A(n_3507),
.Y(n_3639)
);

NAND2xp33_ASAP7_75t_SL g3640 ( 
.A(n_3455),
.B(n_3493),
.Y(n_3640)
);

AND2x2_ASAP7_75t_L g3641 ( 
.A(n_3538),
.B(n_3244),
.Y(n_3641)
);

HB1xp67_ASAP7_75t_L g3642 ( 
.A(n_3440),
.Y(n_3642)
);

INVx1_ASAP7_75t_L g3643 ( 
.A(n_3392),
.Y(n_3643)
);

INVx1_ASAP7_75t_L g3644 ( 
.A(n_3405),
.Y(n_3644)
);

NAND2xp5_ASAP7_75t_SL g3645 ( 
.A(n_3447),
.B(n_3355),
.Y(n_3645)
);

INVx2_ASAP7_75t_L g3646 ( 
.A(n_3441),
.Y(n_3646)
);

AND2x4_ASAP7_75t_SL g3647 ( 
.A(n_3478),
.B(n_3218),
.Y(n_3647)
);

INVx1_ASAP7_75t_L g3648 ( 
.A(n_3406),
.Y(n_3648)
);

AND2x2_ASAP7_75t_L g3649 ( 
.A(n_3539),
.B(n_3244),
.Y(n_3649)
);

AND2x2_ASAP7_75t_L g3650 ( 
.A(n_3528),
.B(n_3277),
.Y(n_3650)
);

INVx1_ASAP7_75t_L g3651 ( 
.A(n_3408),
.Y(n_3651)
);

INVx2_ASAP7_75t_L g3652 ( 
.A(n_3443),
.Y(n_3652)
);

INVx2_ASAP7_75t_L g3653 ( 
.A(n_3573),
.Y(n_3653)
);

AND2x2_ASAP7_75t_L g3654 ( 
.A(n_3617),
.B(n_3503),
.Y(n_3654)
);

NAND2xp5_ASAP7_75t_L g3655 ( 
.A(n_3611),
.B(n_3527),
.Y(n_3655)
);

AOI22xp33_ASAP7_75t_L g3656 ( 
.A1(n_3628),
.A2(n_3467),
.B1(n_3442),
.B2(n_3446),
.Y(n_3656)
);

INVx1_ASAP7_75t_L g3657 ( 
.A(n_3578),
.Y(n_3657)
);

INVx2_ASAP7_75t_L g3658 ( 
.A(n_3573),
.Y(n_3658)
);

AND2x2_ASAP7_75t_L g3659 ( 
.A(n_3568),
.B(n_3464),
.Y(n_3659)
);

NAND2xp5_ASAP7_75t_L g3660 ( 
.A(n_3611),
.B(n_3454),
.Y(n_3660)
);

INVx2_ASAP7_75t_L g3661 ( 
.A(n_3602),
.Y(n_3661)
);

INVx1_ASAP7_75t_L g3662 ( 
.A(n_3578),
.Y(n_3662)
);

NAND2xp5_ASAP7_75t_L g3663 ( 
.A(n_3571),
.B(n_3448),
.Y(n_3663)
);

INVx2_ASAP7_75t_L g3664 ( 
.A(n_3602),
.Y(n_3664)
);

INVx1_ASAP7_75t_SL g3665 ( 
.A(n_3572),
.Y(n_3665)
);

INVx1_ASAP7_75t_L g3666 ( 
.A(n_3585),
.Y(n_3666)
);

NOR2xp33_ASAP7_75t_R g3667 ( 
.A(n_3640),
.B(n_3376),
.Y(n_3667)
);

OR2x2_ASAP7_75t_L g3668 ( 
.A(n_3575),
.B(n_3439),
.Y(n_3668)
);

OR2x2_ASAP7_75t_L g3669 ( 
.A(n_3575),
.B(n_3480),
.Y(n_3669)
);

AND2x2_ASAP7_75t_L g3670 ( 
.A(n_3604),
.B(n_3419),
.Y(n_3670)
);

BUFx3_ASAP7_75t_L g3671 ( 
.A(n_3576),
.Y(n_3671)
);

OR2x2_ASAP7_75t_L g3672 ( 
.A(n_3593),
.B(n_3481),
.Y(n_3672)
);

INVx1_ASAP7_75t_L g3673 ( 
.A(n_3632),
.Y(n_3673)
);

BUFx2_ASAP7_75t_L g3674 ( 
.A(n_3640),
.Y(n_3674)
);

OR2x2_ASAP7_75t_L g3675 ( 
.A(n_3601),
.B(n_3517),
.Y(n_3675)
);

AND2x2_ASAP7_75t_L g3676 ( 
.A(n_3600),
.B(n_3529),
.Y(n_3676)
);

AND2x4_ASAP7_75t_L g3677 ( 
.A(n_3587),
.B(n_3516),
.Y(n_3677)
);

AND2x2_ASAP7_75t_L g3678 ( 
.A(n_3580),
.B(n_3509),
.Y(n_3678)
);

INVx2_ASAP7_75t_L g3679 ( 
.A(n_3646),
.Y(n_3679)
);

NOR2x1_ASAP7_75t_L g3680 ( 
.A(n_3581),
.B(n_3407),
.Y(n_3680)
);

INVx1_ASAP7_75t_L g3681 ( 
.A(n_3635),
.Y(n_3681)
);

INVx1_ASAP7_75t_L g3682 ( 
.A(n_3637),
.Y(n_3682)
);

AND2x4_ASAP7_75t_L g3683 ( 
.A(n_3587),
.B(n_3515),
.Y(n_3683)
);

AND2x2_ASAP7_75t_L g3684 ( 
.A(n_3570),
.B(n_3624),
.Y(n_3684)
);

NAND2xp5_ASAP7_75t_L g3685 ( 
.A(n_3574),
.B(n_3534),
.Y(n_3685)
);

NAND2xp5_ASAP7_75t_L g3686 ( 
.A(n_3614),
.B(n_3505),
.Y(n_3686)
);

BUFx2_ASAP7_75t_L g3687 ( 
.A(n_3636),
.Y(n_3687)
);

AND2x2_ASAP7_75t_L g3688 ( 
.A(n_3605),
.B(n_3483),
.Y(n_3688)
);

INVx2_ASAP7_75t_L g3689 ( 
.A(n_3646),
.Y(n_3689)
);

HB1xp67_ASAP7_75t_L g3690 ( 
.A(n_3615),
.Y(n_3690)
);

AND2x2_ASAP7_75t_L g3691 ( 
.A(n_3622),
.B(n_3559),
.Y(n_3691)
);

OR2x2_ASAP7_75t_L g3692 ( 
.A(n_3615),
.B(n_3561),
.Y(n_3692)
);

NAND2xp5_ASAP7_75t_L g3693 ( 
.A(n_3630),
.B(n_3505),
.Y(n_3693)
);

INVxp67_ASAP7_75t_SL g3694 ( 
.A(n_3631),
.Y(n_3694)
);

AND2x4_ASAP7_75t_L g3695 ( 
.A(n_3623),
.B(n_3515),
.Y(n_3695)
);

OR2x2_ASAP7_75t_L g3696 ( 
.A(n_3631),
.B(n_3536),
.Y(n_3696)
);

INVx1_ASAP7_75t_L g3697 ( 
.A(n_3639),
.Y(n_3697)
);

NAND2xp5_ASAP7_75t_L g3698 ( 
.A(n_3584),
.B(n_3490),
.Y(n_3698)
);

AND2x2_ASAP7_75t_L g3699 ( 
.A(n_3577),
.B(n_3556),
.Y(n_3699)
);

INVxp67_ASAP7_75t_L g3700 ( 
.A(n_3642),
.Y(n_3700)
);

AND2x2_ASAP7_75t_L g3701 ( 
.A(n_3650),
.B(n_3485),
.Y(n_3701)
);

NAND2xp5_ASAP7_75t_L g3702 ( 
.A(n_3584),
.B(n_3492),
.Y(n_3702)
);

INVx2_ASAP7_75t_L g3703 ( 
.A(n_3652),
.Y(n_3703)
);

INVx2_ASAP7_75t_L g3704 ( 
.A(n_3652),
.Y(n_3704)
);

HB1xp67_ASAP7_75t_L g3705 ( 
.A(n_3642),
.Y(n_3705)
);

AND2x2_ASAP7_75t_L g3706 ( 
.A(n_3579),
.B(n_3494),
.Y(n_3706)
);

CKINVDCx5p33_ASAP7_75t_R g3707 ( 
.A(n_3576),
.Y(n_3707)
);

INVx2_ASAP7_75t_L g3708 ( 
.A(n_3619),
.Y(n_3708)
);

INVx1_ASAP7_75t_L g3709 ( 
.A(n_3608),
.Y(n_3709)
);

AND2x2_ASAP7_75t_L g3710 ( 
.A(n_3588),
.B(n_3498),
.Y(n_3710)
);

AND2x2_ASAP7_75t_L g3711 ( 
.A(n_3616),
.B(n_3502),
.Y(n_3711)
);

AND2x2_ASAP7_75t_L g3712 ( 
.A(n_3641),
.B(n_3649),
.Y(n_3712)
);

INVx2_ASAP7_75t_L g3713 ( 
.A(n_3621),
.Y(n_3713)
);

AND2x2_ASAP7_75t_L g3714 ( 
.A(n_3612),
.B(n_3523),
.Y(n_3714)
);

INVx1_ASAP7_75t_L g3715 ( 
.A(n_3643),
.Y(n_3715)
);

AND2x2_ASAP7_75t_L g3716 ( 
.A(n_3638),
.B(n_3543),
.Y(n_3716)
);

NAND2xp5_ASAP7_75t_L g3717 ( 
.A(n_3598),
.B(n_3496),
.Y(n_3717)
);

AND2x4_ASAP7_75t_L g3718 ( 
.A(n_3623),
.B(n_3501),
.Y(n_3718)
);

OR2x2_ASAP7_75t_L g3719 ( 
.A(n_3566),
.B(n_3499),
.Y(n_3719)
);

NAND2xp5_ASAP7_75t_L g3720 ( 
.A(n_3598),
.B(n_3513),
.Y(n_3720)
);

INVx1_ASAP7_75t_L g3721 ( 
.A(n_3644),
.Y(n_3721)
);

AND2x2_ASAP7_75t_L g3722 ( 
.A(n_3595),
.B(n_3545),
.Y(n_3722)
);

INVx3_ASAP7_75t_L g3723 ( 
.A(n_3671),
.Y(n_3723)
);

NAND2xp5_ASAP7_75t_L g3724 ( 
.A(n_3686),
.B(n_3693),
.Y(n_3724)
);

INVx2_ASAP7_75t_L g3725 ( 
.A(n_3705),
.Y(n_3725)
);

INVx1_ASAP7_75t_L g3726 ( 
.A(n_3705),
.Y(n_3726)
);

INVx1_ASAP7_75t_L g3727 ( 
.A(n_3692),
.Y(n_3727)
);

INVx2_ASAP7_75t_L g3728 ( 
.A(n_3700),
.Y(n_3728)
);

OR2x2_ASAP7_75t_L g3729 ( 
.A(n_3696),
.B(n_3583),
.Y(n_3729)
);

INVx2_ASAP7_75t_L g3730 ( 
.A(n_3700),
.Y(n_3730)
);

HB1xp67_ASAP7_75t_L g3731 ( 
.A(n_3694),
.Y(n_3731)
);

AOI22xp5_ASAP7_75t_L g3732 ( 
.A1(n_3656),
.A2(n_3628),
.B1(n_3626),
.B2(n_3569),
.Y(n_3732)
);

INVx1_ASAP7_75t_L g3733 ( 
.A(n_3717),
.Y(n_3733)
);

NAND2xp5_ASAP7_75t_L g3734 ( 
.A(n_3720),
.B(n_3607),
.Y(n_3734)
);

NAND2xp5_ASAP7_75t_L g3735 ( 
.A(n_3655),
.B(n_3607),
.Y(n_3735)
);

NOR2xp33_ASAP7_75t_SL g3736 ( 
.A(n_3707),
.B(n_3599),
.Y(n_3736)
);

INVx1_ASAP7_75t_L g3737 ( 
.A(n_3657),
.Y(n_3737)
);

OR2x2_ASAP7_75t_L g3738 ( 
.A(n_3694),
.B(n_3672),
.Y(n_3738)
);

NAND2x1p5_ASAP7_75t_L g3739 ( 
.A(n_3671),
.B(n_3411),
.Y(n_3739)
);

INVx1_ASAP7_75t_L g3740 ( 
.A(n_3662),
.Y(n_3740)
);

XNOR2xp5_ASAP7_75t_L g3741 ( 
.A(n_3707),
.B(n_3307),
.Y(n_3741)
);

OAI322xp33_ASAP7_75t_L g3742 ( 
.A1(n_3660),
.A2(n_3567),
.A3(n_3569),
.B1(n_3645),
.B2(n_3606),
.C1(n_3395),
.C2(n_3589),
.Y(n_3742)
);

OR2x6_ASAP7_75t_L g3743 ( 
.A(n_3680),
.B(n_3623),
.Y(n_3743)
);

AND2x2_ASAP7_75t_L g3744 ( 
.A(n_3687),
.B(n_3670),
.Y(n_3744)
);

INVx1_ASAP7_75t_L g3745 ( 
.A(n_3690),
.Y(n_3745)
);

NOR4xp25_ASAP7_75t_L g3746 ( 
.A(n_3656),
.B(n_3589),
.C(n_3645),
.D(n_3486),
.Y(n_3746)
);

AND2x4_ASAP7_75t_L g3747 ( 
.A(n_3695),
.B(n_3563),
.Y(n_3747)
);

INVx3_ASAP7_75t_SL g3748 ( 
.A(n_3716),
.Y(n_3748)
);

AOI22xp5_ASAP7_75t_L g3749 ( 
.A1(n_3674),
.A2(n_3590),
.B1(n_3484),
.B2(n_3333),
.Y(n_3749)
);

INVx1_ASAP7_75t_L g3750 ( 
.A(n_3666),
.Y(n_3750)
);

INVx2_ASAP7_75t_L g3751 ( 
.A(n_3690),
.Y(n_3751)
);

INVx1_ASAP7_75t_L g3752 ( 
.A(n_3673),
.Y(n_3752)
);

INVx1_ASAP7_75t_L g3753 ( 
.A(n_3681),
.Y(n_3753)
);

OR2x6_ASAP7_75t_L g3754 ( 
.A(n_3695),
.B(n_3514),
.Y(n_3754)
);

INVx1_ASAP7_75t_L g3755 ( 
.A(n_3682),
.Y(n_3755)
);

HB1xp67_ASAP7_75t_L g3756 ( 
.A(n_3668),
.Y(n_3756)
);

INVx1_ASAP7_75t_L g3757 ( 
.A(n_3653),
.Y(n_3757)
);

AOI22xp5_ASAP7_75t_L g3758 ( 
.A1(n_3665),
.A2(n_3590),
.B1(n_3484),
.B2(n_3343),
.Y(n_3758)
);

INVx2_ASAP7_75t_L g3759 ( 
.A(n_3653),
.Y(n_3759)
);

INVx2_ASAP7_75t_L g3760 ( 
.A(n_3658),
.Y(n_3760)
);

INVx4_ASAP7_75t_L g3761 ( 
.A(n_3695),
.Y(n_3761)
);

OAI22xp5_ASAP7_75t_L g3762 ( 
.A1(n_3683),
.A2(n_3563),
.B1(n_3647),
.B2(n_3625),
.Y(n_3762)
);

NAND2xp5_ASAP7_75t_L g3763 ( 
.A(n_3688),
.B(n_3698),
.Y(n_3763)
);

HB1xp67_ASAP7_75t_L g3764 ( 
.A(n_3669),
.Y(n_3764)
);

AND2x2_ASAP7_75t_L g3765 ( 
.A(n_3677),
.B(n_3591),
.Y(n_3765)
);

AND2x2_ASAP7_75t_L g3766 ( 
.A(n_3677),
.B(n_3592),
.Y(n_3766)
);

BUFx3_ASAP7_75t_L g3767 ( 
.A(n_3714),
.Y(n_3767)
);

XOR2x2_ASAP7_75t_L g3768 ( 
.A(n_3699),
.B(n_3197),
.Y(n_3768)
);

INVx1_ASAP7_75t_L g3769 ( 
.A(n_3697),
.Y(n_3769)
);

OAI33xp33_ASAP7_75t_L g3770 ( 
.A1(n_3685),
.A2(n_3663),
.A3(n_3675),
.B1(n_3702),
.B2(n_3395),
.B3(n_3709),
.Y(n_3770)
);

INVx1_ASAP7_75t_L g3771 ( 
.A(n_3715),
.Y(n_3771)
);

AND2x2_ASAP7_75t_L g3772 ( 
.A(n_3677),
.B(n_3603),
.Y(n_3772)
);

INVx1_ASAP7_75t_L g3773 ( 
.A(n_3658),
.Y(n_3773)
);

OR2x2_ASAP7_75t_L g3774 ( 
.A(n_3719),
.B(n_3594),
.Y(n_3774)
);

AND2x2_ASAP7_75t_L g3775 ( 
.A(n_3678),
.B(n_3618),
.Y(n_3775)
);

INVx1_ASAP7_75t_SL g3776 ( 
.A(n_3659),
.Y(n_3776)
);

OA222x2_ASAP7_75t_L g3777 ( 
.A1(n_3667),
.A2(n_3453),
.B1(n_3413),
.B2(n_3544),
.C1(n_3478),
.C2(n_3491),
.Y(n_3777)
);

INVx1_ASAP7_75t_L g3778 ( 
.A(n_3721),
.Y(n_3778)
);

OR2x2_ASAP7_75t_L g3779 ( 
.A(n_3688),
.B(n_3654),
.Y(n_3779)
);

INVxp67_ASAP7_75t_SL g3780 ( 
.A(n_3661),
.Y(n_3780)
);

INVxp67_ASAP7_75t_L g3781 ( 
.A(n_3684),
.Y(n_3781)
);

OR2x2_ASAP7_75t_L g3782 ( 
.A(n_3654),
.B(n_3678),
.Y(n_3782)
);

INVx2_ASAP7_75t_L g3783 ( 
.A(n_3661),
.Y(n_3783)
);

NOR2xp33_ASAP7_75t_L g3784 ( 
.A(n_3710),
.B(n_3225),
.Y(n_3784)
);

HB1xp67_ASAP7_75t_L g3785 ( 
.A(n_3731),
.Y(n_3785)
);

AND2x2_ASAP7_75t_L g3786 ( 
.A(n_3723),
.B(n_3683),
.Y(n_3786)
);

INVx1_ASAP7_75t_L g3787 ( 
.A(n_3764),
.Y(n_3787)
);

INVx1_ASAP7_75t_L g3788 ( 
.A(n_3756),
.Y(n_3788)
);

NAND2xp5_ASAP7_75t_L g3789 ( 
.A(n_3724),
.B(n_3722),
.Y(n_3789)
);

INVx1_ASAP7_75t_SL g3790 ( 
.A(n_3748),
.Y(n_3790)
);

INVxp67_ASAP7_75t_L g3791 ( 
.A(n_3736),
.Y(n_3791)
);

O2A1O1Ixp33_ASAP7_75t_L g3792 ( 
.A1(n_3770),
.A2(n_3442),
.B(n_3309),
.C(n_3526),
.Y(n_3792)
);

INVx1_ASAP7_75t_L g3793 ( 
.A(n_3738),
.Y(n_3793)
);

INVx1_ASAP7_75t_L g3794 ( 
.A(n_3733),
.Y(n_3794)
);

OAI22xp33_ASAP7_75t_L g3795 ( 
.A1(n_3743),
.A2(n_3564),
.B1(n_3718),
.B2(n_3683),
.Y(n_3795)
);

AOI21xp5_ASAP7_75t_SL g3796 ( 
.A1(n_3743),
.A2(n_3718),
.B(n_3636),
.Y(n_3796)
);

AOI22xp5_ASAP7_75t_L g3797 ( 
.A1(n_3732),
.A2(n_3718),
.B1(n_3722),
.B2(n_3370),
.Y(n_3797)
);

OAI22xp33_ASAP7_75t_L g3798 ( 
.A1(n_3754),
.A2(n_3564),
.B1(n_3150),
.B2(n_3533),
.Y(n_3798)
);

AOI21xp33_ASAP7_75t_SL g3799 ( 
.A1(n_3739),
.A2(n_3151),
.B(n_3542),
.Y(n_3799)
);

OAI31xp33_ASAP7_75t_L g3800 ( 
.A1(n_3723),
.A2(n_3647),
.A3(n_3433),
.B(n_3610),
.Y(n_3800)
);

OAI31xp33_ASAP7_75t_L g3801 ( 
.A1(n_3762),
.A2(n_3468),
.A3(n_3469),
.B(n_3445),
.Y(n_3801)
);

OAI22xp33_ASAP7_75t_L g3802 ( 
.A1(n_3754),
.A2(n_3610),
.B1(n_3625),
.B2(n_3567),
.Y(n_3802)
);

INVx2_ASAP7_75t_L g3803 ( 
.A(n_3779),
.Y(n_3803)
);

XOR2x2_ASAP7_75t_L g3804 ( 
.A(n_3741),
.B(n_3334),
.Y(n_3804)
);

OAI21xp5_ASAP7_75t_L g3805 ( 
.A1(n_3746),
.A2(n_3418),
.B(n_3446),
.Y(n_3805)
);

INVx2_ASAP7_75t_L g3806 ( 
.A(n_3782),
.Y(n_3806)
);

INVxp67_ASAP7_75t_L g3807 ( 
.A(n_3758),
.Y(n_3807)
);

XOR2x2_ASAP7_75t_L g3808 ( 
.A(n_3768),
.B(n_3399),
.Y(n_3808)
);

NAND3xp33_ASAP7_75t_L g3809 ( 
.A(n_3749),
.B(n_3542),
.C(n_3126),
.Y(n_3809)
);

AOI22xp5_ASAP7_75t_L g3810 ( 
.A1(n_3735),
.A2(n_3609),
.B1(n_3711),
.B2(n_3317),
.Y(n_3810)
);

INVx1_ASAP7_75t_L g3811 ( 
.A(n_3737),
.Y(n_3811)
);

INVxp67_ASAP7_75t_L g3812 ( 
.A(n_3784),
.Y(n_3812)
);

AOI21xp33_ASAP7_75t_L g3813 ( 
.A1(n_3734),
.A2(n_3154),
.B(n_3562),
.Y(n_3813)
);

INVx1_ASAP7_75t_L g3814 ( 
.A(n_3740),
.Y(n_3814)
);

AOI22xp5_ASAP7_75t_L g3815 ( 
.A1(n_3727),
.A2(n_3606),
.B1(n_3468),
.B2(n_3706),
.Y(n_3815)
);

INVx1_ASAP7_75t_SL g3816 ( 
.A(n_3767),
.Y(n_3816)
);

XOR2xp5_ASAP7_75t_L g3817 ( 
.A(n_3747),
.B(n_3124),
.Y(n_3817)
);

INVx1_ASAP7_75t_L g3818 ( 
.A(n_3750),
.Y(n_3818)
);

INVx1_ASAP7_75t_L g3819 ( 
.A(n_3752),
.Y(n_3819)
);

AOI21xp5_ASAP7_75t_L g3820 ( 
.A1(n_3742),
.A2(n_3586),
.B(n_3565),
.Y(n_3820)
);

A2O1A1Ixp33_ASAP7_75t_L g3821 ( 
.A1(n_3747),
.A2(n_3522),
.B(n_3489),
.C(n_3565),
.Y(n_3821)
);

XOR2x2_ASAP7_75t_L g3822 ( 
.A(n_3776),
.B(n_3260),
.Y(n_3822)
);

NAND4xp25_ASAP7_75t_SL g3823 ( 
.A(n_3777),
.B(n_3667),
.C(n_3532),
.D(n_3676),
.Y(n_3823)
);

INVx1_ASAP7_75t_L g3824 ( 
.A(n_3753),
.Y(n_3824)
);

INVx1_ASAP7_75t_SL g3825 ( 
.A(n_3790),
.Y(n_3825)
);

O2A1O1Ixp33_ASAP7_75t_L g3826 ( 
.A1(n_3807),
.A2(n_3526),
.B(n_3190),
.C(n_3745),
.Y(n_3826)
);

NAND3xp33_ASAP7_75t_L g3827 ( 
.A(n_3805),
.B(n_3745),
.C(n_3726),
.Y(n_3827)
);

NAND2xp5_ASAP7_75t_L g3828 ( 
.A(n_3815),
.B(n_3781),
.Y(n_3828)
);

OAI31xp33_ASAP7_75t_L g3829 ( 
.A1(n_3809),
.A2(n_3548),
.A3(n_3456),
.B(n_3416),
.Y(n_3829)
);

AOI21xp5_ASAP7_75t_L g3830 ( 
.A1(n_3796),
.A2(n_3761),
.B(n_3780),
.Y(n_3830)
);

AOI222xp33_ASAP7_75t_L g3831 ( 
.A1(n_3809),
.A2(n_3726),
.B1(n_3596),
.B2(n_3361),
.C1(n_3321),
.C2(n_3335),
.Y(n_3831)
);

INVx1_ASAP7_75t_SL g3832 ( 
.A(n_3816),
.Y(n_3832)
);

HB1xp67_ASAP7_75t_L g3833 ( 
.A(n_3785),
.Y(n_3833)
);

INVx1_ASAP7_75t_L g3834 ( 
.A(n_3793),
.Y(n_3834)
);

INVx1_ASAP7_75t_L g3835 ( 
.A(n_3787),
.Y(n_3835)
);

AOI322xp5_ASAP7_75t_L g3836 ( 
.A1(n_3791),
.A2(n_3744),
.A3(n_3763),
.B1(n_3772),
.B2(n_3775),
.C1(n_3766),
.C2(n_3765),
.Y(n_3836)
);

NAND2xp5_ASAP7_75t_L g3837 ( 
.A(n_3788),
.B(n_3728),
.Y(n_3837)
);

NAND2xp5_ASAP7_75t_L g3838 ( 
.A(n_3794),
.B(n_3730),
.Y(n_3838)
);

OR2x2_ASAP7_75t_L g3839 ( 
.A(n_3789),
.B(n_3729),
.Y(n_3839)
);

INVx1_ASAP7_75t_L g3840 ( 
.A(n_3818),
.Y(n_3840)
);

NAND2xp5_ASAP7_75t_L g3841 ( 
.A(n_3797),
.B(n_3792),
.Y(n_3841)
);

OAI21xp33_ASAP7_75t_L g3842 ( 
.A1(n_3823),
.A2(n_3820),
.B(n_3799),
.Y(n_3842)
);

AOI21xp33_ASAP7_75t_L g3843 ( 
.A1(n_3801),
.A2(n_3562),
.B(n_3755),
.Y(n_3843)
);

OAI221xp5_ASAP7_75t_L g3844 ( 
.A1(n_3800),
.A2(n_3761),
.B1(n_3418),
.B2(n_3771),
.C(n_3769),
.Y(n_3844)
);

INVx1_ASAP7_75t_L g3845 ( 
.A(n_3819),
.Y(n_3845)
);

INVx1_ASAP7_75t_L g3846 ( 
.A(n_3824),
.Y(n_3846)
);

INVx2_ASAP7_75t_L g3847 ( 
.A(n_3803),
.Y(n_3847)
);

AND2x2_ASAP7_75t_L g3848 ( 
.A(n_3786),
.B(n_3712),
.Y(n_3848)
);

BUFx2_ASAP7_75t_L g3849 ( 
.A(n_3821),
.Y(n_3849)
);

OAI22xp33_ASAP7_75t_L g3850 ( 
.A1(n_3795),
.A2(n_3774),
.B1(n_3725),
.B2(n_3487),
.Y(n_3850)
);

OAI22xp33_ASAP7_75t_L g3851 ( 
.A1(n_3798),
.A2(n_3487),
.B1(n_3504),
.B2(n_3491),
.Y(n_3851)
);

INVx1_ASAP7_75t_L g3852 ( 
.A(n_3811),
.Y(n_3852)
);

AND2x2_ASAP7_75t_L g3853 ( 
.A(n_3800),
.B(n_3676),
.Y(n_3853)
);

INVx1_ASAP7_75t_L g3854 ( 
.A(n_3814),
.Y(n_3854)
);

OR2x2_ASAP7_75t_L g3855 ( 
.A(n_3806),
.B(n_3751),
.Y(n_3855)
);

INVx2_ASAP7_75t_L g3856 ( 
.A(n_3822),
.Y(n_3856)
);

NAND2xp5_ASAP7_75t_SL g3857 ( 
.A(n_3802),
.B(n_3586),
.Y(n_3857)
);

NAND2xp5_ASAP7_75t_L g3858 ( 
.A(n_3810),
.B(n_3778),
.Y(n_3858)
);

AND2x2_ASAP7_75t_L g3859 ( 
.A(n_3812),
.B(n_3701),
.Y(n_3859)
);

INVx1_ASAP7_75t_L g3860 ( 
.A(n_3817),
.Y(n_3860)
);

AOI21xp33_ASAP7_75t_L g3861 ( 
.A1(n_3813),
.A2(n_3374),
.B(n_3613),
.Y(n_3861)
);

INVx1_ASAP7_75t_L g3862 ( 
.A(n_3808),
.Y(n_3862)
);

NAND2xp5_ASAP7_75t_L g3863 ( 
.A(n_3804),
.B(n_3757),
.Y(n_3863)
);

AND2x2_ASAP7_75t_SL g3864 ( 
.A(n_3797),
.B(n_3187),
.Y(n_3864)
);

AOI222xp33_ASAP7_75t_L g3865 ( 
.A1(n_3809),
.A2(n_3596),
.B1(n_3414),
.B2(n_3648),
.C1(n_3651),
.C2(n_3757),
.Y(n_3865)
);

NAND2xp5_ASAP7_75t_L g3866 ( 
.A(n_3807),
.B(n_3773),
.Y(n_3866)
);

INVx1_ASAP7_75t_L g3867 ( 
.A(n_3833),
.Y(n_3867)
);

AOI221xp5_ASAP7_75t_L g3868 ( 
.A1(n_3841),
.A2(n_3773),
.B1(n_3257),
.B2(n_3414),
.C(n_3240),
.Y(n_3868)
);

AOI221x1_ASAP7_75t_L g3869 ( 
.A1(n_3862),
.A2(n_3241),
.B1(n_3547),
.B2(n_3278),
.C(n_3379),
.Y(n_3869)
);

AOI221xp5_ASAP7_75t_L g3870 ( 
.A1(n_3842),
.A2(n_3783),
.B1(n_3760),
.B2(n_3759),
.C(n_3279),
.Y(n_3870)
);

NAND2xp5_ASAP7_75t_SL g3871 ( 
.A(n_3829),
.B(n_3135),
.Y(n_3871)
);

NAND2xp5_ASAP7_75t_L g3872 ( 
.A(n_3865),
.B(n_3691),
.Y(n_3872)
);

INVx1_ASAP7_75t_L g3873 ( 
.A(n_3832),
.Y(n_3873)
);

INVx1_ASAP7_75t_L g3874 ( 
.A(n_3832),
.Y(n_3874)
);

NOR2xp33_ASAP7_75t_L g3875 ( 
.A(n_3825),
.B(n_3212),
.Y(n_3875)
);

NAND2xp5_ASAP7_75t_SL g3876 ( 
.A(n_3829),
.B(n_3230),
.Y(n_3876)
);

OAI21xp33_ASAP7_75t_SL g3877 ( 
.A1(n_3836),
.A2(n_3501),
.B(n_3427),
.Y(n_3877)
);

INVx2_ASAP7_75t_L g3878 ( 
.A(n_3825),
.Y(n_3878)
);

INVx1_ASAP7_75t_L g3879 ( 
.A(n_3866),
.Y(n_3879)
);

OAI21xp5_ASAP7_75t_L g3880 ( 
.A1(n_3831),
.A2(n_3532),
.B(n_3170),
.Y(n_3880)
);

INVx1_ASAP7_75t_L g3881 ( 
.A(n_3837),
.Y(n_3881)
);

OAI21xp5_ASAP7_75t_L g3882 ( 
.A1(n_3831),
.A2(n_3292),
.B(n_3155),
.Y(n_3882)
);

NAND2xp5_ASAP7_75t_L g3883 ( 
.A(n_3835),
.B(n_3597),
.Y(n_3883)
);

NAND3xp33_ASAP7_75t_SL g3884 ( 
.A(n_3826),
.B(n_3166),
.C(n_3161),
.Y(n_3884)
);

NOR3x1_ASAP7_75t_L g3885 ( 
.A(n_3849),
.B(n_3844),
.C(n_3827),
.Y(n_3885)
);

AOI221xp5_ASAP7_75t_L g3886 ( 
.A1(n_3850),
.A2(n_3520),
.B1(n_3547),
.B2(n_3427),
.C(n_3627),
.Y(n_3886)
);

NAND2xp5_ASAP7_75t_L g3887 ( 
.A(n_3834),
.B(n_3708),
.Y(n_3887)
);

AND2x2_ASAP7_75t_L g3888 ( 
.A(n_3856),
.B(n_3620),
.Y(n_3888)
);

NOR2x1_ASAP7_75t_SL g3889 ( 
.A(n_3857),
.B(n_3260),
.Y(n_3889)
);

NAND2xp5_ASAP7_75t_L g3890 ( 
.A(n_3863),
.B(n_3708),
.Y(n_3890)
);

INVx2_ASAP7_75t_SL g3891 ( 
.A(n_3860),
.Y(n_3891)
);

NOR2xp33_ASAP7_75t_L g3892 ( 
.A(n_3828),
.B(n_3504),
.Y(n_3892)
);

NAND2xp5_ASAP7_75t_L g3893 ( 
.A(n_3858),
.B(n_3713),
.Y(n_3893)
);

NOR3xp33_ASAP7_75t_L g3894 ( 
.A(n_3851),
.B(n_3520),
.C(n_2947),
.Y(n_3894)
);

NAND2xp5_ASAP7_75t_L g3895 ( 
.A(n_3859),
.B(n_3713),
.Y(n_3895)
);

AOI21xp5_ASAP7_75t_L g3896 ( 
.A1(n_3876),
.A2(n_3864),
.B(n_3830),
.Y(n_3896)
);

OAI211xp5_ASAP7_75t_L g3897 ( 
.A1(n_3870),
.A2(n_3861),
.B(n_3843),
.C(n_3853),
.Y(n_3897)
);

AOI21xp5_ASAP7_75t_L g3898 ( 
.A1(n_3871),
.A2(n_3884),
.B(n_3880),
.Y(n_3898)
);

OA22x2_ASAP7_75t_L g3899 ( 
.A1(n_3880),
.A2(n_3847),
.B1(n_3838),
.B2(n_3845),
.Y(n_3899)
);

INVxp67_ASAP7_75t_L g3900 ( 
.A(n_3875),
.Y(n_3900)
);

INVx1_ASAP7_75t_L g3901 ( 
.A(n_3878),
.Y(n_3901)
);

OAI22xp5_ASAP7_75t_L g3902 ( 
.A1(n_3872),
.A2(n_3839),
.B1(n_3855),
.B2(n_3846),
.Y(n_3902)
);

NAND2xp5_ASAP7_75t_L g3903 ( 
.A(n_3873),
.B(n_3854),
.Y(n_3903)
);

OA22x2_ASAP7_75t_L g3904 ( 
.A1(n_3874),
.A2(n_3891),
.B1(n_3867),
.B2(n_3882),
.Y(n_3904)
);

NOR4xp25_ASAP7_75t_L g3905 ( 
.A(n_3877),
.B(n_3852),
.C(n_3840),
.D(n_3848),
.Y(n_3905)
);

NAND2xp5_ASAP7_75t_L g3906 ( 
.A(n_3881),
.B(n_3634),
.Y(n_3906)
);

OAI21xp5_ASAP7_75t_L g3907 ( 
.A1(n_3869),
.A2(n_3495),
.B(n_3331),
.Y(n_3907)
);

AOI22xp5_ASAP7_75t_L g3908 ( 
.A1(n_3868),
.A2(n_3544),
.B1(n_3495),
.B2(n_3545),
.Y(n_3908)
);

A2O1A1Ixp33_ASAP7_75t_L g3909 ( 
.A1(n_3882),
.A2(n_3429),
.B(n_3388),
.C(n_3358),
.Y(n_3909)
);

NOR3x1_ASAP7_75t_L g3910 ( 
.A(n_3879),
.B(n_3266),
.C(n_3582),
.Y(n_3910)
);

AND4x1_ASAP7_75t_L g3911 ( 
.A(n_3885),
.B(n_3429),
.C(n_3380),
.D(n_3311),
.Y(n_3911)
);

INVx1_ASAP7_75t_L g3912 ( 
.A(n_3890),
.Y(n_3912)
);

AOI22xp5_ASAP7_75t_L g3913 ( 
.A1(n_3894),
.A2(n_3627),
.B1(n_3331),
.B2(n_3404),
.Y(n_3913)
);

OAI211xp5_ASAP7_75t_SL g3914 ( 
.A1(n_3886),
.A2(n_3342),
.B(n_3404),
.C(n_3402),
.Y(n_3914)
);

NAND3xp33_ASAP7_75t_SL g3915 ( 
.A(n_3892),
.B(n_3367),
.C(n_3080),
.Y(n_3915)
);

NOR2x1_ASAP7_75t_L g3916 ( 
.A(n_3888),
.B(n_2757),
.Y(n_3916)
);

AO22x2_ASAP7_75t_L g3917 ( 
.A1(n_3893),
.A2(n_3402),
.B1(n_3553),
.B2(n_3552),
.Y(n_3917)
);

NAND4xp25_ASAP7_75t_SL g3918 ( 
.A(n_3898),
.B(n_3889),
.C(n_3895),
.D(n_3883),
.Y(n_3918)
);

NOR2x1_ASAP7_75t_L g3919 ( 
.A(n_3901),
.B(n_3887),
.Y(n_3919)
);

AOI221xp5_ASAP7_75t_L g3920 ( 
.A1(n_3905),
.A2(n_3444),
.B1(n_3449),
.B2(n_3438),
.C(n_3451),
.Y(n_3920)
);

OAI211xp5_ASAP7_75t_SL g3921 ( 
.A1(n_3896),
.A2(n_3582),
.B(n_3221),
.C(n_3294),
.Y(n_3921)
);

OAI322xp33_ASAP7_75t_L g3922 ( 
.A1(n_3904),
.A2(n_2833),
.A3(n_3432),
.B1(n_3435),
.B2(n_3412),
.C1(n_3417),
.C2(n_3422),
.Y(n_3922)
);

NOR2xp33_ASAP7_75t_R g3923 ( 
.A(n_3900),
.B(n_608),
.Y(n_3923)
);

HB1xp67_ASAP7_75t_L g3924 ( 
.A(n_3903),
.Y(n_3924)
);

OAI211xp5_ASAP7_75t_L g3925 ( 
.A1(n_3908),
.A2(n_3897),
.B(n_3909),
.C(n_3907),
.Y(n_3925)
);

OA22x2_ASAP7_75t_L g3926 ( 
.A1(n_3902),
.A2(n_3704),
.B1(n_3703),
.B2(n_3689),
.Y(n_3926)
);

AND2x2_ASAP7_75t_L g3927 ( 
.A(n_3912),
.B(n_3664),
.Y(n_3927)
);

OAI221xp5_ASAP7_75t_L g3928 ( 
.A1(n_3911),
.A2(n_3554),
.B1(n_3382),
.B2(n_3541),
.C(n_3518),
.Y(n_3928)
);

NAND2xp5_ASAP7_75t_SL g3929 ( 
.A(n_3899),
.B(n_3207),
.Y(n_3929)
);

NAND3xp33_ASAP7_75t_L g3930 ( 
.A(n_3913),
.B(n_3315),
.C(n_3299),
.Y(n_3930)
);

AOI221xp5_ASAP7_75t_L g3931 ( 
.A1(n_3915),
.A2(n_3914),
.B1(n_3917),
.B2(n_3906),
.C(n_3910),
.Y(n_3931)
);

AND3x1_ASAP7_75t_L g3932 ( 
.A(n_3916),
.B(n_3294),
.C(n_3277),
.Y(n_3932)
);

NAND4xp25_ASAP7_75t_L g3933 ( 
.A(n_3898),
.B(n_2890),
.C(n_3352),
.D(n_3462),
.Y(n_3933)
);

AOI321xp33_ASAP7_75t_L g3934 ( 
.A1(n_3905),
.A2(n_3541),
.A3(n_3459),
.B1(n_3462),
.B2(n_3463),
.C(n_3436),
.Y(n_3934)
);

INVxp67_ASAP7_75t_L g3935 ( 
.A(n_3901),
.Y(n_3935)
);

AND2x2_ASAP7_75t_L g3936 ( 
.A(n_3924),
.B(n_3664),
.Y(n_3936)
);

INVx1_ASAP7_75t_L g3937 ( 
.A(n_3919),
.Y(n_3937)
);

NOR2xp33_ASAP7_75t_L g3938 ( 
.A(n_3922),
.B(n_608),
.Y(n_3938)
);

OAI22xp33_ASAP7_75t_L g3939 ( 
.A1(n_3928),
.A2(n_3207),
.B1(n_3216),
.B2(n_3382),
.Y(n_3939)
);

AOI22xp5_ASAP7_75t_L g3940 ( 
.A1(n_3925),
.A2(n_2926),
.B1(n_3042),
.B2(n_3689),
.Y(n_3940)
);

INVx1_ASAP7_75t_L g3941 ( 
.A(n_3935),
.Y(n_3941)
);

INVxp67_ASAP7_75t_L g3942 ( 
.A(n_3929),
.Y(n_3942)
);

AOI22xp5_ASAP7_75t_L g3943 ( 
.A1(n_3918),
.A2(n_3704),
.B1(n_3703),
.B2(n_3679),
.Y(n_3943)
);

INVx1_ASAP7_75t_L g3944 ( 
.A(n_3927),
.Y(n_3944)
);

OR2x2_ASAP7_75t_L g3945 ( 
.A(n_3933),
.B(n_3679),
.Y(n_3945)
);

AND3x4_ASAP7_75t_L g3946 ( 
.A(n_3921),
.B(n_3511),
.C(n_3629),
.Y(n_3946)
);

AOI22xp5_ASAP7_75t_L g3947 ( 
.A1(n_3931),
.A2(n_3511),
.B1(n_2529),
.B2(n_2552),
.Y(n_3947)
);

NAND2x1_ASAP7_75t_L g3948 ( 
.A(n_3926),
.B(n_3207),
.Y(n_3948)
);

HB1xp67_ASAP7_75t_L g3949 ( 
.A(n_3941),
.Y(n_3949)
);

NAND2xp5_ASAP7_75t_SL g3950 ( 
.A(n_3942),
.B(n_3923),
.Y(n_3950)
);

NOR2x1_ASAP7_75t_L g3951 ( 
.A(n_3937),
.B(n_3930),
.Y(n_3951)
);

AOI211xp5_ASAP7_75t_L g3952 ( 
.A1(n_3938),
.A2(n_3920),
.B(n_3934),
.C(n_3932),
.Y(n_3952)
);

INVxp67_ASAP7_75t_SL g3953 ( 
.A(n_3947),
.Y(n_3953)
);

AND3x4_ASAP7_75t_L g3954 ( 
.A(n_3946),
.B(n_3318),
.C(n_3633),
.Y(n_3954)
);

INVx1_ASAP7_75t_L g3955 ( 
.A(n_3936),
.Y(n_3955)
);

OR2x2_ASAP7_75t_L g3956 ( 
.A(n_3944),
.B(n_609),
.Y(n_3956)
);

NAND2xp5_ASAP7_75t_SL g3957 ( 
.A(n_3939),
.B(n_3216),
.Y(n_3957)
);

AND2x4_ASAP7_75t_L g3958 ( 
.A(n_3945),
.B(n_3216),
.Y(n_3958)
);

AND3x1_ASAP7_75t_L g3959 ( 
.A(n_3940),
.B(n_3352),
.C(n_3032),
.Y(n_3959)
);

INVx1_ASAP7_75t_SL g3960 ( 
.A(n_3956),
.Y(n_3960)
);

HB1xp67_ASAP7_75t_L g3961 ( 
.A(n_3949),
.Y(n_3961)
);

NAND2xp33_ASAP7_75t_R g3962 ( 
.A(n_3955),
.B(n_610),
.Y(n_3962)
);

NAND2xp5_ASAP7_75t_L g3963 ( 
.A(n_3952),
.B(n_3943),
.Y(n_3963)
);

CKINVDCx5p33_ASAP7_75t_R g3964 ( 
.A(n_3950),
.Y(n_3964)
);

NAND3xp33_ASAP7_75t_L g3965 ( 
.A(n_3951),
.B(n_3948),
.C(n_610),
.Y(n_3965)
);

INVx1_ASAP7_75t_L g3966 ( 
.A(n_3958),
.Y(n_3966)
);

INVx1_ASAP7_75t_L g3967 ( 
.A(n_3961),
.Y(n_3967)
);

INVx1_ASAP7_75t_L g3968 ( 
.A(n_3963),
.Y(n_3968)
);

INVx1_ASAP7_75t_L g3969 ( 
.A(n_3966),
.Y(n_3969)
);

HB1xp67_ASAP7_75t_L g3970 ( 
.A(n_3969),
.Y(n_3970)
);

INVx1_ASAP7_75t_L g3971 ( 
.A(n_3967),
.Y(n_3971)
);

INVx1_ASAP7_75t_L g3972 ( 
.A(n_3970),
.Y(n_3972)
);

OAI22xp5_ASAP7_75t_SL g3973 ( 
.A1(n_3972),
.A2(n_3964),
.B1(n_3968),
.B2(n_3971),
.Y(n_3973)
);

NAND3xp33_ASAP7_75t_SL g3974 ( 
.A(n_3973),
.B(n_3960),
.C(n_3965),
.Y(n_3974)
);

AOI22xp33_ASAP7_75t_L g3975 ( 
.A1(n_3974),
.A2(n_3953),
.B1(n_3954),
.B2(n_3957),
.Y(n_3975)
);

NAND2xp5_ASAP7_75t_L g3976 ( 
.A(n_3975),
.B(n_3959),
.Y(n_3976)
);

AOI22xp5_ASAP7_75t_L g3977 ( 
.A1(n_3976),
.A2(n_3962),
.B1(n_2746),
.B2(n_2637),
.Y(n_3977)
);


endmodule