module fake_jpeg_30689_n_47 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_47);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_47;

wire n_21;
wire n_33;
wire n_45;
wire n_23;
wire n_27;
wire n_22;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_32;

INVx2_ASAP7_75t_SL g16 ( 
.A(n_4),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_SL g17 ( 
.A(n_0),
.B(n_11),
.Y(n_17)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_17),
.B(n_0),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_22),
.B(n_25),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_17),
.B(n_1),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_23),
.B(n_26),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g24 ( 
.A1(n_16),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_24),
.A2(n_19),
.B1(n_18),
.B2(n_20),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_16),
.B(n_2),
.Y(n_25)
);

INVx1_ASAP7_75t_SL g26 ( 
.A(n_16),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_18),
.B(n_21),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_27),
.B(n_20),
.Y(n_29)
);

BUFx2_ASAP7_75t_L g28 ( 
.A(n_24),
.Y(n_28)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_29),
.B(n_8),
.Y(n_38)
);

BUFx24_ASAP7_75t_SL g31 ( 
.A(n_22),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_31),
.B(n_3),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g35 ( 
.A1(n_33),
.A2(n_19),
.B1(n_20),
.B2(n_21),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_35),
.A2(n_36),
.B1(n_30),
.B2(n_14),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_28),
.A2(n_19),
.B1(n_12),
.B2(n_13),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_37),
.B(n_5),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_38),
.B(n_32),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_39),
.B(n_40),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_41),
.A2(n_42),
.B1(n_5),
.B2(n_6),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_34),
.B(n_35),
.C(n_36),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_44),
.A2(n_7),
.B1(n_42),
.B2(n_15),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_45),
.B(n_44),
.Y(n_46)
);

AOI21xp5_ASAP7_75t_L g47 ( 
.A1(n_46),
.A2(n_43),
.B(n_7),
.Y(n_47)
);


endmodule