module fake_jpeg_25253_n_411 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_411);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_411;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_3),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_3),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx6f_ASAP7_75t_SL g31 ( 
.A(n_9),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_14),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_10),
.Y(n_34)
);

CKINVDCx16_ASAP7_75t_R g35 ( 
.A(n_7),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_11),
.B(n_8),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_9),
.B(n_1),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_6),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

BUFx12_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_46),
.Y(n_90)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_47),
.Y(n_91)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_25),
.Y(n_48)
);

INVx1_ASAP7_75t_SL g134 ( 
.A(n_48),
.Y(n_134)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_49),
.B(n_53),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_50),
.Y(n_93)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_25),
.Y(n_51)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_51),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_30),
.Y(n_52)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_52),
.Y(n_97)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_25),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_30),
.Y(n_54)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_54),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_30),
.Y(n_55)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_55),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_41),
.B(n_15),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_56),
.B(n_59),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_25),
.Y(n_57)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_57),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_29),
.Y(n_58)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_58),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_38),
.B(n_15),
.Y(n_59)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_31),
.Y(n_60)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_60),
.Y(n_110)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_31),
.Y(n_61)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_61),
.Y(n_120)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_29),
.Y(n_62)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_62),
.Y(n_92)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_29),
.Y(n_63)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_63),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_64),
.Y(n_122)
);

INVx13_ASAP7_75t_L g65 ( 
.A(n_18),
.Y(n_65)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_65),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_38),
.B(n_8),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_66),
.B(n_69),
.Y(n_128)
);

INVx2_ASAP7_75t_SL g67 ( 
.A(n_27),
.Y(n_67)
);

INVx2_ASAP7_75t_SL g104 ( 
.A(n_67),
.Y(n_104)
);

INVx2_ASAP7_75t_SL g68 ( 
.A(n_27),
.Y(n_68)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_68),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_33),
.Y(n_69)
);

BUFx24_ASAP7_75t_L g70 ( 
.A(n_18),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_70),
.Y(n_88)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_28),
.Y(n_71)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_71),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_72),
.Y(n_130)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_37),
.Y(n_73)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_73),
.Y(n_98)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_40),
.Y(n_74)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_74),
.Y(n_111)
);

INVx3_ASAP7_75t_SL g75 ( 
.A(n_40),
.Y(n_75)
);

BUFx4f_ASAP7_75t_L g123 ( 
.A(n_75),
.Y(n_123)
);

INVx11_ASAP7_75t_L g76 ( 
.A(n_44),
.Y(n_76)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_76),
.Y(n_133)
);

AOI21xp33_ASAP7_75t_L g77 ( 
.A1(n_33),
.A2(n_13),
.B(n_12),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_77),
.B(n_35),
.C(n_26),
.Y(n_101)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_34),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_78),
.B(n_22),
.Y(n_117)
);

BUFx5_ASAP7_75t_L g79 ( 
.A(n_44),
.Y(n_79)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_79),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_34),
.Y(n_80)
);

OR2x2_ASAP7_75t_SL g96 ( 
.A(n_80),
.B(n_78),
.Y(n_96)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_19),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_81),
.Y(n_113)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_19),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_82),
.Y(n_118)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_19),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_83),
.Y(n_119)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_36),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_84),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_45),
.Y(n_85)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_85),
.Y(n_106)
);

INVx11_ASAP7_75t_L g86 ( 
.A(n_28),
.Y(n_86)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_86),
.Y(n_112)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_21),
.Y(n_87)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_87),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_96),
.B(n_126),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_87),
.A2(n_37),
.B1(n_16),
.B2(n_26),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_99),
.A2(n_127),
.B1(n_35),
.B2(n_32),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_101),
.B(n_117),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_75),
.A2(n_16),
.B1(n_23),
.B2(n_20),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_108),
.A2(n_22),
.B1(n_32),
.B2(n_65),
.Y(n_147)
);

BUFx16f_ASAP7_75t_L g116 ( 
.A(n_70),
.Y(n_116)
);

INVx5_ASAP7_75t_L g172 ( 
.A(n_116),
.Y(n_172)
);

INVx11_ASAP7_75t_L g121 ( 
.A(n_62),
.Y(n_121)
);

INVx8_ASAP7_75t_L g140 ( 
.A(n_121),
.Y(n_140)
);

INVx11_ASAP7_75t_L g125 ( 
.A(n_62),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_125),
.Y(n_161)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_81),
.Y(n_126)
);

OAI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_46),
.A2(n_20),
.B1(n_23),
.B2(n_43),
.Y(n_127)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_82),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_132),
.B(n_55),
.Y(n_145)
);

BUFx8_ASAP7_75t_L g135 ( 
.A(n_116),
.Y(n_135)
);

INVx11_ASAP7_75t_L g181 ( 
.A(n_135),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_108),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_136),
.B(n_143),
.Y(n_184)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_90),
.Y(n_138)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_138),
.Y(n_197)
);

CKINVDCx12_ASAP7_75t_R g139 ( 
.A(n_134),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_139),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_L g141 ( 
.A1(n_127),
.A2(n_83),
.B1(n_47),
.B2(n_84),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_141),
.A2(n_147),
.B1(n_148),
.B2(n_149),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_91),
.B(n_63),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_142),
.A2(n_165),
.B(n_120),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_128),
.B(n_49),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_109),
.A2(n_68),
.B1(n_67),
.B2(n_61),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_144),
.A2(n_150),
.B1(n_151),
.B2(n_166),
.Y(n_180)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_145),
.Y(n_200)
);

BUFx2_ASAP7_75t_L g146 ( 
.A(n_88),
.Y(n_146)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_146),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_115),
.A2(n_60),
.B1(n_51),
.B2(n_86),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_L g150 ( 
.A1(n_97),
.A2(n_76),
.B1(n_42),
.B2(n_39),
.Y(n_150)
);

OAI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_97),
.A2(n_42),
.B1(n_39),
.B2(n_43),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_117),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_152),
.B(n_156),
.Y(n_177)
);

BUFx2_ASAP7_75t_L g153 ( 
.A(n_88),
.Y(n_153)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_153),
.Y(n_182)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_121),
.Y(n_154)
);

INVx11_ASAP7_75t_L g196 ( 
.A(n_154),
.Y(n_196)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_131),
.Y(n_155)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_155),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_100),
.Y(n_156)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_94),
.Y(n_157)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_157),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_124),
.B(n_36),
.Y(n_158)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_158),
.Y(n_201)
);

BUFx2_ASAP7_75t_L g159 ( 
.A(n_131),
.Y(n_159)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_159),
.Y(n_186)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_105),
.Y(n_160)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_160),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_100),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_162),
.B(n_163),
.Y(n_178)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_110),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_98),
.B(n_36),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_164),
.B(n_167),
.Y(n_189)
);

NAND2xp33_ASAP7_75t_SL g165 ( 
.A(n_113),
.B(n_53),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_L g166 ( 
.A1(n_106),
.A2(n_42),
.B1(n_39),
.B2(n_43),
.Y(n_166)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_110),
.Y(n_167)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_102),
.Y(n_168)
);

BUFx3_ASAP7_75t_L g212 ( 
.A(n_168),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_113),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_169),
.B(n_171),
.Y(n_191)
);

BUFx12f_ASAP7_75t_L g170 ( 
.A(n_92),
.Y(n_170)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_170),
.Y(n_188)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_118),
.Y(n_171)
);

CKINVDCx12_ASAP7_75t_R g174 ( 
.A(n_129),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_174),
.B(n_175),
.Y(n_203)
);

INVx1_ASAP7_75t_SL g175 ( 
.A(n_123),
.Y(n_175)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_122),
.Y(n_176)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_176),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_162),
.B(n_118),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_183),
.B(n_194),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_136),
.A2(n_103),
.B1(n_130),
.B2(n_89),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_185),
.A2(n_195),
.B1(n_199),
.B2(n_206),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_187),
.A2(n_209),
.B(n_208),
.Y(n_220)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_159),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_192),
.B(n_205),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_173),
.B(n_119),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_144),
.A2(n_112),
.B1(n_133),
.B2(n_104),
.Y(n_195)
);

OAI22xp33_ASAP7_75t_L g199 ( 
.A1(n_165),
.A2(n_155),
.B1(n_167),
.B2(n_163),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_142),
.B(n_57),
.C(n_119),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_204),
.B(n_213),
.Y(n_231)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_140),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_142),
.A2(n_112),
.B1(n_104),
.B2(n_93),
.Y(n_206)
);

AOI22x1_ASAP7_75t_L g208 ( 
.A1(n_148),
.A2(n_123),
.B1(n_48),
.B2(n_58),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_208),
.A2(n_185),
.B1(n_180),
.B2(n_210),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_175),
.A2(n_149),
.B(n_2),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_137),
.A2(n_114),
.B1(n_111),
.B2(n_95),
.Y(n_210)
);

INVx1_ASAP7_75t_SL g225 ( 
.A(n_210),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_157),
.B(n_24),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_191),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_214),
.B(n_215),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_189),
.B(n_170),
.Y(n_215)
);

INVxp67_ASAP7_75t_SL g217 ( 
.A(n_181),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_217),
.B(n_229),
.Y(n_262)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_213),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_218),
.B(n_235),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_200),
.B(n_170),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_219),
.B(n_221),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_L g275 ( 
.A1(n_220),
.A2(n_226),
.B(n_202),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_183),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_194),
.B(n_11),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_222),
.B(n_233),
.Y(n_247)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_181),
.Y(n_223)
);

INVx4_ASAP7_75t_L g270 ( 
.A(n_223),
.Y(n_270)
);

OA21x2_ASAP7_75t_L g226 ( 
.A1(n_209),
.A2(n_168),
.B(n_63),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g227 ( 
.A(n_203),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_227),
.B(n_234),
.Y(n_274)
);

INVx6_ASAP7_75t_L g229 ( 
.A(n_188),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_208),
.A2(n_140),
.B1(n_154),
.B2(n_172),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_230),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_178),
.B(n_160),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_232),
.B(n_241),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_184),
.B(n_13),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_177),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_201),
.B(n_161),
.Y(n_235)
);

AND2x6_ASAP7_75t_L g236 ( 
.A(n_187),
.B(n_14),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_236),
.A2(n_237),
.B(n_244),
.Y(n_260)
);

INVx1_ASAP7_75t_SL g237 ( 
.A(n_212),
.Y(n_237)
);

CKINVDCx14_ASAP7_75t_R g238 ( 
.A(n_206),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_238),
.B(n_240),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_198),
.A2(n_107),
.B1(n_54),
.B2(n_52),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_239),
.A2(n_180),
.B1(n_186),
.B2(n_192),
.Y(n_256)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_195),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_204),
.B(n_21),
.Y(n_241)
);

OAI22xp33_ASAP7_75t_SL g264 ( 
.A1(n_242),
.A2(n_190),
.B1(n_202),
.B2(n_197),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_207),
.B(n_21),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_243),
.B(n_245),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_197),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_211),
.Y(n_245)
);

CKINVDCx12_ASAP7_75t_R g246 ( 
.A(n_193),
.Y(n_246)
);

CKINVDCx16_ASAP7_75t_R g248 ( 
.A(n_246),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_228),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_249),
.B(n_254),
.Y(n_280)
);

INVx5_ASAP7_75t_L g250 ( 
.A(n_246),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_L g279 ( 
.A1(n_250),
.A2(n_264),
.B1(n_275),
.B2(n_225),
.Y(n_279)
);

O2A1O1Ixp33_ASAP7_75t_L g253 ( 
.A1(n_220),
.A2(n_221),
.B(n_240),
.C(n_226),
.Y(n_253)
);

OA22x2_ASAP7_75t_L g285 ( 
.A1(n_253),
.A2(n_271),
.B1(n_244),
.B2(n_239),
.Y(n_285)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_228),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_243),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_255),
.B(n_245),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_256),
.A2(n_257),
.B1(n_182),
.B2(n_179),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_224),
.A2(n_199),
.B1(n_190),
.B2(n_211),
.Y(n_257)
);

AND2x2_ASAP7_75t_SL g258 ( 
.A(n_218),
.B(n_226),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_258),
.B(n_71),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_SL g261 ( 
.A(n_224),
.B(n_193),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_261),
.B(n_234),
.Y(n_289)
);

BUFx3_ASAP7_75t_L g265 ( 
.A(n_229),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_265),
.B(n_223),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_222),
.B(n_205),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_268),
.B(n_269),
.Y(n_276)
);

OR2x2_ASAP7_75t_L g269 ( 
.A(n_242),
.B(n_212),
.Y(n_269)
);

AO22x1_ASAP7_75t_L g271 ( 
.A1(n_216),
.A2(n_188),
.B1(n_207),
.B2(n_186),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_231),
.B(n_241),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_272),
.B(n_231),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_277),
.B(n_281),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_272),
.B(n_216),
.C(n_225),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_278),
.B(n_289),
.C(n_282),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g317 ( 
.A1(n_279),
.A2(n_297),
.B1(n_258),
.B2(n_271),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_274),
.B(n_214),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_269),
.A2(n_253),
.B1(n_275),
.B2(n_266),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_282),
.A2(n_299),
.B1(n_258),
.B2(n_257),
.Y(n_309)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_267),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_283),
.B(n_288),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_267),
.B(n_232),
.Y(n_284)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_284),
.Y(n_313)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_285),
.Y(n_316)
);

OAI21xp33_ASAP7_75t_L g286 ( 
.A1(n_252),
.A2(n_233),
.B(n_236),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_286),
.A2(n_301),
.B(n_260),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_252),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_287),
.Y(n_302)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_262),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_289),
.B(n_260),
.Y(n_318)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_273),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_290),
.B(n_291),
.Y(n_311)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_273),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_251),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_292),
.B(n_295),
.Y(n_315)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_293),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_294),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_249),
.B(n_227),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_SL g296 ( 
.A(n_268),
.B(n_13),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_296),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_274),
.B(n_251),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g304 ( 
.A(n_298),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_269),
.A2(n_237),
.B1(n_179),
.B2(n_182),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_265),
.B(n_223),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_300),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_303),
.B(n_318),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_L g306 ( 
.A1(n_276),
.A2(n_253),
.B(n_259),
.Y(n_306)
);

CKINVDCx14_ASAP7_75t_R g337 ( 
.A(n_306),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_277),
.B(n_261),
.C(n_263),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_308),
.B(n_314),
.C(n_322),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_309),
.A2(n_297),
.B1(n_285),
.B2(n_284),
.Y(n_326)
);

AOI21xp33_ASAP7_75t_L g333 ( 
.A1(n_310),
.A2(n_321),
.B(n_306),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_SL g312 ( 
.A1(n_276),
.A2(n_258),
.B(n_266),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g331 ( 
.A(n_312),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_278),
.B(n_263),
.C(n_254),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_317),
.A2(n_285),
.B1(n_287),
.B2(n_280),
.Y(n_335)
);

AND2x4_ASAP7_75t_SL g319 ( 
.A(n_301),
.B(n_271),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_319),
.B(n_299),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_L g321 ( 
.A1(n_290),
.A2(n_255),
.B(n_248),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_283),
.B(n_256),
.C(n_248),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_326),
.A2(n_344),
.B1(n_337),
.B2(n_313),
.Y(n_359)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_327),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_303),
.B(n_291),
.C(n_292),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_329),
.B(n_332),
.C(n_338),
.Y(n_345)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_311),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_330),
.B(n_339),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_314),
.B(n_293),
.C(n_295),
.Y(n_332)
);

XNOR2x1_ASAP7_75t_L g358 ( 
.A(n_333),
.B(n_307),
.Y(n_358)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_335),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_316),
.A2(n_285),
.B1(n_280),
.B2(n_288),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_336),
.A2(n_341),
.B1(n_319),
.B2(n_324),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_318),
.B(n_281),
.C(n_285),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_315),
.Y(n_339)
);

BUFx6f_ASAP7_75t_L g340 ( 
.A(n_304),
.Y(n_340)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_340),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_316),
.A2(n_296),
.B1(n_270),
.B2(n_250),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_302),
.B(n_247),
.Y(n_342)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_342),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_308),
.B(n_270),
.C(n_247),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_343),
.B(n_322),
.C(n_321),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_309),
.A2(n_196),
.B1(n_172),
.B2(n_24),
.Y(n_344)
);

BUFx24_ASAP7_75t_SL g346 ( 
.A(n_334),
.Y(n_346)
);

NOR3xp33_ASAP7_75t_L g363 ( 
.A(n_346),
.B(n_343),
.C(n_328),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_348),
.A2(n_351),
.B1(n_196),
.B2(n_24),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_349),
.B(n_354),
.C(n_360),
.Y(n_366)
);

OAI21xp5_ASAP7_75t_SL g350 ( 
.A1(n_331),
.A2(n_310),
.B(n_304),
.Y(n_350)
);

OAI21xp5_ASAP7_75t_SL g369 ( 
.A1(n_350),
.A2(n_358),
.B(n_320),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_331),
.A2(n_319),
.B1(n_324),
.B2(n_313),
.Y(n_351)
);

XOR2xp5_ASAP7_75t_L g354 ( 
.A(n_334),
.B(n_312),
.Y(n_354)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_336),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_356),
.B(n_348),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_L g368 ( 
.A1(n_359),
.A2(n_341),
.B1(n_323),
.B2(n_305),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_329),
.B(n_323),
.C(n_325),
.Y(n_360)
);

INVx13_ASAP7_75t_L g361 ( 
.A(n_358),
.Y(n_361)
);

AOI22xp33_ASAP7_75t_SL g374 ( 
.A1(n_361),
.A2(n_364),
.B1(n_349),
.B2(n_354),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_352),
.A2(n_335),
.B1(n_338),
.B2(n_325),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_SL g377 ( 
.A1(n_362),
.A2(n_360),
.B1(n_14),
.B2(n_12),
.Y(n_377)
);

OAI21xp5_ASAP7_75t_SL g376 ( 
.A1(n_363),
.A2(n_355),
.B(n_357),
.Y(n_376)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_351),
.Y(n_364)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_365),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_345),
.B(n_328),
.C(n_332),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_367),
.B(n_370),
.C(n_64),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_368),
.A2(n_371),
.B1(n_373),
.B2(n_74),
.Y(n_380)
);

AOI21xp5_ASAP7_75t_L g379 ( 
.A1(n_369),
.A2(n_372),
.B(n_2),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_345),
.B(n_340),
.C(n_305),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_353),
.B(n_1),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_SL g373 ( 
.A1(n_347),
.A2(n_153),
.B1(n_146),
.B2(n_161),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_374),
.B(n_377),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_376),
.B(n_378),
.Y(n_385)
);

AOI21xp5_ASAP7_75t_SL g378 ( 
.A1(n_369),
.A2(n_9),
.B(n_4),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_SL g386 ( 
.A(n_379),
.B(n_384),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_380),
.B(n_381),
.C(n_382),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_370),
.B(n_85),
.C(n_72),
.Y(n_382)
);

OAI21xp5_ASAP7_75t_SL g383 ( 
.A1(n_362),
.A2(n_2),
.B(n_4),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_383),
.B(n_372),
.C(n_371),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g384 ( 
.A(n_366),
.B(n_79),
.Y(n_384)
);

INVx1_ASAP7_75t_SL g388 ( 
.A(n_378),
.Y(n_388)
);

AOI21xp5_ASAP7_75t_L g394 ( 
.A1(n_388),
.A2(n_392),
.B(n_375),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_L g399 ( 
.A1(n_390),
.A2(n_135),
.B1(n_71),
.B2(n_50),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_381),
.B(n_367),
.C(n_366),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_391),
.B(n_393),
.Y(n_395)
);

AND2x2_ASAP7_75t_L g392 ( 
.A(n_384),
.B(n_361),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_SL g393 ( 
.A(n_374),
.B(n_368),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_394),
.B(n_398),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_389),
.B(n_382),
.C(n_364),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_396),
.B(n_397),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_385),
.B(n_365),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_386),
.B(n_373),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_399),
.B(n_387),
.Y(n_402)
);

AOI21xp5_ASAP7_75t_L g405 ( 
.A1(n_402),
.A2(n_403),
.B(n_4),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_395),
.B(n_387),
.Y(n_403)
);

AOI21xp5_ASAP7_75t_SL g404 ( 
.A1(n_400),
.A2(n_396),
.B(n_135),
.Y(n_404)
);

OR2x2_ASAP7_75t_L g406 ( 
.A(n_404),
.B(n_405),
.Y(n_406)
);

AOI21xp5_ASAP7_75t_L g407 ( 
.A1(n_406),
.A2(n_400),
.B(n_401),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_407),
.Y(n_408)
);

AOI21xp5_ASAP7_75t_L g409 ( 
.A1(n_408),
.A2(n_5),
.B(n_6),
.Y(n_409)
);

AOI21xp5_ASAP7_75t_L g410 ( 
.A1(n_409),
.A2(n_5),
.B(n_7),
.Y(n_410)
);

AO21x1_ASAP7_75t_L g411 ( 
.A1(n_410),
.A2(n_5),
.B(n_70),
.Y(n_411)
);


endmodule