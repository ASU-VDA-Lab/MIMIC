module fake_jpeg_28985_n_410 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_410);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_410;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_1),
.B(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx16_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_3),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_14),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_5),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_0),
.B(n_8),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_7),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_11),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_16),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_2),
.Y(n_45)
);

BUFx12_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_7),
.Y(n_47)
);

BUFx2_ASAP7_75t_R g48 ( 
.A(n_14),
.Y(n_48)
);

BUFx16f_ASAP7_75t_L g49 ( 
.A(n_10),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_4),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_51),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_23),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_52),
.B(n_56),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_19),
.B(n_0),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_53),
.B(n_64),
.Y(n_111)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_32),
.Y(n_54)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_54),
.Y(n_113)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_55),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_23),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_23),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_57),
.B(n_68),
.Y(n_108)
);

INVx1_ASAP7_75t_SL g58 ( 
.A(n_48),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_58),
.B(n_59),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_19),
.B(n_17),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_27),
.Y(n_60)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_60),
.Y(n_100)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_61),
.Y(n_118)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_22),
.Y(n_62)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_62),
.Y(n_131)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_49),
.Y(n_63)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_63),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_40),
.B(n_0),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_27),
.Y(n_65)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_65),
.Y(n_142)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_28),
.Y(n_66)
);

INVx5_ASAP7_75t_L g145 ( 
.A(n_66),
.Y(n_145)
);

INVx2_ASAP7_75t_R g67 ( 
.A(n_48),
.Y(n_67)
);

OR2x2_ASAP7_75t_L g135 ( 
.A(n_67),
.B(n_86),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_39),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_33),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_69),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_33),
.Y(n_70)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_70),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_35),
.Y(n_71)
);

INVx6_ASAP7_75t_L g144 ( 
.A(n_71),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_39),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_72),
.B(n_73),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_40),
.B(n_10),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_22),
.Y(n_74)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_74),
.Y(n_148)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_35),
.Y(n_75)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_75),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_32),
.Y(n_76)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_76),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_35),
.Y(n_77)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_77),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_26),
.Y(n_78)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_78),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_18),
.B(n_17),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_79),
.B(n_85),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_26),
.Y(n_80)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_80),
.Y(n_112)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_39),
.Y(n_81)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_81),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_26),
.Y(n_82)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_82),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_38),
.Y(n_83)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_83),
.Y(n_143)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_29),
.Y(n_84)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_84),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_18),
.B(n_44),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_49),
.B(n_1),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_49),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_87),
.B(n_93),
.Y(n_147)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_38),
.Y(n_88)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_88),
.Y(n_122)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_34),
.Y(n_89)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_89),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_38),
.Y(n_90)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_90),
.Y(n_128)
);

BUFx16f_ASAP7_75t_L g91 ( 
.A(n_49),
.Y(n_91)
);

BUFx10_ASAP7_75t_L g140 ( 
.A(n_91),
.Y(n_140)
);

BUFx5_ASAP7_75t_L g92 ( 
.A(n_28),
.Y(n_92)
);

HB1xp67_ASAP7_75t_L g125 ( 
.A(n_92),
.Y(n_125)
);

INVx1_ASAP7_75t_SL g93 ( 
.A(n_45),
.Y(n_93)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_34),
.Y(n_94)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_94),
.Y(n_134)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_45),
.Y(n_95)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_95),
.Y(n_136)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_50),
.Y(n_96)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_96),
.Y(n_151)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_50),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_97),
.B(n_99),
.Y(n_123)
);

BUFx2_ASAP7_75t_L g98 ( 
.A(n_42),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_98),
.B(n_21),
.Y(n_101)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_42),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_101),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_71),
.A2(n_29),
.B1(n_37),
.B2(n_28),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_110),
.A2(n_119),
.B1(n_137),
.B2(n_141),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_53),
.B(n_47),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_114),
.B(n_129),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_51),
.A2(n_47),
.B1(n_44),
.B2(n_41),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_67),
.A2(n_37),
.B1(n_29),
.B2(n_28),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_120),
.A2(n_121),
.B1(n_146),
.B2(n_150),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_58),
.A2(n_37),
.B1(n_29),
.B2(n_30),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_64),
.B(n_30),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_124),
.B(n_126),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_62),
.B(n_41),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_97),
.B(n_20),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_86),
.A2(n_20),
.B1(n_36),
.B2(n_31),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_93),
.B(n_36),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_138),
.B(n_84),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_77),
.A2(n_70),
.B1(n_69),
.B2(n_75),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_98),
.A2(n_37),
.B1(n_25),
.B2(n_31),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_99),
.A2(n_25),
.B1(n_21),
.B2(n_24),
.Y(n_150)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_100),
.Y(n_153)
);

INVx4_ASAP7_75t_L g220 ( 
.A(n_153),
.Y(n_220)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_131),
.Y(n_154)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_154),
.Y(n_197)
);

OAI32xp33_ASAP7_75t_L g156 ( 
.A1(n_111),
.A2(n_60),
.A3(n_96),
.B1(n_81),
.B2(n_86),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_156),
.B(n_176),
.Y(n_195)
);

BUFx3_ASAP7_75t_L g157 ( 
.A(n_145),
.Y(n_157)
);

BUFx3_ASAP7_75t_L g205 ( 
.A(n_157),
.Y(n_205)
);

BUFx3_ASAP7_75t_L g158 ( 
.A(n_145),
.Y(n_158)
);

INVx4_ASAP7_75t_L g224 ( 
.A(n_158),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_117),
.B(n_24),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_160),
.B(n_164),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_123),
.B(n_55),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_161),
.B(n_167),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_149),
.B(n_91),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_163),
.B(n_186),
.C(n_190),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_107),
.A2(n_94),
.B1(n_88),
.B2(n_76),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_165),
.A2(n_168),
.B1(n_187),
.B2(n_191),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_135),
.B(n_91),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_142),
.A2(n_54),
.B1(n_89),
.B2(n_90),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_135),
.B(n_83),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_169),
.B(n_173),
.Y(n_198)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_130),
.Y(n_170)
);

INVx8_ASAP7_75t_L g208 ( 
.A(n_170),
.Y(n_208)
);

BUFx3_ASAP7_75t_L g171 ( 
.A(n_133),
.Y(n_171)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_171),
.Y(n_218)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_151),
.Y(n_172)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_172),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_148),
.B(n_82),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_149),
.A2(n_24),
.B1(n_11),
.B2(n_12),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_174),
.Y(n_200)
);

INVx8_ASAP7_75t_L g175 ( 
.A(n_139),
.Y(n_175)
);

INVx8_ASAP7_75t_L g226 ( 
.A(n_175),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_116),
.B(n_24),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_102),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_177),
.B(n_182),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_118),
.B(n_80),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_178),
.B(n_184),
.Y(n_206)
);

INVx1_ASAP7_75t_SL g179 ( 
.A(n_103),
.Y(n_179)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_179),
.Y(n_204)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_152),
.Y(n_180)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_180),
.Y(n_210)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_136),
.Y(n_181)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_181),
.Y(n_213)
);

INVx5_ASAP7_75t_L g182 ( 
.A(n_133),
.Y(n_182)
);

INVx1_ASAP7_75t_SL g183 ( 
.A(n_103),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g214 ( 
.A(n_183),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_147),
.B(n_78),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_108),
.B(n_63),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_185),
.B(n_188),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_SL g186 ( 
.A(n_120),
.B(n_2),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_104),
.A2(n_122),
.B1(n_134),
.B2(n_128),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_150),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_109),
.B(n_92),
.C(n_66),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_104),
.A2(n_46),
.B1(n_9),
.B2(n_13),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_105),
.B(n_2),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_192),
.B(n_132),
.Y(n_217)
);

BUFx12f_ASAP7_75t_L g193 ( 
.A(n_140),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_193),
.B(n_46),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_159),
.A2(n_110),
.B1(n_146),
.B2(n_121),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_201),
.A2(n_202),
.B1(n_212),
.B2(n_219),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_188),
.A2(n_105),
.B1(n_127),
.B2(n_144),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_163),
.B(n_167),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_207),
.B(n_222),
.C(n_223),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_161),
.A2(n_127),
.B1(n_144),
.B2(n_132),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_164),
.B(n_130),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_216),
.B(n_217),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_173),
.A2(n_143),
.B1(n_106),
.B2(n_112),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_169),
.B(n_143),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_221),
.B(n_192),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_162),
.B(n_125),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_162),
.B(n_139),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_225),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g227 ( 
.A(n_204),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g257 ( 
.A(n_227),
.Y(n_257)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_197),
.Y(n_229)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_229),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_211),
.A2(n_186),
.B(n_178),
.Y(n_230)
);

A2O1A1Ixp33_ASAP7_75t_L g259 ( 
.A1(n_230),
.A2(n_194),
.B(n_221),
.C(n_217),
.Y(n_259)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_197),
.Y(n_231)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_231),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_234),
.B(n_237),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_201),
.A2(n_190),
.B(n_184),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_235),
.A2(n_238),
.B(n_194),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_195),
.A2(n_189),
.B1(n_156),
.B2(n_166),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_236),
.A2(n_240),
.B1(n_245),
.B2(n_214),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_215),
.B(n_155),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_211),
.A2(n_154),
.B(n_183),
.Y(n_238)
);

BUFx2_ASAP7_75t_L g239 ( 
.A(n_226),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_239),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_206),
.A2(n_189),
.B1(n_166),
.B2(n_174),
.Y(n_240)
);

FAx1_ASAP7_75t_SL g241 ( 
.A(n_198),
.B(n_172),
.CI(n_153),
.CON(n_241),
.SN(n_241)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_241),
.B(n_251),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_215),
.B(n_177),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_242),
.B(n_246),
.Y(n_269)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_220),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_SL g270 ( 
.A1(n_243),
.A2(n_244),
.B1(n_247),
.B2(n_250),
.Y(n_270)
);

INVx8_ASAP7_75t_L g244 ( 
.A(n_226),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_206),
.A2(n_115),
.B1(n_112),
.B2(n_106),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_198),
.B(n_180),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_199),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_207),
.B(n_181),
.C(n_179),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_249),
.B(n_223),
.C(n_222),
.Y(n_255)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_199),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_196),
.B(n_170),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_212),
.A2(n_115),
.B1(n_175),
.B2(n_113),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_252),
.A2(n_209),
.B1(n_216),
.B2(n_214),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_253),
.A2(n_261),
.B1(n_236),
.B2(n_240),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_SL g294 ( 
.A(n_255),
.B(n_256),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_SL g276 ( 
.A1(n_259),
.A2(n_262),
.B(n_232),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_233),
.A2(n_203),
.B1(n_200),
.B2(n_219),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_261),
.A2(n_230),
.B1(n_246),
.B2(n_249),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_235),
.A2(n_202),
.B(n_200),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_263),
.A2(n_267),
.B1(n_271),
.B2(n_252),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_251),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_264),
.B(n_265),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_239),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_248),
.B(n_213),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_266),
.B(n_268),
.Y(n_278)
);

AOI22xp33_ASAP7_75t_L g267 ( 
.A1(n_233),
.A2(n_226),
.B1(n_204),
.B2(n_213),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_SL g268 ( 
.A(n_248),
.B(n_230),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_L g271 ( 
.A1(n_252),
.A2(n_224),
.B1(n_218),
.B2(n_208),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_248),
.B(n_210),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_272),
.B(n_275),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_232),
.A2(n_210),
.B1(n_220),
.B2(n_113),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_276),
.B(n_268),
.Y(n_303)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_254),
.Y(n_277)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_277),
.Y(n_299)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_254),
.Y(n_279)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_279),
.Y(n_301)
);

AOI22xp33_ASAP7_75t_SL g280 ( 
.A1(n_264),
.A2(n_239),
.B1(n_244),
.B2(n_224),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_280),
.A2(n_297),
.B1(n_258),
.B2(n_265),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_281),
.A2(n_291),
.B1(n_295),
.B2(n_259),
.Y(n_316)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_273),
.Y(n_282)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_282),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_SL g283 ( 
.A(n_260),
.B(n_237),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g308 ( 
.A(n_283),
.B(n_296),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_269),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_284),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_285),
.A2(n_297),
.B1(n_288),
.B2(n_284),
.Y(n_317)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_273),
.Y(n_286)
);

INVx1_ASAP7_75t_SL g298 ( 
.A(n_286),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_269),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_287),
.B(n_290),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_270),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_260),
.B(n_241),
.Y(n_292)
);

CKINVDCx16_ASAP7_75t_R g305 ( 
.A(n_292),
.Y(n_305)
);

INVx1_ASAP7_75t_SL g293 ( 
.A(n_253),
.Y(n_293)
);

CKINVDCx16_ASAP7_75t_R g314 ( 
.A(n_293),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_263),
.A2(n_242),
.B1(n_241),
.B2(n_234),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_257),
.B(n_229),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_275),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_278),
.B(n_272),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_300),
.B(n_245),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_L g302 ( 
.A1(n_276),
.A2(n_290),
.B(n_293),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_SL g336 ( 
.A1(n_302),
.A2(n_315),
.B(n_271),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_SL g331 ( 
.A(n_303),
.B(n_277),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_L g304 ( 
.A1(n_293),
.A2(n_274),
.B(n_256),
.Y(n_304)
);

AND2x2_ASAP7_75t_L g337 ( 
.A(n_304),
.B(n_250),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_307),
.A2(n_317),
.B1(n_281),
.B2(n_295),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_SL g309 ( 
.A(n_283),
.B(n_228),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_309),
.B(n_241),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_285),
.A2(n_274),
.B1(n_262),
.B2(n_257),
.Y(n_312)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_312),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_294),
.B(n_268),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_313),
.B(n_319),
.Y(n_332)
);

AOI21xp5_ASAP7_75t_L g315 ( 
.A1(n_289),
.A2(n_238),
.B(n_266),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_L g327 ( 
.A1(n_316),
.A2(n_305),
.B1(n_304),
.B2(n_306),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_294),
.B(n_255),
.C(n_249),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_318),
.B(n_291),
.C(n_288),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_278),
.B(n_259),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_306),
.B(n_287),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_320),
.B(n_324),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_321),
.B(n_335),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_323),
.A2(n_325),
.B1(n_334),
.B2(n_322),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_308),
.B(n_292),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_314),
.A2(n_289),
.B1(n_296),
.B2(n_286),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_L g352 ( 
.A1(n_326),
.A2(n_310),
.B1(n_300),
.B2(n_244),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_327),
.B(n_329),
.Y(n_349)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_328),
.B(n_331),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_316),
.B(n_282),
.Y(n_329)
);

NAND2xp33_ASAP7_75t_R g330 ( 
.A(n_303),
.B(n_279),
.Y(n_330)
);

OAI21xp33_ASAP7_75t_L g340 ( 
.A1(n_330),
.A2(n_315),
.B(n_319),
.Y(n_340)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_298),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_333),
.B(n_334),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_311),
.B(n_231),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_318),
.B(n_227),
.C(n_247),
.Y(n_335)
);

AOI21xp5_ASAP7_75t_L g339 ( 
.A1(n_336),
.A2(n_337),
.B(n_302),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_311),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_SL g342 ( 
.A(n_338),
.B(n_298),
.Y(n_342)
);

O2A1O1Ixp33_ASAP7_75t_L g359 ( 
.A1(n_339),
.A2(n_345),
.B(n_328),
.C(n_332),
.Y(n_359)
);

XOR2xp5_ASAP7_75t_L g358 ( 
.A(n_340),
.B(n_344),
.Y(n_358)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_342),
.Y(n_356)
);

BUFx2_ASAP7_75t_L g343 ( 
.A(n_325),
.Y(n_343)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_343),
.Y(n_360)
);

AOI21xp5_ASAP7_75t_L g345 ( 
.A1(n_336),
.A2(n_317),
.B(n_313),
.Y(n_345)
);

OAI21xp5_ASAP7_75t_SL g347 ( 
.A1(n_337),
.A2(n_301),
.B(n_299),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_347),
.B(n_193),
.Y(n_364)
);

AO221x1_ASAP7_75t_L g348 ( 
.A1(n_320),
.A2(n_310),
.B1(n_301),
.B2(n_299),
.C(n_258),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_348),
.B(n_352),
.Y(n_361)
);

XOR2xp5_ASAP7_75t_L g353 ( 
.A(n_332),
.B(n_321),
.Y(n_353)
);

XOR2xp5_ASAP7_75t_L g366 ( 
.A(n_353),
.B(n_140),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_323),
.A2(n_218),
.B1(n_205),
.B2(n_243),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_354),
.B(n_335),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_L g355 ( 
.A1(n_337),
.A2(n_205),
.B1(n_208),
.B2(n_157),
.Y(n_355)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_355),
.Y(n_368)
);

NAND2x1_ASAP7_75t_L g357 ( 
.A(n_339),
.B(n_331),
.Y(n_357)
);

AND2x2_ASAP7_75t_L g377 ( 
.A(n_357),
.B(n_343),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_359),
.B(n_362),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_350),
.B(n_208),
.C(n_158),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_363),
.B(n_353),
.C(n_350),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_364),
.B(n_365),
.Y(n_375)
);

BUFx6f_ASAP7_75t_L g365 ( 
.A(n_346),
.Y(n_365)
);

XOR2xp5_ASAP7_75t_L g374 ( 
.A(n_366),
.B(n_341),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_342),
.B(n_351),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_367),
.B(n_369),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_349),
.B(n_15),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_370),
.B(n_371),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_362),
.B(n_344),
.C(n_341),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_368),
.A2(n_343),
.B1(n_354),
.B2(n_345),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_372),
.A2(n_361),
.B1(n_359),
.B2(n_358),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_366),
.B(n_363),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_SL g388 ( 
.A(n_373),
.B(n_376),
.Y(n_388)
);

XOR2xp5_ASAP7_75t_L g391 ( 
.A(n_374),
.B(n_377),
.Y(n_391)
);

AOI21xp5_ASAP7_75t_L g376 ( 
.A1(n_356),
.A2(n_348),
.B(n_347),
.Y(n_376)
);

AND2x2_ASAP7_75t_L g380 ( 
.A(n_365),
.B(n_367),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_380),
.B(n_358),
.Y(n_385)
);

NOR2xp67_ASAP7_75t_L g381 ( 
.A(n_357),
.B(n_15),
.Y(n_381)
);

AOI21x1_ASAP7_75t_L g387 ( 
.A1(n_381),
.A2(n_14),
.B(n_17),
.Y(n_387)
);

AOI21xp5_ASAP7_75t_SL g382 ( 
.A1(n_379),
.A2(n_360),
.B(n_361),
.Y(n_382)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_382),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_384),
.B(n_385),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_380),
.A2(n_369),
.B1(n_182),
.B2(n_171),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_386),
.B(n_387),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_378),
.B(n_13),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_389),
.B(n_390),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_SL g390 ( 
.A(n_378),
.B(n_375),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_382),
.B(n_375),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_393),
.B(n_397),
.Y(n_403)
);

OAI21xp5_ASAP7_75t_SL g394 ( 
.A1(n_383),
.A2(n_377),
.B(n_193),
.Y(n_394)
);

XOR2xp5_ASAP7_75t_L g399 ( 
.A(n_394),
.B(n_391),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_388),
.B(n_193),
.C(n_13),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_SL g405 ( 
.A(n_399),
.B(n_401),
.Y(n_405)
);

OAI21xp5_ASAP7_75t_SL g400 ( 
.A1(n_392),
.A2(n_391),
.B(n_140),
.Y(n_400)
);

AOI21xp5_ASAP7_75t_L g404 ( 
.A1(n_400),
.A2(n_402),
.B(n_395),
.Y(n_404)
);

BUFx24_ASAP7_75t_SL g401 ( 
.A(n_396),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_SL g402 ( 
.A1(n_393),
.A2(n_7),
.B1(n_4),
.B2(n_6),
.Y(n_402)
);

OAI21xp5_ASAP7_75t_L g407 ( 
.A1(n_404),
.A2(n_406),
.B(n_3),
.Y(n_407)
);

A2O1A1O1Ixp25_ASAP7_75t_L g406 ( 
.A1(n_403),
.A2(n_398),
.B(n_6),
.C(n_3),
.D(n_46),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_407),
.B(n_6),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_408),
.B(n_405),
.C(n_6),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_SL g410 ( 
.A(n_409),
.B(n_46),
.Y(n_410)
);


endmodule