module real_jpeg_24409_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_0),
.B(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_0),
.B(n_33),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_0),
.B(n_17),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_0),
.B(n_54),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_0),
.B(n_51),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_0),
.B(n_49),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_0),
.B(n_68),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_0),
.B(n_27),
.Y(n_274)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_1),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_2),
.Y(n_52)
);

INVx1_ASAP7_75t_SL g55 ( 
.A(n_3),
.Y(n_55)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_4),
.B(n_54),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_4),
.B(n_49),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

INVx8_ASAP7_75t_SL g28 ( 
.A(n_6),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_7),
.B(n_33),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_7),
.B(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_7),
.B(n_51),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_7),
.B(n_49),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_7),
.B(n_68),
.Y(n_121)
);

CKINVDCx14_ASAP7_75t_R g293 ( 
.A(n_7),
.Y(n_293)
);

CKINVDCx14_ASAP7_75t_R g60 ( 
.A(n_8),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_8),
.B(n_72),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_8),
.B(n_150),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_8),
.B(n_33),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_8),
.B(n_54),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_8),
.B(n_51),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_8),
.B(n_49),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_8),
.B(n_68),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_9),
.B(n_51),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_9),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_9),
.B(n_33),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_9),
.B(n_49),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_9),
.B(n_68),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_9),
.B(n_27),
.Y(n_228)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_10),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_11),
.B(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_11),
.B(n_49),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_11),
.B(n_68),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_11),
.B(n_27),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_11),
.B(n_37),
.Y(n_252)
);

CKINVDCx14_ASAP7_75t_R g291 ( 
.A(n_11),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_11),
.B(n_54),
.Y(n_317)
);

INVx13_ASAP7_75t_L g46 ( 
.A(n_12),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_13),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_13),
.B(n_68),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_13),
.B(n_27),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_13),
.B(n_45),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_13),
.B(n_17),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_13),
.B(n_33),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_13),
.B(n_54),
.Y(n_260)
);

CKINVDCx14_ASAP7_75t_R g25 ( 
.A(n_14),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_14),
.B(n_45),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_14),
.B(n_37),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_14),
.B(n_33),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_14),
.B(n_54),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_14),
.B(n_51),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_14),
.B(n_49),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_14),
.B(n_68),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_15),
.B(n_49),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_15),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_15),
.B(n_68),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_15),
.B(n_127),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_15),
.B(n_216),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_15),
.B(n_33),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_15),
.B(n_54),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_16),
.B(n_54),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_16),
.B(n_33),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_16),
.B(n_170),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_16),
.B(n_51),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_16),
.B(n_49),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_16),
.B(n_68),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_16),
.B(n_27),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_16),
.B(n_295),
.Y(n_294)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_17),
.Y(n_171)
);

INVx6_ASAP7_75t_L g217 ( 
.A(n_17),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_136),
.Y(n_18)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_114),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_79),
.C(n_97),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_21),
.B(n_347),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_56),
.C(n_73),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_SL g342 ( 
.A(n_22),
.B(n_343),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_41),
.C(n_47),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_23),
.B(n_328),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_29),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_24),
.B(n_30),
.C(n_39),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_26),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_26),
.B(n_60),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_26),
.B(n_62),
.Y(n_83)
);

CKINVDCx5p33_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_35),
.B1(n_39),
.B2(n_40),
.Y(n_29)
);

CKINVDCx14_ASAP7_75t_R g40 ( 
.A(n_30),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_SL g95 ( 
.A(n_30),
.B(n_86),
.C(n_96),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_30),
.A2(n_40),
.B1(n_85),
.B2(n_86),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_32),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_31),
.B(n_36),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_31),
.B(n_63),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_32),
.B(n_291),
.Y(n_290)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_35),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_35),
.A2(n_39),
.B1(n_42),
.B2(n_310),
.Y(n_309)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx5_ASAP7_75t_L g150 ( 
.A(n_38),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_39),
.B(n_42),
.C(n_43),
.Y(n_41)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_41),
.B(n_47),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_42),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_43),
.A2(n_44),
.B1(n_308),
.B2(n_309),
.Y(n_307)
);

CKINVDCx16_ASAP7_75t_R g43 ( 
.A(n_44),
.Y(n_43)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

INVx8_ASAP7_75t_L g127 ( 
.A(n_46),
.Y(n_127)
);

INVx6_ASAP7_75t_L g297 ( 
.A(n_46),
.Y(n_297)
);

BUFx24_ASAP7_75t_SL g353 ( 
.A(n_47),
.Y(n_353)
);

FAx1_ASAP7_75t_SL g47 ( 
.A(n_48),
.B(n_50),
.CI(n_53),
.CON(n_47),
.SN(n_47)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_48),
.B(n_50),
.C(n_53),
.Y(n_101)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_51),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx3_ASAP7_75t_SL g54 ( 
.A(n_55),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_55),
.B(n_166),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_56),
.B(n_73),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_67),
.C(n_71),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_57),
.A2(n_58),
.B1(n_333),
.B2(n_335),
.Y(n_332)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_61),
.C(n_64),
.Y(n_58)
);

FAx1_ASAP7_75t_SL g304 ( 
.A(n_59),
.B(n_61),
.CI(n_64),
.CON(n_304),
.SN(n_304)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_63),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_63),
.B(n_65),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_66),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_67),
.A2(n_75),
.B1(n_76),
.B2(n_77),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_67),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_67),
.B(n_76),
.C(n_78),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_67),
.A2(n_71),
.B1(n_77),
.B2(n_334),
.Y(n_333)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_71),
.Y(n_334)
);

INVx8_ASAP7_75t_L g257 ( 
.A(n_72),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_78),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_75),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_79),
.A2(n_80),
.B1(n_97),
.B2(n_348),
.Y(n_347)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_82),
.B1(n_89),
.B2(n_90),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_81),
.B(n_91),
.C(n_95),
.Y(n_116)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

XOR2xp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_84),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_SL g124 ( 
.A(n_83),
.B(n_86),
.C(n_87),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_86),
.B1(n_87),
.B2(n_88),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_86),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_87),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g128 ( 
.A1(n_87),
.A2(n_88),
.B1(n_129),
.B2(n_130),
.Y(n_128)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

XOR2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_95),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_93),
.C(n_94),
.Y(n_91)
);

FAx1_ASAP7_75t_SL g102 ( 
.A(n_92),
.B(n_93),
.CI(n_94),
.CON(n_102),
.SN(n_102)
);

XOR2xp5_ASAP7_75t_L g99 ( 
.A(n_96),
.B(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_97),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_103),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_98),
.B(n_104),
.C(n_107),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_101),
.C(n_102),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g340 ( 
.A(n_99),
.B(n_341),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_101),
.B(n_102),
.Y(n_341)
);

BUFx24_ASAP7_75t_SL g349 ( 
.A(n_102),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_104),
.A2(n_105),
.B1(n_106),
.B2(n_107),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_109),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_108),
.B(n_110),
.C(n_113),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_110),
.A2(n_111),
.B1(n_112),
.B2(n_113),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_111),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_112),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_115),
.A2(n_133),
.B1(n_134),
.B2(n_135),
.Y(n_114)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_115),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_SL g115 ( 
.A(n_116),
.B(n_117),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_123),
.Y(n_117)
);

CKINVDCx5p33_ASAP7_75t_R g118 ( 
.A(n_119),
.Y(n_118)
);

BUFx24_ASAP7_75t_SL g356 ( 
.A(n_119),
.Y(n_356)
);

FAx1_ASAP7_75t_SL g119 ( 
.A(n_120),
.B(n_121),
.CI(n_122),
.CON(n_119),
.SN(n_119)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_125),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_126),
.A2(n_128),
.B1(n_131),
.B2(n_132),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_126),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_128),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_133),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_345),
.C(n_346),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_337),
.C(n_338),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_322),
.C(n_323),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_299),
.C(n_300),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_263),
.C(n_264),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_232),
.C(n_233),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_210),
.C(n_211),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_192),
.C(n_193),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_172),
.C(n_173),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_158),
.C(n_163),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_147),
.A2(n_148),
.B1(n_154),
.B2(n_155),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_147),
.B(n_156),
.C(n_157),
.Y(n_172)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_149),
.A2(n_151),
.B1(n_152),
.B2(n_153),
.Y(n_148)
);

CKINVDCx14_ASAP7_75t_R g153 ( 
.A(n_149),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_151),
.B(n_153),
.Y(n_176)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_SL g155 ( 
.A(n_156),
.B(n_157),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_159),
.B(n_161),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_159),
.A2(n_160),
.B1(n_161),
.B2(n_162),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_160),
.Y(n_159)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_165),
.C(n_167),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_166),
.B(n_257),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_169),
.Y(n_167)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_171),
.B(n_293),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_183),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_175),
.A2(n_176),
.B1(n_177),
.B2(n_178),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_175),
.B(n_178),
.C(n_183),
.Y(n_192)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_179),
.A2(n_180),
.B1(n_181),
.B2(n_182),
.Y(n_178)
);

CKINVDCx14_ASAP7_75t_R g182 ( 
.A(n_179),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_180),
.B(n_182),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_181),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_185),
.B1(n_186),
.B2(n_191),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_184),
.Y(n_191)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_187),
.A2(n_188),
.B1(n_189),
.B2(n_190),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g190 ( 
.A(n_187),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_188),
.B(n_190),
.C(n_191),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_189),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_SL g193 ( 
.A(n_194),
.B(n_201),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_196),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_195),
.B(n_196),
.C(n_201),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_198),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_197),
.B(n_199),
.C(n_200),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_200),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_SL g201 ( 
.A(n_202),
.B(n_203),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_202),
.B(n_204),
.C(n_205),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_205),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_206),
.A2(n_207),
.B1(n_208),
.B2(n_209),
.Y(n_205)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_206),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_207),
.B(n_209),
.Y(n_230)
);

CKINVDCx14_ASAP7_75t_R g207 ( 
.A(n_208),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_226),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_212),
.B(n_227),
.C(n_231),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_SL g212 ( 
.A(n_213),
.B(n_222),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_221),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_214),
.B(n_221),
.C(n_222),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_215),
.A2(n_218),
.B1(n_219),
.B2(n_220),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_215),
.Y(n_220)
);

INVx5_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_218),
.B(n_220),
.Y(n_245)
);

CKINVDCx16_ASAP7_75t_R g218 ( 
.A(n_219),
.Y(n_218)
);

BUFx24_ASAP7_75t_SL g351 ( 
.A(n_222),
.Y(n_351)
);

FAx1_ASAP7_75t_SL g222 ( 
.A(n_223),
.B(n_224),
.CI(n_225),
.CON(n_222),
.SN(n_222)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_223),
.B(n_224),
.C(n_225),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_231),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_227),
.Y(n_249)
);

FAx1_ASAP7_75t_SL g227 ( 
.A(n_228),
.B(n_229),
.CI(n_230),
.CON(n_227),
.SN(n_227)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_248),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_235),
.A2(n_236),
.B1(n_237),
.B2(n_238),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_236),
.B(n_237),
.C(n_248),
.Y(n_263)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_SL g238 ( 
.A(n_239),
.B(n_243),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_239),
.B(n_244),
.C(n_247),
.Y(n_267)
);

BUFx24_ASAP7_75t_SL g350 ( 
.A(n_239),
.Y(n_350)
);

FAx1_ASAP7_75t_SL g239 ( 
.A(n_240),
.B(n_241),
.CI(n_242),
.CON(n_239),
.SN(n_239)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_240),
.B(n_241),
.C(n_242),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_244),
.A2(n_245),
.B1(n_246),
.B2(n_247),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

CKINVDCx16_ASAP7_75t_R g246 ( 
.A(n_247),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_SL g248 ( 
.A(n_249),
.B(n_250),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_249),
.B(n_255),
.C(n_261),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_251),
.A2(n_255),
.B1(n_261),
.B2(n_262),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_251),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_252),
.A2(n_253),
.B(n_254),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_252),
.B(n_253),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_254),
.B(n_287),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_254),
.B(n_287),
.C(n_288),
.Y(n_312)
);

CKINVDCx14_ASAP7_75t_R g262 ( 
.A(n_255),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_258),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_256),
.B(n_259),
.C(n_260),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_260),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_265),
.A2(n_266),
.B1(n_283),
.B2(n_298),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_265),
.B(n_284),
.C(n_285),
.Y(n_299)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_SL g266 ( 
.A(n_267),
.B(n_268),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_267),
.B(n_269),
.C(n_276),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_276),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_271),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_270),
.B(n_272),
.C(n_275),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_272),
.A2(n_273),
.B1(n_274),
.B2(n_275),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_273),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_274),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_282),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_278),
.A2(n_279),
.B1(n_280),
.B2(n_281),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_278),
.B(n_281),
.C(n_282),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_279),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_280),
.Y(n_281)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_283),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_SL g283 ( 
.A(n_284),
.B(n_285),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_288),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_SL g288 ( 
.A(n_289),
.B(n_294),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_292),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_290),
.B(n_292),
.C(n_294),
.Y(n_319)
);

INVx8_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx8_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_301),
.A2(n_302),
.B1(n_320),
.B2(n_321),
.Y(n_300)
);

CKINVDCx16_ASAP7_75t_R g320 ( 
.A(n_301),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_302),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_SL g302 ( 
.A(n_303),
.B(n_311),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_303),
.B(n_311),
.C(n_320),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_305),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_304),
.B(n_306),
.C(n_307),
.Y(n_330)
);

BUFx24_ASAP7_75t_SL g355 ( 
.A(n_304),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_307),
.Y(n_305)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_313),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_312),
.B(n_314),
.C(n_315),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_315),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_319),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_318),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_317),
.B(n_318),
.C(n_319),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_325),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_324),
.B(n_326),
.C(n_336),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_326),
.A2(n_327),
.B1(n_329),
.B2(n_336),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_329),
.Y(n_336)
);

BUFx24_ASAP7_75t_SL g352 ( 
.A(n_329),
.Y(n_352)
);

FAx1_ASAP7_75t_SL g329 ( 
.A(n_330),
.B(n_331),
.CI(n_332),
.CON(n_329),
.SN(n_329)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_330),
.B(n_331),
.C(n_332),
.Y(n_344)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_333),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_339),
.B(n_344),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_340),
.B(n_342),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_340),
.B(n_342),
.C(n_344),
.Y(n_345)
);


endmodule