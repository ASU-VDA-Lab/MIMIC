module fake_jpeg_13374_n_75 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_75);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_75;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_40;
wire n_73;
wire n_59;
wire n_71;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_65;
wire n_63;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_72;
wire n_44;
wire n_28;
wire n_38;
wire n_26;
wire n_36;
wire n_74;
wire n_62;
wire n_25;
wire n_31;
wire n_56;
wire n_67;
wire n_29;
wire n_37;
wire n_50;
wire n_43;
wire n_32;
wire n_70;
wire n_66;

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_22),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_13),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_20),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_23),
.B(n_12),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_29),
.B(n_0),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_33),
.B(n_34),
.Y(n_40)
);

CKINVDCx14_ASAP7_75t_R g34 ( 
.A(n_25),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_36),
.B(n_0),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_38),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_39),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_39),
.B(n_26),
.C(n_31),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_44),
.B(n_48),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_38),
.A2(n_27),
.B1(n_32),
.B2(n_10),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_46),
.A2(n_47),
.B1(n_11),
.B2(n_21),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_35),
.A2(n_32),
.B1(n_27),
.B2(n_37),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_46),
.A2(n_37),
.B1(n_2),
.B2(n_3),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_49),
.A2(n_41),
.B1(n_5),
.B2(n_6),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_50),
.B(n_56),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_52),
.B(n_55),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_44),
.B(n_1),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_53),
.B(n_54),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_43),
.B(n_3),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_L g55 ( 
.A1(n_43),
.A2(n_4),
.B(n_5),
.Y(n_55)
);

INVxp33_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_57),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_51),
.A2(n_41),
.B1(n_42),
.B2(n_57),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_58),
.A2(n_60),
.B1(n_64),
.B2(n_7),
.Y(n_67)
);

XNOR2xp5_ASAP7_75t_L g59 ( 
.A(n_56),
.B(n_42),
.Y(n_59)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_59),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_54),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_62),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_66)
);

AOI21xp5_ASAP7_75t_L g70 ( 
.A1(n_66),
.A2(n_67),
.B(n_69),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_61),
.A2(n_8),
.B1(n_9),
.B2(n_14),
.Y(n_69)
);

AOI21xp5_ASAP7_75t_L g71 ( 
.A1(n_70),
.A2(n_68),
.B(n_65),
.Y(n_71)
);

AOI21x1_ASAP7_75t_SL g72 ( 
.A1(n_71),
.A2(n_68),
.B(n_58),
.Y(n_72)
);

A2O1A1Ixp33_ASAP7_75t_SL g73 ( 
.A1(n_72),
.A2(n_66),
.B(n_59),
.C(n_63),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_73),
.A2(n_24),
.B1(n_17),
.B2(n_18),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_74),
.B(n_16),
.Y(n_75)
);


endmodule