module fake_netlist_5_1593_n_1673 (n_137, n_294, n_318, n_82, n_194, n_316, n_248, n_124, n_86, n_136, n_146, n_315, n_268, n_61, n_127, n_75, n_235, n_226, n_74, n_57, n_353, n_351, n_111, n_155, n_43, n_116, n_22, n_284, n_46, n_245, n_21, n_139, n_38, n_105, n_280, n_4, n_17, n_254, n_33, n_23, n_302, n_265, n_293, n_244, n_47, n_173, n_198, n_247, n_314, n_8, n_321, n_292, n_100, n_212, n_119, n_275, n_252, n_26, n_295, n_133, n_330, n_2, n_6, n_39, n_147, n_67, n_307, n_87, n_150, n_106, n_209, n_259, n_301, n_68, n_93, n_186, n_134, n_191, n_51, n_63, n_171, n_153, n_341, n_204, n_250, n_260, n_298, n_320, n_286, n_122, n_282, n_331, n_10, n_24, n_325, n_132, n_90, n_101, n_281, n_240, n_189, n_220, n_291, n_231, n_257, n_31, n_13, n_152, n_317, n_9, n_323, n_195, n_42, n_356, n_227, n_45, n_271, n_94, n_335, n_123, n_167, n_234, n_343, n_308, n_267, n_297, n_156, n_5, n_225, n_219, n_157, n_131, n_192, n_223, n_158, n_138, n_264, n_109, n_163, n_276, n_339, n_95, n_183, n_185, n_243, n_347, n_169, n_59, n_255, n_215, n_350, n_196, n_211, n_218, n_181, n_3, n_290, n_221, n_178, n_287, n_344, n_72, n_104, n_41, n_56, n_141, n_355, n_15, n_336, n_145, n_48, n_50, n_337, n_313, n_88, n_216, n_168, n_164, n_311, n_208, n_142, n_214, n_328, n_140, n_299, n_303, n_296, n_241, n_357, n_184, n_65, n_78, n_144, n_114, n_96, n_165, n_213, n_129, n_342, n_98, n_361, n_363, n_197, n_107, n_69, n_236, n_1, n_249, n_304, n_329, n_203, n_274, n_80, n_35, n_73, n_277, n_92, n_19, n_338, n_149, n_333, n_309, n_30, n_14, n_84, n_130, n_322, n_258, n_29, n_79, n_151, n_25, n_306, n_288, n_188, n_190, n_201, n_263, n_44, n_224, n_40, n_34, n_228, n_283, n_112, n_85, n_239, n_55, n_49, n_310, n_54, n_12, n_76, n_358, n_362, n_170, n_332, n_27, n_77, n_102, n_161, n_273, n_349, n_270, n_230, n_81, n_118, n_279, n_70, n_253, n_261, n_174, n_289, n_172, n_206, n_217, n_312, n_345, n_210, n_365, n_91, n_176, n_182, n_143, n_83, n_354, n_237, n_180, n_340, n_207, n_37, n_346, n_229, n_108, n_66, n_177, n_60, n_16, n_0, n_58, n_18, n_359, n_117, n_326, n_233, n_205, n_366, n_113, n_246, n_179, n_125, n_269, n_128, n_285, n_120, n_232, n_327, n_135, n_126, n_202, n_266, n_272, n_193, n_251, n_352, n_53, n_160, n_154, n_62, n_148, n_71, n_300, n_159, n_334, n_175, n_262, n_238, n_99, n_319, n_364, n_20, n_121, n_242, n_360, n_36, n_200, n_162, n_64, n_222, n_28, n_89, n_115, n_324, n_199, n_187, n_32, n_103, n_348, n_97, n_166, n_11, n_7, n_256, n_305, n_52, n_278, n_110, n_1673);

input n_137;
input n_294;
input n_318;
input n_82;
input n_194;
input n_316;
input n_248;
input n_124;
input n_86;
input n_136;
input n_146;
input n_315;
input n_268;
input n_61;
input n_127;
input n_75;
input n_235;
input n_226;
input n_74;
input n_57;
input n_353;
input n_351;
input n_111;
input n_155;
input n_43;
input n_116;
input n_22;
input n_284;
input n_46;
input n_245;
input n_21;
input n_139;
input n_38;
input n_105;
input n_280;
input n_4;
input n_17;
input n_254;
input n_33;
input n_23;
input n_302;
input n_265;
input n_293;
input n_244;
input n_47;
input n_173;
input n_198;
input n_247;
input n_314;
input n_8;
input n_321;
input n_292;
input n_100;
input n_212;
input n_119;
input n_275;
input n_252;
input n_26;
input n_295;
input n_133;
input n_330;
input n_2;
input n_6;
input n_39;
input n_147;
input n_67;
input n_307;
input n_87;
input n_150;
input n_106;
input n_209;
input n_259;
input n_301;
input n_68;
input n_93;
input n_186;
input n_134;
input n_191;
input n_51;
input n_63;
input n_171;
input n_153;
input n_341;
input n_204;
input n_250;
input n_260;
input n_298;
input n_320;
input n_286;
input n_122;
input n_282;
input n_331;
input n_10;
input n_24;
input n_325;
input n_132;
input n_90;
input n_101;
input n_281;
input n_240;
input n_189;
input n_220;
input n_291;
input n_231;
input n_257;
input n_31;
input n_13;
input n_152;
input n_317;
input n_9;
input n_323;
input n_195;
input n_42;
input n_356;
input n_227;
input n_45;
input n_271;
input n_94;
input n_335;
input n_123;
input n_167;
input n_234;
input n_343;
input n_308;
input n_267;
input n_297;
input n_156;
input n_5;
input n_225;
input n_219;
input n_157;
input n_131;
input n_192;
input n_223;
input n_158;
input n_138;
input n_264;
input n_109;
input n_163;
input n_276;
input n_339;
input n_95;
input n_183;
input n_185;
input n_243;
input n_347;
input n_169;
input n_59;
input n_255;
input n_215;
input n_350;
input n_196;
input n_211;
input n_218;
input n_181;
input n_3;
input n_290;
input n_221;
input n_178;
input n_287;
input n_344;
input n_72;
input n_104;
input n_41;
input n_56;
input n_141;
input n_355;
input n_15;
input n_336;
input n_145;
input n_48;
input n_50;
input n_337;
input n_313;
input n_88;
input n_216;
input n_168;
input n_164;
input n_311;
input n_208;
input n_142;
input n_214;
input n_328;
input n_140;
input n_299;
input n_303;
input n_296;
input n_241;
input n_357;
input n_184;
input n_65;
input n_78;
input n_144;
input n_114;
input n_96;
input n_165;
input n_213;
input n_129;
input n_342;
input n_98;
input n_361;
input n_363;
input n_197;
input n_107;
input n_69;
input n_236;
input n_1;
input n_249;
input n_304;
input n_329;
input n_203;
input n_274;
input n_80;
input n_35;
input n_73;
input n_277;
input n_92;
input n_19;
input n_338;
input n_149;
input n_333;
input n_309;
input n_30;
input n_14;
input n_84;
input n_130;
input n_322;
input n_258;
input n_29;
input n_79;
input n_151;
input n_25;
input n_306;
input n_288;
input n_188;
input n_190;
input n_201;
input n_263;
input n_44;
input n_224;
input n_40;
input n_34;
input n_228;
input n_283;
input n_112;
input n_85;
input n_239;
input n_55;
input n_49;
input n_310;
input n_54;
input n_12;
input n_76;
input n_358;
input n_362;
input n_170;
input n_332;
input n_27;
input n_77;
input n_102;
input n_161;
input n_273;
input n_349;
input n_270;
input n_230;
input n_81;
input n_118;
input n_279;
input n_70;
input n_253;
input n_261;
input n_174;
input n_289;
input n_172;
input n_206;
input n_217;
input n_312;
input n_345;
input n_210;
input n_365;
input n_91;
input n_176;
input n_182;
input n_143;
input n_83;
input n_354;
input n_237;
input n_180;
input n_340;
input n_207;
input n_37;
input n_346;
input n_229;
input n_108;
input n_66;
input n_177;
input n_60;
input n_16;
input n_0;
input n_58;
input n_18;
input n_359;
input n_117;
input n_326;
input n_233;
input n_205;
input n_366;
input n_113;
input n_246;
input n_179;
input n_125;
input n_269;
input n_128;
input n_285;
input n_120;
input n_232;
input n_327;
input n_135;
input n_126;
input n_202;
input n_266;
input n_272;
input n_193;
input n_251;
input n_352;
input n_53;
input n_160;
input n_154;
input n_62;
input n_148;
input n_71;
input n_300;
input n_159;
input n_334;
input n_175;
input n_262;
input n_238;
input n_99;
input n_319;
input n_364;
input n_20;
input n_121;
input n_242;
input n_360;
input n_36;
input n_200;
input n_162;
input n_64;
input n_222;
input n_28;
input n_89;
input n_115;
input n_324;
input n_199;
input n_187;
input n_32;
input n_103;
input n_348;
input n_97;
input n_166;
input n_11;
input n_7;
input n_256;
input n_305;
input n_52;
input n_278;
input n_110;

output n_1673;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1166;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1150;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_1494;
wire n_625;
wire n_854;
wire n_1462;
wire n_1580;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1607;
wire n_1563;
wire n_606;
wire n_877;
wire n_1118;
wire n_755;
wire n_947;
wire n_1285;
wire n_373;
wire n_1359;
wire n_530;
wire n_1107;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_929;
wire n_1124;
wire n_902;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1261;
wire n_938;
wire n_1098;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_519;
wire n_406;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_1236;
wire n_1633;
wire n_569;
wire n_920;
wire n_1289;
wire n_1517;
wire n_1669;
wire n_370;
wire n_976;
wire n_1449;
wire n_1566;
wire n_1078;
wire n_1670;
wire n_775;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_1598;
wire n_955;
wire n_1146;
wire n_882;
wire n_1036;
wire n_1097;
wire n_550;
wire n_696;
wire n_897;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_845;
wire n_663;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_1672;
wire n_675;
wire n_888;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1556;
wire n_1384;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_468;
wire n_464;
wire n_1582;
wire n_1069;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_989;
wire n_1039;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1581;
wire n_1463;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_1053;
wire n_1224;
wire n_1248;
wire n_1331;
wire n_953;
wire n_1014;
wire n_1241;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_944;
wire n_1623;
wire n_1565;
wire n_647;
wire n_407;
wire n_1072;
wire n_857;
wire n_832;
wire n_561;
wire n_1319;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_728;
wire n_1162;
wire n_1538;
wire n_1199;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1660;
wire n_887;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1662;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_935;
wire n_817;
wire n_1175;
wire n_1479;
wire n_759;
wire n_806;
wire n_1477;
wire n_1635;
wire n_1571;
wire n_1189;
wire n_1259;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_843;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_776;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1647;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1128;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_372;
wire n_677;
wire n_1333;
wire n_1121;
wire n_368;
wire n_604;
wire n_433;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_624;
wire n_1380;
wire n_1617;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_448;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1614;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1009;
wire n_1148;
wire n_750;
wire n_742;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_396;
wire n_1383;
wire n_1073;
wire n_662;
wire n_459;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_486;
wire n_1548;
wire n_614;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_743;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1568;
wire n_1006;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_512;
wire n_1591;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_1031;
wire n_609;
wire n_1041;
wire n_1265;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_572;
wire n_815;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_960;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_1252;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_950;
wire n_1553;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_389;
wire n_418;
wire n_912;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1288;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1363;
wire n_1301;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_992;
wire n_543;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_1643;
wire n_883;
wire n_470;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_894;
wire n_1636;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_1575;
wire n_833;
wire n_1646;
wire n_1307;
wire n_988;
wire n_814;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_1219;
wire n_1204;
wire n_1035;
wire n_783;
wire n_555;
wire n_1188;
wire n_661;
wire n_849;
wire n_681;
wire n_584;
wire n_1638;
wire n_430;
wire n_510;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_875;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1637;
wire n_1419;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_917;
wire n_601;
wire n_966;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_818;
wire n_861;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1440;
wire n_421;
wire n_1356;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_1109;
wire n_895;
wire n_1310;
wire n_427;
wire n_1543;
wire n_1399;
wire n_791;
wire n_732;
wire n_1533;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_1291;
wire n_1297;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_676;
wire n_653;
wire n_642;
wire n_1602;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_664;
wire n_503;
wire n_1372;
wire n_605;
wire n_1273;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_980;
wire n_698;
wire n_703;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1013;
wire n_1452;
wire n_718;
wire n_1120;
wire n_719;
wire n_443;
wire n_714;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_1564;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_518;
wire n_505;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_390;
wire n_1330;
wire n_481;
wire n_1554;
wire n_769;
wire n_1046;
wire n_934;
wire n_1618;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_961;
wire n_771;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_1411;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1344;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_432;
wire n_839;
wire n_1210;
wire n_1364;
wire n_1250;
wire n_369;
wire n_871;
wire n_685;
wire n_598;
wire n_608;
wire n_928;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1619;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_740;
wire n_384;
wire n_1404;
wire n_1315;
wire n_1061;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1255;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_844;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_465;
wire n_1321;
wire n_585;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1540;
wire n_437;
wire n_1642;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_712;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_666;
wire n_1433;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_1018;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_178),
.Y(n_367)
);

BUFx5_ASAP7_75t_L g368 ( 
.A(n_302),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_349),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_75),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_358),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_345),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_232),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_68),
.Y(n_374)
);

BUFx3_ASAP7_75t_L g375 ( 
.A(n_8),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_334),
.Y(n_376)
);

BUFx8_ASAP7_75t_SL g377 ( 
.A(n_129),
.Y(n_377)
);

INVx2_ASAP7_75t_SL g378 ( 
.A(n_266),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_131),
.Y(n_379)
);

CKINVDCx16_ASAP7_75t_R g380 ( 
.A(n_170),
.Y(n_380)
);

CKINVDCx16_ASAP7_75t_R g381 ( 
.A(n_114),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_143),
.Y(n_382)
);

BUFx10_ASAP7_75t_L g383 ( 
.A(n_247),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_32),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_268),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_364),
.Y(n_386)
);

BUFx3_ASAP7_75t_L g387 ( 
.A(n_304),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_50),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_324),
.Y(n_389)
);

BUFx2_ASAP7_75t_L g390 ( 
.A(n_46),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_322),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_205),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_79),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_238),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_233),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_299),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_111),
.Y(n_397)
);

HB1xp67_ASAP7_75t_L g398 ( 
.A(n_267),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_138),
.Y(n_399)
);

BUFx2_ASAP7_75t_L g400 ( 
.A(n_119),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_72),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_46),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_265),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_339),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_213),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_189),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_91),
.Y(n_407)
);

INVxp67_ASAP7_75t_L g408 ( 
.A(n_100),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_353),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_321),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_359),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_126),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_365),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_37),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_209),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_274),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_35),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_89),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_120),
.Y(n_419)
);

BUFx6f_ASAP7_75t_L g420 ( 
.A(n_354),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_229),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_18),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_71),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_43),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_332),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_137),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_201),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_328),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_180),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_179),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_307),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_235),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_296),
.Y(n_433)
);

BUFx2_ASAP7_75t_L g434 ( 
.A(n_47),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_20),
.Y(n_435)
);

BUFx10_ASAP7_75t_L g436 ( 
.A(n_35),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_133),
.Y(n_437)
);

BUFx3_ASAP7_75t_L g438 ( 
.A(n_156),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_363),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_224),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_331),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_330),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_206),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_336),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_31),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_169),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_161),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_74),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_195),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_168),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_153),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_277),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_182),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_59),
.Y(n_454)
);

BUFx3_ASAP7_75t_L g455 ( 
.A(n_65),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_306),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_264),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_40),
.Y(n_458)
);

NOR2xp67_ASAP7_75t_L g459 ( 
.A(n_211),
.B(n_340),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_262),
.Y(n_460)
);

NOR2xp67_ASAP7_75t_L g461 ( 
.A(n_37),
.B(n_38),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_269),
.Y(n_462)
);

HB1xp67_ASAP7_75t_L g463 ( 
.A(n_256),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_29),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_62),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_22),
.Y(n_466)
);

BUFx3_ASAP7_75t_L g467 ( 
.A(n_17),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_124),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_355),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_239),
.Y(n_470)
);

BUFx6f_ASAP7_75t_L g471 ( 
.A(n_30),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_176),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_226),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_313),
.Y(n_474)
);

CKINVDCx20_ASAP7_75t_R g475 ( 
.A(n_9),
.Y(n_475)
);

BUFx3_ASAP7_75t_L g476 ( 
.A(n_34),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_149),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_16),
.Y(n_478)
);

BUFx2_ASAP7_75t_L g479 ( 
.A(n_48),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_54),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_291),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_192),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_155),
.Y(n_483)
);

NOR2xp67_ASAP7_75t_L g484 ( 
.A(n_152),
.B(n_202),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_66),
.Y(n_485)
);

BUFx10_ASAP7_75t_L g486 ( 
.A(n_132),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_312),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_245),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_309),
.Y(n_489)
);

BUFx3_ASAP7_75t_L g490 ( 
.A(n_236),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_320),
.Y(n_491)
);

CKINVDCx20_ASAP7_75t_R g492 ( 
.A(n_341),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_188),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_343),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_284),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_150),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_94),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_12),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_301),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_80),
.Y(n_500)
);

BUFx10_ASAP7_75t_L g501 ( 
.A(n_151),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_69),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_342),
.Y(n_503)
);

HB1xp67_ASAP7_75t_L g504 ( 
.A(n_146),
.Y(n_504)
);

BUFx3_ASAP7_75t_L g505 ( 
.A(n_70),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_250),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_142),
.Y(n_507)
);

NOR2xp67_ASAP7_75t_L g508 ( 
.A(n_110),
.B(n_338),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_337),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_11),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_348),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_293),
.Y(n_512)
);

BUFx2_ASAP7_75t_L g513 ( 
.A(n_171),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_30),
.Y(n_514)
);

CKINVDCx20_ASAP7_75t_R g515 ( 
.A(n_7),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_145),
.Y(n_516)
);

INVx1_ASAP7_75t_SL g517 ( 
.A(n_207),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_3),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_15),
.Y(n_519)
);

INVx1_ASAP7_75t_SL g520 ( 
.A(n_162),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_198),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_57),
.Y(n_522)
);

CKINVDCx20_ASAP7_75t_R g523 ( 
.A(n_215),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_362),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_63),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_254),
.Y(n_526)
);

CKINVDCx14_ASAP7_75t_R g527 ( 
.A(n_159),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_272),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_298),
.Y(n_529)
);

BUFx2_ASAP7_75t_SL g530 ( 
.A(n_67),
.Y(n_530)
);

BUFx2_ASAP7_75t_L g531 ( 
.A(n_219),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_112),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_241),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_96),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_288),
.Y(n_535)
);

BUFx2_ASAP7_75t_L g536 ( 
.A(n_344),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_319),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_212),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_360),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_86),
.Y(n_540)
);

CKINVDCx20_ASAP7_75t_R g541 ( 
.A(n_109),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_276),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_286),
.Y(n_543)
);

CKINVDCx16_ASAP7_75t_R g544 ( 
.A(n_115),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_88),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_253),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_148),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_329),
.Y(n_548)
);

CKINVDCx16_ASAP7_75t_R g549 ( 
.A(n_134),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_18),
.Y(n_550)
);

CKINVDCx20_ASAP7_75t_R g551 ( 
.A(n_76),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_273),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_23),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_234),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_52),
.Y(n_555)
);

BUFx6f_ASAP7_75t_L g556 ( 
.A(n_107),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_290),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_130),
.Y(n_558)
);

BUFx3_ASAP7_75t_L g559 ( 
.A(n_90),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_9),
.Y(n_560)
);

BUFx3_ASAP7_75t_L g561 ( 
.A(n_333),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_102),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_186),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_15),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_103),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_221),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_228),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_83),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_318),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_208),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_135),
.Y(n_571)
);

BUFx3_ASAP7_75t_L g572 ( 
.A(n_242),
.Y(n_572)
);

CKINVDCx20_ASAP7_75t_R g573 ( 
.A(n_199),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_217),
.Y(n_574)
);

INVx2_ASAP7_75t_SL g575 ( 
.A(n_45),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_294),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_214),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_27),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_325),
.Y(n_579)
);

BUFx2_ASAP7_75t_L g580 ( 
.A(n_12),
.Y(n_580)
);

BUFx10_ASAP7_75t_L g581 ( 
.A(n_45),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_13),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_305),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_73),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_157),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_244),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_243),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_237),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_230),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_352),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_297),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_53),
.Y(n_592)
);

INVx2_ASAP7_75t_SL g593 ( 
.A(n_13),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_177),
.Y(n_594)
);

INVx1_ASAP7_75t_SL g595 ( 
.A(n_147),
.Y(n_595)
);

INVx1_ASAP7_75t_SL g596 ( 
.A(n_193),
.Y(n_596)
);

BUFx10_ASAP7_75t_L g597 ( 
.A(n_121),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_55),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_127),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_20),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_210),
.Y(n_601)
);

BUFx10_ASAP7_75t_L g602 ( 
.A(n_60),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_471),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_375),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_375),
.Y(n_605)
);

BUFx8_ASAP7_75t_SL g606 ( 
.A(n_390),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_471),
.Y(n_607)
);

AND2x4_ASAP7_75t_L g608 ( 
.A(n_387),
.B(n_0),
.Y(n_608)
);

HB1xp67_ASAP7_75t_L g609 ( 
.A(n_434),
.Y(n_609)
);

INVx3_ASAP7_75t_L g610 ( 
.A(n_471),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_467),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_398),
.B(n_0),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_471),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_467),
.Y(n_614)
);

BUFx6f_ASAP7_75t_L g615 ( 
.A(n_420),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_398),
.B(n_1),
.Y(n_616)
);

BUFx2_ASAP7_75t_L g617 ( 
.A(n_479),
.Y(n_617)
);

BUFx2_ASAP7_75t_L g618 ( 
.A(n_580),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_476),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_463),
.B(n_1),
.Y(n_620)
);

AND2x2_ASAP7_75t_L g621 ( 
.A(n_527),
.B(n_2),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_463),
.B(n_2),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_476),
.Y(n_623)
);

AOI22xp5_ASAP7_75t_L g624 ( 
.A1(n_527),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_624)
);

BUFx8_ASAP7_75t_SL g625 ( 
.A(n_377),
.Y(n_625)
);

HB1xp67_ASAP7_75t_L g626 ( 
.A(n_414),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_368),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_368),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_368),
.Y(n_629)
);

AND2x2_ASAP7_75t_L g630 ( 
.A(n_400),
.B(n_4),
.Y(n_630)
);

BUFx6f_ASAP7_75t_L g631 ( 
.A(n_420),
.Y(n_631)
);

INVx3_ASAP7_75t_L g632 ( 
.A(n_436),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_384),
.Y(n_633)
);

NOR2x1_ASAP7_75t_L g634 ( 
.A(n_387),
.B(n_49),
.Y(n_634)
);

INVx5_ASAP7_75t_L g635 ( 
.A(n_420),
.Y(n_635)
);

HB1xp67_ASAP7_75t_L g636 ( 
.A(n_417),
.Y(n_636)
);

INVx5_ASAP7_75t_L g637 ( 
.A(n_420),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_504),
.B(n_5),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_445),
.Y(n_639)
);

BUFx6f_ASAP7_75t_L g640 ( 
.A(n_556),
.Y(n_640)
);

BUFx12f_ASAP7_75t_L g641 ( 
.A(n_436),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_458),
.Y(n_642)
);

AOI22xp5_ASAP7_75t_L g643 ( 
.A1(n_380),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_368),
.Y(n_644)
);

BUFx6f_ASAP7_75t_L g645 ( 
.A(n_556),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_368),
.Y(n_646)
);

NOR2xp33_ASAP7_75t_L g647 ( 
.A(n_504),
.B(n_6),
.Y(n_647)
);

INVx3_ASAP7_75t_L g648 ( 
.A(n_581),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_464),
.Y(n_649)
);

OAI21x1_ASAP7_75t_L g650 ( 
.A1(n_373),
.A2(n_56),
.B(n_51),
.Y(n_650)
);

BUFx2_ASAP7_75t_L g651 ( 
.A(n_422),
.Y(n_651)
);

CKINVDCx20_ASAP7_75t_R g652 ( 
.A(n_370),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_519),
.Y(n_653)
);

INVx3_ASAP7_75t_L g654 ( 
.A(n_581),
.Y(n_654)
);

AND2x4_ASAP7_75t_L g655 ( 
.A(n_438),
.B(n_10),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_513),
.B(n_10),
.Y(n_656)
);

AND2x4_ASAP7_75t_L g657 ( 
.A(n_438),
.B(n_455),
.Y(n_657)
);

BUFx6f_ASAP7_75t_L g658 ( 
.A(n_556),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_550),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_560),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_368),
.Y(n_661)
);

HB1xp67_ASAP7_75t_L g662 ( 
.A(n_424),
.Y(n_662)
);

AOI22xp5_ASAP7_75t_L g663 ( 
.A1(n_381),
.A2(n_11),
.B1(n_14),
.B2(n_16),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_564),
.Y(n_664)
);

AND2x4_ASAP7_75t_L g665 ( 
.A(n_455),
.B(n_14),
.Y(n_665)
);

INVx4_ASAP7_75t_L g666 ( 
.A(n_556),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_600),
.Y(n_667)
);

BUFx3_ASAP7_75t_L g668 ( 
.A(n_383),
.Y(n_668)
);

INVx5_ASAP7_75t_L g669 ( 
.A(n_383),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_382),
.Y(n_670)
);

INVx2_ASAP7_75t_SL g671 ( 
.A(n_602),
.Y(n_671)
);

BUFx6f_ASAP7_75t_L g672 ( 
.A(n_490),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_490),
.Y(n_673)
);

BUFx12f_ASAP7_75t_L g674 ( 
.A(n_486),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_367),
.Y(n_675)
);

BUFx6f_ASAP7_75t_L g676 ( 
.A(n_505),
.Y(n_676)
);

HB1xp67_ASAP7_75t_L g677 ( 
.A(n_435),
.Y(n_677)
);

BUFx12f_ASAP7_75t_L g678 ( 
.A(n_486),
.Y(n_678)
);

AND2x4_ASAP7_75t_L g679 ( 
.A(n_505),
.B(n_17),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_559),
.Y(n_680)
);

INVx5_ASAP7_75t_L g681 ( 
.A(n_501),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_531),
.B(n_19),
.Y(n_682)
);

OA21x2_ASAP7_75t_L g683 ( 
.A1(n_382),
.A2(n_19),
.B(n_21),
.Y(n_683)
);

AND2x4_ASAP7_75t_L g684 ( 
.A(n_559),
.B(n_21),
.Y(n_684)
);

BUFx6f_ASAP7_75t_L g685 ( 
.A(n_561),
.Y(n_685)
);

BUFx6f_ASAP7_75t_L g686 ( 
.A(n_561),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_572),
.Y(n_687)
);

BUFx12f_ASAP7_75t_L g688 ( 
.A(n_501),
.Y(n_688)
);

BUFx6f_ASAP7_75t_L g689 ( 
.A(n_572),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_369),
.Y(n_690)
);

BUFx12f_ASAP7_75t_L g691 ( 
.A(n_597),
.Y(n_691)
);

BUFx2_ASAP7_75t_L g692 ( 
.A(n_466),
.Y(n_692)
);

BUFx2_ASAP7_75t_L g693 ( 
.A(n_478),
.Y(n_693)
);

INVx5_ASAP7_75t_L g694 ( 
.A(n_597),
.Y(n_694)
);

BUFx6f_ASAP7_75t_L g695 ( 
.A(n_591),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_374),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_371),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_372),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_376),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_536),
.B(n_22),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_591),
.Y(n_701)
);

BUFx2_ASAP7_75t_L g702 ( 
.A(n_498),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_386),
.Y(n_703)
);

AND2x4_ASAP7_75t_L g704 ( 
.A(n_378),
.B(n_23),
.Y(n_704)
);

OAI22xp5_ASAP7_75t_R g705 ( 
.A1(n_510),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_393),
.B(n_24),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_441),
.B(n_25),
.Y(n_707)
);

OAI21x1_ASAP7_75t_L g708 ( 
.A1(n_488),
.A2(n_61),
.B(n_58),
.Y(n_708)
);

BUFx6f_ASAP7_75t_L g709 ( 
.A(n_552),
.Y(n_709)
);

INVx3_ASAP7_75t_L g710 ( 
.A(n_602),
.Y(n_710)
);

BUFx6f_ASAP7_75t_L g711 ( 
.A(n_565),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_587),
.B(n_26),
.Y(n_712)
);

BUFx6f_ASAP7_75t_L g713 ( 
.A(n_395),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_401),
.Y(n_714)
);

BUFx2_ASAP7_75t_L g715 ( 
.A(n_514),
.Y(n_715)
);

NOR2xp33_ASAP7_75t_L g716 ( 
.A(n_408),
.B(n_27),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_544),
.B(n_28),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_403),
.Y(n_718)
);

BUFx12f_ASAP7_75t_L g719 ( 
.A(n_518),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_379),
.Y(n_720)
);

BUFx2_ASAP7_75t_L g721 ( 
.A(n_553),
.Y(n_721)
);

BUFx12f_ASAP7_75t_L g722 ( 
.A(n_578),
.Y(n_722)
);

HB1xp67_ASAP7_75t_L g723 ( 
.A(n_582),
.Y(n_723)
);

INVx3_ASAP7_75t_L g724 ( 
.A(n_575),
.Y(n_724)
);

INVx3_ASAP7_75t_L g725 ( 
.A(n_593),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_405),
.Y(n_726)
);

BUFx2_ASAP7_75t_L g727 ( 
.A(n_402),
.Y(n_727)
);

BUFx12f_ASAP7_75t_L g728 ( 
.A(n_385),
.Y(n_728)
);

OAI21x1_ASAP7_75t_L g729 ( 
.A1(n_406),
.A2(n_410),
.B(n_407),
.Y(n_729)
);

BUFx6f_ASAP7_75t_L g730 ( 
.A(n_411),
.Y(n_730)
);

BUFx8_ASAP7_75t_SL g731 ( 
.A(n_475),
.Y(n_731)
);

BUFx3_ASAP7_75t_L g732 ( 
.A(n_388),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_413),
.Y(n_733)
);

AND2x4_ASAP7_75t_L g734 ( 
.A(n_416),
.B(n_28),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_423),
.Y(n_735)
);

INVx5_ASAP7_75t_L g736 ( 
.A(n_549),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_425),
.Y(n_737)
);

HB1xp67_ASAP7_75t_L g738 ( 
.A(n_461),
.Y(n_738)
);

BUFx2_ASAP7_75t_L g739 ( 
.A(n_515),
.Y(n_739)
);

INVx3_ASAP7_75t_L g740 ( 
.A(n_427),
.Y(n_740)
);

HB1xp67_ASAP7_75t_L g741 ( 
.A(n_431),
.Y(n_741)
);

AOI22x1_ASAP7_75t_SL g742 ( 
.A1(n_432),
.A2(n_29),
.B1(n_31),
.B2(n_32),
.Y(n_742)
);

AND2x2_ASAP7_75t_L g743 ( 
.A(n_517),
.B(n_33),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_437),
.B(n_33),
.Y(n_744)
);

INVx4_ASAP7_75t_L g745 ( 
.A(n_389),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_440),
.Y(n_746)
);

BUFx3_ASAP7_75t_L g747 ( 
.A(n_391),
.Y(n_747)
);

HB1xp67_ASAP7_75t_L g748 ( 
.A(n_442),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_443),
.Y(n_749)
);

OA21x2_ASAP7_75t_L g750 ( 
.A1(n_447),
.A2(n_34),
.B(n_36),
.Y(n_750)
);

BUFx6f_ASAP7_75t_L g751 ( 
.A(n_448),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_452),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_465),
.Y(n_753)
);

BUFx8_ASAP7_75t_SL g754 ( 
.A(n_492),
.Y(n_754)
);

BUFx6f_ASAP7_75t_L g755 ( 
.A(n_469),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_483),
.B(n_36),
.Y(n_756)
);

BUFx2_ASAP7_75t_L g757 ( 
.A(n_523),
.Y(n_757)
);

INVx5_ASAP7_75t_L g758 ( 
.A(n_530),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_487),
.Y(n_759)
);

BUFx3_ASAP7_75t_L g760 ( 
.A(n_392),
.Y(n_760)
);

BUFx6f_ASAP7_75t_L g761 ( 
.A(n_491),
.Y(n_761)
);

BUFx8_ASAP7_75t_SL g762 ( 
.A(n_541),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_625),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_607),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_754),
.Y(n_765)
);

CKINVDCx16_ASAP7_75t_R g766 ( 
.A(n_652),
.Y(n_766)
);

CKINVDCx5p33_ASAP7_75t_R g767 ( 
.A(n_762),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_613),
.Y(n_768)
);

CKINVDCx5p33_ASAP7_75t_R g769 ( 
.A(n_675),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_690),
.Y(n_770)
);

CKINVDCx5p33_ASAP7_75t_R g771 ( 
.A(n_696),
.Y(n_771)
);

INVx3_ASAP7_75t_L g772 ( 
.A(n_610),
.Y(n_772)
);

CKINVDCx5p33_ASAP7_75t_R g773 ( 
.A(n_720),
.Y(n_773)
);

CKINVDCx5p33_ASAP7_75t_R g774 ( 
.A(n_728),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_603),
.Y(n_775)
);

NOR2xp33_ASAP7_75t_R g776 ( 
.A(n_710),
.B(n_551),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_731),
.Y(n_777)
);

BUFx6f_ASAP7_75t_L g778 ( 
.A(n_615),
.Y(n_778)
);

CKINVDCx16_ASAP7_75t_R g779 ( 
.A(n_641),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_732),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_747),
.Y(n_781)
);

CKINVDCx20_ASAP7_75t_R g782 ( 
.A(n_757),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_760),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_606),
.Y(n_784)
);

NOR2xp33_ASAP7_75t_R g785 ( 
.A(n_710),
.B(n_573),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_603),
.Y(n_786)
);

CKINVDCx20_ASAP7_75t_R g787 ( 
.A(n_727),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_674),
.Y(n_788)
);

OR2x2_ASAP7_75t_L g789 ( 
.A(n_632),
.B(n_38),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_695),
.Y(n_790)
);

CKINVDCx5p33_ASAP7_75t_R g791 ( 
.A(n_678),
.Y(n_791)
);

CKINVDCx5p33_ASAP7_75t_R g792 ( 
.A(n_688),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_695),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_695),
.Y(n_794)
);

CKINVDCx20_ASAP7_75t_R g795 ( 
.A(n_739),
.Y(n_795)
);

CKINVDCx20_ASAP7_75t_R g796 ( 
.A(n_651),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_610),
.Y(n_797)
);

CKINVDCx5p33_ASAP7_75t_R g798 ( 
.A(n_691),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_615),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_719),
.Y(n_800)
);

AND2x2_ASAP7_75t_L g801 ( 
.A(n_736),
.B(n_520),
.Y(n_801)
);

AOI21x1_ASAP7_75t_L g802 ( 
.A1(n_670),
.A2(n_495),
.B(n_493),
.Y(n_802)
);

CKINVDCx16_ASAP7_75t_R g803 ( 
.A(n_722),
.Y(n_803)
);

CKINVDCx5p33_ASAP7_75t_R g804 ( 
.A(n_745),
.Y(n_804)
);

NOR2x1p5_ASAP7_75t_L g805 ( 
.A(n_668),
.B(n_394),
.Y(n_805)
);

CKINVDCx20_ASAP7_75t_R g806 ( 
.A(n_692),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_672),
.Y(n_807)
);

CKINVDCx5p33_ASAP7_75t_R g808 ( 
.A(n_745),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_615),
.Y(n_809)
);

CKINVDCx5p33_ASAP7_75t_R g810 ( 
.A(n_736),
.Y(n_810)
);

BUFx2_ASAP7_75t_L g811 ( 
.A(n_693),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_672),
.Y(n_812)
);

NOR2xp33_ASAP7_75t_R g813 ( 
.A(n_632),
.B(n_396),
.Y(n_813)
);

CKINVDCx5p33_ASAP7_75t_R g814 ( 
.A(n_736),
.Y(n_814)
);

CKINVDCx5p33_ASAP7_75t_R g815 ( 
.A(n_702),
.Y(n_815)
);

BUFx3_ASAP7_75t_L g816 ( 
.A(n_672),
.Y(n_816)
);

BUFx6f_ASAP7_75t_L g817 ( 
.A(n_631),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_676),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_715),
.Y(n_819)
);

NOR2xp33_ASAP7_75t_L g820 ( 
.A(n_656),
.B(n_595),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_631),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_676),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_676),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_721),
.Y(n_824)
);

BUFx6f_ASAP7_75t_L g825 ( 
.A(n_631),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_685),
.Y(n_826)
);

CKINVDCx5p33_ASAP7_75t_R g827 ( 
.A(n_669),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_685),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_640),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_685),
.Y(n_830)
);

NOR2xp33_ASAP7_75t_R g831 ( 
.A(n_648),
.B(n_397),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_686),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_640),
.Y(n_833)
);

CKINVDCx5p33_ASAP7_75t_R g834 ( 
.A(n_669),
.Y(n_834)
);

BUFx10_ASAP7_75t_L g835 ( 
.A(n_671),
.Y(n_835)
);

CKINVDCx20_ASAP7_75t_R g836 ( 
.A(n_626),
.Y(n_836)
);

CKINVDCx5p33_ASAP7_75t_R g837 ( 
.A(n_669),
.Y(n_837)
);

CKINVDCx5p33_ASAP7_75t_R g838 ( 
.A(n_681),
.Y(n_838)
);

CKINVDCx5p33_ASAP7_75t_R g839 ( 
.A(n_681),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_686),
.Y(n_840)
);

CKINVDCx5p33_ASAP7_75t_R g841 ( 
.A(n_681),
.Y(n_841)
);

CKINVDCx20_ASAP7_75t_R g842 ( 
.A(n_636),
.Y(n_842)
);

CKINVDCx5p33_ASAP7_75t_R g843 ( 
.A(n_694),
.Y(n_843)
);

CKINVDCx5p33_ASAP7_75t_R g844 ( 
.A(n_694),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_640),
.Y(n_845)
);

CKINVDCx20_ASAP7_75t_R g846 ( 
.A(n_662),
.Y(n_846)
);

INVx3_ASAP7_75t_L g847 ( 
.A(n_645),
.Y(n_847)
);

BUFx2_ASAP7_75t_L g848 ( 
.A(n_694),
.Y(n_848)
);

CKINVDCx5p33_ASAP7_75t_R g849 ( 
.A(n_677),
.Y(n_849)
);

CKINVDCx5p33_ASAP7_75t_R g850 ( 
.A(n_723),
.Y(n_850)
);

CKINVDCx5p33_ASAP7_75t_R g851 ( 
.A(n_617),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_686),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_689),
.Y(n_853)
);

BUFx10_ASAP7_75t_L g854 ( 
.A(n_647),
.Y(n_854)
);

NOR2xp67_ASAP7_75t_L g855 ( 
.A(n_758),
.B(n_497),
.Y(n_855)
);

CKINVDCx5p33_ASAP7_75t_R g856 ( 
.A(n_618),
.Y(n_856)
);

HB1xp67_ASAP7_75t_L g857 ( 
.A(n_609),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_689),
.Y(n_858)
);

CKINVDCx20_ASAP7_75t_R g859 ( 
.A(n_717),
.Y(n_859)
);

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_689),
.Y(n_860)
);

CKINVDCx5p33_ASAP7_75t_R g861 ( 
.A(n_758),
.Y(n_861)
);

HB1xp67_ASAP7_75t_L g862 ( 
.A(n_648),
.Y(n_862)
);

NOR2xp33_ASAP7_75t_R g863 ( 
.A(n_654),
.B(n_399),
.Y(n_863)
);

OAI22xp33_ASAP7_75t_SL g864 ( 
.A1(n_682),
.A2(n_503),
.B1(n_506),
.B2(n_499),
.Y(n_864)
);

CKINVDCx20_ASAP7_75t_R g865 ( 
.A(n_741),
.Y(n_865)
);

CKINVDCx5p33_ASAP7_75t_R g866 ( 
.A(n_758),
.Y(n_866)
);

NOR2xp67_ASAP7_75t_L g867 ( 
.A(n_635),
.B(n_507),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_SL g868 ( 
.A(n_820),
.B(n_630),
.Y(n_868)
);

INVxp67_ASAP7_75t_SL g869 ( 
.A(n_816),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_801),
.B(n_621),
.Y(n_870)
);

INVx3_ASAP7_75t_L g871 ( 
.A(n_778),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_790),
.B(n_793),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_794),
.B(n_799),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_847),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_809),
.B(n_635),
.Y(n_875)
);

NOR2xp33_ASAP7_75t_L g876 ( 
.A(n_862),
.B(n_700),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_821),
.B(n_635),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_847),
.Y(n_878)
);

BUFx8_ASAP7_75t_L g879 ( 
.A(n_811),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_829),
.Y(n_880)
);

NOR2xp33_ASAP7_75t_L g881 ( 
.A(n_862),
.B(n_743),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_833),
.B(n_637),
.Y(n_882)
);

NAND2xp33_ASAP7_75t_L g883 ( 
.A(n_860),
.B(n_612),
.Y(n_883)
);

NAND2xp33_ASAP7_75t_L g884 ( 
.A(n_813),
.B(n_616),
.Y(n_884)
);

NOR2xp33_ASAP7_75t_L g885 ( 
.A(n_804),
.B(n_620),
.Y(n_885)
);

NOR2xp33_ASAP7_75t_L g886 ( 
.A(n_808),
.B(n_622),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_845),
.B(n_637),
.Y(n_887)
);

NOR2xp33_ASAP7_75t_L g888 ( 
.A(n_769),
.B(n_638),
.Y(n_888)
);

BUFx6f_ASAP7_75t_L g889 ( 
.A(n_778),
.Y(n_889)
);

NOR2xp33_ASAP7_75t_L g890 ( 
.A(n_770),
.B(n_654),
.Y(n_890)
);

BUFx6f_ASAP7_75t_L g891 ( 
.A(n_778),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_SL g892 ( 
.A(n_776),
.B(n_704),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_768),
.B(n_637),
.Y(n_893)
);

NAND2xp33_ASAP7_75t_L g894 ( 
.A(n_831),
.B(n_706),
.Y(n_894)
);

AND2x2_ASAP7_75t_L g895 ( 
.A(n_848),
.B(n_657),
.Y(n_895)
);

INVx3_ASAP7_75t_L g896 ( 
.A(n_778),
.Y(n_896)
);

INVx2_ASAP7_75t_L g897 ( 
.A(n_817),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_807),
.Y(n_898)
);

CKINVDCx5p33_ASAP7_75t_R g899 ( 
.A(n_771),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_812),
.Y(n_900)
);

NOR2xp33_ASAP7_75t_L g901 ( 
.A(n_773),
.B(n_657),
.Y(n_901)
);

NOR2xp67_ASAP7_75t_L g902 ( 
.A(n_772),
.B(n_666),
.Y(n_902)
);

NAND2xp33_ASAP7_75t_L g903 ( 
.A(n_863),
.B(n_707),
.Y(n_903)
);

INVx2_ASAP7_75t_L g904 ( 
.A(n_817),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_772),
.B(n_666),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_775),
.B(n_704),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_786),
.B(n_734),
.Y(n_907)
);

NAND3xp33_ASAP7_75t_L g908 ( 
.A(n_849),
.B(n_748),
.C(n_716),
.Y(n_908)
);

INVx8_ASAP7_75t_L g909 ( 
.A(n_763),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_SL g910 ( 
.A(n_785),
.B(n_608),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_818),
.B(n_822),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_823),
.B(n_734),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_826),
.B(n_709),
.Y(n_913)
);

AND2x2_ASAP7_75t_L g914 ( 
.A(n_835),
.B(n_680),
.Y(n_914)
);

NOR3xp33_ASAP7_75t_L g915 ( 
.A(n_864),
.B(n_756),
.C(n_744),
.Y(n_915)
);

AND2x2_ASAP7_75t_L g916 ( 
.A(n_835),
.B(n_687),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_817),
.Y(n_917)
);

INVxp67_ASAP7_75t_L g918 ( 
.A(n_857),
.Y(n_918)
);

INVx2_ASAP7_75t_SL g919 ( 
.A(n_805),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_828),
.B(n_830),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_832),
.Y(n_921)
);

INVxp67_ASAP7_75t_SL g922 ( 
.A(n_817),
.Y(n_922)
);

BUFx6f_ASAP7_75t_SL g923 ( 
.A(n_854),
.Y(n_923)
);

AOI22xp5_ASAP7_75t_L g924 ( 
.A1(n_859),
.A2(n_624),
.B1(n_663),
.B2(n_643),
.Y(n_924)
);

AOI22xp33_ASAP7_75t_L g925 ( 
.A1(n_789),
.A2(n_655),
.B1(n_665),
.B2(n_608),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_SL g926 ( 
.A(n_815),
.B(n_655),
.Y(n_926)
);

BUFx3_ASAP7_75t_L g927 ( 
.A(n_840),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_SL g928 ( 
.A(n_819),
.B(n_665),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_825),
.Y(n_929)
);

INVxp33_ASAP7_75t_L g930 ( 
.A(n_857),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_SL g931 ( 
.A(n_824),
.B(n_679),
.Y(n_931)
);

INVx2_ASAP7_75t_L g932 ( 
.A(n_825),
.Y(n_932)
);

AND2x4_ASAP7_75t_L g933 ( 
.A(n_852),
.B(n_679),
.Y(n_933)
);

NOR2xp33_ASAP7_75t_L g934 ( 
.A(n_780),
.B(n_673),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_853),
.B(n_709),
.Y(n_935)
);

INVx2_ASAP7_75t_L g936 ( 
.A(n_825),
.Y(n_936)
);

AND2x2_ASAP7_75t_L g937 ( 
.A(n_861),
.B(n_738),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_858),
.B(n_825),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_SL g939 ( 
.A(n_850),
.B(n_684),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_764),
.B(n_797),
.Y(n_940)
);

INVx3_ASAP7_75t_L g941 ( 
.A(n_802),
.Y(n_941)
);

BUFx6f_ASAP7_75t_L g942 ( 
.A(n_854),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_855),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_SL g944 ( 
.A(n_781),
.B(n_684),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_867),
.Y(n_945)
);

BUFx6f_ASAP7_75t_L g946 ( 
.A(n_866),
.Y(n_946)
);

AND2x4_ASAP7_75t_L g947 ( 
.A(n_783),
.B(n_604),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_810),
.B(n_709),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_814),
.Y(n_949)
);

BUFx5_ASAP7_75t_L g950 ( 
.A(n_827),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_834),
.B(n_711),
.Y(n_951)
);

NOR2xp33_ASAP7_75t_L g952 ( 
.A(n_851),
.B(n_856),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_837),
.Y(n_953)
);

INVx2_ASAP7_75t_L g954 ( 
.A(n_838),
.Y(n_954)
);

INVx2_ASAP7_75t_L g955 ( 
.A(n_839),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_841),
.B(n_711),
.Y(n_956)
);

OR2x2_ASAP7_75t_L g957 ( 
.A(n_766),
.B(n_605),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_843),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_844),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_865),
.Y(n_960)
);

BUFx3_ASAP7_75t_L g961 ( 
.A(n_909),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_885),
.B(n_886),
.Y(n_962)
);

INVx2_ASAP7_75t_L g963 ( 
.A(n_874),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_870),
.B(n_711),
.Y(n_964)
);

NAND2xp33_ASAP7_75t_SL g965 ( 
.A(n_942),
.B(n_892),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_881),
.B(n_729),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_868),
.B(n_511),
.Y(n_967)
);

INVx2_ASAP7_75t_SL g968 ( 
.A(n_914),
.Y(n_968)
);

AO22x1_ASAP7_75t_L g969 ( 
.A1(n_915),
.A2(n_705),
.B1(n_634),
.B2(n_619),
.Y(n_969)
);

AOI21xp5_ASAP7_75t_L g970 ( 
.A1(n_941),
.A2(n_628),
.B(n_627),
.Y(n_970)
);

NOR3xp33_ASAP7_75t_L g971 ( 
.A(n_888),
.B(n_803),
.C(n_779),
.Y(n_971)
);

NOR2xp33_ASAP7_75t_L g972 ( 
.A(n_934),
.B(n_796),
.Y(n_972)
);

OAI21xp5_ASAP7_75t_L g973 ( 
.A1(n_941),
.A2(n_708),
.B(n_650),
.Y(n_973)
);

INVx2_ASAP7_75t_L g974 ( 
.A(n_878),
.Y(n_974)
);

HB1xp67_ASAP7_75t_L g975 ( 
.A(n_918),
.Y(n_975)
);

INVx2_ASAP7_75t_L g976 ( 
.A(n_880),
.Y(n_976)
);

AOI22xp5_ASAP7_75t_L g977 ( 
.A1(n_876),
.A2(n_806),
.B1(n_842),
.B2(n_836),
.Y(n_977)
);

AOI22xp33_ASAP7_75t_L g978 ( 
.A1(n_925),
.A2(n_750),
.B1(n_683),
.B2(n_712),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_940),
.Y(n_979)
);

AOI22xp5_ASAP7_75t_L g980 ( 
.A1(n_884),
.A2(n_846),
.B1(n_596),
.B2(n_409),
.Y(n_980)
);

OAI21xp5_ASAP7_75t_L g981 ( 
.A1(n_907),
.A2(n_750),
.B(n_683),
.Y(n_981)
);

INVx2_ASAP7_75t_SL g982 ( 
.A(n_916),
.Y(n_982)
);

NOR3xp33_ASAP7_75t_SL g983 ( 
.A(n_908),
.B(n_800),
.C(n_784),
.Y(n_983)
);

INVx2_ASAP7_75t_SL g984 ( 
.A(n_895),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_913),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_935),
.Y(n_986)
);

INVx5_ASAP7_75t_L g987 ( 
.A(n_946),
.Y(n_987)
);

INVxp67_ASAP7_75t_SL g988 ( 
.A(n_902),
.Y(n_988)
);

AND2x4_ASAP7_75t_L g989 ( 
.A(n_869),
.B(n_933),
.Y(n_989)
);

NOR2xp67_ASAP7_75t_L g990 ( 
.A(n_952),
.B(n_765),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_SL g991 ( 
.A(n_947),
.B(n_890),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_873),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_906),
.B(n_933),
.Y(n_993)
);

BUFx4f_ASAP7_75t_L g994 ( 
.A(n_942),
.Y(n_994)
);

INVx8_ASAP7_75t_L g995 ( 
.A(n_909),
.Y(n_995)
);

AND2x4_ASAP7_75t_L g996 ( 
.A(n_927),
.B(n_633),
.Y(n_996)
);

NOR2x1p5_ASAP7_75t_L g997 ( 
.A(n_942),
.B(n_788),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_SL g998 ( 
.A(n_947),
.B(n_774),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_872),
.Y(n_999)
);

INVxp67_ASAP7_75t_SL g1000 ( 
.A(n_902),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_SL g1001 ( 
.A(n_901),
.B(n_791),
.Y(n_1001)
);

CKINVDCx5p33_ASAP7_75t_R g1002 ( 
.A(n_899),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_912),
.B(n_522),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_911),
.Y(n_1004)
);

BUFx3_ASAP7_75t_L g1005 ( 
.A(n_946),
.Y(n_1005)
);

BUFx6f_ASAP7_75t_L g1006 ( 
.A(n_889),
.Y(n_1006)
);

OAI22xp33_ASAP7_75t_L g1007 ( 
.A1(n_924),
.A2(n_930),
.B1(n_919),
.B2(n_910),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_950),
.B(n_524),
.Y(n_1008)
);

NOR2xp33_ASAP7_75t_L g1009 ( 
.A(n_939),
.B(n_782),
.Y(n_1009)
);

AND2x4_ASAP7_75t_L g1010 ( 
.A(n_898),
.B(n_900),
.Y(n_1010)
);

INVx2_ASAP7_75t_L g1011 ( 
.A(n_871),
.Y(n_1011)
);

INVx3_ASAP7_75t_L g1012 ( 
.A(n_957),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_920),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_921),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_950),
.B(n_534),
.Y(n_1015)
);

OAI21xp33_ASAP7_75t_L g1016 ( 
.A1(n_926),
.A2(n_623),
.B(n_611),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_938),
.Y(n_1017)
);

INVx2_ASAP7_75t_L g1018 ( 
.A(n_871),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_905),
.Y(n_1019)
);

AND2x4_ASAP7_75t_L g1020 ( 
.A(n_948),
.B(n_951),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_897),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_SL g1022 ( 
.A(n_946),
.B(n_798),
.Y(n_1022)
);

CKINVDCx5p33_ASAP7_75t_R g1023 ( 
.A(n_923),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_950),
.B(n_535),
.Y(n_1024)
);

INVx4_ASAP7_75t_L g1025 ( 
.A(n_889),
.Y(n_1025)
);

AOI22xp5_ASAP7_75t_L g1026 ( 
.A1(n_894),
.A2(n_412),
.B1(n_415),
.B2(n_404),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_950),
.B(n_545),
.Y(n_1027)
);

BUFx6f_ASAP7_75t_L g1028 ( 
.A(n_889),
.Y(n_1028)
);

INVx2_ASAP7_75t_L g1029 ( 
.A(n_896),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_904),
.Y(n_1030)
);

INVxp67_ASAP7_75t_L g1031 ( 
.A(n_937),
.Y(n_1031)
);

AND2x4_ASAP7_75t_L g1032 ( 
.A(n_956),
.B(n_639),
.Y(n_1032)
);

BUFx2_ASAP7_75t_L g1033 ( 
.A(n_960),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_917),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_950),
.B(n_548),
.Y(n_1035)
);

INVx2_ASAP7_75t_L g1036 ( 
.A(n_896),
.Y(n_1036)
);

INVx4_ASAP7_75t_L g1037 ( 
.A(n_891),
.Y(n_1037)
);

NOR2xp33_ASAP7_75t_L g1038 ( 
.A(n_944),
.B(n_787),
.Y(n_1038)
);

INVx2_ASAP7_75t_L g1039 ( 
.A(n_891),
.Y(n_1039)
);

AND2x2_ASAP7_75t_L g1040 ( 
.A(n_928),
.B(n_614),
.Y(n_1040)
);

AND2x4_ASAP7_75t_L g1041 ( 
.A(n_953),
.B(n_954),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_929),
.Y(n_1042)
);

INVxp67_ASAP7_75t_L g1043 ( 
.A(n_931),
.Y(n_1043)
);

AOI22xp5_ASAP7_75t_L g1044 ( 
.A1(n_903),
.A2(n_883),
.B1(n_949),
.B2(n_958),
.Y(n_1044)
);

INVx2_ASAP7_75t_L g1045 ( 
.A(n_891),
.Y(n_1045)
);

A2O1A1Ixp33_ASAP7_75t_L g1046 ( 
.A1(n_959),
.A2(n_484),
.B(n_508),
.C(n_459),
.Y(n_1046)
);

INVx2_ASAP7_75t_SL g1047 ( 
.A(n_955),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_SL g1048 ( 
.A(n_943),
.B(n_792),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_932),
.B(n_558),
.Y(n_1049)
);

INVx3_ASAP7_75t_L g1050 ( 
.A(n_936),
.Y(n_1050)
);

INVx2_ASAP7_75t_SL g1051 ( 
.A(n_879),
.Y(n_1051)
);

BUFx3_ASAP7_75t_L g1052 ( 
.A(n_879),
.Y(n_1052)
);

AOI22xp5_ASAP7_75t_L g1053 ( 
.A1(n_945),
.A2(n_419),
.B1(n_421),
.B2(n_418),
.Y(n_1053)
);

AOI22xp5_ASAP7_75t_L g1054 ( 
.A1(n_923),
.A2(n_428),
.B1(n_429),
.B2(n_426),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_922),
.B(n_563),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_893),
.B(n_567),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_SL g1057 ( 
.A(n_875),
.B(n_430),
.Y(n_1057)
);

AOI22xp5_ASAP7_75t_L g1058 ( 
.A1(n_877),
.A2(n_439),
.B1(n_444),
.B2(n_433),
.Y(n_1058)
);

BUFx4f_ASAP7_75t_L g1059 ( 
.A(n_882),
.Y(n_1059)
);

NOR2xp33_ASAP7_75t_R g1060 ( 
.A(n_887),
.B(n_767),
.Y(n_1060)
);

NOR2xp33_ASAP7_75t_SL g1061 ( 
.A(n_1002),
.B(n_777),
.Y(n_1061)
);

OA21x2_ASAP7_75t_L g1062 ( 
.A1(n_981),
.A2(n_973),
.B(n_966),
.Y(n_1062)
);

CKINVDCx5p33_ASAP7_75t_R g1063 ( 
.A(n_995),
.Y(n_1063)
);

CKINVDCx5p33_ASAP7_75t_R g1064 ( 
.A(n_995),
.Y(n_1064)
);

OAI22xp5_ASAP7_75t_L g1065 ( 
.A1(n_962),
.A2(n_571),
.B1(n_579),
.B2(n_569),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_979),
.B(n_583),
.Y(n_1066)
);

BUFx12f_ASAP7_75t_L g1067 ( 
.A(n_997),
.Y(n_1067)
);

NOR2xp33_ASAP7_75t_L g1068 ( 
.A(n_1031),
.B(n_795),
.Y(n_1068)
);

NAND3xp33_ASAP7_75t_SL g1069 ( 
.A(n_977),
.B(n_449),
.C(n_446),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_SL g1070 ( 
.A(n_987),
.B(n_993),
.Y(n_1070)
);

INVx4_ASAP7_75t_L g1071 ( 
.A(n_987),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_1014),
.Y(n_1072)
);

BUFx2_ASAP7_75t_L g1073 ( 
.A(n_1012),
.Y(n_1073)
);

AOI21xp5_ASAP7_75t_L g1074 ( 
.A1(n_988),
.A2(n_658),
.B(n_645),
.Y(n_1074)
);

INVx5_ASAP7_75t_L g1075 ( 
.A(n_987),
.Y(n_1075)
);

AOI21xp5_ASAP7_75t_L g1076 ( 
.A1(n_1000),
.A2(n_658),
.B(n_645),
.Y(n_1076)
);

AOI21xp5_ASAP7_75t_L g1077 ( 
.A1(n_964),
.A2(n_658),
.B(n_586),
.Y(n_1077)
);

CKINVDCx14_ASAP7_75t_R g1078 ( 
.A(n_961),
.Y(n_1078)
);

AO22x1_ASAP7_75t_L g1079 ( 
.A1(n_972),
.A2(n_742),
.B1(n_614),
.B2(n_590),
.Y(n_1079)
);

INVx3_ASAP7_75t_L g1080 ( 
.A(n_1050),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_SL g1081 ( 
.A(n_994),
.B(n_450),
.Y(n_1081)
);

INVx2_ASAP7_75t_L g1082 ( 
.A(n_1050),
.Y(n_1082)
);

NOR2xp33_ASAP7_75t_R g1083 ( 
.A(n_965),
.B(n_451),
.Y(n_1083)
);

BUFx8_ASAP7_75t_L g1084 ( 
.A(n_1051),
.Y(n_1084)
);

HB1xp67_ASAP7_75t_L g1085 ( 
.A(n_975),
.Y(n_1085)
);

AO21x1_ASAP7_75t_L g1086 ( 
.A1(n_1008),
.A2(n_585),
.B(n_670),
.Y(n_1086)
);

BUFx3_ASAP7_75t_L g1087 ( 
.A(n_1005),
.Y(n_1087)
);

AOI21xp5_ASAP7_75t_L g1088 ( 
.A1(n_978),
.A2(n_644),
.B(n_629),
.Y(n_1088)
);

A2O1A1Ixp33_ASAP7_75t_L g1089 ( 
.A1(n_1019),
.A2(n_699),
.B(n_714),
.C(n_697),
.Y(n_1089)
);

OAI22xp5_ASAP7_75t_L g1090 ( 
.A1(n_1044),
.A2(n_454),
.B1(n_456),
.B2(n_453),
.Y(n_1090)
);

INVx2_ASAP7_75t_L g1091 ( 
.A(n_976),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_1021),
.Y(n_1092)
);

NOR2xp33_ASAP7_75t_L g1093 ( 
.A(n_1007),
.B(n_742),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_1030),
.Y(n_1094)
);

AOI22xp33_ASAP7_75t_SL g1095 ( 
.A1(n_1009),
.A2(n_725),
.B1(n_724),
.B2(n_460),
.Y(n_1095)
);

AOI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_1015),
.A2(n_661),
.B(n_646),
.Y(n_1096)
);

AND2x2_ASAP7_75t_SL g1097 ( 
.A(n_971),
.B(n_724),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_SL g1098 ( 
.A(n_989),
.B(n_457),
.Y(n_1098)
);

AOI22xp5_ASAP7_75t_L g1099 ( 
.A1(n_999),
.A2(n_468),
.B1(n_470),
.B2(n_462),
.Y(n_1099)
);

NAND2xp33_ASAP7_75t_SL g1100 ( 
.A(n_983),
.B(n_472),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_SL g1101 ( 
.A(n_989),
.B(n_473),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_1034),
.Y(n_1102)
);

NAND3xp33_ASAP7_75t_SL g1103 ( 
.A(n_980),
.B(n_477),
.C(n_474),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_1004),
.B(n_698),
.Y(n_1104)
);

INVx2_ASAP7_75t_L g1105 ( 
.A(n_963),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_SL g1106 ( 
.A(n_968),
.B(n_480),
.Y(n_1106)
);

NAND3xp33_ASAP7_75t_L g1107 ( 
.A(n_1043),
.B(n_726),
.C(n_718),
.Y(n_1107)
);

HB1xp67_ASAP7_75t_L g1108 ( 
.A(n_1033),
.Y(n_1108)
);

HB1xp67_ASAP7_75t_L g1109 ( 
.A(n_982),
.Y(n_1109)
);

BUFx6f_ASAP7_75t_L g1110 ( 
.A(n_1006),
.Y(n_1110)
);

AOI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_1024),
.A2(n_482),
.B(n_481),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_1042),
.Y(n_1112)
);

AOI21x1_ASAP7_75t_L g1113 ( 
.A1(n_1027),
.A2(n_1035),
.B(n_970),
.Y(n_1113)
);

OA21x2_ASAP7_75t_L g1114 ( 
.A1(n_1049),
.A2(n_701),
.B(n_703),
.Y(n_1114)
);

NOR2xp33_ASAP7_75t_R g1115 ( 
.A(n_1023),
.B(n_485),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_1013),
.B(n_733),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_SL g1117 ( 
.A(n_1020),
.B(n_489),
.Y(n_1117)
);

OAI22xp5_ASAP7_75t_L g1118 ( 
.A1(n_967),
.A2(n_577),
.B1(n_496),
.B2(n_500),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_992),
.B(n_752),
.Y(n_1119)
);

BUFx3_ASAP7_75t_L g1120 ( 
.A(n_996),
.Y(n_1120)
);

O2A1O1Ixp33_ASAP7_75t_L g1121 ( 
.A1(n_1046),
.A2(n_737),
.B(n_749),
.C(n_735),
.Y(n_1121)
);

OAI22xp5_ASAP7_75t_L g1122 ( 
.A1(n_1017),
.A2(n_574),
.B1(n_502),
.B2(n_509),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_985),
.B(n_759),
.Y(n_1123)
);

HB1xp67_ASAP7_75t_L g1124 ( 
.A(n_984),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_986),
.B(n_494),
.Y(n_1125)
);

OAI21x1_ASAP7_75t_L g1126 ( 
.A1(n_1011),
.A2(n_701),
.B(n_740),
.Y(n_1126)
);

NOR2xp33_ASAP7_75t_L g1127 ( 
.A(n_991),
.B(n_1038),
.Y(n_1127)
);

OAI22xp5_ASAP7_75t_L g1128 ( 
.A1(n_1020),
.A2(n_576),
.B1(n_516),
.B2(n_521),
.Y(n_1128)
);

INVx2_ASAP7_75t_L g1129 ( 
.A(n_974),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_1003),
.B(n_512),
.Y(n_1130)
);

AOI21xp5_ASAP7_75t_L g1131 ( 
.A1(n_1025),
.A2(n_526),
.B(n_525),
.Y(n_1131)
);

NOR2xp33_ASAP7_75t_R g1132 ( 
.A(n_1047),
.B(n_528),
.Y(n_1132)
);

OR2x6_ASAP7_75t_SL g1133 ( 
.A(n_1056),
.B(n_529),
.Y(n_1133)
);

AOI21xp5_ASAP7_75t_L g1134 ( 
.A1(n_1025),
.A2(n_533),
.B(n_532),
.Y(n_1134)
);

A2O1A1Ixp33_ASAP7_75t_L g1135 ( 
.A1(n_1040),
.A2(n_753),
.B(n_703),
.C(n_746),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_1018),
.Y(n_1136)
);

BUFx2_ASAP7_75t_L g1137 ( 
.A(n_996),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_SL g1138 ( 
.A(n_1032),
.B(n_1041),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_1032),
.B(n_537),
.Y(n_1139)
);

OAI21xp33_ASAP7_75t_SL g1140 ( 
.A1(n_1055),
.A2(n_746),
.B(n_649),
.Y(n_1140)
);

OAI21xp33_ASAP7_75t_L g1141 ( 
.A1(n_1016),
.A2(n_653),
.B(n_642),
.Y(n_1141)
);

O2A1O1Ixp33_ASAP7_75t_L g1142 ( 
.A1(n_1057),
.A2(n_740),
.B(n_660),
.C(n_664),
.Y(n_1142)
);

INVx3_ASAP7_75t_L g1143 ( 
.A(n_1039),
.Y(n_1143)
);

AOI21xp5_ASAP7_75t_L g1144 ( 
.A1(n_1037),
.A2(n_1028),
.B(n_1006),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_1072),
.Y(n_1145)
);

HB1xp67_ASAP7_75t_L g1146 ( 
.A(n_1085),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_1092),
.Y(n_1147)
);

OAI21x1_ASAP7_75t_L g1148 ( 
.A1(n_1113),
.A2(n_1036),
.B(n_1029),
.Y(n_1148)
);

INVx1_ASAP7_75t_SL g1149 ( 
.A(n_1108),
.Y(n_1149)
);

AND2x2_ASAP7_75t_L g1150 ( 
.A(n_1127),
.B(n_990),
.Y(n_1150)
);

AND2x2_ASAP7_75t_L g1151 ( 
.A(n_1137),
.B(n_1041),
.Y(n_1151)
);

NAND2x1p5_ASAP7_75t_L g1152 ( 
.A(n_1075),
.B(n_1071),
.Y(n_1152)
);

BUFx2_ASAP7_75t_L g1153 ( 
.A(n_1073),
.Y(n_1153)
);

NOR2xp33_ASAP7_75t_L g1154 ( 
.A(n_1093),
.B(n_1001),
.Y(n_1154)
);

INVx3_ASAP7_75t_L g1155 ( 
.A(n_1110),
.Y(n_1155)
);

OAI21x1_ASAP7_75t_L g1156 ( 
.A1(n_1126),
.A2(n_1045),
.B(n_1048),
.Y(n_1156)
);

NAND2x1p5_ASAP7_75t_L g1157 ( 
.A(n_1075),
.B(n_1037),
.Y(n_1157)
);

AND2x2_ASAP7_75t_L g1158 ( 
.A(n_1124),
.B(n_969),
.Y(n_1158)
);

BUFx2_ASAP7_75t_SL g1159 ( 
.A(n_1075),
.Y(n_1159)
);

BUFx2_ASAP7_75t_L g1160 ( 
.A(n_1087),
.Y(n_1160)
);

OR2x2_ASAP7_75t_L g1161 ( 
.A(n_1068),
.B(n_998),
.Y(n_1161)
);

OAI21x1_ASAP7_75t_L g1162 ( 
.A1(n_1088),
.A2(n_1026),
.B(n_1053),
.Y(n_1162)
);

BUFx3_ASAP7_75t_L g1163 ( 
.A(n_1063),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_1094),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_1102),
.Y(n_1165)
);

AO21x2_ASAP7_75t_L g1166 ( 
.A1(n_1086),
.A2(n_1010),
.B(n_1058),
.Y(n_1166)
);

BUFx2_ASAP7_75t_R g1167 ( 
.A(n_1064),
.Y(n_1167)
);

INVx4_ASAP7_75t_L g1168 ( 
.A(n_1110),
.Y(n_1168)
);

BUFx3_ASAP7_75t_L g1169 ( 
.A(n_1120),
.Y(n_1169)
);

BUFx6f_ASAP7_75t_L g1170 ( 
.A(n_1110),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_1112),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1091),
.Y(n_1172)
);

OAI21x1_ASAP7_75t_SL g1173 ( 
.A1(n_1144),
.A2(n_1054),
.B(n_667),
.Y(n_1173)
);

AND2x4_ASAP7_75t_L g1174 ( 
.A(n_1138),
.B(n_1010),
.Y(n_1174)
);

OAI21xp5_ASAP7_75t_L g1175 ( 
.A1(n_1062),
.A2(n_1059),
.B(n_1022),
.Y(n_1175)
);

AO21x2_ASAP7_75t_L g1176 ( 
.A1(n_1066),
.A2(n_1060),
.B(n_659),
.Y(n_1176)
);

OAI21xp5_ASAP7_75t_L g1177 ( 
.A1(n_1062),
.A2(n_539),
.B(n_538),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_1105),
.Y(n_1178)
);

OAI21x1_ASAP7_75t_L g1179 ( 
.A1(n_1143),
.A2(n_1028),
.B(n_1006),
.Y(n_1179)
);

NAND2x1p5_ASAP7_75t_L g1180 ( 
.A(n_1071),
.B(n_1028),
.Y(n_1180)
);

NAND2x1p5_ASAP7_75t_L g1181 ( 
.A(n_1080),
.B(n_1052),
.Y(n_1181)
);

INVx3_ASAP7_75t_L g1182 ( 
.A(n_1080),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_1104),
.B(n_540),
.Y(n_1183)
);

AND2x4_ASAP7_75t_L g1184 ( 
.A(n_1129),
.B(n_64),
.Y(n_1184)
);

AO21x2_ASAP7_75t_L g1185 ( 
.A1(n_1103),
.A2(n_1077),
.B(n_1130),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_1136),
.Y(n_1186)
);

INVx4_ASAP7_75t_SL g1187 ( 
.A(n_1067),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_1082),
.Y(n_1188)
);

AO21x2_ASAP7_75t_L g1189 ( 
.A1(n_1123),
.A2(n_730),
.B(n_713),
.Y(n_1189)
);

INVx2_ASAP7_75t_L g1190 ( 
.A(n_1114),
.Y(n_1190)
);

AO21x2_ASAP7_75t_L g1191 ( 
.A1(n_1119),
.A2(n_1070),
.B(n_1116),
.Y(n_1191)
);

INVx2_ASAP7_75t_L g1192 ( 
.A(n_1114),
.Y(n_1192)
);

BUFx10_ASAP7_75t_L g1193 ( 
.A(n_1097),
.Y(n_1193)
);

INVx3_ASAP7_75t_L g1194 ( 
.A(n_1143),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_1125),
.B(n_542),
.Y(n_1195)
);

OAI21x1_ASAP7_75t_L g1196 ( 
.A1(n_1096),
.A2(n_725),
.B(n_78),
.Y(n_1196)
);

BUFx3_ASAP7_75t_L g1197 ( 
.A(n_1084),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_1107),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_1089),
.Y(n_1199)
);

INVx2_ASAP7_75t_L g1200 ( 
.A(n_1109),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1135),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_1139),
.B(n_543),
.Y(n_1202)
);

INVx3_ASAP7_75t_L g1203 ( 
.A(n_1084),
.Y(n_1203)
);

AO21x2_ASAP7_75t_L g1204 ( 
.A1(n_1111),
.A2(n_730),
.B(n_713),
.Y(n_1204)
);

AO21x2_ASAP7_75t_L g1205 ( 
.A1(n_1069),
.A2(n_730),
.B(n_713),
.Y(n_1205)
);

INVx2_ASAP7_75t_L g1206 ( 
.A(n_1117),
.Y(n_1206)
);

OAI21x1_ASAP7_75t_L g1207 ( 
.A1(n_1074),
.A2(n_81),
.B(n_77),
.Y(n_1207)
);

INVx5_ASAP7_75t_L g1208 ( 
.A(n_1078),
.Y(n_1208)
);

BUFx6f_ASAP7_75t_L g1209 ( 
.A(n_1098),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1141),
.Y(n_1210)
);

AND2x4_ASAP7_75t_L g1211 ( 
.A(n_1101),
.B(n_82),
.Y(n_1211)
);

INVx8_ASAP7_75t_L g1212 ( 
.A(n_1061),
.Y(n_1212)
);

BUFx6f_ASAP7_75t_L g1213 ( 
.A(n_1106),
.Y(n_1213)
);

OR3x4_ASAP7_75t_SL g1214 ( 
.A(n_1079),
.B(n_39),
.C(n_40),
.Y(n_1214)
);

OAI21xp5_ASAP7_75t_L g1215 ( 
.A1(n_1065),
.A2(n_547),
.B(n_546),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_1140),
.Y(n_1216)
);

INVx2_ASAP7_75t_L g1217 ( 
.A(n_1145),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1147),
.Y(n_1218)
);

BUFx12f_ASAP7_75t_L g1219 ( 
.A(n_1208),
.Y(n_1219)
);

INVx2_ASAP7_75t_L g1220 ( 
.A(n_1164),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_L g1221 ( 
.A(n_1150),
.B(n_1210),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1165),
.Y(n_1222)
);

INVx2_ASAP7_75t_L g1223 ( 
.A(n_1171),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1186),
.Y(n_1224)
);

AO21x1_ASAP7_75t_SL g1225 ( 
.A1(n_1175),
.A2(n_1099),
.B(n_1133),
.Y(n_1225)
);

NAND2x1p5_ASAP7_75t_L g1226 ( 
.A(n_1168),
.B(n_1081),
.Y(n_1226)
);

OAI22xp5_ASAP7_75t_L g1227 ( 
.A1(n_1154),
.A2(n_1095),
.B1(n_1090),
.B2(n_1121),
.Y(n_1227)
);

INVx2_ASAP7_75t_L g1228 ( 
.A(n_1172),
.Y(n_1228)
);

BUFx12f_ASAP7_75t_L g1229 ( 
.A(n_1208),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1178),
.Y(n_1230)
);

OAI21x1_ASAP7_75t_L g1231 ( 
.A1(n_1148),
.A2(n_1156),
.B(n_1179),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1188),
.Y(n_1232)
);

HB1xp67_ASAP7_75t_L g1233 ( 
.A(n_1146),
.Y(n_1233)
);

INVxp67_ASAP7_75t_SL g1234 ( 
.A(n_1146),
.Y(n_1234)
);

INVx2_ASAP7_75t_L g1235 ( 
.A(n_1194),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1216),
.Y(n_1236)
);

AOI22xp33_ASAP7_75t_SL g1237 ( 
.A1(n_1154),
.A2(n_1083),
.B1(n_1115),
.B2(n_1132),
.Y(n_1237)
);

NAND2x1_ASAP7_75t_L g1238 ( 
.A(n_1168),
.B(n_1076),
.Y(n_1238)
);

HB1xp67_ASAP7_75t_L g1239 ( 
.A(n_1149),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_1182),
.B(n_1122),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_1194),
.Y(n_1241)
);

AO21x1_ASAP7_75t_L g1242 ( 
.A1(n_1177),
.A2(n_1100),
.B(n_1118),
.Y(n_1242)
);

INVx3_ASAP7_75t_L g1243 ( 
.A(n_1182),
.Y(n_1243)
);

OAI22xp5_ASAP7_75t_L g1244 ( 
.A1(n_1211),
.A2(n_1128),
.B1(n_1142),
.B2(n_1131),
.Y(n_1244)
);

OAI21x1_ASAP7_75t_L g1245 ( 
.A1(n_1196),
.A2(n_1134),
.B(n_85),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1198),
.Y(n_1246)
);

AOI22xp33_ASAP7_75t_SL g1247 ( 
.A1(n_1212),
.A2(n_588),
.B1(n_555),
.B2(n_557),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1184),
.Y(n_1248)
);

OAI22xp33_ASAP7_75t_L g1249 ( 
.A1(n_1161),
.A2(n_1212),
.B1(n_1214),
.B2(n_1206),
.Y(n_1249)
);

NAND2x1p5_ASAP7_75t_L g1250 ( 
.A(n_1170),
.B(n_751),
.Y(n_1250)
);

BUFx12f_ASAP7_75t_L g1251 ( 
.A(n_1208),
.Y(n_1251)
);

AND2x2_ASAP7_75t_L g1252 ( 
.A(n_1151),
.B(n_554),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1184),
.Y(n_1253)
);

INVx2_ASAP7_75t_L g1254 ( 
.A(n_1190),
.Y(n_1254)
);

BUFx10_ASAP7_75t_L g1255 ( 
.A(n_1209),
.Y(n_1255)
);

OAI21x1_ASAP7_75t_SL g1256 ( 
.A1(n_1175),
.A2(n_87),
.B(n_84),
.Y(n_1256)
);

BUFx12f_ASAP7_75t_L g1257 ( 
.A(n_1208),
.Y(n_1257)
);

BUFx4f_ASAP7_75t_L g1258 ( 
.A(n_1212),
.Y(n_1258)
);

AOI22xp33_ASAP7_75t_SL g1259 ( 
.A1(n_1214),
.A2(n_592),
.B1(n_566),
.B2(n_568),
.Y(n_1259)
);

BUFx3_ASAP7_75t_L g1260 ( 
.A(n_1160),
.Y(n_1260)
);

INVx2_ASAP7_75t_L g1261 ( 
.A(n_1190),
.Y(n_1261)
);

BUFx4f_ASAP7_75t_SL g1262 ( 
.A(n_1163),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1199),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1201),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1174),
.Y(n_1265)
);

AOI21x1_ASAP7_75t_L g1266 ( 
.A1(n_1192),
.A2(n_755),
.B(n_751),
.Y(n_1266)
);

AOI22xp33_ASAP7_75t_L g1267 ( 
.A1(n_1215),
.A2(n_598),
.B1(n_570),
.B2(n_584),
.Y(n_1267)
);

AOI22xp33_ASAP7_75t_L g1268 ( 
.A1(n_1215),
.A2(n_599),
.B1(n_589),
.B2(n_594),
.Y(n_1268)
);

INVx2_ASAP7_75t_SL g1269 ( 
.A(n_1169),
.Y(n_1269)
);

OAI21xp5_ASAP7_75t_L g1270 ( 
.A1(n_1162),
.A2(n_601),
.B(n_562),
.Y(n_1270)
);

NAND2x1p5_ASAP7_75t_L g1271 ( 
.A(n_1170),
.B(n_751),
.Y(n_1271)
);

OR2x2_ASAP7_75t_L g1272 ( 
.A(n_1149),
.B(n_761),
.Y(n_1272)
);

AND2x2_ASAP7_75t_L g1273 ( 
.A(n_1158),
.B(n_755),
.Y(n_1273)
);

INVx2_ASAP7_75t_L g1274 ( 
.A(n_1192),
.Y(n_1274)
);

NAND2x1p5_ASAP7_75t_L g1275 ( 
.A(n_1170),
.B(n_1155),
.Y(n_1275)
);

AND2x4_ASAP7_75t_L g1276 ( 
.A(n_1174),
.B(n_92),
.Y(n_1276)
);

INVx3_ASAP7_75t_L g1277 ( 
.A(n_1180),
.Y(n_1277)
);

CKINVDCx14_ASAP7_75t_R g1278 ( 
.A(n_1163),
.Y(n_1278)
);

OAI21x1_ASAP7_75t_SL g1279 ( 
.A1(n_1173),
.A2(n_1177),
.B(n_1202),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_L g1280 ( 
.A(n_1195),
.B(n_755),
.Y(n_1280)
);

AOI22xp33_ASAP7_75t_L g1281 ( 
.A1(n_1211),
.A2(n_761),
.B1(n_41),
.B2(n_42),
.Y(n_1281)
);

INVx2_ASAP7_75t_L g1282 ( 
.A(n_1155),
.Y(n_1282)
);

AOI21xp5_ASAP7_75t_SL g1283 ( 
.A1(n_1157),
.A2(n_761),
.B(n_222),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1200),
.Y(n_1284)
);

NAND2x1p5_ASAP7_75t_L g1285 ( 
.A(n_1213),
.B(n_93),
.Y(n_1285)
);

OAI22xp5_ASAP7_75t_L g1286 ( 
.A1(n_1202),
.A2(n_39),
.B1(n_41),
.B2(n_42),
.Y(n_1286)
);

AND2x2_ASAP7_75t_L g1287 ( 
.A(n_1153),
.B(n_43),
.Y(n_1287)
);

INVx2_ASAP7_75t_L g1288 ( 
.A(n_1180),
.Y(n_1288)
);

INVx2_ASAP7_75t_L g1289 ( 
.A(n_1191),
.Y(n_1289)
);

NAND2xp33_ASAP7_75t_R g1290 ( 
.A(n_1276),
.B(n_1203),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1236),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1254),
.Y(n_1292)
);

INVx2_ASAP7_75t_L g1293 ( 
.A(n_1217),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1220),
.Y(n_1294)
);

BUFx6f_ASAP7_75t_L g1295 ( 
.A(n_1219),
.Y(n_1295)
);

INVx2_ASAP7_75t_L g1296 ( 
.A(n_1223),
.Y(n_1296)
);

BUFx3_ASAP7_75t_L g1297 ( 
.A(n_1262),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_L g1298 ( 
.A(n_1221),
.B(n_1195),
.Y(n_1298)
);

CKINVDCx5p33_ASAP7_75t_R g1299 ( 
.A(n_1278),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_L g1300 ( 
.A(n_1221),
.B(n_1183),
.Y(n_1300)
);

CKINVDCx12_ASAP7_75t_R g1301 ( 
.A(n_1287),
.Y(n_1301)
);

OR2x4_ASAP7_75t_L g1302 ( 
.A(n_1272),
.B(n_1209),
.Y(n_1302)
);

INVx2_ASAP7_75t_L g1303 ( 
.A(n_1228),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1218),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1222),
.Y(n_1305)
);

NAND2x1p5_ASAP7_75t_L g1306 ( 
.A(n_1260),
.B(n_1169),
.Y(n_1306)
);

NOR2xp33_ASAP7_75t_L g1307 ( 
.A(n_1249),
.B(n_1237),
.Y(n_1307)
);

AOI22xp33_ASAP7_75t_L g1308 ( 
.A1(n_1227),
.A2(n_1259),
.B1(n_1249),
.B2(n_1237),
.Y(n_1308)
);

NAND2xp33_ASAP7_75t_R g1309 ( 
.A(n_1276),
.B(n_1203),
.Y(n_1309)
);

BUFx2_ASAP7_75t_L g1310 ( 
.A(n_1239),
.Y(n_1310)
);

CKINVDCx5p33_ASAP7_75t_R g1311 ( 
.A(n_1229),
.Y(n_1311)
);

OR2x6_ASAP7_75t_L g1312 ( 
.A(n_1251),
.B(n_1159),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1224),
.Y(n_1313)
);

AOI22xp33_ASAP7_75t_L g1314 ( 
.A1(n_1227),
.A2(n_1209),
.B1(n_1213),
.B2(n_1193),
.Y(n_1314)
);

AOI22xp33_ASAP7_75t_SL g1315 ( 
.A1(n_1286),
.A2(n_1213),
.B1(n_1193),
.B2(n_1176),
.Y(n_1315)
);

AND2x2_ASAP7_75t_L g1316 ( 
.A(n_1273),
.B(n_1183),
.Y(n_1316)
);

CKINVDCx5p33_ASAP7_75t_R g1317 ( 
.A(n_1257),
.Y(n_1317)
);

AND2x2_ASAP7_75t_SL g1318 ( 
.A(n_1258),
.B(n_1167),
.Y(n_1318)
);

BUFx3_ASAP7_75t_L g1319 ( 
.A(n_1255),
.Y(n_1319)
);

INVxp67_ASAP7_75t_SL g1320 ( 
.A(n_1239),
.Y(n_1320)
);

HB1xp67_ASAP7_75t_L g1321 ( 
.A(n_1233),
.Y(n_1321)
);

INVx4_ASAP7_75t_L g1322 ( 
.A(n_1258),
.Y(n_1322)
);

INVx2_ASAP7_75t_L g1323 ( 
.A(n_1230),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1232),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_L g1325 ( 
.A(n_1246),
.B(n_1176),
.Y(n_1325)
);

CKINVDCx5p33_ASAP7_75t_R g1326 ( 
.A(n_1255),
.Y(n_1326)
);

OAI22xp5_ASAP7_75t_L g1327 ( 
.A1(n_1259),
.A2(n_1181),
.B1(n_1167),
.B2(n_1152),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1263),
.Y(n_1328)
);

O2A1O1Ixp33_ASAP7_75t_SL g1329 ( 
.A1(n_1240),
.A2(n_1166),
.B(n_1152),
.C(n_1157),
.Y(n_1329)
);

INVx3_ASAP7_75t_L g1330 ( 
.A(n_1277),
.Y(n_1330)
);

CKINVDCx5p33_ASAP7_75t_R g1331 ( 
.A(n_1269),
.Y(n_1331)
);

CKINVDCx16_ASAP7_75t_R g1332 ( 
.A(n_1252),
.Y(n_1332)
);

CKINVDCx5p33_ASAP7_75t_R g1333 ( 
.A(n_1233),
.Y(n_1333)
);

OR2x6_ASAP7_75t_L g1334 ( 
.A(n_1285),
.B(n_1197),
.Y(n_1334)
);

NOR2x1_ASAP7_75t_L g1335 ( 
.A(n_1277),
.B(n_1197),
.Y(n_1335)
);

AOI22xp33_ASAP7_75t_L g1336 ( 
.A1(n_1281),
.A2(n_1166),
.B1(n_1191),
.B2(n_1205),
.Y(n_1336)
);

INVxp67_ASAP7_75t_L g1337 ( 
.A(n_1234),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_L g1338 ( 
.A(n_1284),
.B(n_1181),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1264),
.Y(n_1339)
);

NAND2xp33_ASAP7_75t_SL g1340 ( 
.A(n_1248),
.B(n_1187),
.Y(n_1340)
);

NOR2xp33_ASAP7_75t_R g1341 ( 
.A(n_1265),
.B(n_1187),
.Y(n_1341)
);

AND2x2_ASAP7_75t_L g1342 ( 
.A(n_1234),
.B(n_1205),
.Y(n_1342)
);

INVx8_ASAP7_75t_L g1343 ( 
.A(n_1243),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1261),
.Y(n_1344)
);

AND2x2_ASAP7_75t_L g1345 ( 
.A(n_1247),
.B(n_1187),
.Y(n_1345)
);

AND2x2_ASAP7_75t_L g1346 ( 
.A(n_1247),
.B(n_1189),
.Y(n_1346)
);

INVx2_ASAP7_75t_L g1347 ( 
.A(n_1274),
.Y(n_1347)
);

AO31x2_ASAP7_75t_L g1348 ( 
.A1(n_1242),
.A2(n_1189),
.A3(n_1204),
.B(n_1185),
.Y(n_1348)
);

NOR2xp33_ASAP7_75t_R g1349 ( 
.A(n_1253),
.B(n_95),
.Y(n_1349)
);

AO32x2_ASAP7_75t_L g1350 ( 
.A1(n_1286),
.A2(n_1185),
.A3(n_1207),
.B1(n_1204),
.B2(n_44),
.Y(n_1350)
);

AND2x2_ASAP7_75t_L g1351 ( 
.A(n_1225),
.B(n_44),
.Y(n_1351)
);

AO31x2_ASAP7_75t_L g1352 ( 
.A1(n_1289),
.A2(n_47),
.A3(n_48),
.B(n_97),
.Y(n_1352)
);

NAND2xp33_ASAP7_75t_R g1353 ( 
.A(n_1240),
.B(n_98),
.Y(n_1353)
);

AND3x1_ASAP7_75t_L g1354 ( 
.A(n_1282),
.B(n_1235),
.C(n_1267),
.Y(n_1354)
);

AND2x2_ASAP7_75t_L g1355 ( 
.A(n_1243),
.B(n_1241),
.Y(n_1355)
);

NAND2xp33_ASAP7_75t_R g1356 ( 
.A(n_1288),
.B(n_99),
.Y(n_1356)
);

NOR2xp33_ASAP7_75t_R g1357 ( 
.A(n_1280),
.B(n_101),
.Y(n_1357)
);

O2A1O1Ixp33_ASAP7_75t_SL g1358 ( 
.A1(n_1244),
.A2(n_104),
.B(n_105),
.C(n_106),
.Y(n_1358)
);

OAI21xp5_ASAP7_75t_L g1359 ( 
.A1(n_1268),
.A2(n_108),
.B(n_113),
.Y(n_1359)
);

BUFx12f_ASAP7_75t_L g1360 ( 
.A(n_1285),
.Y(n_1360)
);

AND2x2_ASAP7_75t_L g1361 ( 
.A(n_1280),
.B(n_116),
.Y(n_1361)
);

BUFx3_ASAP7_75t_L g1362 ( 
.A(n_1275),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1231),
.Y(n_1363)
);

INVx2_ASAP7_75t_L g1364 ( 
.A(n_1291),
.Y(n_1364)
);

AND2x2_ASAP7_75t_L g1365 ( 
.A(n_1342),
.B(n_1270),
.Y(n_1365)
);

INVx2_ASAP7_75t_L g1366 ( 
.A(n_1291),
.Y(n_1366)
);

NAND2xp5_ASAP7_75t_L g1367 ( 
.A(n_1298),
.B(n_1226),
.Y(n_1367)
);

INVx2_ASAP7_75t_R g1368 ( 
.A(n_1363),
.Y(n_1368)
);

AND2x2_ASAP7_75t_L g1369 ( 
.A(n_1328),
.B(n_1270),
.Y(n_1369)
);

AND2x2_ASAP7_75t_L g1370 ( 
.A(n_1339),
.B(n_1275),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1304),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1305),
.Y(n_1372)
);

OAI321xp33_ASAP7_75t_L g1373 ( 
.A1(n_1308),
.A2(n_1244),
.A3(n_1226),
.B1(n_1271),
.B2(n_1250),
.C(n_1266),
.Y(n_1373)
);

AND2x2_ASAP7_75t_L g1374 ( 
.A(n_1313),
.B(n_1250),
.Y(n_1374)
);

INVx3_ASAP7_75t_L g1375 ( 
.A(n_1292),
.Y(n_1375)
);

INVx2_ASAP7_75t_L g1376 ( 
.A(n_1292),
.Y(n_1376)
);

INVx3_ASAP7_75t_L g1377 ( 
.A(n_1330),
.Y(n_1377)
);

INVx2_ASAP7_75t_L g1378 ( 
.A(n_1344),
.Y(n_1378)
);

AND2x2_ASAP7_75t_L g1379 ( 
.A(n_1323),
.B(n_1271),
.Y(n_1379)
);

OR2x2_ASAP7_75t_L g1380 ( 
.A(n_1320),
.B(n_1245),
.Y(n_1380)
);

BUFx2_ASAP7_75t_L g1381 ( 
.A(n_1333),
.Y(n_1381)
);

AND2x2_ASAP7_75t_L g1382 ( 
.A(n_1324),
.B(n_1355),
.Y(n_1382)
);

INVx1_ASAP7_75t_SL g1383 ( 
.A(n_1310),
.Y(n_1383)
);

AND2x4_ASAP7_75t_L g1384 ( 
.A(n_1330),
.B(n_1238),
.Y(n_1384)
);

AND2x2_ASAP7_75t_L g1385 ( 
.A(n_1325),
.B(n_117),
.Y(n_1385)
);

AND2x2_ASAP7_75t_L g1386 ( 
.A(n_1346),
.B(n_118),
.Y(n_1386)
);

OR2x2_ASAP7_75t_L g1387 ( 
.A(n_1321),
.B(n_1283),
.Y(n_1387)
);

AND2x2_ASAP7_75t_L g1388 ( 
.A(n_1352),
.B(n_122),
.Y(n_1388)
);

AND2x2_ASAP7_75t_L g1389 ( 
.A(n_1352),
.B(n_123),
.Y(n_1389)
);

INVx2_ASAP7_75t_L g1390 ( 
.A(n_1347),
.Y(n_1390)
);

AND2x2_ASAP7_75t_L g1391 ( 
.A(n_1352),
.B(n_125),
.Y(n_1391)
);

OR2x6_ASAP7_75t_L g1392 ( 
.A(n_1334),
.B(n_1279),
.Y(n_1392)
);

AND2x2_ASAP7_75t_L g1393 ( 
.A(n_1294),
.B(n_128),
.Y(n_1393)
);

AOI22xp5_ASAP7_75t_L g1394 ( 
.A1(n_1307),
.A2(n_1256),
.B1(n_139),
.B2(n_140),
.Y(n_1394)
);

INVxp33_ASAP7_75t_L g1395 ( 
.A(n_1306),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1337),
.Y(n_1396)
);

AND2x4_ASAP7_75t_L g1397 ( 
.A(n_1293),
.B(n_136),
.Y(n_1397)
);

HB1xp67_ASAP7_75t_L g1398 ( 
.A(n_1296),
.Y(n_1398)
);

AND2x4_ASAP7_75t_L g1399 ( 
.A(n_1334),
.B(n_141),
.Y(n_1399)
);

AND2x2_ASAP7_75t_L g1400 ( 
.A(n_1303),
.B(n_1316),
.Y(n_1400)
);

OR2x2_ASAP7_75t_L g1401 ( 
.A(n_1300),
.B(n_144),
.Y(n_1401)
);

INVxp67_ASAP7_75t_SL g1402 ( 
.A(n_1338),
.Y(n_1402)
);

BUFx2_ASAP7_75t_L g1403 ( 
.A(n_1302),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1363),
.Y(n_1404)
);

OA21x2_ASAP7_75t_L g1405 ( 
.A1(n_1336),
.A2(n_154),
.B(n_158),
.Y(n_1405)
);

AND2x2_ASAP7_75t_L g1406 ( 
.A(n_1351),
.B(n_366),
.Y(n_1406)
);

INVx2_ASAP7_75t_L g1407 ( 
.A(n_1348),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1350),
.Y(n_1408)
);

AND2x2_ASAP7_75t_L g1409 ( 
.A(n_1350),
.B(n_160),
.Y(n_1409)
);

INVx2_ASAP7_75t_L g1410 ( 
.A(n_1348),
.Y(n_1410)
);

AND2x2_ASAP7_75t_L g1411 ( 
.A(n_1350),
.B(n_361),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1329),
.Y(n_1412)
);

AND2x2_ASAP7_75t_L g1413 ( 
.A(n_1315),
.B(n_163),
.Y(n_1413)
);

INVx2_ASAP7_75t_L g1414 ( 
.A(n_1348),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1362),
.Y(n_1415)
);

AOI22xp33_ASAP7_75t_SL g1416 ( 
.A1(n_1359),
.A2(n_164),
.B1(n_165),
.B2(n_166),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1354),
.Y(n_1417)
);

BUFx6f_ASAP7_75t_L g1418 ( 
.A(n_1360),
.Y(n_1418)
);

INVx2_ASAP7_75t_L g1419 ( 
.A(n_1361),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1335),
.Y(n_1420)
);

AND2x2_ASAP7_75t_L g1421 ( 
.A(n_1314),
.B(n_167),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_L g1422 ( 
.A(n_1332),
.B(n_1345),
.Y(n_1422)
);

OR2x2_ASAP7_75t_L g1423 ( 
.A(n_1327),
.B(n_357),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1343),
.Y(n_1424)
);

INVx2_ASAP7_75t_L g1425 ( 
.A(n_1343),
.Y(n_1425)
);

NAND2x1_ASAP7_75t_L g1426 ( 
.A(n_1322),
.B(n_172),
.Y(n_1426)
);

INVx2_ASAP7_75t_L g1427 ( 
.A(n_1319),
.Y(n_1427)
);

AOI22xp33_ASAP7_75t_L g1428 ( 
.A1(n_1357),
.A2(n_173),
.B1(n_174),
.B2(n_175),
.Y(n_1428)
);

INVxp33_ASAP7_75t_L g1429 ( 
.A(n_1341),
.Y(n_1429)
);

AND2x2_ASAP7_75t_L g1430 ( 
.A(n_1318),
.B(n_181),
.Y(n_1430)
);

INVx2_ASAP7_75t_L g1431 ( 
.A(n_1322),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1358),
.Y(n_1432)
);

INVx2_ASAP7_75t_L g1433 ( 
.A(n_1331),
.Y(n_1433)
);

OR2x2_ASAP7_75t_L g1434 ( 
.A(n_1340),
.B(n_356),
.Y(n_1434)
);

AND2x2_ASAP7_75t_L g1435 ( 
.A(n_1400),
.B(n_1312),
.Y(n_1435)
);

OR2x2_ASAP7_75t_L g1436 ( 
.A(n_1365),
.B(n_1312),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1364),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_L g1438 ( 
.A(n_1402),
.B(n_1349),
.Y(n_1438)
);

NAND2x1p5_ASAP7_75t_L g1439 ( 
.A(n_1405),
.B(n_1295),
.Y(n_1439)
);

INVx2_ASAP7_75t_L g1440 ( 
.A(n_1382),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1364),
.Y(n_1441)
);

INVx2_ASAP7_75t_L g1442 ( 
.A(n_1382),
.Y(n_1442)
);

AND2x2_ASAP7_75t_L g1443 ( 
.A(n_1400),
.B(n_1295),
.Y(n_1443)
);

AND2x4_ASAP7_75t_L g1444 ( 
.A(n_1366),
.B(n_1295),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1366),
.Y(n_1445)
);

AND2x2_ASAP7_75t_L g1446 ( 
.A(n_1386),
.B(n_1299),
.Y(n_1446)
);

NAND2xp5_ASAP7_75t_L g1447 ( 
.A(n_1369),
.B(n_1326),
.Y(n_1447)
);

AND2x4_ASAP7_75t_L g1448 ( 
.A(n_1375),
.B(n_1297),
.Y(n_1448)
);

AOI221xp5_ASAP7_75t_L g1449 ( 
.A1(n_1409),
.A2(n_1353),
.B1(n_1317),
.B2(n_1311),
.C(n_1356),
.Y(n_1449)
);

AND2x2_ASAP7_75t_L g1450 ( 
.A(n_1386),
.B(n_1422),
.Y(n_1450)
);

NAND2xp5_ASAP7_75t_L g1451 ( 
.A(n_1369),
.B(n_1290),
.Y(n_1451)
);

INVx2_ASAP7_75t_SL g1452 ( 
.A(n_1433),
.Y(n_1452)
);

AOI21xp5_ASAP7_75t_L g1453 ( 
.A1(n_1405),
.A2(n_1309),
.B(n_1301),
.Y(n_1453)
);

BUFx2_ASAP7_75t_L g1454 ( 
.A(n_1403),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1371),
.Y(n_1455)
);

INVxp67_ASAP7_75t_SL g1456 ( 
.A(n_1412),
.Y(n_1456)
);

NAND2xp5_ASAP7_75t_L g1457 ( 
.A(n_1396),
.B(n_183),
.Y(n_1457)
);

AND2x2_ASAP7_75t_L g1458 ( 
.A(n_1365),
.B(n_351),
.Y(n_1458)
);

INVx2_ASAP7_75t_L g1459 ( 
.A(n_1378),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_L g1460 ( 
.A(n_1372),
.B(n_184),
.Y(n_1460)
);

INVx2_ASAP7_75t_L g1461 ( 
.A(n_1378),
.Y(n_1461)
);

NAND2xp5_ASAP7_75t_L g1462 ( 
.A(n_1376),
.B(n_185),
.Y(n_1462)
);

AND2x4_ASAP7_75t_SL g1463 ( 
.A(n_1433),
.B(n_187),
.Y(n_1463)
);

HB1xp67_ASAP7_75t_L g1464 ( 
.A(n_1383),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1404),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1376),
.Y(n_1466)
);

NAND2xp5_ASAP7_75t_L g1467 ( 
.A(n_1408),
.B(n_190),
.Y(n_1467)
);

HB1xp67_ASAP7_75t_L g1468 ( 
.A(n_1398),
.Y(n_1468)
);

AND2x2_ASAP7_75t_L g1469 ( 
.A(n_1417),
.B(n_191),
.Y(n_1469)
);

AND2x4_ASAP7_75t_L g1470 ( 
.A(n_1375),
.B(n_350),
.Y(n_1470)
);

AND2x2_ASAP7_75t_L g1471 ( 
.A(n_1370),
.B(n_194),
.Y(n_1471)
);

INVxp33_ASAP7_75t_L g1472 ( 
.A(n_1381),
.Y(n_1472)
);

NAND2xp5_ASAP7_75t_L g1473 ( 
.A(n_1367),
.B(n_1375),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1390),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1390),
.Y(n_1475)
);

AND2x4_ASAP7_75t_L g1476 ( 
.A(n_1392),
.B(n_347),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_L g1477 ( 
.A(n_1409),
.B(n_196),
.Y(n_1477)
);

OR2x2_ASAP7_75t_L g1478 ( 
.A(n_1380),
.B(n_197),
.Y(n_1478)
);

AND2x2_ASAP7_75t_L g1479 ( 
.A(n_1370),
.B(n_200),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1407),
.Y(n_1480)
);

AND2x2_ASAP7_75t_L g1481 ( 
.A(n_1419),
.B(n_346),
.Y(n_1481)
);

INVxp67_ASAP7_75t_SL g1482 ( 
.A(n_1387),
.Y(n_1482)
);

AND2x2_ASAP7_75t_L g1483 ( 
.A(n_1419),
.B(n_203),
.Y(n_1483)
);

NAND2xp5_ASAP7_75t_L g1484 ( 
.A(n_1411),
.B(n_204),
.Y(n_1484)
);

OR2x2_ASAP7_75t_L g1485 ( 
.A(n_1401),
.B(n_216),
.Y(n_1485)
);

INVx3_ASAP7_75t_L g1486 ( 
.A(n_1377),
.Y(n_1486)
);

AND2x4_ASAP7_75t_SL g1487 ( 
.A(n_1418),
.B(n_218),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_L g1488 ( 
.A(n_1411),
.B(n_220),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1407),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1410),
.Y(n_1490)
);

BUFx3_ASAP7_75t_L g1491 ( 
.A(n_1427),
.Y(n_1491)
);

INVx3_ASAP7_75t_L g1492 ( 
.A(n_1377),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1410),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1455),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_1468),
.B(n_1385),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1465),
.Y(n_1496)
);

INVx4_ASAP7_75t_L g1497 ( 
.A(n_1476),
.Y(n_1497)
);

AND2x2_ASAP7_75t_L g1498 ( 
.A(n_1450),
.B(n_1427),
.Y(n_1498)
);

HB1xp67_ASAP7_75t_L g1499 ( 
.A(n_1456),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1440),
.B(n_1392),
.Y(n_1500)
);

INVx2_ASAP7_75t_L g1501 ( 
.A(n_1459),
.Y(n_1501)
);

OR2x2_ASAP7_75t_L g1502 ( 
.A(n_1482),
.B(n_1473),
.Y(n_1502)
);

AND2x2_ASAP7_75t_L g1503 ( 
.A(n_1442),
.B(n_1368),
.Y(n_1503)
);

NAND2x1p5_ASAP7_75t_L g1504 ( 
.A(n_1453),
.B(n_1405),
.Y(n_1504)
);

AND2x2_ASAP7_75t_L g1505 ( 
.A(n_1464),
.B(n_1392),
.Y(n_1505)
);

NOR2x1_ASAP7_75t_L g1506 ( 
.A(n_1447),
.B(n_1438),
.Y(n_1506)
);

AND2x4_ASAP7_75t_SL g1507 ( 
.A(n_1448),
.B(n_1392),
.Y(n_1507)
);

AND2x4_ASAP7_75t_L g1508 ( 
.A(n_1436),
.B(n_1415),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_SL g1509 ( 
.A(n_1453),
.B(n_1387),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1437),
.Y(n_1510)
);

AND2x2_ASAP7_75t_L g1511 ( 
.A(n_1435),
.B(n_1406),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_L g1512 ( 
.A(n_1473),
.B(n_1385),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1441),
.Y(n_1513)
);

AND2x4_ASAP7_75t_L g1514 ( 
.A(n_1461),
.B(n_1420),
.Y(n_1514)
);

INVx2_ASAP7_75t_L g1515 ( 
.A(n_1445),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1466),
.Y(n_1516)
);

AND2x2_ASAP7_75t_L g1517 ( 
.A(n_1454),
.B(n_1406),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1474),
.Y(n_1518)
);

INVx4_ASAP7_75t_L g1519 ( 
.A(n_1476),
.Y(n_1519)
);

INVx3_ASAP7_75t_L g1520 ( 
.A(n_1444),
.Y(n_1520)
);

NOR2xp33_ASAP7_75t_L g1521 ( 
.A(n_1451),
.B(n_1423),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1443),
.B(n_1374),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_L g1523 ( 
.A(n_1451),
.B(n_1374),
.Y(n_1523)
);

AND2x2_ASAP7_75t_L g1524 ( 
.A(n_1472),
.B(n_1491),
.Y(n_1524)
);

OR2x2_ASAP7_75t_L g1525 ( 
.A(n_1447),
.B(n_1368),
.Y(n_1525)
);

AND2x4_ASAP7_75t_L g1526 ( 
.A(n_1486),
.B(n_1414),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1475),
.Y(n_1527)
);

OR2x2_ASAP7_75t_L g1528 ( 
.A(n_1452),
.B(n_1480),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1456),
.Y(n_1529)
);

INVx2_ASAP7_75t_L g1530 ( 
.A(n_1489),
.Y(n_1530)
);

INVx3_ASAP7_75t_L g1531 ( 
.A(n_1444),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1490),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1496),
.Y(n_1533)
);

INVx2_ASAP7_75t_L g1534 ( 
.A(n_1515),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1494),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1515),
.Y(n_1536)
);

OAI32xp33_ASAP7_75t_L g1537 ( 
.A1(n_1504),
.A2(n_1423),
.A3(n_1488),
.B1(n_1477),
.B2(n_1484),
.Y(n_1537)
);

HB1xp67_ASAP7_75t_L g1538 ( 
.A(n_1499),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1510),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1513),
.Y(n_1540)
);

AOI22xp5_ASAP7_75t_L g1541 ( 
.A1(n_1506),
.A2(n_1449),
.B1(n_1413),
.B2(n_1438),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_L g1542 ( 
.A(n_1523),
.B(n_1486),
.Y(n_1542)
);

AND2x2_ASAP7_75t_L g1543 ( 
.A(n_1505),
.B(n_1524),
.Y(n_1543)
);

NAND2x2_ASAP7_75t_L g1544 ( 
.A(n_1495),
.B(n_1485),
.Y(n_1544)
);

NAND2x1p5_ASAP7_75t_L g1545 ( 
.A(n_1497),
.B(n_1492),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1530),
.Y(n_1546)
);

NAND4xp75_ASAP7_75t_L g1547 ( 
.A(n_1509),
.B(n_1449),
.C(n_1413),
.D(n_1488),
.Y(n_1547)
);

OAI322xp33_ASAP7_75t_L g1548 ( 
.A1(n_1521),
.A2(n_1484),
.A3(n_1477),
.B1(n_1467),
.B2(n_1457),
.C1(n_1401),
.C2(n_1460),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1516),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1518),
.Y(n_1550)
);

OR2x2_ASAP7_75t_L g1551 ( 
.A(n_1502),
.B(n_1493),
.Y(n_1551)
);

OR2x2_ASAP7_75t_L g1552 ( 
.A(n_1525),
.B(n_1414),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1527),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1512),
.B(n_1492),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1501),
.Y(n_1555)
);

HB1xp67_ASAP7_75t_L g1556 ( 
.A(n_1499),
.Y(n_1556)
);

AND2x4_ASAP7_75t_L g1557 ( 
.A(n_1520),
.B(n_1448),
.Y(n_1557)
);

INVx2_ASAP7_75t_SL g1558 ( 
.A(n_1508),
.Y(n_1558)
);

AOI32xp33_ASAP7_75t_L g1559 ( 
.A1(n_1521),
.A2(n_1469),
.A3(n_1421),
.B1(n_1416),
.B2(n_1429),
.Y(n_1559)
);

INVx2_ASAP7_75t_SL g1560 ( 
.A(n_1543),
.Y(n_1560)
);

INVx2_ASAP7_75t_L g1561 ( 
.A(n_1534),
.Y(n_1561)
);

AOI22xp5_ASAP7_75t_L g1562 ( 
.A1(n_1547),
.A2(n_1509),
.B1(n_1497),
.B2(n_1519),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1557),
.B(n_1508),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1539),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1540),
.Y(n_1565)
);

INVxp67_ASAP7_75t_SL g1566 ( 
.A(n_1538),
.Y(n_1566)
);

INVx1_ASAP7_75t_SL g1567 ( 
.A(n_1557),
.Y(n_1567)
);

XOR2x2_ASAP7_75t_L g1568 ( 
.A(n_1541),
.B(n_1446),
.Y(n_1568)
);

NAND2xp5_ASAP7_75t_L g1569 ( 
.A(n_1556),
.B(n_1529),
.Y(n_1569)
);

NOR3xp33_ASAP7_75t_L g1570 ( 
.A(n_1548),
.B(n_1457),
.C(n_1467),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1549),
.Y(n_1571)
);

AND2x2_ASAP7_75t_L g1572 ( 
.A(n_1558),
.B(n_1508),
.Y(n_1572)
);

AOI211xp5_ASAP7_75t_L g1573 ( 
.A1(n_1537),
.A2(n_1430),
.B(n_1517),
.C(n_1429),
.Y(n_1573)
);

AND2x2_ASAP7_75t_L g1574 ( 
.A(n_1545),
.B(n_1522),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1550),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1553),
.Y(n_1576)
);

OR2x2_ASAP7_75t_L g1577 ( 
.A(n_1542),
.B(n_1554),
.Y(n_1577)
);

INVx2_ASAP7_75t_L g1578 ( 
.A(n_1546),
.Y(n_1578)
);

OAI221xp5_ASAP7_75t_L g1579 ( 
.A1(n_1559),
.A2(n_1504),
.B1(n_1394),
.B2(n_1428),
.C(n_1439),
.Y(n_1579)
);

NOR3xp33_ASAP7_75t_L g1580 ( 
.A(n_1537),
.B(n_1460),
.C(n_1430),
.Y(n_1580)
);

OAI221xp5_ASAP7_75t_L g1581 ( 
.A1(n_1544),
.A2(n_1439),
.B1(n_1421),
.B2(n_1519),
.C(n_1497),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1570),
.B(n_1533),
.Y(n_1582)
);

NOR2xp33_ASAP7_75t_L g1583 ( 
.A(n_1581),
.B(n_1511),
.Y(n_1583)
);

OAI211xp5_ASAP7_75t_SL g1584 ( 
.A1(n_1573),
.A2(n_1535),
.B(n_1555),
.C(n_1551),
.Y(n_1584)
);

NAND3xp33_ASAP7_75t_L g1585 ( 
.A(n_1580),
.B(n_1389),
.C(n_1391),
.Y(n_1585)
);

NOR3xp33_ASAP7_75t_SL g1586 ( 
.A(n_1581),
.B(n_1579),
.C(n_1566),
.Y(n_1586)
);

OAI221xp5_ASAP7_75t_L g1587 ( 
.A1(n_1580),
.A2(n_1519),
.B1(n_1552),
.B2(n_1536),
.C(n_1531),
.Y(n_1587)
);

OAI22xp5_ASAP7_75t_L g1588 ( 
.A1(n_1579),
.A2(n_1507),
.B1(n_1531),
.B2(n_1520),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_L g1589 ( 
.A(n_1570),
.B(n_1498),
.Y(n_1589)
);

AND2x2_ASAP7_75t_L g1590 ( 
.A(n_1563),
.B(n_1520),
.Y(n_1590)
);

OR2x2_ASAP7_75t_L g1591 ( 
.A(n_1577),
.B(n_1528),
.Y(n_1591)
);

INVxp67_ASAP7_75t_SL g1592 ( 
.A(n_1562),
.Y(n_1592)
);

OAI21xp5_ASAP7_75t_SL g1593 ( 
.A1(n_1568),
.A2(n_1463),
.B(n_1507),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1564),
.Y(n_1594)
);

XOR2x2_ASAP7_75t_L g1595 ( 
.A(n_1560),
.B(n_1399),
.Y(n_1595)
);

OAI22xp33_ASAP7_75t_L g1596 ( 
.A1(n_1567),
.A2(n_1531),
.B1(n_1478),
.B2(n_1546),
.Y(n_1596)
);

AOI332xp33_ASAP7_75t_L g1597 ( 
.A1(n_1565),
.A2(n_1532),
.A3(n_1501),
.B1(n_1530),
.B2(n_1514),
.B3(n_1503),
.C1(n_1500),
.C2(n_1424),
.Y(n_1597)
);

NOR4xp25_ASAP7_75t_SL g1598 ( 
.A(n_1571),
.B(n_1373),
.C(n_1432),
.D(n_1514),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1575),
.Y(n_1599)
);

XNOR2xp5_ASAP7_75t_L g1600 ( 
.A(n_1574),
.B(n_1395),
.Y(n_1600)
);

AND2x2_ASAP7_75t_L g1601 ( 
.A(n_1572),
.B(n_1514),
.Y(n_1601)
);

INVxp67_ASAP7_75t_L g1602 ( 
.A(n_1576),
.Y(n_1602)
);

NOR2xp33_ASAP7_75t_SL g1603 ( 
.A(n_1585),
.B(n_1418),
.Y(n_1603)
);

NOR2xp67_ASAP7_75t_SL g1604 ( 
.A(n_1585),
.B(n_1418),
.Y(n_1604)
);

AOI211xp5_ASAP7_75t_L g1605 ( 
.A1(n_1592),
.A2(n_1391),
.B(n_1389),
.C(n_1388),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_L g1606 ( 
.A(n_1582),
.B(n_1569),
.Y(n_1606)
);

AOI221x1_ASAP7_75t_L g1607 ( 
.A1(n_1584),
.A2(n_1569),
.B1(n_1561),
.B2(n_1578),
.C(n_1462),
.Y(n_1607)
);

HB1xp67_ASAP7_75t_L g1608 ( 
.A(n_1602),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1594),
.Y(n_1609)
);

AOI21xp5_ASAP7_75t_L g1610 ( 
.A1(n_1593),
.A2(n_1395),
.B(n_1399),
.Y(n_1610)
);

AND2x2_ASAP7_75t_L g1611 ( 
.A(n_1590),
.B(n_1503),
.Y(n_1611)
);

NOR2xp33_ASAP7_75t_L g1612 ( 
.A(n_1600),
.B(n_1418),
.Y(n_1612)
);

NOR3x1_ASAP7_75t_L g1613 ( 
.A(n_1588),
.B(n_1587),
.C(n_1589),
.Y(n_1613)
);

NAND3xp33_ASAP7_75t_L g1614 ( 
.A(n_1586),
.B(n_1598),
.C(n_1599),
.Y(n_1614)
);

NOR2x1_ASAP7_75t_L g1615 ( 
.A(n_1583),
.B(n_1399),
.Y(n_1615)
);

O2A1O1Ixp33_ASAP7_75t_L g1616 ( 
.A1(n_1614),
.A2(n_1596),
.B(n_1388),
.C(n_1434),
.Y(n_1616)
);

NOR3xp33_ASAP7_75t_SL g1617 ( 
.A(n_1612),
.B(n_1462),
.C(n_1597),
.Y(n_1617)
);

INVxp33_ASAP7_75t_L g1618 ( 
.A(n_1615),
.Y(n_1618)
);

XNOR2x1_ASAP7_75t_L g1619 ( 
.A(n_1608),
.B(n_1595),
.Y(n_1619)
);

OR3x1_ASAP7_75t_L g1620 ( 
.A(n_1609),
.B(n_1487),
.C(n_1591),
.Y(n_1620)
);

AOI22xp33_ASAP7_75t_L g1621 ( 
.A1(n_1604),
.A2(n_1601),
.B1(n_1458),
.B2(n_1431),
.Y(n_1621)
);

AOI211xp5_ASAP7_75t_L g1622 ( 
.A1(n_1603),
.A2(n_1471),
.B(n_1479),
.C(n_1431),
.Y(n_1622)
);

AOI21xp5_ASAP7_75t_L g1623 ( 
.A1(n_1606),
.A2(n_1426),
.B(n_1425),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_L g1624 ( 
.A(n_1607),
.B(n_1425),
.Y(n_1624)
);

AND2x2_ASAP7_75t_L g1625 ( 
.A(n_1618),
.B(n_1613),
.Y(n_1625)
);

NOR2xp33_ASAP7_75t_L g1626 ( 
.A(n_1619),
.B(n_1610),
.Y(n_1626)
);

AOI221x1_ASAP7_75t_L g1627 ( 
.A1(n_1623),
.A2(n_1611),
.B1(n_1470),
.B2(n_1483),
.C(n_1481),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1624),
.Y(n_1628)
);

AOI22xp5_ASAP7_75t_L g1629 ( 
.A1(n_1620),
.A2(n_1605),
.B1(n_1526),
.B2(n_1470),
.Y(n_1629)
);

NAND3xp33_ASAP7_75t_L g1630 ( 
.A(n_1616),
.B(n_1434),
.C(n_1379),
.Y(n_1630)
);

NOR3xp33_ASAP7_75t_L g1631 ( 
.A(n_1622),
.B(n_1393),
.C(n_1397),
.Y(n_1631)
);

XNOR2xp5_ASAP7_75t_L g1632 ( 
.A(n_1617),
.B(n_1393),
.Y(n_1632)
);

OAI221xp5_ASAP7_75t_L g1633 ( 
.A1(n_1621),
.A2(n_1377),
.B1(n_1379),
.B2(n_1397),
.C(n_231),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1628),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_L g1635 ( 
.A(n_1625),
.B(n_1626),
.Y(n_1635)
);

AND2x2_ASAP7_75t_L g1636 ( 
.A(n_1632),
.B(n_1526),
.Y(n_1636)
);

AND3x4_ASAP7_75t_L g1637 ( 
.A(n_1631),
.B(n_1397),
.C(n_1526),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1630),
.Y(n_1638)
);

INVx3_ASAP7_75t_L g1639 ( 
.A(n_1627),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1629),
.Y(n_1640)
);

INVxp33_ASAP7_75t_SL g1641 ( 
.A(n_1635),
.Y(n_1641)
);

OAI22xp5_ASAP7_75t_L g1642 ( 
.A1(n_1639),
.A2(n_1633),
.B1(n_1384),
.B2(n_227),
.Y(n_1642)
);

NAND4xp25_ASAP7_75t_L g1643 ( 
.A(n_1640),
.B(n_1384),
.C(n_225),
.D(n_240),
.Y(n_1643)
);

OAI22xp5_ASAP7_75t_L g1644 ( 
.A1(n_1639),
.A2(n_1384),
.B1(n_246),
.B2(n_248),
.Y(n_1644)
);

XOR2x1_ASAP7_75t_L g1645 ( 
.A(n_1644),
.B(n_1634),
.Y(n_1645)
);

NOR2xp33_ASAP7_75t_L g1646 ( 
.A(n_1641),
.B(n_1638),
.Y(n_1646)
);

INVx1_ASAP7_75t_SL g1647 ( 
.A(n_1642),
.Y(n_1647)
);

OAI22xp33_ASAP7_75t_L g1648 ( 
.A1(n_1643),
.A2(n_1636),
.B1(n_1637),
.B2(n_251),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1646),
.Y(n_1649)
);

OAI22xp5_ASAP7_75t_L g1650 ( 
.A1(n_1647),
.A2(n_223),
.B1(n_249),
.B2(n_252),
.Y(n_1650)
);

AOI22xp33_ASAP7_75t_L g1651 ( 
.A1(n_1648),
.A2(n_255),
.B1(n_257),
.B2(n_258),
.Y(n_1651)
);

AOI22xp33_ASAP7_75t_L g1652 ( 
.A1(n_1649),
.A2(n_1651),
.B1(n_1650),
.B2(n_1645),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1649),
.Y(n_1653)
);

OAI22xp5_ASAP7_75t_L g1654 ( 
.A1(n_1651),
.A2(n_259),
.B1(n_260),
.B2(n_261),
.Y(n_1654)
);

OAI22xp5_ASAP7_75t_L g1655 ( 
.A1(n_1652),
.A2(n_263),
.B1(n_270),
.B2(n_271),
.Y(n_1655)
);

CKINVDCx20_ASAP7_75t_R g1656 ( 
.A(n_1653),
.Y(n_1656)
);

INVx2_ASAP7_75t_SL g1657 ( 
.A(n_1654),
.Y(n_1657)
);

BUFx2_ASAP7_75t_L g1658 ( 
.A(n_1653),
.Y(n_1658)
);

OAI221xp5_ASAP7_75t_L g1659 ( 
.A1(n_1658),
.A2(n_275),
.B1(n_278),
.B2(n_279),
.C(n_280),
.Y(n_1659)
);

AOI22xp33_ASAP7_75t_L g1660 ( 
.A1(n_1656),
.A2(n_281),
.B1(n_282),
.B2(n_283),
.Y(n_1660)
);

O2A1O1Ixp33_ASAP7_75t_L g1661 ( 
.A1(n_1655),
.A2(n_285),
.B(n_287),
.C(n_289),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1657),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1658),
.Y(n_1663)
);

OAI21xp5_ASAP7_75t_L g1664 ( 
.A1(n_1663),
.A2(n_292),
.B(n_295),
.Y(n_1664)
);

AOI21xp5_ASAP7_75t_L g1665 ( 
.A1(n_1662),
.A2(n_300),
.B(n_303),
.Y(n_1665)
);

XNOR2x1_ASAP7_75t_L g1666 ( 
.A(n_1661),
.B(n_1659),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_L g1667 ( 
.A(n_1660),
.B(n_308),
.Y(n_1667)
);

AOI21xp5_ASAP7_75t_L g1668 ( 
.A1(n_1663),
.A2(n_310),
.B(n_311),
.Y(n_1668)
);

AOI22xp5_ASAP7_75t_SL g1669 ( 
.A1(n_1665),
.A2(n_314),
.B1(n_315),
.B2(n_316),
.Y(n_1669)
);

AOI21x1_ASAP7_75t_L g1670 ( 
.A1(n_1668),
.A2(n_317),
.B(n_323),
.Y(n_1670)
);

AOI22xp5_ASAP7_75t_L g1671 ( 
.A1(n_1667),
.A2(n_326),
.B1(n_327),
.B2(n_335),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1669),
.B(n_1666),
.Y(n_1672)
);

AOI22xp33_ASAP7_75t_L g1673 ( 
.A1(n_1672),
.A2(n_1664),
.B1(n_1671),
.B2(n_1670),
.Y(n_1673)
);


endmodule