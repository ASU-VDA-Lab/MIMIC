module fake_jpeg_26745_n_131 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_131);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_131;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx13_ASAP7_75t_L g13 ( 
.A(n_11),
.Y(n_13)
);

BUFx3_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

INVx4_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_5),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_11),
.Y(n_24)
);

INVx2_ASAP7_75t_SL g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_25),
.B(n_0),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_28),
.B(n_25),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_27),
.Y(n_29)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_14),
.B(n_0),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_30),
.B(n_14),
.Y(n_41)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_31),
.B(n_36),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_32),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_35),
.Y(n_39)
);

CKINVDCx16_ASAP7_75t_R g36 ( 
.A(n_25),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_43),
.Y(n_51)
);

XOR2xp5_ASAP7_75t_L g62 ( 
.A(n_41),
.B(n_17),
.Y(n_62)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_30),
.B(n_14),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_31),
.A2(n_27),
.B1(n_25),
.B2(n_13),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_44),
.A2(n_17),
.B1(n_15),
.B2(n_18),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_35),
.A2(n_27),
.B1(n_13),
.B2(n_21),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_45),
.A2(n_17),
.B1(n_15),
.B2(n_23),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_36),
.A2(n_21),
.B1(n_22),
.B2(n_23),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_53),
.A2(n_58),
.B1(n_15),
.B2(n_20),
.Y(n_78)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_54),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_55),
.B(n_59),
.Y(n_66)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_57),
.Y(n_73)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_50),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_60),
.B(n_63),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_62),
.B(n_41),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_40),
.B(n_24),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_42),
.B(n_24),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_64),
.B(n_26),
.Y(n_76)
);

XOR2xp5_ASAP7_75t_L g88 ( 
.A(n_65),
.B(n_69),
.Y(n_88)
);

OAI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_56),
.A2(n_50),
.B1(n_22),
.B2(n_44),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_67),
.B(n_70),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_SL g68 ( 
.A1(n_56),
.A2(n_37),
.B(n_43),
.Y(n_68)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_68),
.A2(n_39),
.B(n_18),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_62),
.B(n_37),
.C(n_47),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_69),
.B(n_77),
.C(n_60),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_51),
.B(n_32),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_L g71 ( 
.A1(n_52),
.A2(n_61),
.B(n_58),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_L g86 ( 
.A1(n_71),
.A2(n_54),
.B(n_49),
.Y(n_86)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_61),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_75),
.B(n_76),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_52),
.B(n_33),
.C(n_39),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_78),
.B(n_26),
.Y(n_89)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_71),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_79),
.B(n_80),
.Y(n_91)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_74),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_70),
.B(n_66),
.Y(n_82)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_82),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_77),
.B(n_57),
.Y(n_84)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_84),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_72),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_85),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_86),
.A2(n_90),
.B(n_20),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_87),
.B(n_88),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_89),
.B(n_26),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_79),
.A2(n_68),
.B(n_75),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_93),
.A2(n_95),
.B(n_97),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_86),
.A2(n_65),
.B(n_78),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_81),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_98),
.B(n_80),
.Y(n_102)
);

AOI221xp5_ASAP7_75t_L g99 ( 
.A1(n_90),
.A2(n_73),
.B1(n_26),
.B2(n_19),
.C(n_10),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_99),
.B(n_9),
.Y(n_108)
);

OAI21xp33_ASAP7_75t_SL g103 ( 
.A1(n_100),
.A2(n_83),
.B(n_85),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_102),
.B(n_104),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_103),
.B(n_108),
.Y(n_112)
);

HB1xp67_ASAP7_75t_L g104 ( 
.A(n_94),
.Y(n_104)
);

OR2x2_ASAP7_75t_L g105 ( 
.A(n_91),
.B(n_83),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_105),
.B(n_106),
.Y(n_113)
);

AOI31xp67_ASAP7_75t_L g106 ( 
.A1(n_97),
.A2(n_89),
.A3(n_87),
.B(n_88),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_92),
.B(n_89),
.C(n_33),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_107),
.B(n_92),
.C(n_101),
.Y(n_111)
);

A2O1A1O1Ixp25_ASAP7_75t_L g109 ( 
.A1(n_93),
.A2(n_19),
.B(n_55),
.C(n_34),
.D(n_10),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_109),
.A2(n_98),
.B(n_96),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_111),
.B(n_113),
.C(n_112),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_114),
.B(n_116),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_110),
.A2(n_1),
.B(n_2),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_104),
.A2(n_1),
.B(n_3),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_117),
.B(n_1),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_118),
.B(n_120),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_113),
.B(n_103),
.C(n_33),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_121),
.A2(n_122),
.B(n_3),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_115),
.B(n_7),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_119),
.A2(n_8),
.B(n_12),
.Y(n_123)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_123),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_124),
.B(n_125),
.Y(n_128)
);

A2O1A1Ixp33_ASAP7_75t_L g125 ( 
.A1(n_121),
.A2(n_8),
.B(n_12),
.C(n_4),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_127),
.B(n_126),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_129),
.B(n_130),
.Y(n_131)
);

AO21x1_ASAP7_75t_L g130 ( 
.A1(n_128),
.A2(n_6),
.B(n_29),
.Y(n_130)
);


endmodule