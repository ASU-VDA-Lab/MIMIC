module fake_jpeg_1754_n_371 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_371);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_371;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_14),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

BUFx16f_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx4f_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx24_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_11),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_7),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_2),
.B(n_1),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_7),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_41),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

INVx1_ASAP7_75t_SL g95 ( 
.A(n_42),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_43),
.Y(n_98)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_44),
.Y(n_77)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_45),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_21),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_46),
.Y(n_108)
);

AND2x2_ASAP7_75t_SL g47 ( 
.A(n_17),
.B(n_0),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_47),
.B(n_48),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_35),
.B(n_1),
.Y(n_48)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_26),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_49),
.Y(n_92)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_18),
.Y(n_50)
);

HB1xp67_ASAP7_75t_L g107 ( 
.A(n_50),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_21),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_51),
.Y(n_109)
);

INVx2_ASAP7_75t_SL g52 ( 
.A(n_28),
.Y(n_52)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_52),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_15),
.B(n_2),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_53),
.B(n_67),
.Y(n_86)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_26),
.Y(n_54)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_54),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_21),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_55),
.Y(n_128)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_17),
.Y(n_56)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_56),
.Y(n_120)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_17),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_57),
.Y(n_79)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_29),
.Y(n_58)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_58),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_59),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_35),
.B(n_2),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_60),
.B(n_74),
.Y(n_85)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_16),
.Y(n_61)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_61),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_33),
.Y(n_62)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_62),
.Y(n_81)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_19),
.Y(n_63)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_63),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_26),
.Y(n_64)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_64),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_33),
.Y(n_65)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_65),
.Y(n_102)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_16),
.Y(n_66)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_66),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_15),
.B(n_13),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_33),
.Y(n_68)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_68),
.Y(n_103)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_20),
.Y(n_69)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_69),
.Y(n_124)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_29),
.Y(n_70)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_70),
.Y(n_118)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_37),
.Y(n_71)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_71),
.Y(n_111)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_37),
.Y(n_72)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_72),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_37),
.Y(n_73)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_73),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_39),
.Y(n_74)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_23),
.Y(n_75)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_75),
.Y(n_125)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_19),
.Y(n_76)
);

NAND2xp33_ASAP7_75t_SL g110 ( 
.A(n_76),
.B(n_28),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_48),
.B(n_19),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_84),
.B(n_88),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_60),
.B(n_30),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_43),
.A2(n_19),
.B1(n_46),
.B2(n_55),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_91),
.A2(n_99),
.B1(n_113),
.B2(n_127),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_42),
.B(n_40),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_94),
.B(n_96),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_42),
.B(n_40),
.Y(n_96)
);

HAxp5_ASAP7_75t_SL g97 ( 
.A(n_47),
.B(n_28),
.CON(n_97),
.SN(n_97)
);

AOI21xp33_ASAP7_75t_L g138 ( 
.A1(n_97),
.A2(n_100),
.B(n_101),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_51),
.A2(n_39),
.B1(n_34),
.B2(n_32),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_59),
.B(n_30),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_62),
.B(n_31),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_58),
.B(n_32),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_106),
.B(n_116),
.Y(n_162)
);

OR2x2_ASAP7_75t_L g174 ( 
.A(n_110),
.B(n_112),
.Y(n_174)
);

AOI21xp33_ASAP7_75t_L g112 ( 
.A1(n_52),
.A2(n_20),
.B(n_36),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_75),
.A2(n_29),
.B1(n_24),
.B2(n_36),
.Y(n_113)
);

OA22x2_ASAP7_75t_L g132 ( 
.A1(n_113),
.A2(n_119),
.B1(n_28),
.B2(n_22),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_65),
.B(n_31),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_115),
.B(n_2),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_54),
.B(n_34),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_54),
.B(n_27),
.Y(n_117)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_117),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_64),
.A2(n_29),
.B1(n_24),
.B2(n_27),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_71),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_121),
.Y(n_139)
);

NAND2xp33_ASAP7_75t_SL g126 ( 
.A(n_49),
.B(n_24),
.Y(n_126)
);

BUFx5_ASAP7_75t_L g141 ( 
.A(n_126),
.Y(n_141)
);

INVx6_ASAP7_75t_L g127 ( 
.A(n_68),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_127),
.Y(n_172)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_123),
.Y(n_129)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_129),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_85),
.A2(n_73),
.B1(n_22),
.B2(n_39),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_130),
.A2(n_135),
.B1(n_145),
.B2(n_149),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_132),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_82),
.B(n_72),
.Y(n_133)
);

MAJx2_ASAP7_75t_L g197 ( 
.A(n_133),
.B(n_152),
.C(n_156),
.Y(n_197)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_104),
.Y(n_134)
);

INVx1_ASAP7_75t_SL g206 ( 
.A(n_134),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_97),
.A2(n_72),
.B1(n_28),
.B2(n_29),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_123),
.A2(n_38),
.B1(n_25),
.B2(n_23),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_136),
.Y(n_191)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_80),
.Y(n_137)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_137),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_120),
.A2(n_38),
.B1(n_25),
.B2(n_23),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_140),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_142),
.B(n_144),
.Y(n_182)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_95),
.Y(n_143)
);

HB1xp67_ASAP7_75t_L g187 ( 
.A(n_143),
.Y(n_187)
);

OA22x2_ASAP7_75t_L g144 ( 
.A1(n_119),
.A2(n_38),
.B1(n_25),
.B2(n_5),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_86),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_120),
.A2(n_124),
.B1(n_105),
.B2(n_95),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_146),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_87),
.B(n_3),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_147),
.B(n_175),
.Y(n_193)
);

FAx1_ASAP7_75t_SL g148 ( 
.A(n_107),
.B(n_3),
.CI(n_6),
.CON(n_148),
.SN(n_148)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_148),
.B(n_165),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_L g149 ( 
.A1(n_111),
.A2(n_3),
.B1(n_6),
.B2(n_8),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_150),
.A2(n_161),
.B1(n_170),
.B2(n_171),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_L g151 ( 
.A1(n_111),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_151),
.A2(n_166),
.B1(n_160),
.B2(n_179),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_118),
.B(n_6),
.C(n_8),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_125),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_154),
.Y(n_222)
);

INVx5_ASAP7_75t_SL g155 ( 
.A(n_77),
.Y(n_155)
);

OR2x2_ASAP7_75t_L g183 ( 
.A(n_155),
.B(n_179),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_83),
.B(n_93),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_90),
.Y(n_157)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_157),
.Y(n_216)
);

INVx11_ASAP7_75t_L g158 ( 
.A(n_79),
.Y(n_158)
);

INVx8_ASAP7_75t_L g208 ( 
.A(n_158),
.Y(n_208)
);

HB1xp67_ASAP7_75t_L g159 ( 
.A(n_90),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_159),
.Y(n_203)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_78),
.Y(n_160)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_160),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_78),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_93),
.A2(n_92),
.B1(n_77),
.B2(n_79),
.Y(n_163)
);

OAI22xp33_ASAP7_75t_L g213 ( 
.A1(n_163),
.A2(n_169),
.B1(n_144),
.B2(n_158),
.Y(n_213)
);

MAJx2_ASAP7_75t_L g164 ( 
.A(n_98),
.B(n_11),
.C(n_12),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_164),
.B(n_173),
.Y(n_192)
);

FAx1_ASAP7_75t_SL g165 ( 
.A(n_122),
.B(n_12),
.CI(n_13),
.CON(n_165),
.SN(n_165)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_98),
.A2(n_128),
.B1(n_109),
.B2(n_108),
.Y(n_166)
);

AO22x1_ASAP7_75t_L g167 ( 
.A1(n_92),
.A2(n_12),
.B1(n_89),
.B2(n_79),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_167),
.B(n_177),
.Y(n_184)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_114),
.Y(n_168)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_168),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_89),
.A2(n_108),
.B1(n_109),
.B2(n_128),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_81),
.A2(n_102),
.B1(n_103),
.B2(n_114),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_81),
.A2(n_85),
.B1(n_82),
.B2(n_86),
.Y(n_171)
);

MAJx2_ASAP7_75t_L g173 ( 
.A(n_102),
.B(n_88),
.C(n_84),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_103),
.B(n_82),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_82),
.B(n_112),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_176),
.B(n_174),
.Y(n_195)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_104),
.Y(n_177)
);

INVx2_ASAP7_75t_SL g179 ( 
.A(n_123),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_142),
.B(n_176),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_181),
.B(n_186),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_174),
.A2(n_175),
.B1(n_130),
.B2(n_173),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_185),
.A2(n_199),
.B1(n_209),
.B2(n_212),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_139),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_178),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_188),
.B(n_190),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_178),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_195),
.B(n_207),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_172),
.Y(n_196)
);

CKINVDCx14_ASAP7_75t_R g255 ( 
.A(n_196),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_138),
.A2(n_135),
.B1(n_141),
.B2(n_131),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_141),
.A2(n_156),
.B(n_133),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_201),
.A2(n_221),
.B(n_192),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_147),
.B(n_164),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_204),
.B(n_219),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_162),
.B(n_153),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_166),
.A2(n_145),
.B1(n_132),
.B2(n_144),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_213),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_152),
.B(n_148),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_214),
.B(n_204),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_172),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_215),
.B(n_196),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_132),
.A2(n_144),
.B1(n_165),
.B2(n_137),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_218),
.A2(n_220),
.B1(n_201),
.B2(n_185),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_165),
.B(n_148),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_132),
.A2(n_174),
.B1(n_176),
.B2(n_175),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_167),
.A2(n_174),
.B(n_141),
.Y(n_221)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_183),
.Y(n_223)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_223),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_183),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_224),
.B(n_228),
.Y(n_267)
);

OAI22x1_ASAP7_75t_SL g225 ( 
.A1(n_189),
.A2(n_167),
.B1(n_179),
.B2(n_211),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_225),
.A2(n_246),
.B1(n_223),
.B2(n_249),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_227),
.A2(n_248),
.B(n_200),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_183),
.Y(n_228)
);

INVx13_ASAP7_75t_L g230 ( 
.A(n_208),
.Y(n_230)
);

CKINVDCx14_ASAP7_75t_R g261 ( 
.A(n_230),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_187),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_231),
.B(n_237),
.Y(n_273)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_232),
.Y(n_282)
);

INVx2_ASAP7_75t_SL g233 ( 
.A(n_210),
.Y(n_233)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_233),
.Y(n_278)
);

INVx5_ASAP7_75t_L g234 ( 
.A(n_208),
.Y(n_234)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_234),
.Y(n_288)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_210),
.Y(n_235)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_235),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_236),
.B(n_226),
.Y(n_279)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_216),
.Y(n_237)
);

O2A1O1Ixp33_ASAP7_75t_L g238 ( 
.A1(n_189),
.A2(n_221),
.B(n_219),
.C(n_217),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g259 ( 
.A1(n_238),
.A2(n_191),
.B(n_222),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_240),
.B(n_239),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_209),
.A2(n_182),
.B1(n_218),
.B2(n_211),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_241),
.A2(n_243),
.B1(n_254),
.B2(n_206),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_182),
.A2(n_220),
.B1(n_205),
.B2(n_184),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_182),
.A2(n_184),
.B1(n_193),
.B2(n_195),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_186),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_247),
.B(n_249),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_184),
.A2(n_199),
.B1(n_194),
.B2(n_198),
.Y(n_248)
);

CKINVDCx16_ASAP7_75t_R g249 ( 
.A(n_207),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_193),
.B(n_197),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_250),
.B(n_203),
.Y(n_264)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_216),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_251),
.B(n_253),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_197),
.B(n_181),
.C(n_188),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_252),
.B(n_257),
.C(n_227),
.Y(n_262)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_202),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_205),
.A2(n_214),
.B1(n_212),
.B2(n_194),
.Y(n_254)
);

HB1xp67_ASAP7_75t_L g256 ( 
.A(n_202),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_256),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_197),
.B(n_190),
.C(n_203),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_200),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_258),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_259),
.A2(n_265),
.B(n_272),
.Y(n_295)
);

NOR2xp67_ASAP7_75t_R g260 ( 
.A(n_224),
.B(n_180),
.Y(n_260)
);

OAI322xp33_ASAP7_75t_L g291 ( 
.A1(n_260),
.A2(n_244),
.A3(n_246),
.B1(n_225),
.B2(n_231),
.C1(n_235),
.C2(n_237),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_262),
.B(n_251),
.C(n_233),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_263),
.A2(n_277),
.B1(n_279),
.B2(n_284),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_SL g304 ( 
.A(n_264),
.B(n_285),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_L g265 ( 
.A1(n_238),
.A2(n_208),
.B(n_215),
.Y(n_265)
);

CKINVDCx16_ASAP7_75t_R g266 ( 
.A(n_245),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_266),
.B(n_274),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_270),
.B(n_244),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_255),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_242),
.B(n_180),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_275),
.B(n_286),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_SL g276 ( 
.A1(n_248),
.A2(n_236),
.B(n_254),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_L g290 ( 
.A1(n_276),
.A2(n_259),
.B(n_272),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_241),
.A2(n_226),
.B1(n_243),
.B2(n_229),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_229),
.A2(n_250),
.B1(n_239),
.B2(n_240),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_252),
.B(n_257),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_247),
.B(n_228),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_287),
.A2(n_269),
.B1(n_264),
.B2(n_275),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_SL g326 ( 
.A(n_290),
.B(n_302),
.Y(n_326)
);

NOR3xp33_ASAP7_75t_L g315 ( 
.A(n_291),
.B(n_283),
.C(n_278),
.Y(n_315)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_286),
.Y(n_292)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_292),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_281),
.Y(n_293)
);

AOI22xp33_ASAP7_75t_L g325 ( 
.A1(n_293),
.A2(n_297),
.B1(n_301),
.B2(n_303),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_285),
.B(n_262),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_294),
.B(n_298),
.C(n_300),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_SL g329 ( 
.A(n_296),
.B(n_309),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_281),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_262),
.B(n_233),
.C(n_253),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_283),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_L g302 ( 
.A1(n_267),
.A2(n_287),
.B(n_276),
.Y(n_302)
);

INVxp33_ASAP7_75t_L g303 ( 
.A(n_280),
.Y(n_303)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_273),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_305),
.B(n_307),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_284),
.B(n_258),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_306),
.B(n_304),
.C(n_298),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_280),
.B(n_234),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_274),
.B(n_230),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_279),
.A2(n_277),
.B1(n_267),
.B2(n_263),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_310),
.B(n_271),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_265),
.A2(n_230),
.B(n_269),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_311),
.B(n_278),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_L g321 ( 
.A1(n_312),
.A2(n_268),
.B1(n_288),
.B2(n_261),
.Y(n_321)
);

OA21x2_ASAP7_75t_SL g313 ( 
.A1(n_292),
.A2(n_282),
.B(n_260),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_294),
.B(n_273),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_314),
.B(n_327),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_315),
.B(n_295),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_317),
.B(n_324),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_320),
.A2(n_321),
.B1(n_323),
.B2(n_310),
.Y(n_332)
);

BUFx6f_ASAP7_75t_L g322 ( 
.A(n_305),
.Y(n_322)
);

HB1xp67_ASAP7_75t_L g331 ( 
.A(n_322),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_308),
.A2(n_261),
.B1(n_288),
.B2(n_312),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_293),
.B(n_297),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_299),
.B(n_300),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_328),
.B(n_330),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_299),
.B(n_289),
.Y(n_330)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_332),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_316),
.B(n_304),
.C(n_306),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_334),
.B(n_313),
.C(n_325),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_316),
.B(n_302),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_335),
.B(n_344),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_323),
.A2(n_308),
.B1(n_290),
.B2(n_289),
.Y(n_337)
);

OR2x2_ASAP7_75t_L g351 ( 
.A(n_337),
.B(n_340),
.Y(n_351)
);

OAI21xp5_ASAP7_75t_SL g338 ( 
.A1(n_324),
.A2(n_295),
.B(n_307),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_338),
.B(n_329),
.Y(n_352)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_327),
.B(n_311),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g342 ( 
.A(n_314),
.B(n_291),
.Y(n_342)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_326),
.B(n_309),
.Y(n_343)
);

XOR2xp5_ASAP7_75t_L g344 ( 
.A(n_326),
.B(n_319),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_333),
.A2(n_320),
.B1(n_318),
.B2(n_319),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_345),
.B(n_350),
.Y(n_354)
);

INVx11_ASAP7_75t_L g348 ( 
.A(n_331),
.Y(n_348)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_348),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_339),
.Y(n_350)
);

AOI31xp33_ASAP7_75t_L g357 ( 
.A1(n_352),
.A2(n_334),
.A3(n_341),
.B(n_322),
.Y(n_357)
);

OAI21xp5_ASAP7_75t_L g353 ( 
.A1(n_344),
.A2(n_329),
.B(n_318),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_353),
.B(n_336),
.Y(n_359)
);

OA21x2_ASAP7_75t_L g355 ( 
.A1(n_353),
.A2(n_343),
.B(n_342),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_355),
.B(n_356),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_346),
.B(n_335),
.C(n_336),
.Y(n_356)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_357),
.Y(n_361)
);

XOR2xp5_ASAP7_75t_L g360 ( 
.A(n_359),
.B(n_349),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_L g364 ( 
.A1(n_360),
.A2(n_351),
.B(n_354),
.Y(n_364)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_358),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_363),
.B(n_345),
.Y(n_366)
);

XOR2xp5_ASAP7_75t_L g367 ( 
.A(n_364),
.B(n_366),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_361),
.A2(n_350),
.B1(n_347),
.B2(n_351),
.Y(n_365)
);

INVxp67_ASAP7_75t_L g368 ( 
.A(n_365),
.Y(n_368)
);

INVxp67_ASAP7_75t_L g369 ( 
.A(n_367),
.Y(n_369)
);

O2A1O1Ixp33_ASAP7_75t_L g370 ( 
.A1(n_369),
.A2(n_362),
.B(n_368),
.C(n_356),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_370),
.B(n_362),
.Y(n_371)
);


endmodule