module real_jpeg_29591_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_312;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_0),
.A2(n_64),
.B1(n_65),
.B2(n_66),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_0),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_0),
.A2(n_48),
.B1(n_49),
.B2(n_66),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_0),
.A2(n_28),
.B1(n_29),
.B2(n_66),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_0),
.A2(n_34),
.B1(n_37),
.B2(n_66),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_1),
.A2(n_28),
.B1(n_29),
.B2(n_40),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_1),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_1),
.A2(n_34),
.B1(n_37),
.B2(n_40),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_1),
.A2(n_40),
.B1(n_64),
.B2(n_65),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_1),
.A2(n_40),
.B1(n_48),
.B2(n_49),
.Y(n_112)
);

INVx11_ASAP7_75t_L g90 ( 
.A(n_2),
.Y(n_90)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_2),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_3),
.A2(n_48),
.B1(n_49),
.B2(n_57),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_3),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_3),
.A2(n_57),
.B1(n_64),
.B2(n_65),
.Y(n_71)
);

OAI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_3),
.A2(n_28),
.B1(n_29),
.B2(n_57),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g132 ( 
.A1(n_3),
.A2(n_34),
.B1(n_37),
.B2(n_57),
.Y(n_132)
);

BUFx12_ASAP7_75t_L g62 ( 
.A(n_4),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_5),
.A2(n_48),
.B1(n_49),
.B2(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_5),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_5),
.A2(n_28),
.B1(n_29),
.B2(n_54),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_5),
.A2(n_54),
.B1(n_64),
.B2(n_65),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_5),
.A2(n_34),
.B1(n_37),
.B2(n_54),
.Y(n_159)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

INVx13_ASAP7_75t_L g64 ( 
.A(n_7),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_8),
.A2(n_64),
.B1(n_65),
.B2(n_168),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_8),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_8),
.A2(n_48),
.B1(n_49),
.B2(n_168),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g233 ( 
.A1(n_8),
.A2(n_28),
.B1(n_29),
.B2(n_168),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_SL g266 ( 
.A1(n_8),
.A2(n_34),
.B1(n_37),
.B2(n_168),
.Y(n_266)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_9),
.A2(n_64),
.B1(n_65),
.B2(n_141),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_9),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_9),
.A2(n_48),
.B1(n_49),
.B2(n_141),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_9),
.A2(n_28),
.B1(n_29),
.B2(n_141),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_SL g261 ( 
.A1(n_9),
.A2(n_34),
.B1(n_37),
.B2(n_141),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_10),
.A2(n_64),
.B1(n_65),
.B2(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_10),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_10),
.A2(n_48),
.B1(n_49),
.B2(n_189),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_10),
.A2(n_28),
.B1(n_29),
.B2(n_189),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_SL g274 ( 
.A1(n_10),
.A2(n_34),
.B1(n_37),
.B2(n_189),
.Y(n_274)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_12),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_12),
.B(n_60),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_12),
.B(n_48),
.Y(n_226)
);

AOI21xp33_ASAP7_75t_L g230 ( 
.A1(n_12),
.A2(n_48),
.B(n_226),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_SL g250 ( 
.A1(n_12),
.A2(n_28),
.B1(n_29),
.B2(n_187),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_12),
.A2(n_31),
.B(n_34),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_12),
.B(n_137),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_12),
.A2(n_87),
.B1(n_91),
.B2(n_274),
.Y(n_276)
);

BUFx24_ASAP7_75t_L g50 ( 
.A(n_13),
.Y(n_50)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_14),
.Y(n_47)
);

INVx11_ASAP7_75t_SL g36 ( 
.A(n_15),
.Y(n_36)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_118),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_117),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_101),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_20),
.B(n_101),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_74),
.C(n_84),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_21),
.A2(n_22),
.B1(n_74),
.B2(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_58),
.B1(n_72),
.B2(n_73),
.Y(n_22)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_23),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_41),
.B2(n_42),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_24),
.A2(n_25),
.B1(n_109),
.B2(n_110),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_24),
.B(n_42),
.C(n_58),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

AOI21xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_33),
.B(n_38),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_26),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_26),
.A2(n_96),
.B(n_97),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_26),
.A2(n_33),
.B1(n_96),
.B2(n_135),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_26),
.A2(n_38),
.B(n_97),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_26),
.A2(n_33),
.B1(n_233),
.B2(n_234),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_26),
.A2(n_79),
.B(n_234),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_26),
.A2(n_33),
.B1(n_250),
.B2(n_251),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_26),
.A2(n_33),
.B1(n_233),
.B2(n_251),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_33),
.Y(n_26)
);

OAI22xp33_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_29),
.B1(n_31),
.B2(n_32),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_28),
.A2(n_29),
.B1(n_46),
.B2(n_47),
.Y(n_51)
);

AOI32xp33_ASAP7_75t_L g224 ( 
.A1(n_28),
.A2(n_49),
.A3(n_225),
.B1(n_226),
.B2(n_227),
.Y(n_224)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NAND2xp33_ASAP7_75t_SL g227 ( 
.A(n_29),
.B(n_46),
.Y(n_227)
);

A2O1A1Ixp33_ASAP7_75t_L g252 ( 
.A1(n_29),
.A2(n_32),
.B(n_187),
.C(n_253),
.Y(n_252)
);

BUFx10_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

OA22x2_ASAP7_75t_L g33 ( 
.A1(n_31),
.A2(n_32),
.B1(n_34),
.B2(n_37),
.Y(n_33)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_33),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_33),
.A2(n_81),
.B(n_135),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g272 ( 
.A(n_33),
.B(n_187),
.Y(n_272)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_34),
.Y(n_37)
);

BUFx4f_ASAP7_75t_SL g34 ( 
.A(n_35),
.Y(n_34)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_37),
.B(n_89),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_37),
.B(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_39),
.B(n_80),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

AOI21xp5_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_52),
.B(n_55),
.Y(n_42)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_43),
.A2(n_55),
.B(n_164),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_43),
.A2(n_111),
.B(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_44),
.A2(n_51),
.B1(n_53),
.B2(n_76),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_44),
.B(n_56),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_44),
.A2(n_51),
.B1(n_183),
.B2(n_184),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_44),
.A2(n_51),
.B1(n_183),
.B2(n_211),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_44),
.A2(n_51),
.B1(n_211),
.B2(n_230),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_51),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_46),
.A2(n_47),
.B1(n_48),
.B2(n_49),
.Y(n_45)
);

INVx6_ASAP7_75t_L g225 ( 
.A(n_46),
.Y(n_225)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_48),
.A2(n_49),
.B1(n_61),
.B2(n_62),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_48),
.B(n_61),
.Y(n_200)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_49),
.A2(n_69),
.B1(n_186),
.B2(n_200),
.Y(n_199)
);

BUFx4f_ASAP7_75t_SL g49 ( 
.A(n_50),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_51),
.B(n_56),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_51),
.B(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_51),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_53),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_58),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_58),
.A2(n_73),
.B1(n_103),
.B2(n_115),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_63),
.B(n_67),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_59),
.B(n_71),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_59),
.A2(n_63),
.B1(n_105),
.B2(n_106),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_59),
.A2(n_105),
.B1(n_140),
.B2(n_167),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_59),
.A2(n_105),
.B1(n_167),
.B2(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

O2A1O1Ixp33_ASAP7_75t_L g68 ( 
.A1(n_60),
.A2(n_61),
.B(n_65),
.C(n_69),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_60),
.B(n_99),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_60),
.A2(n_68),
.B1(n_186),
.B2(n_188),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_61),
.B(n_65),
.Y(n_69)
);

CKINVDCx14_ASAP7_75t_R g61 ( 
.A(n_62),
.Y(n_61)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_64),
.Y(n_65)
);

HAxp5_ASAP7_75t_SL g186 ( 
.A(n_65),
.B(n_187),
.CON(n_186),
.SN(n_186)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_68),
.B(n_70),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_68),
.A2(n_99),
.B(n_100),
.Y(n_98)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_68),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_74),
.A2(n_75),
.B(n_78),
.Y(n_125)
);

CKINVDCx14_ASAP7_75t_R g146 ( 
.A(n_74),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_78),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_77),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_77),
.A2(n_113),
.B(n_137),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_81),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_80),
.B(n_83),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_82),
.B(n_83),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_84),
.A2(n_85),
.B1(n_144),
.B2(n_145),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_85),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_94),
.B(n_98),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_86),
.B(n_95),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_86),
.A2(n_98),
.B1(n_123),
.B2(n_124),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_86),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_86),
.A2(n_95),
.B1(n_124),
.B2(n_155),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_91),
.B(n_92),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_87),
.A2(n_159),
.B(n_160),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_87),
.A2(n_90),
.B1(n_159),
.B2(n_202),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g260 ( 
.A1(n_87),
.A2(n_133),
.B(n_261),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_87),
.A2(n_215),
.B1(n_266),
.B2(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_88),
.B(n_131),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_88),
.A2(n_93),
.B(n_161),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_88),
.A2(n_89),
.B1(n_265),
.B2(n_267),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_89),
.B(n_93),
.Y(n_133)
);

INVx11_ASAP7_75t_L g215 ( 
.A(n_89),
.Y(n_215)
);

INVx11_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_91),
.B(n_132),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_91),
.B(n_187),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_94),
.B(n_122),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_95),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_98),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_116),
.Y(n_101)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_103),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_104),
.A2(n_107),
.B1(n_108),
.B2(n_114),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_104),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_105),
.A2(n_140),
.B(n_142),
.Y(n_139)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_110),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_113),
.Y(n_110)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_112),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_119),
.A2(n_147),
.B(n_318),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_143),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_120),
.B(n_143),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_125),
.C(n_126),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_121),
.B(n_125),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_126),
.A2(n_127),
.B1(n_170),
.B2(n_171),
.Y(n_169)
);

CKINVDCx14_ASAP7_75t_R g126 ( 
.A(n_127),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_136),
.C(n_138),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_128),
.B(n_152),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_134),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_129),
.B(n_134),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_133),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_130),
.A2(n_202),
.B(n_215),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_136),
.A2(n_138),
.B1(n_139),
.B2(n_153),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_136),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_148),
.A2(n_172),
.B(n_317),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_169),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g317 ( 
.A(n_149),
.B(n_169),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_154),
.C(n_156),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_150),
.A2(n_151),
.B1(n_154),
.B2(n_315),
.Y(n_314)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_154),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_156),
.B(n_314),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_163),
.C(n_165),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_157),
.B(n_306),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_162),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_158),
.B(n_162),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_161),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_163),
.A2(n_165),
.B1(n_166),
.B2(n_307),
.Y(n_306)
);

CKINVDCx16_ASAP7_75t_R g307 ( 
.A(n_163),
.Y(n_307)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_173),
.A2(n_311),
.B(n_316),
.Y(n_172)
);

O2A1O1Ixp33_ASAP7_75t_SL g173 ( 
.A1(n_174),
.A2(n_216),
.B(n_297),
.C(n_310),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_203),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_175),
.B(n_203),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_190),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_178),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_177),
.B(n_178),
.C(n_190),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_181),
.C(n_185),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_179),
.A2(n_180),
.B1(n_181),
.B2(n_182),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_180),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_182),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_184),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_SL g205 ( 
.A(n_185),
.B(n_206),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_188),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_SL g190 ( 
.A(n_191),
.B(n_198),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_192),
.A2(n_193),
.B1(n_195),
.B2(n_196),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_192),
.B(n_196),
.C(n_198),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_193),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_196),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_201),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_199),
.B(n_201),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_207),
.C(n_209),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_204),
.A2(n_205),
.B1(n_292),
.B2(n_294),
.Y(n_291)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_207),
.A2(n_208),
.B1(n_209),
.B2(n_293),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_209),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_212),
.C(n_214),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_210),
.B(n_238),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_212),
.A2(n_213),
.B1(n_214),
.B2(n_239),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_213),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_214),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_217),
.B(n_296),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_218),
.A2(n_289),
.B(n_295),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_219),
.A2(n_244),
.B(n_288),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_235),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_220),
.B(n_235),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_228),
.C(n_231),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_221),
.A2(n_222),
.B1(n_285),
.B2(n_286),
.Y(n_284)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_224),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_223),
.B(n_224),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_228),
.A2(n_229),
.B1(n_231),
.B2(n_232),
.Y(n_286)
);

CKINVDCx16_ASAP7_75t_R g228 ( 
.A(n_229),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_232),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_236),
.A2(n_237),
.B1(n_240),
.B2(n_241),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_236),
.B(n_242),
.C(n_243),
.Y(n_290)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_243),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_245),
.A2(n_282),
.B(n_287),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_L g245 ( 
.A1(n_246),
.A2(n_262),
.B(n_281),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_254),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_247),
.B(n_254),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_248),
.B(n_252),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_248),
.A2(n_249),
.B1(n_252),
.B2(n_269),
.Y(n_268)
);

CKINVDCx16_ASAP7_75t_R g248 ( 
.A(n_249),
.Y(n_248)
);

CKINVDCx16_ASAP7_75t_R g269 ( 
.A(n_252),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_260),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_256),
.A2(n_257),
.B1(n_258),
.B2(n_259),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_256),
.B(n_259),
.C(n_260),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_257),
.Y(n_256)
);

CKINVDCx16_ASAP7_75t_R g258 ( 
.A(n_259),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_261),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_263),
.A2(n_270),
.B(n_280),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_268),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g280 ( 
.A(n_264),
.B(n_268),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_271),
.A2(n_275),
.B(n_279),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_273),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_272),
.B(n_273),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_276),
.B(n_277),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_284),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_SL g287 ( 
.A(n_283),
.B(n_284),
.Y(n_287)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_291),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_SL g295 ( 
.A(n_290),
.B(n_291),
.Y(n_295)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_292),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_299),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_SL g310 ( 
.A(n_298),
.B(n_299),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_300),
.A2(n_301),
.B1(n_308),
.B2(n_309),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_302),
.A2(n_303),
.B1(n_304),
.B2(n_305),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_302),
.B(n_305),
.C(n_309),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_303),
.Y(n_302)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_308),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_313),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_312),
.B(n_313),
.Y(n_316)
);


endmodule