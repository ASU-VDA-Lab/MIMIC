module real_jpeg_14865_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_380, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_380;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_366;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_373;
wire n_375;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_0),
.Y(n_68)
);

BUFx4f_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_2),
.Y(n_44)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_3),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_3),
.B(n_40),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_3),
.B(n_25),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_3),
.B(n_88),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_3),
.B(n_68),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_3),
.B(n_34),
.Y(n_285)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_5),
.B(n_88),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_5),
.B(n_54),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_5),
.B(n_25),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_5),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_5),
.B(n_40),
.Y(n_266)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_6),
.B(n_31),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_6),
.B(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_6),
.B(n_40),
.Y(n_39)
);

AND2x2_ASAP7_75t_SL g67 ( 
.A(n_6),
.B(n_68),
.Y(n_67)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_6),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_6),
.B(n_25),
.Y(n_91)
);

AND2x2_ASAP7_75t_SL g140 ( 
.A(n_6),
.B(n_88),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_6),
.B(n_54),
.Y(n_164)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_7),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_8),
.B(n_43),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_8),
.B(n_31),
.Y(n_181)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_8),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_8),
.B(n_68),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_8),
.B(n_88),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_8),
.B(n_40),
.Y(n_311)
);

AND2x2_ASAP7_75t_L g24 ( 
.A(n_9),
.B(n_25),
.Y(n_24)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_9),
.B(n_40),
.Y(n_49)
);

CKINVDCx14_ASAP7_75t_R g71 ( 
.A(n_9),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_9),
.B(n_54),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_9),
.B(n_88),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_9),
.B(n_34),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_9),
.B(n_68),
.Y(n_210)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_10),
.B(n_40),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_10),
.B(n_34),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_10),
.B(n_31),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_10),
.B(n_88),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_10),
.B(n_54),
.Y(n_318)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_11),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_13),
.B(n_25),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_13),
.B(n_88),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_13),
.B(n_34),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_13),
.B(n_31),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_13),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_13),
.B(n_54),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_13),
.B(n_40),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_13),
.B(n_43),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_14),
.B(n_25),
.Y(n_46)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_14),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_14),
.B(n_54),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_14),
.B(n_31),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_14),
.B(n_34),
.Y(n_326)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_147),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_146),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_122),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_20),
.B(n_122),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_20),
.B(n_149),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g376 ( 
.A(n_20),
.B(n_149),
.Y(n_376)
);

FAx1_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_61),
.CI(n_96),
.CON(n_20),
.SN(n_20)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_38),
.C(n_47),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_22),
.A2(n_23),
.B1(n_38),
.B2(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_27),
.B1(n_28),
.B2(n_37),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_24),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_24),
.B(n_30),
.C(n_32),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_24),
.A2(n_37),
.B1(n_309),
.B2(n_310),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_24),
.B(n_140),
.C(n_312),
.Y(n_340)
);

INVx5_ASAP7_75t_SL g198 ( 
.A(n_25),
.Y(n_198)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_30),
.B1(n_32),
.B2(n_33),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_29),
.A2(n_30),
.B1(n_91),
.B2(n_92),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_29),
.A2(n_30),
.B1(n_252),
.B2(n_253),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_30),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_30),
.B(n_87),
.C(n_91),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_30),
.B(n_250),
.C(n_252),
.Y(n_290)
);

INVx13_ASAP7_75t_L g72 ( 
.A(n_31),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_32),
.B(n_65),
.C(n_74),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_32),
.A2(n_33),
.B1(n_74),
.B2(n_116),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_32),
.A2(n_33),
.B1(n_121),
.B2(n_158),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_32),
.A2(n_33),
.B1(n_210),
.B2(n_211),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_33),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_33),
.B(n_118),
.C(n_121),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_33),
.B(n_210),
.Y(n_264)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_35),
.B(n_186),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_35),
.B(n_229),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_38),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_41),
.C(n_46),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_39),
.A2(n_41),
.B1(n_102),
.B2(n_103),
.Y(n_101)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_39),
.Y(n_103)
);

INVx1_ASAP7_75t_SL g131 ( 
.A(n_40),
.Y(n_131)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_41),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_45),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_42),
.B(n_75),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_42),
.B(n_71),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_42),
.B(n_56),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_42),
.B(n_229),
.Y(n_300)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_45),
.B(n_188),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_45),
.B(n_198),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g100 ( 
.A(n_46),
.B(n_101),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_47),
.A2(n_48),
.B1(n_166),
.B2(n_167),
.Y(n_165)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_49),
.A2(n_50),
.B1(n_51),
.B2(n_60),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_49),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_49),
.B(n_52),
.C(n_57),
.Y(n_94)
);

CKINVDCx14_ASAP7_75t_R g50 ( 
.A(n_51),
.Y(n_50)
);

XOR2xp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_57),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_56),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_53),
.B(n_186),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_54),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_56),
.B(n_72),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_59),
.Y(n_57)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_58),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_59),
.B(n_131),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_59),
.B(n_188),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_84),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_63),
.A2(n_64),
.B1(n_76),
.B2(n_77),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_63),
.B(n_77),
.C(n_84),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_64),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_65),
.A2(n_66),
.B1(n_114),
.B2(n_115),
.Y(n_113)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_69),
.C(n_73),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_67),
.A2(n_69),
.B1(n_70),
.B2(n_111),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_67),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_67),
.B(n_119),
.C(n_120),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_67),
.A2(n_111),
.B1(n_119),
.B2(n_162),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_67),
.A2(n_111),
.B1(n_190),
.B2(n_191),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_67),
.B(n_190),
.Y(n_206)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_68),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_69),
.A2(n_70),
.B1(n_91),
.B2(n_92),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_69),
.B(n_91),
.C(n_300),
.Y(n_319)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_71),
.B(n_72),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_72),
.B(n_229),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_73),
.A2(n_109),
.B1(n_110),
.B2(n_112),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_73),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_73),
.A2(n_109),
.B1(n_137),
.B2(n_138),
.Y(n_136)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_74),
.Y(n_116)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_79),
.B1(n_80),
.B2(n_83),
.Y(n_77)
);

CKINVDCx14_ASAP7_75t_R g78 ( 
.A(n_79),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_79),
.B(n_81),
.C(n_82),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_80),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_SL g80 ( 
.A(n_81),
.B(n_82),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_SL g84 ( 
.A(n_85),
.B(n_93),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_85),
.B(n_94),
.C(n_95),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_87),
.B1(n_89),
.B2(n_90),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_86),
.A2(n_87),
.B1(n_105),
.B2(n_338),
.Y(n_337)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_87),
.B(n_105),
.C(n_106),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_91),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_91),
.A2(n_92),
.B1(n_139),
.B2(n_140),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_95),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_113),
.C(n_117),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_97),
.A2(n_98),
.B1(n_170),
.B2(n_171),
.Y(n_169)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_104),
.C(n_107),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_99),
.A2(n_100),
.B1(n_153),
.B2(n_154),
.Y(n_152)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_104),
.A2(n_107),
.B1(n_108),
.B2(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_104),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_105),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_106),
.B(n_337),
.Y(n_336)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_110),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_113),
.B(n_117),
.Y(n_171)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_118),
.B(n_157),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_119),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_119),
.A2(n_162),
.B1(n_257),
.B2(n_258),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_119),
.B(n_257),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_120),
.B(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_121),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_145),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_124),
.A2(n_125),
.B1(n_143),
.B2(n_144),
.Y(n_123)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_124),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_125),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_SL g125 ( 
.A(n_126),
.B(n_134),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_128),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_129),
.A2(n_130),
.B1(n_132),
.B2(n_133),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_130),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_133),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_135),
.A2(n_136),
.B1(n_141),
.B2(n_142),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_139),
.A2(n_140),
.B1(n_311),
.B2(n_312),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

OAI21xp33_ASAP7_75t_L g147 ( 
.A1(n_148),
.A2(n_172),
.B(n_376),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_165),
.C(n_169),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g368 ( 
.A(n_150),
.B(n_369),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_156),
.C(n_159),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_151),
.A2(n_152),
.B1(n_363),
.B2(n_364),
.Y(n_362)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g364 ( 
.A(n_156),
.B(n_159),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_163),
.C(n_164),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g346 ( 
.A(n_160),
.B(n_347),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_L g347 ( 
.A1(n_163),
.A2(n_164),
.B1(n_348),
.B2(n_349),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_163),
.Y(n_349)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_164),
.Y(n_348)
);

XOR2xp5_ASAP7_75t_L g369 ( 
.A(n_165),
.B(n_169),
.Y(n_369)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

AOI321xp33_ASAP7_75t_L g172 ( 
.A1(n_173),
.A2(n_356),
.A3(n_366),
.B1(n_370),
.B2(n_375),
.C(n_380),
.Y(n_172)
);

NOR3xp33_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_303),
.C(n_351),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_175),
.A2(n_274),
.B(n_302),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_176),
.A2(n_244),
.B(n_273),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_213),
.B(n_243),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_192),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_178),
.B(n_192),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_183),
.C(n_189),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_179),
.A2(n_195),
.B1(n_196),
.B2(n_204),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_179),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_179),
.B(n_240),
.Y(n_239)
);

FAx1_ASAP7_75t_SL g179 ( 
.A(n_180),
.B(n_181),
.CI(n_182),
.CON(n_179),
.SN(n_179)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_183),
.A2(n_184),
.B1(n_189),
.B2(n_241),
.Y(n_240)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_184),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_187),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_SL g222 ( 
.A(n_185),
.B(n_187),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_186),
.B(n_198),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_188),
.B(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_189),
.Y(n_241)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_193),
.A2(n_194),
.B1(n_205),
.B2(n_212),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_195),
.B(n_204),
.C(n_212),
.Y(n_245)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_196),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_199),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_197),
.B(n_200),
.C(n_203),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_201),
.B1(n_202),
.B2(n_203),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_202),
.Y(n_203)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_205),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_SL g205 ( 
.A(n_206),
.B(n_207),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_206),
.B(n_208),
.C(n_209),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_209),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_210),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_210),
.A2(n_211),
.B1(n_326),
.B2(n_327),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_210),
.B(n_324),
.C(n_327),
.Y(n_341)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_214),
.A2(n_237),
.B(n_242),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_215),
.A2(n_226),
.B(n_236),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_221),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_216),
.B(n_221),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_217),
.B(n_219),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_217),
.A2(n_218),
.B1(n_219),
.B2(n_220),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_218),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_220),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_223),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_222),
.B(n_224),
.C(n_225),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_225),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_227),
.A2(n_231),
.B(n_235),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_230),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_228),
.B(n_230),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_232),
.B(n_234),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_239),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_238),
.B(n_239),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_246),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_245),
.B(n_246),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_247),
.A2(n_248),
.B1(n_259),
.B2(n_260),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_247),
.B(n_261),
.C(n_272),
.Y(n_275)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_254),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_249),
.B(n_255),
.C(n_256),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_SL g249 ( 
.A(n_250),
.B(n_251),
.Y(n_249)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_256),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_258),
.Y(n_257)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_261),
.A2(n_262),
.B1(n_271),
.B2(n_272),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_263),
.A2(n_264),
.B1(n_265),
.B2(n_270),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_263),
.B(n_267),
.C(n_269),
.Y(n_293)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_265),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_266),
.A2(n_267),
.B1(n_268),
.B2(n_269),
.Y(n_265)
);

CKINVDCx14_ASAP7_75t_R g269 ( 
.A(n_266),
.Y(n_269)
);

CKINVDCx14_ASAP7_75t_R g267 ( 
.A(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_276),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_275),
.B(n_276),
.Y(n_302)
);

AOI22xp33_ASAP7_75t_SL g276 ( 
.A1(n_277),
.A2(n_278),
.B1(n_292),
.B2(n_301),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_279),
.A2(n_280),
.B1(n_281),
.B2(n_291),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_279),
.B(n_291),
.C(n_301),
.Y(n_352)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_281),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_282),
.A2(n_283),
.B1(n_287),
.B2(n_288),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_282),
.B(n_289),
.C(n_290),
.Y(n_320)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

BUFx24_ASAP7_75t_SL g379 ( 
.A(n_283),
.Y(n_379)
);

FAx1_ASAP7_75t_SL g283 ( 
.A(n_284),
.B(n_285),
.CI(n_286),
.CON(n_283),
.SN(n_283)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_284),
.B(n_285),
.C(n_286),
.Y(n_329)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_SL g288 ( 
.A(n_289),
.B(n_290),
.Y(n_288)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_292),
.Y(n_301)
);

BUFx24_ASAP7_75t_SL g377 ( 
.A(n_292),
.Y(n_377)
);

FAx1_ASAP7_75t_SL g292 ( 
.A(n_293),
.B(n_294),
.CI(n_298),
.CON(n_292),
.SN(n_292)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_293),
.B(n_294),
.C(n_298),
.Y(n_332)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_295),
.A2(n_296),
.B(n_297),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_295),
.B(n_296),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_297),
.A2(n_329),
.B1(n_330),
.B2(n_331),
.Y(n_328)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_297),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_SL g298 ( 
.A(n_299),
.B(n_300),
.Y(n_298)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

AOI21xp33_ASAP7_75t_L g371 ( 
.A1(n_304),
.A2(n_372),
.B(n_373),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_333),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_305),
.B(n_333),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_321),
.C(n_332),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g353 ( 
.A(n_306),
.B(n_354),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_SL g306 ( 
.A(n_307),
.B(n_320),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_313),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_308),
.B(n_313),
.C(n_320),
.Y(n_350)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

CKINVDCx16_ASAP7_75t_R g312 ( 
.A(n_311),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_319),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_315),
.A2(n_316),
.B1(n_317),
.B2(n_318),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_316),
.B(n_317),
.C(n_319),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_318),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_L g354 ( 
.A1(n_321),
.A2(n_322),
.B1(n_332),
.B2(n_355),
.Y(n_354)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_SL g322 ( 
.A(n_323),
.B(n_328),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_323),
.B(n_329),
.C(n_331),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_SL g323 ( 
.A(n_324),
.B(n_325),
.Y(n_323)
);

CKINVDCx14_ASAP7_75t_R g327 ( 
.A(n_326),
.Y(n_327)
);

CKINVDCx14_ASAP7_75t_R g330 ( 
.A(n_329),
.Y(n_330)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_332),
.Y(n_355)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_334),
.B(n_350),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_335),
.B(n_342),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_335),
.B(n_342),
.C(n_350),
.Y(n_358)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_336),
.B(n_339),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_336),
.B(n_340),
.C(n_341),
.Y(n_361)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_340),
.B(n_341),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_SL g342 ( 
.A(n_343),
.B(n_344),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_343),
.B(n_345),
.C(n_346),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_345),
.B(n_346),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_352),
.B(n_353),
.Y(n_351)
);

AND2x2_ASAP7_75t_L g372 ( 
.A(n_352),
.B(n_353),
.Y(n_372)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

OAI21xp5_ASAP7_75t_SL g370 ( 
.A1(n_357),
.A2(n_371),
.B(n_374),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_358),
.B(n_359),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_SL g374 ( 
.A(n_358),
.B(n_359),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_360),
.B(n_365),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_361),
.B(n_362),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_361),
.B(n_362),
.C(n_365),
.Y(n_367)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_367),
.B(n_368),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_367),
.B(n_368),
.Y(n_375)
);


endmodule