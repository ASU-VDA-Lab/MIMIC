module fake_ariane_1564_n_1083 (n_83, n_8, n_233, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_240, n_167, n_90, n_195, n_38, n_213, n_47, n_110, n_153, n_18, n_197, n_221, n_86, n_269, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_237, n_172, n_69, n_259, n_95, n_175, n_92, n_143, n_183, n_203, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_242, n_260, n_274, n_115, n_272, n_133, n_66, n_205, n_236, n_265, n_71, n_267, n_24, n_7, n_109, n_208, n_245, n_96, n_156, n_209, n_49, n_262, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_210, n_147, n_204, n_225, n_235, n_200, n_51, n_166, n_253, n_76, n_218, n_103, n_79, n_26, n_244, n_226, n_3, n_246, n_271, n_46, n_220, n_0, n_84, n_247, n_261, n_36, n_199, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_217, n_44, n_224, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_263, n_201, n_229, n_70, n_250, n_222, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_256, n_6, n_214, n_227, n_48, n_94, n_101, n_243, n_4, n_134, n_188, n_185, n_2, n_32, n_249, n_37, n_58, n_65, n_123, n_212, n_9, n_138, n_112, n_45, n_162, n_11, n_264, n_129, n_126, n_137, n_255, n_122, n_268, n_257, n_266, n_198, n_148, n_232, n_164, n_52, n_157, n_248, n_184, n_177, n_135, n_258, n_73, n_77, n_171, n_228, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_206, n_13, n_27, n_207, n_241, n_29, n_254, n_238, n_41, n_219, n_140, n_55, n_191, n_151, n_136, n_231, n_192, n_28, n_80, n_146, n_234, n_230, n_211, n_270, n_194, n_97, n_154, n_215, n_252, n_142, n_251, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_202, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_216, n_16, n_5, n_155, n_127, n_239, n_223, n_35, n_273, n_54, n_25, n_1083);

input n_83;
input n_8;
input n_233;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_240;
input n_167;
input n_90;
input n_195;
input n_38;
input n_213;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_221;
input n_86;
input n_269;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_237;
input n_172;
input n_69;
input n_259;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_203;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_242;
input n_260;
input n_274;
input n_115;
input n_272;
input n_133;
input n_66;
input n_205;
input n_236;
input n_265;
input n_71;
input n_267;
input n_24;
input n_7;
input n_109;
input n_208;
input n_245;
input n_96;
input n_156;
input n_209;
input n_49;
input n_262;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_210;
input n_147;
input n_204;
input n_225;
input n_235;
input n_200;
input n_51;
input n_166;
input n_253;
input n_76;
input n_218;
input n_103;
input n_79;
input n_26;
input n_244;
input n_226;
input n_3;
input n_246;
input n_271;
input n_46;
input n_220;
input n_0;
input n_84;
input n_247;
input n_261;
input n_36;
input n_199;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_217;
input n_44;
input n_224;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_263;
input n_201;
input n_229;
input n_70;
input n_250;
input n_222;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_256;
input n_6;
input n_214;
input n_227;
input n_48;
input n_94;
input n_101;
input n_243;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_249;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_264;
input n_129;
input n_126;
input n_137;
input n_255;
input n_122;
input n_268;
input n_257;
input n_266;
input n_198;
input n_148;
input n_232;
input n_164;
input n_52;
input n_157;
input n_248;
input n_184;
input n_177;
input n_135;
input n_258;
input n_73;
input n_77;
input n_171;
input n_228;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_206;
input n_13;
input n_27;
input n_207;
input n_241;
input n_29;
input n_254;
input n_238;
input n_41;
input n_219;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_231;
input n_192;
input n_28;
input n_80;
input n_146;
input n_234;
input n_230;
input n_211;
input n_270;
input n_194;
input n_97;
input n_154;
input n_215;
input n_252;
input n_142;
input n_251;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_202;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_216;
input n_16;
input n_5;
input n_155;
input n_127;
input n_239;
input n_223;
input n_35;
input n_273;
input n_54;
input n_25;

output n_1083;

wire n_295;
wire n_356;
wire n_556;
wire n_698;
wire n_1072;
wire n_695;
wire n_913;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_1008;
wire n_581;
wire n_294;
wire n_1020;
wire n_646;
wire n_640;
wire n_463;
wire n_1024;
wire n_830;
wire n_691;
wire n_404;
wire n_943;
wire n_678;
wire n_1058;
wire n_651;
wire n_987;
wire n_936;
wire n_347;
wire n_423;
wire n_1042;
wire n_961;
wire n_469;
wire n_1046;
wire n_479;
wire n_726;
wire n_603;
wire n_878;
wire n_373;
wire n_299;
wire n_836;
wire n_541;
wire n_499;
wire n_789;
wire n_788;
wire n_850;
wire n_908;
wire n_771;
wire n_1036;
wire n_564;
wire n_610;
wire n_752;
wire n_341;
wire n_1029;
wire n_985;
wire n_421;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_760;
wire n_690;
wire n_906;
wire n_416;
wire n_969;
wire n_283;
wire n_919;
wire n_525;
wire n_806;
wire n_367;
wire n_970;
wire n_713;
wire n_649;
wire n_598;
wire n_345;
wire n_374;
wire n_318;
wire n_817;
wire n_643;
wire n_679;
wire n_924;
wire n_927;
wire n_781;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_717;
wire n_819;
wire n_286;
wire n_443;
wire n_586;
wire n_864;
wire n_952;
wire n_686;
wire n_605;
wire n_776;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_826;
wire n_524;
wire n_391;
wire n_349;
wire n_634;
wire n_466;
wire n_756;
wire n_1016;
wire n_346;
wire n_940;
wire n_764;
wire n_979;
wire n_348;
wire n_552;
wire n_1077;
wire n_462;
wire n_607;
wire n_670;
wire n_897;
wire n_956;
wire n_949;
wire n_410;
wire n_379;
wire n_445;
wire n_515;
wire n_807;
wire n_765;
wire n_891;
wire n_737;
wire n_885;
wire n_441;
wire n_568;
wire n_1032;
wire n_385;
wire n_637;
wire n_917;
wire n_327;
wire n_766;
wire n_372;
wire n_377;
wire n_396;
wire n_802;
wire n_631;
wire n_399;
wire n_554;
wire n_960;
wire n_520;
wire n_980;
wire n_870;
wire n_714;
wire n_279;
wire n_905;
wire n_702;
wire n_958;
wire n_945;
wire n_790;
wire n_857;
wire n_898;
wire n_363;
wire n_720;
wire n_968;
wire n_1067;
wire n_354;
wire n_813;
wire n_926;
wire n_725;
wire n_419;
wire n_1009;
wire n_1064;
wire n_633;
wire n_900;
wire n_883;
wire n_338;
wire n_995;
wire n_285;
wire n_473;
wire n_801;
wire n_733;
wire n_761;
wire n_818;
wire n_500;
wire n_665;
wire n_336;
wire n_731;
wire n_754;
wire n_779;
wire n_871;
wire n_315;
wire n_903;
wire n_1073;
wire n_594;
wire n_311;
wire n_402;
wire n_1052;
wire n_1068;
wire n_829;
wire n_1062;
wire n_668;
wire n_339;
wire n_758;
wire n_738;
wire n_833;
wire n_672;
wire n_487;
wire n_740;
wire n_879;
wire n_422;
wire n_648;
wire n_784;
wire n_597;
wire n_816;
wire n_1018;
wire n_855;
wire n_1047;
wire n_835;
wire n_808;
wire n_953;
wire n_446;
wire n_553;
wire n_1076;
wire n_753;
wire n_1050;
wire n_566;
wire n_814;
wire n_578;
wire n_701;
wire n_1003;
wire n_625;
wire n_405;
wire n_557;
wire n_858;
wire n_645;
wire n_989;
wire n_309;
wire n_331;
wire n_320;
wire n_559;
wire n_401;
wire n_485;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_1035;
wire n_350;
wire n_291;
wire n_822;
wire n_344;
wire n_381;
wire n_795;
wire n_426;
wire n_433;
wire n_481;
wire n_600;
wire n_721;
wire n_840;
wire n_1053;
wire n_398;
wire n_529;
wire n_502;
wire n_561;
wire n_770;
wire n_839;
wire n_821;
wire n_928;
wire n_465;
wire n_486;
wire n_507;
wire n_901;
wire n_759;
wire n_569;
wire n_567;
wire n_825;
wire n_732;
wire n_971;
wire n_369;
wire n_787;
wire n_894;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_478;
wire n_703;
wire n_748;
wire n_786;
wire n_510;
wire n_1061;
wire n_1045;
wire n_831;
wire n_868;
wire n_326;
wire n_681;
wire n_778;
wire n_874;
wire n_323;
wire n_550;
wire n_1023;
wire n_988;
wire n_635;
wire n_707;
wire n_997;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_694;
wire n_884;
wire n_983;
wire n_282;
wire n_328;
wire n_368;
wire n_1034;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_277;
wire n_467;
wire n_432;
wire n_545;
wire n_1015;
wire n_536;
wire n_644;
wire n_293;
wire n_823;
wire n_921;
wire n_620;
wire n_325;
wire n_276;
wire n_688;
wire n_1074;
wire n_859;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_693;
wire n_863;
wire n_303;
wire n_671;
wire n_442;
wire n_777;
wire n_929;
wire n_352;
wire n_538;
wire n_920;
wire n_899;
wire n_576;
wire n_843;
wire n_1080;
wire n_511;
wire n_611;
wire n_365;
wire n_429;
wire n_455;
wire n_654;
wire n_588;
wire n_1013;
wire n_986;
wire n_638;
wire n_334;
wire n_729;
wire n_887;
wire n_661;
wire n_488;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_300;
wire n_533;
wire n_904;
wire n_505;
wire n_869;
wire n_846;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_1059;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_1039;
wire n_305;
wire n_539;
wire n_312;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_977;
wire n_957;
wire n_512;
wire n_715;
wire n_889;
wire n_1066;
wire n_935;
wire n_579;
wire n_844;
wire n_1012;
wire n_459;
wire n_685;
wire n_321;
wire n_911;
wire n_361;
wire n_458;
wire n_383;
wire n_623;
wire n_838;
wire n_861;
wire n_780;
wire n_950;
wire n_1017;
wire n_711;
wire n_877;
wire n_1021;
wire n_1065;
wire n_453;
wire n_734;
wire n_491;
wire n_810;
wire n_723;
wire n_616;
wire n_617;
wire n_658;
wire n_630;
wire n_705;
wire n_570;
wire n_1055;
wire n_362;
wire n_543;
wire n_942;
wire n_310;
wire n_709;
wire n_601;
wire n_683;
wire n_565;
wire n_281;
wire n_628;
wire n_809;
wire n_461;
wire n_490;
wire n_743;
wire n_907;
wire n_1006;
wire n_881;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_1019;
wire n_297;
wire n_962;
wire n_662;
wire n_641;
wire n_1005;
wire n_503;
wire n_941;
wire n_700;
wire n_910;
wire n_290;
wire n_527;
wire n_741;
wire n_747;
wire n_772;
wire n_847;
wire n_939;
wire n_371;
wire n_845;
wire n_888;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_676;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_1038;
wire n_572;
wire n_343;
wire n_865;
wire n_1041;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_993;
wire n_380;
wire n_948;
wire n_582;
wire n_284;
wire n_922;
wire n_1004;
wire n_448;
wire n_593;
wire n_755;
wire n_710;
wire n_860;
wire n_534;
wire n_355;
wire n_444;
wire n_609;
wire n_278;
wire n_851;
wire n_1043;
wire n_560;
wire n_450;
wire n_890;
wire n_842;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_1022;
wire n_1033;
wire n_896;
wire n_409;
wire n_947;
wire n_930;
wire n_519;
wire n_902;
wire n_384;
wire n_1031;
wire n_468;
wire n_1056;
wire n_853;
wire n_526;
wire n_716;
wire n_742;
wire n_696;
wire n_1040;
wire n_674;
wire n_1081;
wire n_482;
wire n_316;
wire n_798;
wire n_769;
wire n_820;
wire n_577;
wire n_407;
wire n_774;
wire n_933;
wire n_872;
wire n_916;
wire n_596;
wire n_954;
wire n_912;
wire n_476;
wire n_460;
wire n_832;
wire n_535;
wire n_366;
wire n_762;
wire n_744;
wire n_656;
wire n_555;
wire n_492;
wire n_574;
wire n_848;
wire n_804;
wire n_280;
wire n_982;
wire n_915;
wire n_629;
wire n_664;
wire n_1075;
wire n_454;
wire n_992;
wire n_966;
wire n_298;
wire n_955;
wire n_532;
wire n_415;
wire n_794;
wire n_763;
wire n_655;
wire n_544;
wire n_540;
wire n_692;
wire n_599;
wire n_768;
wire n_514;
wire n_418;
wire n_984;
wire n_537;
wire n_1063;
wire n_403;
wire n_750;
wire n_834;
wire n_991;
wire n_389;
wire n_1007;
wire n_800;
wire n_657;
wire n_513;
wire n_837;
wire n_288;
wire n_812;
wire n_395;
wire n_621;
wire n_606;
wire n_951;
wire n_1026;
wire n_938;
wire n_862;
wire n_304;
wire n_895;
wire n_659;
wire n_509;
wire n_583;
wire n_1014;
wire n_724;
wire n_306;
wire n_666;
wire n_1000;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_378;
wire n_436;
wire n_946;
wire n_757;
wire n_375;
wire n_324;
wire n_1030;
wire n_585;
wire n_875;
wire n_669;
wire n_785;
wire n_827;
wire n_931;
wire n_619;
wire n_337;
wire n_437;
wire n_622;
wire n_697;
wire n_999;
wire n_998;
wire n_967;
wire n_472;
wire n_937;
wire n_296;
wire n_746;
wire n_456;
wire n_292;
wire n_880;
wire n_793;
wire n_852;
wire n_1079;
wire n_275;
wire n_704;
wire n_1060;
wire n_1044;
wire n_751;
wire n_615;
wire n_1027;
wire n_1070;
wire n_996;
wire n_521;
wire n_963;
wire n_873;
wire n_1082;
wire n_496;
wire n_739;
wire n_1028;
wire n_342;
wire n_866;
wire n_517;
wire n_925;
wire n_530;
wire n_792;
wire n_1001;
wire n_824;
wire n_428;
wire n_1002;
wire n_358;
wire n_580;
wire n_892;
wire n_608;
wire n_959;
wire n_494;
wire n_1051;
wire n_719;
wire n_434;
wire n_360;
wire n_975;
wire n_563;
wire n_394;
wire n_923;
wire n_932;
wire n_773;
wire n_1037;
wire n_981;
wire n_1010;
wire n_882;
wire n_990;
wire n_317;
wire n_867;
wire n_803;
wire n_329;
wire n_718;
wire n_340;
wire n_944;
wire n_749;
wire n_994;
wire n_289;
wire n_548;
wire n_542;
wire n_815;
wire n_973;
wire n_523;
wire n_1078;
wire n_972;
wire n_470;
wire n_457;
wire n_632;
wire n_477;
wire n_364;
wire n_650;
wire n_782;
wire n_856;
wire n_425;
wire n_431;
wire n_811;
wire n_1054;
wire n_508;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1071;
wire n_411;
wire n_484;
wire n_712;
wire n_849;
wire n_909;
wire n_976;
wire n_353;
wire n_736;
wire n_767;
wire n_1025;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_964;
wire n_1057;
wire n_382;
wire n_797;
wire n_489;
wire n_480;
wire n_978;
wire n_642;
wire n_1011;
wire n_408;
wire n_828;
wire n_595;
wire n_322;
wire n_974;
wire n_506;
wire n_893;
wire n_602;
wire n_799;
wire n_558;
wire n_592;
wire n_397;
wire n_841;
wire n_854;
wire n_471;
wire n_351;
wire n_1069;
wire n_965;
wire n_393;
wire n_886;
wire n_474;
wire n_653;
wire n_359;
wire n_573;
wire n_796;
wire n_805;
wire n_531;
wire n_934;
wire n_783;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_242),
.Y(n_275)
);

BUFx3_ASAP7_75t_L g276 ( 
.A(n_75),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_63),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_256),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_149),
.Y(n_279)
);

BUFx4f_ASAP7_75t_SL g280 ( 
.A(n_54),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_204),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_109),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_107),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_103),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_243),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_37),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_81),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_13),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_177),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_186),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_190),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_110),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_119),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_134),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_129),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_180),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_170),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_192),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_7),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_132),
.Y(n_300)
);

BUFx2_ASAP7_75t_L g301 ( 
.A(n_128),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_238),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_66),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_273),
.Y(n_304)
);

HB1xp67_ASAP7_75t_L g305 ( 
.A(n_9),
.Y(n_305)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_199),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_24),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_117),
.Y(n_308)
);

CKINVDCx16_ASAP7_75t_R g309 ( 
.A(n_239),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_162),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_206),
.Y(n_311)
);

BUFx5_ASAP7_75t_L g312 ( 
.A(n_189),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_101),
.Y(n_313)
);

BUFx5_ASAP7_75t_L g314 ( 
.A(n_152),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_262),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_188),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_213),
.Y(n_317)
);

INVx2_ASAP7_75t_SL g318 ( 
.A(n_196),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_155),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_105),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_156),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_145),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_13),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_76),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_227),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_15),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_217),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_267),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_226),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_230),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_253),
.Y(n_331)
);

BUFx2_ASAP7_75t_L g332 ( 
.A(n_157),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_45),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_123),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_96),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_83),
.Y(n_336)
);

CKINVDCx16_ASAP7_75t_R g337 ( 
.A(n_19),
.Y(n_337)
);

BUFx3_ASAP7_75t_L g338 ( 
.A(n_125),
.Y(n_338)
);

BUFx2_ASAP7_75t_SL g339 ( 
.A(n_198),
.Y(n_339)
);

HB1xp67_ASAP7_75t_L g340 ( 
.A(n_305),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_309),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_337),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_305),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_288),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_284),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_301),
.B(n_0),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_303),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_332),
.B(n_0),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_325),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_307),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_326),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_323),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_277),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_285),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_292),
.B(n_1),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_327),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_293),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_294),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_329),
.Y(n_359)
);

NOR2xp67_ASAP7_75t_L g360 ( 
.A(n_299),
.B(n_1),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_296),
.B(n_2),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_297),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_298),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_300),
.Y(n_364)
);

BUFx2_ASAP7_75t_SL g365 ( 
.A(n_276),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_302),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_308),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_275),
.Y(n_368)
);

BUFx2_ASAP7_75t_L g369 ( 
.A(n_276),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_311),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_317),
.Y(n_371)
);

INVxp67_ASAP7_75t_SL g372 ( 
.A(n_338),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_338),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_319),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_278),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_321),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_324),
.B(n_2),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_330),
.Y(n_378)
);

INVxp67_ASAP7_75t_L g379 ( 
.A(n_331),
.Y(n_379)
);

CKINVDCx16_ASAP7_75t_R g380 ( 
.A(n_339),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_335),
.Y(n_381)
);

CKINVDCx16_ASAP7_75t_R g382 ( 
.A(n_318),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_353),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_349),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_345),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_344),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g387 ( 
.A(n_345),
.B(n_3),
.Y(n_387)
);

INVx3_ASAP7_75t_L g388 ( 
.A(n_354),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_357),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_350),
.Y(n_390)
);

NAND2x1_ASAP7_75t_L g391 ( 
.A(n_369),
.B(n_306),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_372),
.B(n_336),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_351),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_347),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_356),
.Y(n_395)
);

AND2x4_ASAP7_75t_L g396 ( 
.A(n_379),
.B(n_306),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_382),
.B(n_316),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_381),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_358),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_362),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_363),
.Y(n_401)
);

HB1xp67_ASAP7_75t_L g402 ( 
.A(n_342),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_347),
.Y(n_403)
);

AND2x2_ASAP7_75t_L g404 ( 
.A(n_380),
.B(n_316),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_364),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_366),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_356),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_367),
.Y(n_408)
);

BUFx6f_ASAP7_75t_L g409 ( 
.A(n_370),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_371),
.Y(n_410)
);

HB1xp67_ASAP7_75t_L g411 ( 
.A(n_342),
.Y(n_411)
);

INVx3_ASAP7_75t_L g412 ( 
.A(n_374),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_359),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_368),
.Y(n_414)
);

AND2x4_ASAP7_75t_L g415 ( 
.A(n_376),
.B(n_378),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_352),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_365),
.B(n_320),
.Y(n_417)
);

HB1xp67_ASAP7_75t_L g418 ( 
.A(n_341),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_359),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_343),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_355),
.Y(n_421)
);

BUFx6f_ASAP7_75t_L g422 ( 
.A(n_361),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_373),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_377),
.Y(n_424)
);

HB1xp67_ASAP7_75t_L g425 ( 
.A(n_341),
.Y(n_425)
);

BUFx6f_ASAP7_75t_L g426 ( 
.A(n_348),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_375),
.B(n_279),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_375),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_373),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_340),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_346),
.Y(n_431)
);

INVx3_ASAP7_75t_L g432 ( 
.A(n_409),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_386),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_427),
.B(n_428),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_416),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_390),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_L g437 ( 
.A1(n_431),
.A2(n_360),
.B1(n_281),
.B2(n_283),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_409),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_409),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_SL g440 ( 
.A(n_428),
.B(n_282),
.Y(n_440)
);

BUFx3_ASAP7_75t_L g441 ( 
.A(n_414),
.Y(n_441)
);

AOI22xp33_ASAP7_75t_L g442 ( 
.A1(n_431),
.A2(n_280),
.B1(n_287),
.B2(n_286),
.Y(n_442)
);

INVx6_ASAP7_75t_L g443 ( 
.A(n_415),
.Y(n_443)
);

HB1xp67_ASAP7_75t_L g444 ( 
.A(n_430),
.Y(n_444)
);

INVx4_ASAP7_75t_L g445 ( 
.A(n_388),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_426),
.B(n_422),
.Y(n_446)
);

INVx2_ASAP7_75t_SL g447 ( 
.A(n_404),
.Y(n_447)
);

BUFx10_ASAP7_75t_L g448 ( 
.A(n_384),
.Y(n_448)
);

BUFx6f_ASAP7_75t_L g449 ( 
.A(n_383),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_393),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_426),
.B(n_289),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_L g452 ( 
.A(n_385),
.B(n_3),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_SL g453 ( 
.A(n_426),
.B(n_422),
.Y(n_453)
);

BUFx10_ASAP7_75t_L g454 ( 
.A(n_384),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_383),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_388),
.B(n_312),
.Y(n_456)
);

AND2x2_ASAP7_75t_L g457 ( 
.A(n_418),
.B(n_290),
.Y(n_457)
);

INVx4_ASAP7_75t_L g458 ( 
.A(n_388),
.Y(n_458)
);

AOI22xp33_ASAP7_75t_L g459 ( 
.A1(n_396),
.A2(n_280),
.B1(n_295),
.B2(n_291),
.Y(n_459)
);

AND3x2_ASAP7_75t_L g460 ( 
.A(n_425),
.B(n_4),
.C(n_5),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_412),
.B(n_312),
.Y(n_461)
);

AND2x2_ASAP7_75t_L g462 ( 
.A(n_396),
.B(n_304),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g463 ( 
.A(n_426),
.B(n_310),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_389),
.Y(n_464)
);

OR2x6_ASAP7_75t_L g465 ( 
.A(n_402),
.B(n_4),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_389),
.Y(n_466)
);

INVx5_ASAP7_75t_L g467 ( 
.A(n_412),
.Y(n_467)
);

OR2x6_ASAP7_75t_L g468 ( 
.A(n_411),
.B(n_5),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_399),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_399),
.Y(n_470)
);

AND2x2_ASAP7_75t_L g471 ( 
.A(n_396),
.B(n_313),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_412),
.B(n_312),
.Y(n_472)
);

AND2x4_ASAP7_75t_L g473 ( 
.A(n_415),
.B(n_6),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_400),
.Y(n_474)
);

AND2x2_ASAP7_75t_SL g475 ( 
.A(n_397),
.B(n_6),
.Y(n_475)
);

BUFx6f_ASAP7_75t_SL g476 ( 
.A(n_415),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_429),
.Y(n_477)
);

INVx4_ASAP7_75t_L g478 ( 
.A(n_422),
.Y(n_478)
);

AND2x2_ASAP7_75t_L g479 ( 
.A(n_421),
.B(n_315),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_424),
.B(n_312),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_419),
.Y(n_481)
);

AOI22xp33_ASAP7_75t_L g482 ( 
.A1(n_422),
.A2(n_314),
.B1(n_312),
.B2(n_322),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_400),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_401),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_401),
.Y(n_485)
);

BUFx8_ASAP7_75t_SL g486 ( 
.A(n_385),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_405),
.Y(n_487)
);

AOI22xp5_ASAP7_75t_L g488 ( 
.A1(n_420),
.A2(n_391),
.B1(n_406),
.B2(n_398),
.Y(n_488)
);

AOI22xp5_ASAP7_75t_L g489 ( 
.A1(n_408),
.A2(n_392),
.B1(n_417),
.B2(n_410),
.Y(n_489)
);

INVx3_ASAP7_75t_L g490 ( 
.A(n_410),
.Y(n_490)
);

INVx5_ASAP7_75t_L g491 ( 
.A(n_395),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_407),
.B(n_312),
.Y(n_492)
);

NAND3xp33_ASAP7_75t_SL g493 ( 
.A(n_407),
.B(n_333),
.C(n_328),
.Y(n_493)
);

INVx4_ASAP7_75t_L g494 ( 
.A(n_387),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_423),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_434),
.B(n_478),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_449),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_478),
.B(n_7),
.Y(n_498)
);

AOI22xp33_ASAP7_75t_L g499 ( 
.A1(n_475),
.A2(n_314),
.B1(n_423),
.B2(n_403),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_SL g500 ( 
.A(n_479),
.B(n_334),
.Y(n_500)
);

BUFx6f_ASAP7_75t_L g501 ( 
.A(n_449),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_445),
.B(n_314),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_449),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_445),
.B(n_314),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_490),
.Y(n_505)
);

INVxp67_ASAP7_75t_L g506 ( 
.A(n_486),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_458),
.B(n_314),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_489),
.B(n_8),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_490),
.Y(n_509)
);

AOI22xp5_ASAP7_75t_L g510 ( 
.A1(n_443),
.A2(n_403),
.B1(n_413),
.B2(n_394),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_433),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_451),
.B(n_8),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_447),
.B(n_9),
.Y(n_513)
);

AND2x2_ASAP7_75t_L g514 ( 
.A(n_441),
.B(n_394),
.Y(n_514)
);

AND2x2_ASAP7_75t_L g515 ( 
.A(n_444),
.B(n_413),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_443),
.B(n_10),
.Y(n_516)
);

AND2x6_ASAP7_75t_SL g517 ( 
.A(n_465),
.B(n_468),
.Y(n_517)
);

AOI22xp33_ASAP7_75t_L g518 ( 
.A1(n_473),
.A2(n_12),
.B1(n_10),
.B2(n_11),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_SL g519 ( 
.A(n_467),
.B(n_11),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_455),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_492),
.B(n_12),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_436),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_492),
.B(n_14),
.Y(n_523)
);

AOI22xp5_ASAP7_75t_L g524 ( 
.A1(n_443),
.A2(n_16),
.B1(n_14),
.B2(n_15),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_480),
.B(n_16),
.Y(n_525)
);

NOR3xp33_ASAP7_75t_L g526 ( 
.A(n_493),
.B(n_17),
.C(n_18),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_SL g527 ( 
.A(n_467),
.B(n_17),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_450),
.Y(n_528)
);

NAND2xp33_ASAP7_75t_SL g529 ( 
.A(n_476),
.B(n_18),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_435),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_SL g531 ( 
.A(n_491),
.B(n_19),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_464),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_480),
.B(n_466),
.Y(n_533)
);

INVx3_ASAP7_75t_L g534 ( 
.A(n_432),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_469),
.Y(n_535)
);

AOI22xp33_ASAP7_75t_L g536 ( 
.A1(n_473),
.A2(n_22),
.B1(n_20),
.B2(n_21),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_446),
.B(n_20),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_470),
.B(n_21),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_474),
.Y(n_539)
);

AND2x2_ASAP7_75t_L g540 ( 
.A(n_444),
.B(n_22),
.Y(n_540)
);

AOI22xp33_ASAP7_75t_L g541 ( 
.A1(n_483),
.A2(n_25),
.B1(n_23),
.B2(n_24),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_453),
.B(n_23),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_484),
.B(n_25),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_485),
.Y(n_544)
);

INVxp67_ASAP7_75t_L g545 ( 
.A(n_481),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_440),
.B(n_26),
.Y(n_546)
);

INVxp67_ASAP7_75t_L g547 ( 
.A(n_477),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_487),
.Y(n_548)
);

BUFx8_ASAP7_75t_L g549 ( 
.A(n_476),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_432),
.Y(n_550)
);

BUFx6f_ASAP7_75t_SL g551 ( 
.A(n_448),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_462),
.B(n_26),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_456),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_456),
.Y(n_554)
);

NAND3xp33_ASAP7_75t_L g555 ( 
.A(n_442),
.B(n_27),
.C(n_28),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_SL g556 ( 
.A(n_467),
.B(n_27),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_471),
.B(n_28),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_461),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_SL g559 ( 
.A(n_467),
.B(n_29),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_461),
.Y(n_560)
);

OAI221xp5_ASAP7_75t_L g561 ( 
.A1(n_459),
.A2(n_29),
.B1(n_30),
.B2(n_31),
.C(n_32),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_438),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_SL g563 ( 
.A(n_491),
.B(n_30),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_437),
.B(n_31),
.Y(n_564)
);

NOR3xp33_ASAP7_75t_L g565 ( 
.A(n_493),
.B(n_32),
.C(n_33),
.Y(n_565)
);

NAND2xp33_ASAP7_75t_L g566 ( 
.A(n_491),
.B(n_33),
.Y(n_566)
);

AOI21xp5_ASAP7_75t_L g567 ( 
.A1(n_496),
.A2(n_463),
.B(n_472),
.Y(n_567)
);

NAND2x1p5_ASAP7_75t_L g568 ( 
.A(n_514),
.B(n_491),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_511),
.B(n_457),
.Y(n_569)
);

AOI21xp5_ASAP7_75t_L g570 ( 
.A1(n_533),
.A2(n_504),
.B(n_502),
.Y(n_570)
);

OAI21xp5_ASAP7_75t_L g571 ( 
.A1(n_553),
.A2(n_482),
.B(n_488),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_522),
.B(n_528),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_516),
.B(n_482),
.Y(n_573)
);

BUFx4f_ASAP7_75t_L g574 ( 
.A(n_515),
.Y(n_574)
);

AOI21xp5_ASAP7_75t_L g575 ( 
.A1(n_507),
.A2(n_439),
.B(n_465),
.Y(n_575)
);

AOI21xp5_ASAP7_75t_L g576 ( 
.A1(n_554),
.A2(n_468),
.B(n_465),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_516),
.B(n_448),
.Y(n_577)
);

AOI21xp5_ASAP7_75t_L g578 ( 
.A1(n_558),
.A2(n_468),
.B(n_495),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_SL g579 ( 
.A(n_545),
.B(n_454),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_540),
.B(n_454),
.Y(n_580)
);

NOR2xp33_ASAP7_75t_L g581 ( 
.A(n_547),
.B(n_494),
.Y(n_581)
);

O2A1O1Ixp33_ASAP7_75t_L g582 ( 
.A1(n_561),
.A2(n_460),
.B(n_34),
.C(n_452),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_L g583 ( 
.A(n_510),
.B(n_494),
.Y(n_583)
);

AOI21xp5_ASAP7_75t_L g584 ( 
.A1(n_560),
.A2(n_460),
.B(n_36),
.Y(n_584)
);

AOI21xp5_ASAP7_75t_L g585 ( 
.A1(n_525),
.A2(n_38),
.B(n_35),
.Y(n_585)
);

AOI21xp5_ASAP7_75t_L g586 ( 
.A1(n_521),
.A2(n_40),
.B(n_39),
.Y(n_586)
);

AO221x2_ASAP7_75t_L g587 ( 
.A1(n_555),
.A2(n_34),
.B1(n_41),
.B2(n_42),
.C(n_43),
.Y(n_587)
);

AOI21xp5_ASAP7_75t_L g588 ( 
.A1(n_523),
.A2(n_44),
.B(n_46),
.Y(n_588)
);

A2O1A1Ixp33_ASAP7_75t_L g589 ( 
.A1(n_546),
.A2(n_47),
.B(n_48),
.C(n_49),
.Y(n_589)
);

A2O1A1Ixp33_ASAP7_75t_L g590 ( 
.A1(n_546),
.A2(n_50),
.B(n_51),
.C(n_52),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_508),
.B(n_53),
.Y(n_591)
);

BUFx6f_ASAP7_75t_L g592 ( 
.A(n_501),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_530),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_539),
.Y(n_594)
);

OR2x2_ASAP7_75t_L g595 ( 
.A(n_499),
.B(n_55),
.Y(n_595)
);

OAI22xp5_ASAP7_75t_L g596 ( 
.A1(n_518),
.A2(n_56),
.B1(n_57),
.B2(n_58),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_498),
.B(n_59),
.Y(n_597)
);

BUFx6f_ASAP7_75t_L g598 ( 
.A(n_501),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_498),
.B(n_60),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_544),
.B(n_61),
.Y(n_600)
);

OAI21x1_ASAP7_75t_L g601 ( 
.A1(n_562),
.A2(n_62),
.B(n_64),
.Y(n_601)
);

HB1xp67_ASAP7_75t_L g602 ( 
.A(n_549),
.Y(n_602)
);

AOI22xp33_ASAP7_75t_L g603 ( 
.A1(n_499),
.A2(n_65),
.B1(n_67),
.B2(n_68),
.Y(n_603)
);

INVx3_ASAP7_75t_L g604 ( 
.A(n_501),
.Y(n_604)
);

INVx1_ASAP7_75t_SL g605 ( 
.A(n_513),
.Y(n_605)
);

AOI22xp5_ASAP7_75t_L g606 ( 
.A1(n_512),
.A2(n_69),
.B1(n_70),
.B2(n_71),
.Y(n_606)
);

NOR2x1_ASAP7_75t_L g607 ( 
.A(n_500),
.B(n_72),
.Y(n_607)
);

NOR2xp67_ASAP7_75t_L g608 ( 
.A(n_506),
.B(n_73),
.Y(n_608)
);

NOR2x1_ASAP7_75t_L g609 ( 
.A(n_564),
.B(n_74),
.Y(n_609)
);

O2A1O1Ixp33_ASAP7_75t_SL g610 ( 
.A1(n_519),
.A2(n_77),
.B(n_78),
.C(n_79),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_548),
.B(n_80),
.Y(n_611)
);

AOI21xp5_ASAP7_75t_L g612 ( 
.A1(n_550),
.A2(n_82),
.B(n_84),
.Y(n_612)
);

NAND2x1p5_ASAP7_75t_L g613 ( 
.A(n_501),
.B(n_85),
.Y(n_613)
);

O2A1O1Ixp33_ASAP7_75t_L g614 ( 
.A1(n_566),
.A2(n_86),
.B(n_87),
.C(n_88),
.Y(n_614)
);

AOI21xp5_ASAP7_75t_L g615 ( 
.A1(n_534),
.A2(n_89),
.B(n_90),
.Y(n_615)
);

AOI21xp5_ASAP7_75t_L g616 ( 
.A1(n_534),
.A2(n_509),
.B(n_505),
.Y(n_616)
);

AOI21xp5_ASAP7_75t_L g617 ( 
.A1(n_497),
.A2(n_91),
.B(n_92),
.Y(n_617)
);

AOI21xp5_ASAP7_75t_L g618 ( 
.A1(n_503),
.A2(n_93),
.B(n_94),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_552),
.B(n_95),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_557),
.B(n_97),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_520),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_532),
.B(n_98),
.Y(n_622)
);

BUFx6f_ASAP7_75t_L g623 ( 
.A(n_535),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_537),
.B(n_99),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_537),
.B(n_100),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_SL g626 ( 
.A(n_518),
.B(n_102),
.Y(n_626)
);

OAI21xp5_ASAP7_75t_L g627 ( 
.A1(n_538),
.A2(n_104),
.B(n_106),
.Y(n_627)
);

OAI21xp5_ASAP7_75t_L g628 ( 
.A1(n_570),
.A2(n_542),
.B(n_543),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_L g629 ( 
.A(n_577),
.B(n_551),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_572),
.B(n_542),
.Y(n_630)
);

AOI21xp5_ASAP7_75t_L g631 ( 
.A1(n_597),
.A2(n_527),
.B(n_519),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_593),
.Y(n_632)
);

OAI21x1_ASAP7_75t_SL g633 ( 
.A1(n_575),
.A2(n_536),
.B(n_541),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_569),
.B(n_536),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_SL g635 ( 
.A(n_574),
.B(n_549),
.Y(n_635)
);

AOI21xp5_ASAP7_75t_L g636 ( 
.A1(n_599),
.A2(n_556),
.B(n_527),
.Y(n_636)
);

AOI21x1_ASAP7_75t_L g637 ( 
.A1(n_624),
.A2(n_559),
.B(n_556),
.Y(n_637)
);

AOI21xp5_ASAP7_75t_L g638 ( 
.A1(n_567),
.A2(n_563),
.B(n_531),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_605),
.B(n_526),
.Y(n_639)
);

OAI21x1_ASAP7_75t_L g640 ( 
.A1(n_601),
.A2(n_541),
.B(n_524),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_594),
.B(n_526),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_SL g642 ( 
.A(n_580),
.B(n_529),
.Y(n_642)
);

NOR2xp33_ASAP7_75t_L g643 ( 
.A(n_583),
.B(n_581),
.Y(n_643)
);

AOI21x1_ASAP7_75t_L g644 ( 
.A1(n_625),
.A2(n_565),
.B(n_517),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_SL g645 ( 
.A(n_576),
.B(n_565),
.Y(n_645)
);

OAI21xp5_ASAP7_75t_L g646 ( 
.A1(n_571),
.A2(n_573),
.B(n_616),
.Y(n_646)
);

OAI21x1_ASAP7_75t_L g647 ( 
.A1(n_622),
.A2(n_108),
.B(n_111),
.Y(n_647)
);

AOI221xp5_ASAP7_75t_L g648 ( 
.A1(n_582),
.A2(n_551),
.B1(n_113),
.B2(n_114),
.C(n_115),
.Y(n_648)
);

AO21x2_ASAP7_75t_L g649 ( 
.A1(n_591),
.A2(n_112),
.B(n_116),
.Y(n_649)
);

AND2x6_ASAP7_75t_L g650 ( 
.A(n_592),
.B(n_118),
.Y(n_650)
);

BUFx2_ASAP7_75t_L g651 ( 
.A(n_602),
.Y(n_651)
);

INVx5_ASAP7_75t_L g652 ( 
.A(n_592),
.Y(n_652)
);

HB1xp67_ASAP7_75t_L g653 ( 
.A(n_623),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_621),
.Y(n_654)
);

AOI21xp5_ASAP7_75t_SL g655 ( 
.A1(n_626),
.A2(n_120),
.B(n_121),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_578),
.B(n_122),
.Y(n_656)
);

BUFx3_ASAP7_75t_L g657 ( 
.A(n_568),
.Y(n_657)
);

A2O1A1Ixp33_ASAP7_75t_L g658 ( 
.A1(n_595),
.A2(n_124),
.B(n_126),
.C(n_127),
.Y(n_658)
);

OAI21x1_ASAP7_75t_L g659 ( 
.A1(n_600),
.A2(n_130),
.B(n_131),
.Y(n_659)
);

AOI21xp5_ASAP7_75t_L g660 ( 
.A1(n_619),
.A2(n_133),
.B(n_135),
.Y(n_660)
);

OAI21xp5_ASAP7_75t_L g661 ( 
.A1(n_611),
.A2(n_136),
.B(n_137),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_623),
.B(n_138),
.Y(n_662)
);

AND2x2_ASAP7_75t_SL g663 ( 
.A(n_603),
.B(n_139),
.Y(n_663)
);

OAI21x1_ASAP7_75t_L g664 ( 
.A1(n_627),
.A2(n_588),
.B(n_586),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_623),
.B(n_604),
.Y(n_665)
);

OAI21x1_ASAP7_75t_L g666 ( 
.A1(n_585),
.A2(n_140),
.B(n_141),
.Y(n_666)
);

OAI21x1_ASAP7_75t_SL g667 ( 
.A1(n_614),
.A2(n_596),
.B(n_584),
.Y(n_667)
);

AOI221x1_ASAP7_75t_L g668 ( 
.A1(n_589),
.A2(n_142),
.B1(n_143),
.B2(n_144),
.C(n_146),
.Y(n_668)
);

AOI21xp5_ASAP7_75t_L g669 ( 
.A1(n_620),
.A2(n_147),
.B(n_148),
.Y(n_669)
);

OR2x2_ASAP7_75t_L g670 ( 
.A(n_579),
.B(n_604),
.Y(n_670)
);

AOI21x1_ASAP7_75t_L g671 ( 
.A1(n_609),
.A2(n_150),
.B(n_151),
.Y(n_671)
);

OR2x2_ASAP7_75t_L g672 ( 
.A(n_592),
.B(n_153),
.Y(n_672)
);

INVx5_ASAP7_75t_L g673 ( 
.A(n_598),
.Y(n_673)
);

A2O1A1Ixp33_ASAP7_75t_L g674 ( 
.A1(n_607),
.A2(n_154),
.B(n_158),
.C(n_159),
.Y(n_674)
);

OAI22xp5_ASAP7_75t_L g675 ( 
.A1(n_598),
.A2(n_160),
.B1(n_161),
.B2(n_163),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_598),
.Y(n_676)
);

OAI21xp5_ASAP7_75t_L g677 ( 
.A1(n_615),
.A2(n_164),
.B(n_165),
.Y(n_677)
);

OAI21x1_ASAP7_75t_L g678 ( 
.A1(n_613),
.A2(n_166),
.B(n_167),
.Y(n_678)
);

A2O1A1Ixp33_ASAP7_75t_L g679 ( 
.A1(n_590),
.A2(n_606),
.B(n_608),
.C(n_612),
.Y(n_679)
);

OAI21xp5_ASAP7_75t_L g680 ( 
.A1(n_617),
.A2(n_168),
.B(n_169),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_587),
.B(n_171),
.Y(n_681)
);

AO31x2_ASAP7_75t_L g682 ( 
.A1(n_618),
.A2(n_172),
.A3(n_173),
.B(n_174),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_587),
.Y(n_683)
);

AOI221x1_ASAP7_75t_L g684 ( 
.A1(n_610),
.A2(n_175),
.B1(n_176),
.B2(n_178),
.C(n_179),
.Y(n_684)
);

AO31x2_ASAP7_75t_L g685 ( 
.A1(n_570),
.A2(n_181),
.A3(n_182),
.B(n_183),
.Y(n_685)
);

A2O1A1Ixp33_ASAP7_75t_L g686 ( 
.A1(n_582),
.A2(n_184),
.B(n_185),
.C(n_187),
.Y(n_686)
);

AND2x4_ASAP7_75t_L g687 ( 
.A(n_657),
.B(n_191),
.Y(n_687)
);

BUFx10_ASAP7_75t_L g688 ( 
.A(n_629),
.Y(n_688)
);

BUFx8_ASAP7_75t_L g689 ( 
.A(n_651),
.Y(n_689)
);

INVx2_ASAP7_75t_SL g690 ( 
.A(n_635),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_654),
.Y(n_691)
);

INVx2_ASAP7_75t_SL g692 ( 
.A(n_670),
.Y(n_692)
);

AOI21xp5_ASAP7_75t_L g693 ( 
.A1(n_628),
.A2(n_193),
.B(n_194),
.Y(n_693)
);

OR2x6_ASAP7_75t_L g694 ( 
.A(n_653),
.B(n_274),
.Y(n_694)
);

AND2x4_ASAP7_75t_L g695 ( 
.A(n_652),
.B(n_195),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_643),
.B(n_272),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_632),
.Y(n_697)
);

BUFx2_ASAP7_75t_L g698 ( 
.A(n_676),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_641),
.Y(n_699)
);

CKINVDCx11_ASAP7_75t_R g700 ( 
.A(n_676),
.Y(n_700)
);

OR2x2_ASAP7_75t_L g701 ( 
.A(n_639),
.B(n_197),
.Y(n_701)
);

AO32x1_ASAP7_75t_L g702 ( 
.A1(n_683),
.A2(n_200),
.A3(n_201),
.B1(n_202),
.B2(n_203),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_634),
.Y(n_703)
);

INVx5_ASAP7_75t_L g704 ( 
.A(n_650),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_665),
.Y(n_705)
);

INVx1_ASAP7_75t_SL g706 ( 
.A(n_672),
.Y(n_706)
);

BUFx6f_ASAP7_75t_L g707 ( 
.A(n_652),
.Y(n_707)
);

INVx3_ASAP7_75t_L g708 ( 
.A(n_652),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_630),
.B(n_271),
.Y(n_709)
);

INVxp67_ASAP7_75t_SL g710 ( 
.A(n_645),
.Y(n_710)
);

AOI21xp5_ASAP7_75t_L g711 ( 
.A1(n_631),
.A2(n_636),
.B(n_679),
.Y(n_711)
);

AND2x2_ASAP7_75t_L g712 ( 
.A(n_644),
.B(n_205),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_642),
.B(n_270),
.Y(n_713)
);

INVx3_ASAP7_75t_L g714 ( 
.A(n_673),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_673),
.B(n_207),
.Y(n_715)
);

NAND2x1p5_ASAP7_75t_L g716 ( 
.A(n_673),
.B(n_208),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_662),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_663),
.B(n_648),
.Y(n_718)
);

NOR2xp67_ASAP7_75t_SL g719 ( 
.A(n_681),
.B(n_209),
.Y(n_719)
);

INVx4_ASAP7_75t_L g720 ( 
.A(n_650),
.Y(n_720)
);

AOI21xp5_ASAP7_75t_L g721 ( 
.A1(n_664),
.A2(n_210),
.B(n_211),
.Y(n_721)
);

INVxp67_ASAP7_75t_L g722 ( 
.A(n_656),
.Y(n_722)
);

BUFx12f_ASAP7_75t_L g723 ( 
.A(n_650),
.Y(n_723)
);

AND2x4_ASAP7_75t_L g724 ( 
.A(n_650),
.B(n_269),
.Y(n_724)
);

INVx3_ASAP7_75t_L g725 ( 
.A(n_671),
.Y(n_725)
);

INVx5_ASAP7_75t_L g726 ( 
.A(n_655),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_633),
.Y(n_727)
);

OAI22xp5_ASAP7_75t_L g728 ( 
.A1(n_638),
.A2(n_212),
.B1(n_214),
.B2(n_215),
.Y(n_728)
);

BUFx3_ASAP7_75t_L g729 ( 
.A(n_678),
.Y(n_729)
);

BUFx6f_ASAP7_75t_L g730 ( 
.A(n_659),
.Y(n_730)
);

AOI21xp5_ASAP7_75t_L g731 ( 
.A1(n_667),
.A2(n_216),
.B(n_218),
.Y(n_731)
);

OR2x6_ASAP7_75t_L g732 ( 
.A(n_686),
.B(n_658),
.Y(n_732)
);

AND2x2_ASAP7_75t_L g733 ( 
.A(n_646),
.B(n_685),
.Y(n_733)
);

BUFx3_ASAP7_75t_L g734 ( 
.A(n_647),
.Y(n_734)
);

AOI21xp5_ASAP7_75t_L g735 ( 
.A1(n_677),
.A2(n_661),
.B(n_680),
.Y(n_735)
);

BUFx6f_ASAP7_75t_L g736 ( 
.A(n_666),
.Y(n_736)
);

OA21x2_ASAP7_75t_L g737 ( 
.A1(n_711),
.A2(n_668),
.B(n_684),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_691),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_697),
.Y(n_739)
);

CKINVDCx11_ASAP7_75t_R g740 ( 
.A(n_688),
.Y(n_740)
);

INVx3_ASAP7_75t_L g741 ( 
.A(n_720),
.Y(n_741)
);

INVx1_ASAP7_75t_SL g742 ( 
.A(n_706),
.Y(n_742)
);

INVx3_ASAP7_75t_L g743 ( 
.A(n_720),
.Y(n_743)
);

BUFx12f_ASAP7_75t_L g744 ( 
.A(n_689),
.Y(n_744)
);

INVx3_ASAP7_75t_L g745 ( 
.A(n_704),
.Y(n_745)
);

INVx1_ASAP7_75t_SL g746 ( 
.A(n_698),
.Y(n_746)
);

INVx3_ASAP7_75t_L g747 ( 
.A(n_704),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_705),
.Y(n_748)
);

CKINVDCx6p67_ASAP7_75t_R g749 ( 
.A(n_700),
.Y(n_749)
);

OR2x6_ASAP7_75t_L g750 ( 
.A(n_723),
.B(n_640),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_692),
.Y(n_751)
);

OAI22xp5_ASAP7_75t_L g752 ( 
.A1(n_718),
.A2(n_637),
.B1(n_674),
.B2(n_669),
.Y(n_752)
);

OAI21x1_ASAP7_75t_SL g753 ( 
.A1(n_735),
.A2(n_660),
.B(n_675),
.Y(n_753)
);

AOI22xp33_ASAP7_75t_L g754 ( 
.A1(n_699),
.A2(n_717),
.B1(n_703),
.B2(n_732),
.Y(n_754)
);

AOI22xp33_ASAP7_75t_L g755 ( 
.A1(n_732),
.A2(n_696),
.B1(n_722),
.B2(n_704),
.Y(n_755)
);

CKINVDCx11_ASAP7_75t_R g756 ( 
.A(n_688),
.Y(n_756)
);

AND2x2_ASAP7_75t_L g757 ( 
.A(n_690),
.B(n_685),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_698),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_710),
.Y(n_759)
);

BUFx6f_ASAP7_75t_L g760 ( 
.A(n_707),
.Y(n_760)
);

INVx3_ASAP7_75t_L g761 ( 
.A(n_707),
.Y(n_761)
);

OAI22xp5_ASAP7_75t_L g762 ( 
.A1(n_701),
.A2(n_685),
.B1(n_682),
.B2(n_649),
.Y(n_762)
);

AO21x2_ASAP7_75t_L g763 ( 
.A1(n_733),
.A2(n_682),
.B(n_220),
.Y(n_763)
);

INVx8_ASAP7_75t_L g764 ( 
.A(n_694),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_727),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_687),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_694),
.Y(n_767)
);

AOI22xp33_ASAP7_75t_L g768 ( 
.A1(n_709),
.A2(n_682),
.B1(n_221),
.B2(n_222),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_707),
.B(n_219),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_712),
.Y(n_770)
);

OAI22xp5_ASAP7_75t_L g771 ( 
.A1(n_724),
.A2(n_223),
.B1(n_224),
.B2(n_225),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_689),
.Y(n_772)
);

AND2x4_ASAP7_75t_L g773 ( 
.A(n_708),
.B(n_228),
.Y(n_773)
);

BUFx6f_ASAP7_75t_L g774 ( 
.A(n_714),
.Y(n_774)
);

INVx3_ASAP7_75t_L g775 ( 
.A(n_695),
.Y(n_775)
);

CKINVDCx20_ASAP7_75t_R g776 ( 
.A(n_715),
.Y(n_776)
);

NAND2x1p5_ASAP7_75t_L g777 ( 
.A(n_724),
.B(n_229),
.Y(n_777)
);

BUFx6f_ASAP7_75t_L g778 ( 
.A(n_695),
.Y(n_778)
);

BUFx8_ASAP7_75t_SL g779 ( 
.A(n_713),
.Y(n_779)
);

AND2x4_ASAP7_75t_L g780 ( 
.A(n_726),
.B(n_231),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_716),
.Y(n_781)
);

HB1xp67_ASAP7_75t_SL g782 ( 
.A(n_729),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_719),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_719),
.Y(n_784)
);

OAI22xp5_ASAP7_75t_L g785 ( 
.A1(n_731),
.A2(n_232),
.B1(n_233),
.B2(n_234),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_725),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_726),
.Y(n_787)
);

AND2x2_ASAP7_75t_L g788 ( 
.A(n_693),
.B(n_235),
.Y(n_788)
);

CKINVDCx5p33_ASAP7_75t_R g789 ( 
.A(n_726),
.Y(n_789)
);

AOI22xp33_ASAP7_75t_L g790 ( 
.A1(n_728),
.A2(n_236),
.B1(n_237),
.B2(n_240),
.Y(n_790)
);

BUFx6f_ASAP7_75t_L g791 ( 
.A(n_734),
.Y(n_791)
);

OA21x2_ASAP7_75t_L g792 ( 
.A1(n_721),
.A2(n_241),
.B(n_244),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_730),
.Y(n_793)
);

CKINVDCx11_ASAP7_75t_R g794 ( 
.A(n_730),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_730),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_746),
.B(n_736),
.Y(n_796)
);

AND2x2_ASAP7_75t_L g797 ( 
.A(n_758),
.B(n_746),
.Y(n_797)
);

HB1xp67_ASAP7_75t_L g798 ( 
.A(n_759),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_765),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_786),
.Y(n_800)
);

INVx3_ASAP7_75t_L g801 ( 
.A(n_791),
.Y(n_801)
);

INVx2_ASAP7_75t_SL g802 ( 
.A(n_791),
.Y(n_802)
);

BUFx3_ASAP7_75t_L g803 ( 
.A(n_794),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_738),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_795),
.Y(n_805)
);

OAI21x1_ASAP7_75t_L g806 ( 
.A1(n_753),
.A2(n_736),
.B(n_702),
.Y(n_806)
);

HB1xp67_ASAP7_75t_L g807 ( 
.A(n_748),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_793),
.Y(n_808)
);

AND2x2_ASAP7_75t_L g809 ( 
.A(n_757),
.B(n_736),
.Y(n_809)
);

OAI21x1_ASAP7_75t_L g810 ( 
.A1(n_762),
.A2(n_702),
.B(n_246),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_791),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_750),
.Y(n_812)
);

INVx2_ASAP7_75t_SL g813 ( 
.A(n_783),
.Y(n_813)
);

BUFx3_ASAP7_75t_L g814 ( 
.A(n_787),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_763),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_750),
.Y(n_816)
);

AO21x2_ASAP7_75t_L g817 ( 
.A1(n_762),
.A2(n_245),
.B(n_247),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_763),
.Y(n_818)
);

OA21x2_ASAP7_75t_L g819 ( 
.A1(n_784),
.A2(n_248),
.B(n_249),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_750),
.Y(n_820)
);

INVx2_ASAP7_75t_SL g821 ( 
.A(n_741),
.Y(n_821)
);

OA21x2_ASAP7_75t_L g822 ( 
.A1(n_770),
.A2(n_250),
.B(n_251),
.Y(n_822)
);

AO21x2_ASAP7_75t_L g823 ( 
.A1(n_752),
.A2(n_252),
.B(n_254),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_739),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_782),
.Y(n_825)
);

INVx2_ASAP7_75t_L g826 ( 
.A(n_737),
.Y(n_826)
);

OAI21xp5_ASAP7_75t_L g827 ( 
.A1(n_752),
.A2(n_255),
.B(n_257),
.Y(n_827)
);

INVxp33_ASAP7_75t_L g828 ( 
.A(n_740),
.Y(n_828)
);

AND2x2_ASAP7_75t_L g829 ( 
.A(n_775),
.B(n_258),
.Y(n_829)
);

INVx3_ASAP7_75t_L g830 ( 
.A(n_741),
.Y(n_830)
);

HB1xp67_ASAP7_75t_L g831 ( 
.A(n_782),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_737),
.Y(n_832)
);

AND2x2_ASAP7_75t_L g833 ( 
.A(n_775),
.B(n_259),
.Y(n_833)
);

INVx3_ASAP7_75t_L g834 ( 
.A(n_743),
.Y(n_834)
);

AND2x4_ASAP7_75t_L g835 ( 
.A(n_745),
.B(n_747),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_792),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_777),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_792),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_745),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_777),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_747),
.Y(n_841)
);

OR2x6_ASAP7_75t_L g842 ( 
.A(n_764),
.B(n_260),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_743),
.Y(n_843)
);

AND2x2_ASAP7_75t_L g844 ( 
.A(n_754),
.B(n_261),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_769),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_799),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_807),
.B(n_742),
.Y(n_847)
);

INVx3_ASAP7_75t_L g848 ( 
.A(n_839),
.Y(n_848)
);

AND2x2_ASAP7_75t_L g849 ( 
.A(n_809),
.B(n_755),
.Y(n_849)
);

AND2x2_ASAP7_75t_L g850 ( 
.A(n_809),
.B(n_742),
.Y(n_850)
);

INVx2_ASAP7_75t_SL g851 ( 
.A(n_811),
.Y(n_851)
);

AND2x4_ASAP7_75t_L g852 ( 
.A(n_825),
.B(n_767),
.Y(n_852)
);

OR2x2_ASAP7_75t_L g853 ( 
.A(n_797),
.B(n_798),
.Y(n_853)
);

AND2x2_ASAP7_75t_L g854 ( 
.A(n_797),
.B(n_749),
.Y(n_854)
);

INVx3_ASAP7_75t_L g855 ( 
.A(n_839),
.Y(n_855)
);

AND2x2_ASAP7_75t_L g856 ( 
.A(n_804),
.B(n_800),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_799),
.Y(n_857)
);

OR2x2_ASAP7_75t_L g858 ( 
.A(n_800),
.B(n_751),
.Y(n_858)
);

NAND3xp33_ASAP7_75t_L g859 ( 
.A(n_827),
.B(n_768),
.C(n_771),
.Y(n_859)
);

OR2x2_ASAP7_75t_L g860 ( 
.A(n_813),
.B(n_764),
.Y(n_860)
);

AND2x2_ASAP7_75t_L g861 ( 
.A(n_804),
.B(n_788),
.Y(n_861)
);

AND2x2_ASAP7_75t_L g862 ( 
.A(n_805),
.B(n_756),
.Y(n_862)
);

HB1xp67_ASAP7_75t_L g863 ( 
.A(n_813),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_813),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_845),
.B(n_776),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_845),
.B(n_764),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_831),
.B(n_825),
.Y(n_867)
);

INVx3_ASAP7_75t_L g868 ( 
.A(n_839),
.Y(n_868)
);

AND2x2_ASAP7_75t_L g869 ( 
.A(n_805),
.B(n_761),
.Y(n_869)
);

CKINVDCx5p33_ASAP7_75t_R g870 ( 
.A(n_803),
.Y(n_870)
);

AND2x2_ASAP7_75t_L g871 ( 
.A(n_808),
.B(n_832),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_824),
.Y(n_872)
);

AND2x2_ASAP7_75t_L g873 ( 
.A(n_808),
.B(n_761),
.Y(n_873)
);

NOR2xp33_ASAP7_75t_L g874 ( 
.A(n_828),
.B(n_772),
.Y(n_874)
);

AND2x2_ASAP7_75t_L g875 ( 
.A(n_832),
.B(n_774),
.Y(n_875)
);

INVx4_ASAP7_75t_L g876 ( 
.A(n_817),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_826),
.Y(n_877)
);

NAND2xp33_ASAP7_75t_L g878 ( 
.A(n_821),
.B(n_789),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_826),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_831),
.B(n_774),
.Y(n_880)
);

AND2x2_ASAP7_75t_L g881 ( 
.A(n_826),
.B(n_774),
.Y(n_881)
);

AND2x2_ASAP7_75t_L g882 ( 
.A(n_796),
.B(n_766),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_802),
.B(n_760),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_836),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_796),
.Y(n_885)
);

INVx2_ASAP7_75t_SL g886 ( 
.A(n_811),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_812),
.Y(n_887)
);

INVx2_ASAP7_75t_L g888 ( 
.A(n_836),
.Y(n_888)
);

AND2x4_ASAP7_75t_L g889 ( 
.A(n_811),
.B(n_778),
.Y(n_889)
);

INVx2_ASAP7_75t_SL g890 ( 
.A(n_802),
.Y(n_890)
);

HB1xp67_ASAP7_75t_L g891 ( 
.A(n_841),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_812),
.Y(n_892)
);

AOI211xp5_ASAP7_75t_L g893 ( 
.A1(n_859),
.A2(n_827),
.B(n_771),
.C(n_785),
.Y(n_893)
);

NAND3xp33_ASAP7_75t_L g894 ( 
.A(n_876),
.B(n_843),
.C(n_840),
.Y(n_894)
);

NOR3xp33_ASAP7_75t_L g895 ( 
.A(n_876),
.B(n_859),
.C(n_867),
.Y(n_895)
);

OA211x2_ASAP7_75t_L g896 ( 
.A1(n_880),
.A2(n_803),
.B(n_823),
.C(n_814),
.Y(n_896)
);

OAI221xp5_ASAP7_75t_L g897 ( 
.A1(n_876),
.A2(n_865),
.B1(n_866),
.B2(n_858),
.C(n_847),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_885),
.B(n_821),
.Y(n_898)
);

AND2x2_ASAP7_75t_L g899 ( 
.A(n_850),
.B(n_803),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_885),
.B(n_821),
.Y(n_900)
);

NOR2xp33_ASAP7_75t_L g901 ( 
.A(n_870),
.B(n_744),
.Y(n_901)
);

AND2x2_ASAP7_75t_L g902 ( 
.A(n_850),
.B(n_814),
.Y(n_902)
);

AND2x2_ASAP7_75t_SL g903 ( 
.A(n_878),
.B(n_840),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_853),
.B(n_801),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_853),
.B(n_801),
.Y(n_905)
);

OAI21xp5_ASAP7_75t_L g906 ( 
.A1(n_876),
.A2(n_810),
.B(n_819),
.Y(n_906)
);

AND2x2_ASAP7_75t_L g907 ( 
.A(n_854),
.B(n_814),
.Y(n_907)
);

OAI221xp5_ASAP7_75t_SL g908 ( 
.A1(n_861),
.A2(n_842),
.B1(n_860),
.B2(n_844),
.C(n_790),
.Y(n_908)
);

OAI21xp5_ASAP7_75t_SL g909 ( 
.A1(n_854),
.A2(n_844),
.B(n_785),
.Y(n_909)
);

AOI211xp5_ASAP7_75t_L g910 ( 
.A1(n_861),
.A2(n_860),
.B(n_862),
.C(n_875),
.Y(n_910)
);

AND2x2_ASAP7_75t_L g911 ( 
.A(n_862),
.B(n_801),
.Y(n_911)
);

OAI221xp5_ASAP7_75t_L g912 ( 
.A1(n_858),
.A2(n_816),
.B1(n_820),
.B2(n_837),
.C(n_842),
.Y(n_912)
);

NOR3xp33_ASAP7_75t_L g913 ( 
.A(n_883),
.B(n_837),
.C(n_801),
.Y(n_913)
);

OAI221xp5_ASAP7_75t_SL g914 ( 
.A1(n_864),
.A2(n_842),
.B1(n_838),
.B2(n_836),
.C(n_823),
.Y(n_914)
);

NAND3xp33_ASAP7_75t_L g915 ( 
.A(n_864),
.B(n_843),
.C(n_816),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_856),
.B(n_843),
.Y(n_916)
);

OAI21xp5_ASAP7_75t_SL g917 ( 
.A1(n_874),
.A2(n_830),
.B(n_834),
.Y(n_917)
);

NAND4xp25_ASAP7_75t_L g918 ( 
.A(n_846),
.B(n_830),
.C(n_834),
.D(n_820),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_SL g919 ( 
.A(n_870),
.B(n_802),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_856),
.B(n_841),
.Y(n_920)
);

AOI221xp5_ASAP7_75t_L g921 ( 
.A1(n_846),
.A2(n_823),
.B1(n_817),
.B2(n_857),
.C(n_871),
.Y(n_921)
);

OAI22xp5_ASAP7_75t_L g922 ( 
.A1(n_852),
.A2(n_842),
.B1(n_781),
.B2(n_778),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_871),
.B(n_830),
.Y(n_923)
);

NAND4xp25_ASAP7_75t_L g924 ( 
.A(n_857),
.B(n_869),
.C(n_873),
.D(n_852),
.Y(n_924)
);

AOI22xp33_ASAP7_75t_L g925 ( 
.A1(n_849),
.A2(n_817),
.B1(n_823),
.B2(n_818),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_869),
.B(n_873),
.Y(n_926)
);

NOR2xp33_ASAP7_75t_L g927 ( 
.A(n_901),
.B(n_779),
.Y(n_927)
);

OR2x2_ASAP7_75t_L g928 ( 
.A(n_920),
.B(n_863),
.Y(n_928)
);

AND2x4_ASAP7_75t_SL g929 ( 
.A(n_907),
.B(n_852),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_898),
.Y(n_930)
);

INVx2_ASAP7_75t_L g931 ( 
.A(n_915),
.Y(n_931)
);

INVx2_ASAP7_75t_L g932 ( 
.A(n_900),
.Y(n_932)
);

AND2x2_ASAP7_75t_L g933 ( 
.A(n_902),
.B(n_899),
.Y(n_933)
);

AND2x2_ASAP7_75t_L g934 ( 
.A(n_910),
.B(n_852),
.Y(n_934)
);

AND2x2_ASAP7_75t_L g935 ( 
.A(n_911),
.B(n_875),
.Y(n_935)
);

INVx2_ASAP7_75t_L g936 ( 
.A(n_916),
.Y(n_936)
);

AND2x2_ASAP7_75t_L g937 ( 
.A(n_895),
.B(n_848),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_904),
.Y(n_938)
);

AND2x2_ASAP7_75t_L g939 ( 
.A(n_926),
.B(n_848),
.Y(n_939)
);

AND2x2_ASAP7_75t_L g940 ( 
.A(n_905),
.B(n_848),
.Y(n_940)
);

AND2x2_ASAP7_75t_L g941 ( 
.A(n_923),
.B(n_906),
.Y(n_941)
);

INVx2_ASAP7_75t_L g942 ( 
.A(n_894),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_913),
.B(n_891),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_924),
.Y(n_944)
);

AND2x2_ASAP7_75t_L g945 ( 
.A(n_917),
.B(n_855),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_SL g946 ( 
.A(n_903),
.B(n_890),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_918),
.Y(n_947)
);

AND2x2_ASAP7_75t_L g948 ( 
.A(n_921),
.B(n_855),
.Y(n_948)
);

AND2x4_ASAP7_75t_SL g949 ( 
.A(n_925),
.B(n_889),
.Y(n_949)
);

INVx2_ASAP7_75t_L g950 ( 
.A(n_897),
.Y(n_950)
);

HB1xp67_ASAP7_75t_L g951 ( 
.A(n_896),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_912),
.Y(n_952)
);

INVx2_ASAP7_75t_SL g953 ( 
.A(n_919),
.Y(n_953)
);

INVx2_ASAP7_75t_L g954 ( 
.A(n_922),
.Y(n_954)
);

NOR2xp33_ASAP7_75t_L g955 ( 
.A(n_931),
.B(n_909),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_931),
.B(n_921),
.Y(n_956)
);

AND2x2_ASAP7_75t_L g957 ( 
.A(n_934),
.B(n_890),
.Y(n_957)
);

INVx2_ASAP7_75t_SL g958 ( 
.A(n_929),
.Y(n_958)
);

AND2x2_ASAP7_75t_L g959 ( 
.A(n_934),
.B(n_868),
.Y(n_959)
);

HB1xp67_ASAP7_75t_L g960 ( 
.A(n_942),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_930),
.B(n_887),
.Y(n_961)
);

INVx2_ASAP7_75t_L g962 ( 
.A(n_932),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_938),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_928),
.Y(n_964)
);

OR2x2_ASAP7_75t_L g965 ( 
.A(n_928),
.B(n_892),
.Y(n_965)
);

AND2x2_ASAP7_75t_L g966 ( 
.A(n_929),
.B(n_881),
.Y(n_966)
);

AND2x2_ASAP7_75t_L g967 ( 
.A(n_933),
.B(n_881),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_947),
.B(n_887),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_936),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_968),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_960),
.Y(n_971)
);

AND2x2_ASAP7_75t_L g972 ( 
.A(n_958),
.B(n_964),
.Y(n_972)
);

INVxp67_ASAP7_75t_L g973 ( 
.A(n_955),
.Y(n_973)
);

AND2x2_ASAP7_75t_L g974 ( 
.A(n_958),
.B(n_941),
.Y(n_974)
);

INVx1_ASAP7_75t_SL g975 ( 
.A(n_960),
.Y(n_975)
);

INVxp67_ASAP7_75t_L g976 ( 
.A(n_955),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_963),
.Y(n_977)
);

AND2x2_ASAP7_75t_L g978 ( 
.A(n_959),
.B(n_941),
.Y(n_978)
);

NOR2x1p5_ASAP7_75t_SL g979 ( 
.A(n_962),
.B(n_942),
.Y(n_979)
);

INVxp67_ASAP7_75t_SL g980 ( 
.A(n_956),
.Y(n_980)
);

INVxp67_ASAP7_75t_L g981 ( 
.A(n_972),
.Y(n_981)
);

INVx2_ASAP7_75t_SL g982 ( 
.A(n_972),
.Y(n_982)
);

HB1xp67_ASAP7_75t_L g983 ( 
.A(n_971),
.Y(n_983)
);

OR2x2_ASAP7_75t_L g984 ( 
.A(n_975),
.B(n_965),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_977),
.Y(n_985)
);

OR2x2_ASAP7_75t_L g986 ( 
.A(n_970),
.B(n_944),
.Y(n_986)
);

NOR2xp33_ASAP7_75t_L g987 ( 
.A(n_973),
.B(n_927),
.Y(n_987)
);

AOI22xp33_ASAP7_75t_L g988 ( 
.A1(n_986),
.A2(n_980),
.B1(n_976),
.B2(n_950),
.Y(n_988)
);

AND2x4_ASAP7_75t_L g989 ( 
.A(n_982),
.B(n_974),
.Y(n_989)
);

NOR2x1_ASAP7_75t_L g990 ( 
.A(n_987),
.B(n_974),
.Y(n_990)
);

AOI22xp5_ASAP7_75t_L g991 ( 
.A1(n_981),
.A2(n_950),
.B1(n_952),
.B2(n_948),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_983),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_990),
.B(n_985),
.Y(n_993)
);

AND2x2_ASAP7_75t_L g994 ( 
.A(n_989),
.B(n_984),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_988),
.B(n_979),
.Y(n_995)
);

OR2x2_ASAP7_75t_L g996 ( 
.A(n_992),
.B(n_978),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_991),
.Y(n_997)
);

AOI21xp5_ASAP7_75t_L g998 ( 
.A1(n_995),
.A2(n_951),
.B(n_893),
.Y(n_998)
);

NOR2xp33_ASAP7_75t_L g999 ( 
.A(n_994),
.B(n_947),
.Y(n_999)
);

AOI221xp5_ASAP7_75t_L g1000 ( 
.A1(n_997),
.A2(n_914),
.B1(n_948),
.B2(n_908),
.C(n_937),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_996),
.Y(n_1001)
);

OAI221xp5_ASAP7_75t_SL g1002 ( 
.A1(n_993),
.A2(n_978),
.B1(n_937),
.B2(n_954),
.C(n_842),
.Y(n_1002)
);

NOR2x1_ASAP7_75t_L g1003 ( 
.A(n_993),
.B(n_842),
.Y(n_1003)
);

AOI221xp5_ASAP7_75t_L g1004 ( 
.A1(n_995),
.A2(n_914),
.B1(n_908),
.B2(n_949),
.C(n_943),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_1001),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_999),
.B(n_959),
.Y(n_1006)
);

AOI211x1_ASAP7_75t_L g1007 ( 
.A1(n_998),
.A2(n_946),
.B(n_957),
.C(n_961),
.Y(n_1007)
);

HB1xp67_ASAP7_75t_L g1008 ( 
.A(n_1003),
.Y(n_1008)
);

INVx1_ASAP7_75t_SL g1009 ( 
.A(n_1002),
.Y(n_1009)
);

NOR3xp33_ASAP7_75t_L g1010 ( 
.A(n_1004),
.B(n_954),
.C(n_962),
.Y(n_1010)
);

OAI211xp5_ASAP7_75t_SL g1011 ( 
.A1(n_1005),
.A2(n_1000),
.B(n_953),
.C(n_932),
.Y(n_1011)
);

AOI22xp5_ASAP7_75t_L g1012 ( 
.A1(n_1009),
.A2(n_817),
.B1(n_949),
.B2(n_953),
.Y(n_1012)
);

INVx3_ASAP7_75t_L g1013 ( 
.A(n_1006),
.Y(n_1013)
);

NOR2xp33_ASAP7_75t_L g1014 ( 
.A(n_1008),
.B(n_969),
.Y(n_1014)
);

AND2x2_ASAP7_75t_L g1015 ( 
.A(n_1010),
.B(n_933),
.Y(n_1015)
);

OAI211xp5_ASAP7_75t_L g1016 ( 
.A1(n_1007),
.A2(n_945),
.B(n_819),
.C(n_966),
.Y(n_1016)
);

NOR2xp33_ASAP7_75t_L g1017 ( 
.A(n_1006),
.B(n_967),
.Y(n_1017)
);

NOR2x1_ASAP7_75t_L g1018 ( 
.A(n_1005),
.B(n_773),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_SL g1019 ( 
.A(n_1013),
.B(n_1018),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_SL g1020 ( 
.A(n_1012),
.B(n_945),
.Y(n_1020)
);

AND2x4_ASAP7_75t_L g1021 ( 
.A(n_1015),
.B(n_935),
.Y(n_1021)
);

INVxp67_ASAP7_75t_SL g1022 ( 
.A(n_1014),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_1017),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_1011),
.Y(n_1024)
);

NOR3xp33_ASAP7_75t_SL g1025 ( 
.A(n_1016),
.B(n_769),
.C(n_892),
.Y(n_1025)
);

HB1xp67_ASAP7_75t_L g1026 ( 
.A(n_1013),
.Y(n_1026)
);

INVx2_ASAP7_75t_L g1027 ( 
.A(n_1013),
.Y(n_1027)
);

AOI22xp5_ASAP7_75t_L g1028 ( 
.A1(n_1012),
.A2(n_936),
.B1(n_778),
.B2(n_819),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_1013),
.Y(n_1029)
);

NOR2x1p5_ASAP7_75t_L g1030 ( 
.A(n_1013),
.B(n_830),
.Y(n_1030)
);

OAI22xp5_ASAP7_75t_L g1031 ( 
.A1(n_1013),
.A2(n_939),
.B1(n_940),
.B2(n_935),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_1013),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_1013),
.Y(n_1033)
);

AND2x4_ASAP7_75t_L g1034 ( 
.A(n_1013),
.B(n_939),
.Y(n_1034)
);

AND2x4_ASAP7_75t_L g1035 ( 
.A(n_1027),
.B(n_940),
.Y(n_1035)
);

NOR4xp25_ASAP7_75t_L g1036 ( 
.A(n_1029),
.B(n_829),
.C(n_833),
.D(n_851),
.Y(n_1036)
);

OR2x2_ASAP7_75t_L g1037 ( 
.A(n_1026),
.B(n_868),
.Y(n_1037)
);

HB1xp67_ASAP7_75t_L g1038 ( 
.A(n_1032),
.Y(n_1038)
);

AND3x2_ASAP7_75t_L g1039 ( 
.A(n_1022),
.B(n_773),
.C(n_780),
.Y(n_1039)
);

NAND3x1_ASAP7_75t_L g1040 ( 
.A(n_1033),
.B(n_834),
.C(n_829),
.Y(n_1040)
);

INVx1_ASAP7_75t_SL g1041 ( 
.A(n_1019),
.Y(n_1041)
);

AND2x4_ASAP7_75t_L g1042 ( 
.A(n_1023),
.B(n_834),
.Y(n_1042)
);

CKINVDCx5p33_ASAP7_75t_R g1043 ( 
.A(n_1024),
.Y(n_1043)
);

OAI322xp33_ASAP7_75t_SL g1044 ( 
.A1(n_1020),
.A2(n_838),
.A3(n_888),
.B1(n_884),
.B2(n_879),
.C1(n_877),
.C2(n_872),
.Y(n_1044)
);

INVx2_ASAP7_75t_L g1045 ( 
.A(n_1034),
.Y(n_1045)
);

AOI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_1021),
.A2(n_819),
.B(n_822),
.Y(n_1046)
);

NOR2xp67_ASAP7_75t_L g1047 ( 
.A(n_1021),
.B(n_1031),
.Y(n_1047)
);

HB1xp67_ASAP7_75t_L g1048 ( 
.A(n_1030),
.Y(n_1048)
);

NAND2x1p5_ASAP7_75t_L g1049 ( 
.A(n_1028),
.B(n_780),
.Y(n_1049)
);

NOR2xp33_ASAP7_75t_SL g1050 ( 
.A(n_1025),
.B(n_760),
.Y(n_1050)
);

XNOR2x1_ASAP7_75t_L g1051 ( 
.A(n_1024),
.B(n_819),
.Y(n_1051)
);

BUFx2_ASAP7_75t_L g1052 ( 
.A(n_1026),
.Y(n_1052)
);

NOR2xp33_ASAP7_75t_L g1053 ( 
.A(n_1052),
.B(n_760),
.Y(n_1053)
);

NOR2xp33_ASAP7_75t_SL g1054 ( 
.A(n_1041),
.B(n_1038),
.Y(n_1054)
);

INVx3_ASAP7_75t_L g1055 ( 
.A(n_1035),
.Y(n_1055)
);

OR2x2_ASAP7_75t_L g1056 ( 
.A(n_1045),
.B(n_810),
.Y(n_1056)
);

HB1xp67_ASAP7_75t_L g1057 ( 
.A(n_1047),
.Y(n_1057)
);

AND2x4_ASAP7_75t_L g1058 ( 
.A(n_1042),
.B(n_835),
.Y(n_1058)
);

AND2x4_ASAP7_75t_L g1059 ( 
.A(n_1042),
.B(n_835),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_1043),
.B(n_851),
.Y(n_1060)
);

AOI22xp33_ASAP7_75t_L g1061 ( 
.A1(n_1051),
.A2(n_815),
.B1(n_818),
.B2(n_822),
.Y(n_1061)
);

NAND2x1p5_ASAP7_75t_L g1062 ( 
.A(n_1037),
.B(n_1048),
.Y(n_1062)
);

AND2x4_ASAP7_75t_L g1063 ( 
.A(n_1039),
.B(n_835),
.Y(n_1063)
);

OA22x2_ASAP7_75t_L g1064 ( 
.A1(n_1057),
.A2(n_1055),
.B1(n_1060),
.B2(n_1059),
.Y(n_1064)
);

AOI22xp5_ASAP7_75t_L g1065 ( 
.A1(n_1054),
.A2(n_1050),
.B1(n_1040),
.B2(n_1049),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_1062),
.Y(n_1066)
);

OAI22xp5_ASAP7_75t_L g1067 ( 
.A1(n_1053),
.A2(n_1046),
.B1(n_1036),
.B2(n_1044),
.Y(n_1067)
);

OR3x1_ASAP7_75t_L g1068 ( 
.A(n_1058),
.B(n_833),
.C(n_822),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_1056),
.Y(n_1069)
);

AOI22xp5_ASAP7_75t_L g1070 ( 
.A1(n_1065),
.A2(n_1063),
.B1(n_1056),
.B2(n_1061),
.Y(n_1070)
);

AOI221xp5_ASAP7_75t_L g1071 ( 
.A1(n_1069),
.A2(n_815),
.B1(n_818),
.B2(n_838),
.C(n_884),
.Y(n_1071)
);

NOR3xp33_ASAP7_75t_L g1072 ( 
.A(n_1066),
.B(n_810),
.C(n_849),
.Y(n_1072)
);

OA22x2_ASAP7_75t_L g1073 ( 
.A1(n_1067),
.A2(n_835),
.B1(n_886),
.B2(n_855),
.Y(n_1073)
);

AOI21xp5_ASAP7_75t_L g1074 ( 
.A1(n_1073),
.A2(n_1064),
.B(n_1068),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_1074),
.Y(n_1075)
);

AOI21xp5_ASAP7_75t_L g1076 ( 
.A1(n_1074),
.A2(n_1070),
.B(n_1072),
.Y(n_1076)
);

AOI21xp5_ASAP7_75t_L g1077 ( 
.A1(n_1076),
.A2(n_1071),
.B(n_822),
.Y(n_1077)
);

OAI22xp33_ASAP7_75t_L g1078 ( 
.A1(n_1075),
.A2(n_822),
.B1(n_815),
.B2(n_886),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_1077),
.B(n_263),
.Y(n_1079)
);

AOI21xp5_ASAP7_75t_L g1080 ( 
.A1(n_1078),
.A2(n_806),
.B(n_265),
.Y(n_1080)
);

OAI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_1079),
.A2(n_806),
.B(n_877),
.Y(n_1081)
);

OAI221xp5_ASAP7_75t_R g1082 ( 
.A1(n_1081),
.A2(n_1080),
.B1(n_266),
.B2(n_268),
.C(n_264),
.Y(n_1082)
);

AOI211xp5_ASAP7_75t_L g1083 ( 
.A1(n_1082),
.A2(n_806),
.B(n_889),
.C(n_882),
.Y(n_1083)
);


endmodule