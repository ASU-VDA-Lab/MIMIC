module fake_ariane_2485_n_1771 (n_83, n_8, n_56, n_60, n_160, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_158, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_52, n_157, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1771);

input n_83;
input n_8;
input n_56;
input n_60;
input n_160;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_158;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_52;
input n_157;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1771;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_1682;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_754;
wire n_665;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_167;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_238;
wire n_365;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1597;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1594;
wire n_680;
wire n_287;
wire n_1716;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_824;
wire n_428;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1163;
wire n_186;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_1726;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_321;
wire n_221;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_888;
wire n_845;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_534;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1753;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1524;
wire n_1476;
wire n_1733;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_169;
wire n_1201;
wire n_1288;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_166;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_168;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_532;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_164;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1735;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_898;
wire n_857;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1727;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1732;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_174;
wire n_275;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_165;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_92),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_63),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_26),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_150),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_137),
.Y(n_168)
);

BUFx8_ASAP7_75t_SL g169 ( 
.A(n_142),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_74),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_83),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_126),
.Y(n_172)
);

INVx1_ASAP7_75t_SL g173 ( 
.A(n_29),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_4),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_55),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_131),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_52),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_94),
.Y(n_178)
);

INVx1_ASAP7_75t_SL g179 ( 
.A(n_134),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_17),
.Y(n_180)
);

INVx1_ASAP7_75t_SL g181 ( 
.A(n_99),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_23),
.Y(n_182)
);

BUFx2_ASAP7_75t_L g183 ( 
.A(n_89),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_22),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_139),
.Y(n_185)
);

BUFx3_ASAP7_75t_L g186 ( 
.A(n_151),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_102),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_138),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_20),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_60),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_118),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_149),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_0),
.Y(n_193)
);

INVx2_ASAP7_75t_SL g194 ( 
.A(n_123),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_24),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_119),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_66),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_114),
.Y(n_198)
);

INVx1_ASAP7_75t_SL g199 ( 
.A(n_29),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_73),
.Y(n_200)
);

BUFx3_ASAP7_75t_L g201 ( 
.A(n_113),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_82),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_79),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_72),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_127),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_11),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_12),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_70),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_24),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_107),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_23),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_64),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_90),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_37),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_62),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_76),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_154),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_110),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_16),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_61),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_141),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_44),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_21),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_160),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_22),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_6),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_4),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_101),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_9),
.Y(n_229)
);

INVx1_ASAP7_75t_SL g230 ( 
.A(n_77),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_117),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_26),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_147),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_12),
.Y(n_234)
);

CKINVDCx14_ASAP7_75t_R g235 ( 
.A(n_140),
.Y(n_235)
);

BUFx3_ASAP7_75t_L g236 ( 
.A(n_38),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_7),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_161),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_157),
.Y(n_239)
);

INVx2_ASAP7_75t_SL g240 ( 
.A(n_34),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_42),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_20),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_125),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_85),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_15),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_42),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_65),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_84),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_124),
.Y(n_249)
);

BUFx10_ASAP7_75t_L g250 ( 
.A(n_155),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_8),
.Y(n_251)
);

INVx2_ASAP7_75t_SL g252 ( 
.A(n_132),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_38),
.Y(n_253)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_93),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_143),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_81),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_55),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_19),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_3),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_43),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_153),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_17),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_69),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_51),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_98),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_16),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_14),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_87),
.Y(n_268)
);

INVx1_ASAP7_75t_SL g269 ( 
.A(n_75),
.Y(n_269)
);

INVx1_ASAP7_75t_SL g270 ( 
.A(n_46),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_39),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_3),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_33),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_162),
.Y(n_274)
);

INVx2_ASAP7_75t_SL g275 ( 
.A(n_34),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_21),
.Y(n_276)
);

BUFx3_ASAP7_75t_L g277 ( 
.A(n_33),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_13),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_32),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_43),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_67),
.Y(n_281)
);

BUFx2_ASAP7_75t_L g282 ( 
.A(n_58),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_128),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_158),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_146),
.Y(n_285)
);

INVx1_ASAP7_75t_SL g286 ( 
.A(n_31),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_6),
.Y(n_287)
);

INVx1_ASAP7_75t_SL g288 ( 
.A(n_145),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_28),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_116),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_68),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_96),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_51),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_144),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_122),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_37),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_133),
.Y(n_297)
);

INVx2_ASAP7_75t_SL g298 ( 
.A(n_15),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_100),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_159),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_53),
.Y(n_301)
);

BUFx8_ASAP7_75t_SL g302 ( 
.A(n_35),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_35),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_58),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_71),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_48),
.Y(n_306)
);

INVxp67_ASAP7_75t_L g307 ( 
.A(n_50),
.Y(n_307)
);

BUFx2_ASAP7_75t_L g308 ( 
.A(n_163),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_2),
.Y(n_309)
);

BUFx3_ASAP7_75t_L g310 ( 
.A(n_57),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_28),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_13),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_106),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_56),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_120),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_111),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_0),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_8),
.Y(n_318)
);

BUFx5_ASAP7_75t_L g319 ( 
.A(n_156),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_129),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_9),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_54),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_50),
.Y(n_323)
);

INVx1_ASAP7_75t_SL g324 ( 
.A(n_130),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_2),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_115),
.Y(n_326)
);

BUFx2_ASAP7_75t_L g327 ( 
.A(n_148),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_49),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_302),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_183),
.B(n_1),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_169),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_180),
.Y(n_332)
);

NOR2xp67_ASAP7_75t_L g333 ( 
.A(n_240),
.B(n_1),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_176),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_180),
.Y(n_335)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_282),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_180),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_185),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_192),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_180),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_308),
.B(n_5),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_217),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_268),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_180),
.Y(n_344)
);

HB1xp67_ASAP7_75t_L g345 ( 
.A(n_177),
.Y(n_345)
);

INVxp67_ASAP7_75t_SL g346 ( 
.A(n_236),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_225),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_225),
.Y(n_348)
);

BUFx2_ASAP7_75t_L g349 ( 
.A(n_236),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_326),
.Y(n_350)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_225),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_225),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_225),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_207),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_242),
.Y(n_355)
);

CKINVDCx16_ASAP7_75t_R g356 ( 
.A(n_164),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_174),
.Y(n_357)
);

INVxp33_ASAP7_75t_SL g358 ( 
.A(n_177),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_242),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_175),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_R g361 ( 
.A(n_235),
.B(n_152),
.Y(n_361)
);

NOR2xp67_ASAP7_75t_L g362 ( 
.A(n_240),
.B(n_5),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_189),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_209),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_242),
.Y(n_365)
);

HB1xp67_ASAP7_75t_L g366 ( 
.A(n_182),
.Y(n_366)
);

HB1xp67_ASAP7_75t_L g367 ( 
.A(n_182),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_245),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_242),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_258),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_271),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_242),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_211),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_214),
.Y(n_374)
);

HB1xp67_ASAP7_75t_L g375 ( 
.A(n_184),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_262),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_219),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_262),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_223),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_312),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_227),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_232),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_234),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_273),
.Y(n_384)
);

HB1xp67_ASAP7_75t_L g385 ( 
.A(n_184),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_237),
.Y(n_386)
);

XNOR2x1_ASAP7_75t_L g387 ( 
.A(n_193),
.B(n_195),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_241),
.Y(n_388)
);

BUFx6f_ASAP7_75t_L g389 ( 
.A(n_238),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_253),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_273),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_254),
.Y(n_392)
);

HB1xp67_ASAP7_75t_L g393 ( 
.A(n_193),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_254),
.Y(n_394)
);

CKINVDCx16_ASAP7_75t_R g395 ( 
.A(n_250),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_325),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_290),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_290),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_260),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_186),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_250),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_166),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_206),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_264),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_250),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_222),
.Y(n_406)
);

BUFx2_ASAP7_75t_L g407 ( 
.A(n_277),
.Y(n_407)
);

BUFx6f_ASAP7_75t_SL g408 ( 
.A(n_186),
.Y(n_408)
);

INVx1_ASAP7_75t_SL g409 ( 
.A(n_173),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_328),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_389),
.Y(n_411)
);

BUFx6f_ASAP7_75t_L g412 ( 
.A(n_389),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_332),
.Y(n_413)
);

HB1xp67_ASAP7_75t_L g414 ( 
.A(n_387),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_389),
.Y(n_415)
);

INVx3_ASAP7_75t_L g416 ( 
.A(n_351),
.Y(n_416)
);

BUFx3_ASAP7_75t_L g417 ( 
.A(n_400),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_338),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_332),
.Y(n_419)
);

BUFx6f_ASAP7_75t_L g420 ( 
.A(n_389),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_342),
.Y(n_421)
);

AND2x6_ASAP7_75t_L g422 ( 
.A(n_389),
.B(n_238),
.Y(n_422)
);

AND2x2_ASAP7_75t_L g423 ( 
.A(n_349),
.B(n_277),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_389),
.Y(n_424)
);

INVxp33_ASAP7_75t_L g425 ( 
.A(n_387),
.Y(n_425)
);

INVxp33_ASAP7_75t_SL g426 ( 
.A(n_331),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_335),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_335),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_337),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_350),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_337),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_340),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_340),
.Y(n_433)
);

BUFx3_ASAP7_75t_L g434 ( 
.A(n_400),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_339),
.Y(n_435)
);

INVx3_ASAP7_75t_L g436 ( 
.A(n_351),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_344),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_343),
.Y(n_438)
);

AND2x4_ASAP7_75t_L g439 ( 
.A(n_346),
.B(n_310),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_329),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_344),
.Y(n_441)
);

NAND2xp33_ASAP7_75t_L g442 ( 
.A(n_354),
.B(n_275),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_347),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_347),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_348),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_348),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_364),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_373),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_352),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_352),
.Y(n_450)
);

AND2x2_ASAP7_75t_L g451 ( 
.A(n_349),
.B(n_310),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_353),
.Y(n_452)
);

AND2x2_ASAP7_75t_L g453 ( 
.A(n_407),
.B(n_402),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_353),
.Y(n_454)
);

BUFx6f_ASAP7_75t_L g455 ( 
.A(n_355),
.Y(n_455)
);

NOR2xp67_ASAP7_75t_L g456 ( 
.A(n_392),
.B(n_194),
.Y(n_456)
);

INVxp67_ASAP7_75t_L g457 ( 
.A(n_409),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_392),
.B(n_327),
.Y(n_458)
);

AND2x4_ASAP7_75t_L g459 ( 
.A(n_394),
.B(n_275),
.Y(n_459)
);

OA21x2_ASAP7_75t_L g460 ( 
.A1(n_355),
.A2(n_168),
.B(n_165),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_374),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_377),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_379),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_359),
.Y(n_464)
);

CKINVDCx20_ASAP7_75t_R g465 ( 
.A(n_357),
.Y(n_465)
);

INVxp67_ASAP7_75t_L g466 ( 
.A(n_345),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_359),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_330),
.B(n_194),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_381),
.Y(n_469)
);

CKINVDCx16_ASAP7_75t_R g470 ( 
.A(n_395),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_382),
.Y(n_471)
);

CKINVDCx20_ASAP7_75t_R g472 ( 
.A(n_360),
.Y(n_472)
);

OAI21x1_ASAP7_75t_L g473 ( 
.A1(n_394),
.A2(n_398),
.B(n_397),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_365),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_397),
.B(n_178),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_398),
.B(n_190),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_383),
.Y(n_477)
);

INVxp67_ASAP7_75t_L g478 ( 
.A(n_366),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_365),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_369),
.Y(n_480)
);

OR2x2_ASAP7_75t_L g481 ( 
.A(n_407),
.B(n_199),
.Y(n_481)
);

INVx1_ASAP7_75t_SL g482 ( 
.A(n_401),
.Y(n_482)
);

HB1xp67_ASAP7_75t_L g483 ( 
.A(n_336),
.Y(n_483)
);

INVxp67_ASAP7_75t_L g484 ( 
.A(n_457),
.Y(n_484)
);

AND2x6_ASAP7_75t_L g485 ( 
.A(n_468),
.B(n_201),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_468),
.B(n_395),
.Y(n_486)
);

OR2x6_ASAP7_75t_L g487 ( 
.A(n_439),
.B(n_341),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_446),
.Y(n_488)
);

INVx3_ASAP7_75t_L g489 ( 
.A(n_473),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_SL g490 ( 
.A(n_447),
.B(n_356),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_466),
.B(n_356),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_417),
.B(n_386),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_417),
.B(n_388),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_SL g494 ( 
.A(n_448),
.B(n_390),
.Y(n_494)
);

AND2x2_ASAP7_75t_L g495 ( 
.A(n_453),
.B(n_402),
.Y(n_495)
);

AOI22xp33_ASAP7_75t_L g496 ( 
.A1(n_439),
.A2(n_459),
.B1(n_434),
.B2(n_417),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_SL g497 ( 
.A(n_461),
.B(n_399),
.Y(n_497)
);

BUFx2_ASAP7_75t_L g498 ( 
.A(n_457),
.Y(n_498)
);

INVx2_ASAP7_75t_SL g499 ( 
.A(n_481),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_434),
.B(n_404),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_434),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_473),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_473),
.Y(n_503)
);

OAI21xp33_ASAP7_75t_SL g504 ( 
.A1(n_453),
.A2(n_362),
.B(n_333),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_446),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_413),
.Y(n_506)
);

INVx4_ASAP7_75t_L g507 ( 
.A(n_422),
.Y(n_507)
);

OR2x2_ASAP7_75t_L g508 ( 
.A(n_481),
.B(n_367),
.Y(n_508)
);

INVx2_ASAP7_75t_SL g509 ( 
.A(n_453),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_413),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_450),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_SL g512 ( 
.A(n_462),
.B(n_410),
.Y(n_512)
);

BUFx2_ASAP7_75t_L g513 ( 
.A(n_463),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_SL g514 ( 
.A(n_426),
.B(n_405),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_439),
.B(n_358),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_450),
.Y(n_516)
);

INVx2_ASAP7_75t_SL g517 ( 
.A(n_423),
.Y(n_517)
);

OR2x6_ASAP7_75t_L g518 ( 
.A(n_439),
.B(n_333),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_419),
.Y(n_519)
);

AND2x2_ASAP7_75t_L g520 ( 
.A(n_439),
.B(n_403),
.Y(n_520)
);

AND2x6_ASAP7_75t_L g521 ( 
.A(n_459),
.B(n_201),
.Y(n_521)
);

CKINVDCx20_ASAP7_75t_R g522 ( 
.A(n_465),
.Y(n_522)
);

INVx1_ASAP7_75t_SL g523 ( 
.A(n_472),
.Y(n_523)
);

BUFx6f_ASAP7_75t_L g524 ( 
.A(n_455),
.Y(n_524)
);

AND2x6_ASAP7_75t_L g525 ( 
.A(n_459),
.B(n_238),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_452),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_452),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_419),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_427),
.Y(n_529)
);

INVx1_ASAP7_75t_SL g530 ( 
.A(n_482),
.Y(n_530)
);

AND2x2_ASAP7_75t_L g531 ( 
.A(n_483),
.B(n_375),
.Y(n_531)
);

AND2x6_ASAP7_75t_L g532 ( 
.A(n_459),
.B(n_238),
.Y(n_532)
);

BUFx3_ASAP7_75t_L g533 ( 
.A(n_469),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_SL g534 ( 
.A(n_470),
.B(n_385),
.Y(n_534)
);

BUFx6f_ASAP7_75t_L g535 ( 
.A(n_455),
.Y(n_535)
);

OR2x2_ASAP7_75t_L g536 ( 
.A(n_483),
.B(n_393),
.Y(n_536)
);

BUFx3_ASAP7_75t_L g537 ( 
.A(n_471),
.Y(n_537)
);

INVx1_ASAP7_75t_SL g538 ( 
.A(n_482),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_452),
.Y(n_539)
);

CKINVDCx20_ASAP7_75t_R g540 ( 
.A(n_470),
.Y(n_540)
);

CKINVDCx20_ASAP7_75t_R g541 ( 
.A(n_414),
.Y(n_541)
);

OAI22xp5_ASAP7_75t_L g542 ( 
.A1(n_466),
.A2(n_362),
.B1(n_307),
.B2(n_321),
.Y(n_542)
);

BUFx4f_ASAP7_75t_L g543 ( 
.A(n_460),
.Y(n_543)
);

OR2x6_ASAP7_75t_L g544 ( 
.A(n_459),
.B(n_298),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_464),
.Y(n_545)
);

BUFx10_ASAP7_75t_L g546 ( 
.A(n_477),
.Y(n_546)
);

NAND2xp33_ASAP7_75t_L g547 ( 
.A(n_422),
.B(n_319),
.Y(n_547)
);

BUFx2_ASAP7_75t_L g548 ( 
.A(n_418),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_427),
.Y(n_549)
);

AOI22xp33_ASAP7_75t_L g550 ( 
.A1(n_460),
.A2(n_361),
.B1(n_298),
.B2(n_408),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_464),
.Y(n_551)
);

NAND2xp33_ASAP7_75t_L g552 ( 
.A(n_422),
.B(n_319),
.Y(n_552)
);

NAND2x1p5_ASAP7_75t_L g553 ( 
.A(n_423),
.B(n_403),
.Y(n_553)
);

INVx3_ASAP7_75t_L g554 ( 
.A(n_455),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_SL g555 ( 
.A(n_478),
.B(n_196),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_SL g556 ( 
.A(n_478),
.B(n_198),
.Y(n_556)
);

BUFx4f_ASAP7_75t_L g557 ( 
.A(n_460),
.Y(n_557)
);

INVx3_ASAP7_75t_L g558 ( 
.A(n_455),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_428),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_442),
.B(n_408),
.Y(n_560)
);

NAND2xp33_ASAP7_75t_L g561 ( 
.A(n_422),
.B(n_319),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_428),
.Y(n_562)
);

AOI22xp33_ASAP7_75t_L g563 ( 
.A1(n_460),
.A2(n_408),
.B1(n_280),
.B2(n_266),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_429),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_458),
.B(n_406),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_429),
.Y(n_566)
);

NAND3xp33_ASAP7_75t_L g567 ( 
.A(n_423),
.B(n_246),
.C(n_195),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_SL g568 ( 
.A(n_458),
.B(n_202),
.Y(n_568)
);

INVx5_ASAP7_75t_L g569 ( 
.A(n_422),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_451),
.B(n_406),
.Y(n_570)
);

AOI22xp33_ASAP7_75t_L g571 ( 
.A1(n_460),
.A2(n_451),
.B1(n_425),
.B2(n_414),
.Y(n_571)
);

BUFx10_ASAP7_75t_L g572 ( 
.A(n_421),
.Y(n_572)
);

BUFx4f_ASAP7_75t_L g573 ( 
.A(n_455),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_464),
.Y(n_574)
);

AND2x6_ASAP7_75t_L g575 ( 
.A(n_451),
.B(n_238),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_431),
.Y(n_576)
);

INVx3_ASAP7_75t_L g577 ( 
.A(n_455),
.Y(n_577)
);

CKINVDCx16_ASAP7_75t_R g578 ( 
.A(n_430),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_SL g579 ( 
.A(n_475),
.B(n_204),
.Y(n_579)
);

BUFx6f_ASAP7_75t_L g580 ( 
.A(n_455),
.Y(n_580)
);

AOI22xp33_ASAP7_75t_L g581 ( 
.A1(n_456),
.A2(n_475),
.B1(n_476),
.B2(n_257),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_SL g582 ( 
.A(n_476),
.B(n_210),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_431),
.B(n_369),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_467),
.Y(n_584)
);

NAND2xp33_ASAP7_75t_L g585 ( 
.A(n_422),
.B(n_319),
.Y(n_585)
);

INVx1_ASAP7_75t_SL g586 ( 
.A(n_435),
.Y(n_586)
);

BUFx3_ASAP7_75t_L g587 ( 
.A(n_432),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_432),
.Y(n_588)
);

INVx3_ASAP7_75t_L g589 ( 
.A(n_467),
.Y(n_589)
);

CKINVDCx20_ASAP7_75t_R g590 ( 
.A(n_438),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_L g591 ( 
.A(n_433),
.B(n_215),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_467),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_SL g593 ( 
.A(n_433),
.B(n_221),
.Y(n_593)
);

BUFx10_ASAP7_75t_L g594 ( 
.A(n_440),
.Y(n_594)
);

INVx3_ASAP7_75t_L g595 ( 
.A(n_416),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_437),
.Y(n_596)
);

INVx6_ASAP7_75t_L g597 ( 
.A(n_412),
.Y(n_597)
);

AND2x2_ASAP7_75t_L g598 ( 
.A(n_437),
.B(n_376),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_441),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_441),
.Y(n_600)
);

OR2x2_ASAP7_75t_L g601 ( 
.A(n_416),
.B(n_270),
.Y(n_601)
);

BUFx2_ASAP7_75t_L g602 ( 
.A(n_443),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_443),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_444),
.Y(n_604)
);

INVx4_ASAP7_75t_L g605 ( 
.A(n_422),
.Y(n_605)
);

AND2x2_ASAP7_75t_L g606 ( 
.A(n_444),
.B(n_376),
.Y(n_606)
);

AND2x2_ASAP7_75t_L g607 ( 
.A(n_445),
.B(n_378),
.Y(n_607)
);

NAND3xp33_ASAP7_75t_L g608 ( 
.A(n_445),
.B(n_276),
.C(n_246),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_449),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_454),
.Y(n_610)
);

AND2x2_ASAP7_75t_L g611 ( 
.A(n_474),
.B(n_378),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_474),
.Y(n_612)
);

OAI22xp5_ASAP7_75t_L g613 ( 
.A1(n_479),
.A2(n_309),
.B1(n_287),
.B2(n_323),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_SL g614 ( 
.A(n_479),
.B(n_228),
.Y(n_614)
);

INVx2_ASAP7_75t_SL g615 ( 
.A(n_416),
.Y(n_615)
);

BUFx6f_ASAP7_75t_L g616 ( 
.A(n_412),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_480),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_480),
.Y(n_618)
);

AOI22xp33_ASAP7_75t_L g619 ( 
.A1(n_416),
.A2(n_317),
.B1(n_272),
.B2(n_293),
.Y(n_619)
);

OR2x6_ASAP7_75t_L g620 ( 
.A(n_436),
.B(n_384),
.Y(n_620)
);

OR2x6_ASAP7_75t_L g621 ( 
.A(n_436),
.B(n_384),
.Y(n_621)
);

AND2x2_ASAP7_75t_L g622 ( 
.A(n_436),
.B(n_391),
.Y(n_622)
);

INVx6_ASAP7_75t_L g623 ( 
.A(n_412),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_SL g624 ( 
.A(n_412),
.B(n_247),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_436),
.Y(n_625)
);

INVx2_ASAP7_75t_SL g626 ( 
.A(n_411),
.Y(n_626)
);

AND2x2_ASAP7_75t_L g627 ( 
.A(n_411),
.B(n_391),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_411),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_424),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_565),
.B(n_179),
.Y(n_630)
);

A2O1A1Ixp33_ASAP7_75t_L g631 ( 
.A1(n_504),
.A2(n_226),
.B(n_229),
.C(n_267),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_587),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_486),
.B(n_181),
.Y(n_633)
);

AOI22xp5_ASAP7_75t_L g634 ( 
.A1(n_487),
.A2(n_252),
.B1(n_291),
.B2(n_292),
.Y(n_634)
);

INVxp67_ASAP7_75t_L g635 ( 
.A(n_498),
.Y(n_635)
);

INVx8_ASAP7_75t_L g636 ( 
.A(n_521),
.Y(n_636)
);

AOI22xp5_ASAP7_75t_L g637 ( 
.A1(n_487),
.A2(n_485),
.B1(n_618),
.B2(n_515),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_520),
.B(n_230),
.Y(n_638)
);

BUFx3_ASAP7_75t_L g639 ( 
.A(n_590),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_587),
.Y(n_640)
);

INVx4_ASAP7_75t_L g641 ( 
.A(n_620),
.Y(n_641)
);

O2A1O1Ixp5_ASAP7_75t_L g642 ( 
.A1(n_489),
.A2(n_249),
.B(n_256),
.C(n_263),
.Y(n_642)
);

NOR2xp33_ASAP7_75t_L g643 ( 
.A(n_517),
.B(n_286),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_SL g644 ( 
.A(n_491),
.B(n_533),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_595),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_622),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_520),
.B(n_269),
.Y(n_647)
);

NOR2xp33_ASAP7_75t_L g648 ( 
.A(n_517),
.B(n_276),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_618),
.B(n_288),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_496),
.B(n_571),
.Y(n_650)
);

AOI22xp5_ASAP7_75t_L g651 ( 
.A1(n_487),
.A2(n_252),
.B1(n_285),
.B2(n_284),
.Y(n_651)
);

O2A1O1Ixp33_ASAP7_75t_L g652 ( 
.A1(n_570),
.A2(n_251),
.B(n_259),
.C(n_311),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_595),
.Y(n_653)
);

AOI22xp33_ASAP7_75t_L g654 ( 
.A1(n_509),
.A2(n_485),
.B1(n_521),
.B2(n_543),
.Y(n_654)
);

INVx2_ASAP7_75t_SL g655 ( 
.A(n_530),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_595),
.Y(n_656)
);

AOI22xp5_ASAP7_75t_L g657 ( 
.A1(n_487),
.A2(n_203),
.B1(n_200),
.B2(n_197),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_589),
.Y(n_658)
);

NOR2xp33_ASAP7_75t_L g659 ( 
.A(n_492),
.B(n_278),
.Y(n_659)
);

AND2x2_ASAP7_75t_L g660 ( 
.A(n_499),
.B(n_363),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_568),
.B(n_324),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_SL g662 ( 
.A(n_489),
.B(n_167),
.Y(n_662)
);

INVx2_ASAP7_75t_SL g663 ( 
.A(n_538),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_SL g664 ( 
.A(n_533),
.B(n_167),
.Y(n_664)
);

INVx8_ASAP7_75t_L g665 ( 
.A(n_521),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_568),
.B(n_170),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_L g667 ( 
.A(n_493),
.B(n_278),
.Y(n_667)
);

BUFx6f_ASAP7_75t_SL g668 ( 
.A(n_594),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_553),
.B(n_170),
.Y(n_669)
);

OAI221xp5_ASAP7_75t_L g670 ( 
.A1(n_509),
.A2(n_289),
.B1(n_314),
.B2(n_323),
.C(n_322),
.Y(n_670)
);

NOR2xp33_ASAP7_75t_L g671 ( 
.A(n_500),
.B(n_279),
.Y(n_671)
);

BUFx3_ASAP7_75t_L g672 ( 
.A(n_590),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_SL g673 ( 
.A(n_537),
.B(n_171),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_SL g674 ( 
.A(n_537),
.B(n_171),
.Y(n_674)
);

INVxp67_ASAP7_75t_L g675 ( 
.A(n_499),
.Y(n_675)
);

AND2x2_ASAP7_75t_L g676 ( 
.A(n_484),
.B(n_368),
.Y(n_676)
);

AOI22xp5_ASAP7_75t_L g677 ( 
.A1(n_485),
.A2(n_285),
.B1(n_203),
.B2(n_200),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_553),
.B(n_172),
.Y(n_678)
);

AOI22xp5_ASAP7_75t_L g679 ( 
.A1(n_485),
.A2(n_291),
.B1(n_197),
.B2(n_191),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_598),
.Y(n_680)
);

BUFx6f_ASAP7_75t_L g681 ( 
.A(n_507),
.Y(n_681)
);

OR2x2_ASAP7_75t_L g682 ( 
.A(n_508),
.B(n_370),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_602),
.B(n_172),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_581),
.B(n_187),
.Y(n_684)
);

OR2x6_ASAP7_75t_L g685 ( 
.A(n_548),
.B(n_371),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_589),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_495),
.B(n_187),
.Y(n_687)
);

OAI22xp5_ASAP7_75t_SL g688 ( 
.A1(n_541),
.A2(n_380),
.B1(n_396),
.B2(n_287),
.Y(n_688)
);

AOI22xp33_ASAP7_75t_L g689 ( 
.A1(n_485),
.A2(n_303),
.B1(n_301),
.B2(n_304),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_495),
.B(n_560),
.Y(n_690)
);

AOI22xp5_ASAP7_75t_L g691 ( 
.A1(n_485),
.A2(n_284),
.B1(n_191),
.B2(n_188),
.Y(n_691)
);

NOR2xp33_ASAP7_75t_L g692 ( 
.A(n_567),
.B(n_279),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_579),
.B(n_292),
.Y(n_693)
);

INVx2_ASAP7_75t_SL g694 ( 
.A(n_601),
.Y(n_694)
);

OAI21xp5_ASAP7_75t_L g695 ( 
.A1(n_543),
.A2(n_557),
.B(n_503),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_579),
.B(n_294),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_SL g697 ( 
.A(n_546),
.B(n_294),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_582),
.B(n_295),
.Y(n_698)
);

AND2x2_ASAP7_75t_L g699 ( 
.A(n_531),
.B(n_296),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_589),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_488),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_488),
.Y(n_702)
);

NOR2xp33_ASAP7_75t_L g703 ( 
.A(n_518),
.B(n_296),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_598),
.Y(n_704)
);

INVx2_ASAP7_75t_SL g705 ( 
.A(n_523),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_505),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_582),
.B(n_295),
.Y(n_707)
);

NOR2xp33_ASAP7_75t_L g708 ( 
.A(n_518),
.B(n_301),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_518),
.B(n_297),
.Y(n_709)
);

BUFx8_ASAP7_75t_L g710 ( 
.A(n_513),
.Y(n_710)
);

INVx2_ASAP7_75t_SL g711 ( 
.A(n_536),
.Y(n_711)
);

INVx4_ASAP7_75t_L g712 ( 
.A(n_620),
.Y(n_712)
);

AOI22xp5_ASAP7_75t_L g713 ( 
.A1(n_518),
.A2(n_297),
.B1(n_320),
.B2(n_305),
.Y(n_713)
);

INVx2_ASAP7_75t_SL g714 ( 
.A(n_546),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_521),
.B(n_299),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_521),
.B(n_299),
.Y(n_716)
);

NAND3xp33_ASAP7_75t_L g717 ( 
.A(n_494),
.B(n_318),
.C(n_306),
.Y(n_717)
);

BUFx5_ASAP7_75t_L g718 ( 
.A(n_502),
.Y(n_718)
);

NOR2xp67_ASAP7_75t_L g719 ( 
.A(n_494),
.B(n_372),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_521),
.B(n_575),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_SL g721 ( 
.A(n_489),
.B(n_300),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_SL g722 ( 
.A(n_543),
.B(n_557),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_575),
.B(n_300),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_SL g724 ( 
.A(n_546),
.B(n_305),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_575),
.B(n_320),
.Y(n_725)
);

AND2x2_ASAP7_75t_L g726 ( 
.A(n_572),
.B(n_303),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_575),
.B(n_304),
.Y(n_727)
);

INVxp67_ASAP7_75t_SL g728 ( 
.A(n_557),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_606),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_606),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_575),
.B(n_306),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_SL g732 ( 
.A(n_497),
.B(n_309),
.Y(n_732)
);

OAI22xp33_ASAP7_75t_L g733 ( 
.A1(n_544),
.A2(n_318),
.B1(n_322),
.B2(n_281),
.Y(n_733)
);

INVxp67_ASAP7_75t_L g734 ( 
.A(n_534),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_575),
.B(n_205),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_SL g736 ( 
.A(n_524),
.B(n_274),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_SL g737 ( 
.A(n_497),
.B(n_208),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_607),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_SL g739 ( 
.A(n_512),
.B(n_212),
.Y(n_739)
);

INVx2_ASAP7_75t_SL g740 ( 
.A(n_572),
.Y(n_740)
);

NOR2xp33_ASAP7_75t_L g741 ( 
.A(n_555),
.B(n_283),
.Y(n_741)
);

AOI22xp5_ASAP7_75t_L g742 ( 
.A1(n_544),
.A2(n_556),
.B1(n_555),
.B2(n_620),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_544),
.B(n_607),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_544),
.B(n_213),
.Y(n_744)
);

INVxp67_ASAP7_75t_L g745 ( 
.A(n_586),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_611),
.B(n_216),
.Y(n_746)
);

OR2x2_ASAP7_75t_L g747 ( 
.A(n_578),
.B(n_7),
.Y(n_747)
);

AND2x2_ASAP7_75t_L g748 ( 
.A(n_572),
.B(n_10),
.Y(n_748)
);

NOR2xp33_ASAP7_75t_L g749 ( 
.A(n_556),
.B(n_313),
.Y(n_749)
);

AOI22xp5_ASAP7_75t_SL g750 ( 
.A1(n_541),
.A2(n_316),
.B1(n_315),
.B2(n_224),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_611),
.B(n_501),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_SL g752 ( 
.A(n_512),
.B(n_248),
.Y(n_752)
);

OR2x6_ASAP7_75t_L g753 ( 
.A(n_490),
.B(n_424),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_506),
.B(n_244),
.Y(n_754)
);

NOR2xp33_ASAP7_75t_L g755 ( 
.A(n_608),
.B(n_10),
.Y(n_755)
);

O2A1O1Ixp5_ASAP7_75t_L g756 ( 
.A1(n_593),
.A2(n_424),
.B(n_415),
.C(n_422),
.Y(n_756)
);

OAI22xp33_ASAP7_75t_L g757 ( 
.A1(n_514),
.A2(n_218),
.B1(n_220),
.B2(n_231),
.Y(n_757)
);

NOR3xp33_ASAP7_75t_L g758 ( 
.A(n_490),
.B(n_233),
.C(n_239),
.Y(n_758)
);

OAI22xp5_ASAP7_75t_SL g759 ( 
.A1(n_522),
.A2(n_243),
.B1(n_255),
.B2(n_261),
.Y(n_759)
);

INVx2_ASAP7_75t_SL g760 ( 
.A(n_594),
.Y(n_760)
);

NOR3xp33_ASAP7_75t_L g761 ( 
.A(n_542),
.B(n_265),
.C(n_415),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_SL g762 ( 
.A(n_550),
.B(n_319),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_511),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_510),
.B(n_415),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_SL g765 ( 
.A(n_613),
.B(n_319),
.Y(n_765)
);

OR2x2_ASAP7_75t_L g766 ( 
.A(n_619),
.B(n_11),
.Y(n_766)
);

NOR2xp33_ASAP7_75t_L g767 ( 
.A(n_519),
.B(n_14),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_SL g768 ( 
.A(n_615),
.B(n_319),
.Y(n_768)
);

AOI22xp5_ASAP7_75t_L g769 ( 
.A1(n_620),
.A2(n_319),
.B1(n_422),
.B2(n_412),
.Y(n_769)
);

AOI22xp33_ASAP7_75t_L g770 ( 
.A1(n_563),
.A2(n_420),
.B1(n_412),
.B2(n_25),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_528),
.B(n_529),
.Y(n_771)
);

AND2x2_ASAP7_75t_L g772 ( 
.A(n_594),
.B(n_540),
.Y(n_772)
);

AND2x6_ASAP7_75t_SL g773 ( 
.A(n_522),
.B(n_18),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_549),
.B(n_18),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_559),
.B(n_19),
.Y(n_775)
);

NOR2xp33_ASAP7_75t_L g776 ( 
.A(n_562),
.B(n_25),
.Y(n_776)
);

NOR2xp67_ASAP7_75t_L g777 ( 
.A(n_615),
.B(n_564),
.Y(n_777)
);

AND2x2_ASAP7_75t_L g778 ( 
.A(n_540),
.B(n_27),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_516),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_566),
.B(n_27),
.Y(n_780)
);

NOR2xp33_ASAP7_75t_L g781 ( 
.A(n_576),
.B(n_30),
.Y(n_781)
);

OAI22xp5_ASAP7_75t_L g782 ( 
.A1(n_588),
.A2(n_30),
.B1(n_31),
.B2(n_32),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_596),
.B(n_36),
.Y(n_783)
);

NOR2xp33_ASAP7_75t_R g784 ( 
.A(n_547),
.B(n_86),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_SL g785 ( 
.A(n_524),
.B(n_420),
.Y(n_785)
);

BUFx6f_ASAP7_75t_L g786 ( 
.A(n_507),
.Y(n_786)
);

INVx8_ASAP7_75t_L g787 ( 
.A(n_525),
.Y(n_787)
);

INVxp67_ASAP7_75t_L g788 ( 
.A(n_621),
.Y(n_788)
);

INVx3_ASAP7_75t_L g789 ( 
.A(n_621),
.Y(n_789)
);

INVx4_ASAP7_75t_L g790 ( 
.A(n_621),
.Y(n_790)
);

OAI22xp5_ASAP7_75t_L g791 ( 
.A1(n_599),
.A2(n_36),
.B1(n_39),
.B2(n_40),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_600),
.B(n_40),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_627),
.Y(n_793)
);

AOI21xp5_ASAP7_75t_L g794 ( 
.A1(n_695),
.A2(n_573),
.B(n_577),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_771),
.Y(n_795)
);

AOI21x1_ASAP7_75t_L g796 ( 
.A1(n_785),
.A2(n_617),
.B(n_604),
.Y(n_796)
);

AOI21xp5_ASAP7_75t_L g797 ( 
.A1(n_722),
.A2(n_573),
.B(n_577),
.Y(n_797)
);

AOI21xp5_ASAP7_75t_L g798 ( 
.A1(n_722),
.A2(n_573),
.B(n_577),
.Y(n_798)
);

OR2x4_ASAP7_75t_L g799 ( 
.A(n_747),
.B(n_591),
.Y(n_799)
);

O2A1O1Ixp33_ASAP7_75t_L g800 ( 
.A1(n_733),
.A2(n_625),
.B(n_614),
.C(n_593),
.Y(n_800)
);

AOI21xp5_ASAP7_75t_L g801 ( 
.A1(n_728),
.A2(n_554),
.B(n_558),
.Y(n_801)
);

AOI21xp5_ASAP7_75t_L g802 ( 
.A1(n_728),
.A2(n_554),
.B(n_558),
.Y(n_802)
);

AOI21xp5_ASAP7_75t_L g803 ( 
.A1(n_764),
.A2(n_554),
.B(n_558),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_751),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_633),
.B(n_627),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_650),
.B(n_603),
.Y(n_806)
);

A2O1A1Ixp33_ASAP7_75t_L g807 ( 
.A1(n_741),
.A2(n_609),
.B(n_610),
.C(n_612),
.Y(n_807)
);

AOI21xp5_ASAP7_75t_L g808 ( 
.A1(n_785),
.A2(n_610),
.B(n_612),
.Y(n_808)
);

NOR2xp67_ASAP7_75t_L g809 ( 
.A(n_745),
.B(n_614),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_646),
.B(n_527),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_701),
.Y(n_811)
);

OR2x6_ASAP7_75t_L g812 ( 
.A(n_685),
.B(n_621),
.Y(n_812)
);

CKINVDCx8_ASAP7_75t_R g813 ( 
.A(n_685),
.Y(n_813)
);

AOI21xp5_ASAP7_75t_L g814 ( 
.A1(n_662),
.A2(n_626),
.B(n_628),
.Y(n_814)
);

BUFx6f_ASAP7_75t_L g815 ( 
.A(n_787),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_659),
.B(n_532),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_702),
.Y(n_817)
);

OR2x2_ASAP7_75t_L g818 ( 
.A(n_682),
.B(n_574),
.Y(n_818)
);

OAI21x1_ASAP7_75t_L g819 ( 
.A1(n_756),
.A2(n_551),
.B(n_539),
.Y(n_819)
);

CKINVDCx5p33_ASAP7_75t_R g820 ( 
.A(n_710),
.Y(n_820)
);

NOR2xp33_ASAP7_75t_L g821 ( 
.A(n_635),
.B(n_626),
.Y(n_821)
);

A2O1A1Ixp33_ASAP7_75t_L g822 ( 
.A1(n_741),
.A2(n_592),
.B(n_551),
.C(n_516),
.Y(n_822)
);

INVxp67_ASAP7_75t_SL g823 ( 
.A(n_681),
.Y(n_823)
);

AOI21xp5_ASAP7_75t_L g824 ( 
.A1(n_662),
.A2(n_629),
.B(n_524),
.Y(n_824)
);

AND2x2_ASAP7_75t_L g825 ( 
.A(n_699),
.B(n_545),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_SL g826 ( 
.A(n_641),
.B(n_580),
.Y(n_826)
);

A2O1A1Ixp33_ASAP7_75t_L g827 ( 
.A1(n_749),
.A2(n_545),
.B(n_584),
.C(n_526),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_659),
.B(n_532),
.Y(n_828)
);

OAI22xp5_ASAP7_75t_L g829 ( 
.A1(n_689),
.A2(n_637),
.B1(n_704),
.B2(n_680),
.Y(n_829)
);

AND2x4_ASAP7_75t_L g830 ( 
.A(n_641),
.B(n_507),
.Y(n_830)
);

AOI21xp5_ASAP7_75t_L g831 ( 
.A1(n_721),
.A2(n_629),
.B(n_535),
.Y(n_831)
);

NOR2x1_ASAP7_75t_L g832 ( 
.A(n_644),
.B(n_717),
.Y(n_832)
);

BUFx6f_ASAP7_75t_L g833 ( 
.A(n_787),
.Y(n_833)
);

NOR2x1_ASAP7_75t_L g834 ( 
.A(n_753),
.B(n_605),
.Y(n_834)
);

OAI321xp33_ASAP7_75t_L g835 ( 
.A1(n_689),
.A2(n_583),
.A3(n_592),
.B1(n_584),
.B2(n_526),
.C(n_527),
.Y(n_835)
);

AOI21xp5_ASAP7_75t_L g836 ( 
.A1(n_721),
.A2(n_686),
.B(n_658),
.Y(n_836)
);

INVx4_ASAP7_75t_L g837 ( 
.A(n_712),
.Y(n_837)
);

AOI21xp5_ASAP7_75t_L g838 ( 
.A1(n_700),
.A2(n_524),
.B(n_535),
.Y(n_838)
);

OAI21xp5_ASAP7_75t_L g839 ( 
.A1(n_642),
.A2(n_539),
.B(n_574),
.Y(n_839)
);

OR2x6_ASAP7_75t_L g840 ( 
.A(n_685),
.B(n_605),
.Y(n_840)
);

AOI22xp5_ASAP7_75t_L g841 ( 
.A1(n_649),
.A2(n_667),
.B1(n_671),
.B2(n_742),
.Y(n_841)
);

AOI21x1_ASAP7_75t_L g842 ( 
.A1(n_762),
.A2(n_768),
.B(n_765),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_667),
.B(n_525),
.Y(n_843)
);

NAND2x1p5_ASAP7_75t_L g844 ( 
.A(n_712),
.B(n_605),
.Y(n_844)
);

OAI22xp5_ASAP7_75t_L g845 ( 
.A1(n_729),
.A2(n_623),
.B1(n_597),
.B2(n_580),
.Y(n_845)
);

INVx2_ASAP7_75t_SL g846 ( 
.A(n_655),
.Y(n_846)
);

AOI21xp5_ASAP7_75t_L g847 ( 
.A1(n_645),
.A2(n_535),
.B(n_580),
.Y(n_847)
);

AOI21xp5_ASAP7_75t_L g848 ( 
.A1(n_653),
.A2(n_656),
.B(n_777),
.Y(n_848)
);

AOI21xp5_ASAP7_75t_L g849 ( 
.A1(n_754),
.A2(n_535),
.B(n_580),
.Y(n_849)
);

BUFx6f_ASAP7_75t_L g850 ( 
.A(n_787),
.Y(n_850)
);

AND2x6_ASAP7_75t_SL g851 ( 
.A(n_772),
.B(n_778),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_671),
.B(n_532),
.Y(n_852)
);

INVx4_ASAP7_75t_L g853 ( 
.A(n_790),
.Y(n_853)
);

OAI22xp5_ASAP7_75t_L g854 ( 
.A1(n_730),
.A2(n_623),
.B1(n_597),
.B2(n_624),
.Y(n_854)
);

INVx1_ASAP7_75t_SL g855 ( 
.A(n_663),
.Y(n_855)
);

AOI21xp33_ASAP7_75t_L g856 ( 
.A1(n_749),
.A2(n_624),
.B(n_585),
.Y(n_856)
);

NAND2xp33_ASAP7_75t_L g857 ( 
.A(n_718),
.B(n_525),
.Y(n_857)
);

NOR2xp33_ASAP7_75t_R g858 ( 
.A(n_714),
.B(n_740),
.Y(n_858)
);

OAI21x1_ASAP7_75t_L g859 ( 
.A1(n_756),
.A2(n_623),
.B(n_597),
.Y(n_859)
);

NOR3xp33_ASAP7_75t_L g860 ( 
.A(n_757),
.B(n_547),
.C(n_552),
.Y(n_860)
);

AOI21x1_ASAP7_75t_L g861 ( 
.A1(n_720),
.A2(n_616),
.B(n_585),
.Y(n_861)
);

A2O1A1Ixp33_ASAP7_75t_L g862 ( 
.A1(n_755),
.A2(n_552),
.B(n_561),
.C(n_616),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_630),
.B(n_532),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_738),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_SL g865 ( 
.A(n_790),
.B(n_616),
.Y(n_865)
);

O2A1O1Ixp33_ASAP7_75t_L g866 ( 
.A1(n_733),
.A2(n_561),
.B(n_44),
.C(n_45),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_SL g867 ( 
.A(n_635),
.B(n_616),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_793),
.B(n_532),
.Y(n_868)
);

BUFx6f_ASAP7_75t_L g869 ( 
.A(n_636),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_SL g870 ( 
.A(n_675),
.B(n_569),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_638),
.B(n_525),
.Y(n_871)
);

A2O1A1Ixp33_ASAP7_75t_L g872 ( 
.A1(n_755),
.A2(n_525),
.B(n_569),
.C(n_420),
.Y(n_872)
);

INVx3_ASAP7_75t_L g873 ( 
.A(n_789),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_632),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_743),
.B(n_525),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_706),
.Y(n_876)
);

NAND3xp33_ASAP7_75t_L g877 ( 
.A(n_675),
.B(n_420),
.C(n_412),
.Y(n_877)
);

A2O1A1Ixp33_ASAP7_75t_L g878 ( 
.A1(n_767),
.A2(n_569),
.B(n_420),
.C(n_46),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_640),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_SL g880 ( 
.A(n_789),
.B(n_569),
.Y(n_880)
);

BUFx6f_ASAP7_75t_L g881 ( 
.A(n_636),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_647),
.B(n_41),
.Y(n_882)
);

OAI21xp5_ASAP7_75t_L g883 ( 
.A1(n_642),
.A2(n_41),
.B(n_45),
.Y(n_883)
);

AO221x2_ASAP7_75t_L g884 ( 
.A1(n_782),
.A2(n_791),
.B1(n_757),
.B2(n_759),
.C(n_688),
.Y(n_884)
);

O2A1O1Ixp5_ASAP7_75t_L g885 ( 
.A1(n_774),
.A2(n_47),
.B(n_48),
.C(n_49),
.Y(n_885)
);

AND2x2_ASAP7_75t_L g886 ( 
.A(n_660),
.B(n_47),
.Y(n_886)
);

INVx3_ASAP7_75t_L g887 ( 
.A(n_681),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_643),
.B(n_52),
.Y(n_888)
);

A2O1A1Ixp33_ASAP7_75t_L g889 ( 
.A1(n_767),
.A2(n_781),
.B(n_776),
.C(n_692),
.Y(n_889)
);

OAI21xp5_ASAP7_75t_L g890 ( 
.A1(n_631),
.A2(n_53),
.B(n_54),
.Y(n_890)
);

OAI21xp33_ASAP7_75t_L g891 ( 
.A1(n_648),
.A2(n_56),
.B(n_57),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_SL g892 ( 
.A(n_788),
.B(n_745),
.Y(n_892)
);

O2A1O1Ixp5_ASAP7_75t_L g893 ( 
.A1(n_775),
.A2(n_59),
.B(n_78),
.C(n_80),
.Y(n_893)
);

AOI21xp5_ASAP7_75t_L g894 ( 
.A1(n_681),
.A2(n_88),
.B(n_91),
.Y(n_894)
);

AOI21xp5_ASAP7_75t_L g895 ( 
.A1(n_786),
.A2(n_95),
.B(n_97),
.Y(n_895)
);

INVx4_ASAP7_75t_L g896 ( 
.A(n_636),
.Y(n_896)
);

AOI21xp5_ASAP7_75t_L g897 ( 
.A1(n_786),
.A2(n_103),
.B(n_104),
.Y(n_897)
);

AOI21xp5_ASAP7_75t_L g898 ( 
.A1(n_786),
.A2(n_105),
.B(n_108),
.Y(n_898)
);

INVxp67_ASAP7_75t_L g899 ( 
.A(n_705),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_643),
.B(n_109),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_687),
.B(n_648),
.Y(n_901)
);

AOI21xp5_ASAP7_75t_L g902 ( 
.A1(n_786),
.A2(n_112),
.B(n_121),
.Y(n_902)
);

NOR3xp33_ASAP7_75t_L g903 ( 
.A(n_711),
.B(n_135),
.C(n_136),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_746),
.B(n_694),
.Y(n_904)
);

AOI21xp5_ASAP7_75t_L g905 ( 
.A1(n_654),
.A2(n_669),
.B(n_678),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_661),
.B(n_703),
.Y(n_906)
);

NOR2xp33_ASAP7_75t_L g907 ( 
.A(n_676),
.B(n_734),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_703),
.B(n_708),
.Y(n_908)
);

BUFx6f_ASAP7_75t_L g909 ( 
.A(n_665),
.Y(n_909)
);

AOI21xp5_ASAP7_75t_L g910 ( 
.A1(n_763),
.A2(n_779),
.B(n_715),
.Y(n_910)
);

AND2x2_ASAP7_75t_L g911 ( 
.A(n_726),
.B(n_734),
.Y(n_911)
);

AOI21x1_ASAP7_75t_L g912 ( 
.A1(n_736),
.A2(n_792),
.B(n_783),
.Y(n_912)
);

O2A1O1Ixp33_ASAP7_75t_L g913 ( 
.A1(n_670),
.A2(n_683),
.B(n_692),
.C(n_780),
.Y(n_913)
);

INVx3_ASAP7_75t_SL g914 ( 
.A(n_639),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_708),
.B(n_781),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_766),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_SL g917 ( 
.A(n_788),
.B(n_758),
.Y(n_917)
);

INVx2_ASAP7_75t_SL g918 ( 
.A(n_672),
.Y(n_918)
);

OAI21xp33_ASAP7_75t_L g919 ( 
.A1(n_657),
.A2(n_634),
.B(n_651),
.Y(n_919)
);

AND2x2_ASAP7_75t_L g920 ( 
.A(n_750),
.B(n_760),
.Y(n_920)
);

INVxp67_ASAP7_75t_L g921 ( 
.A(n_710),
.Y(n_921)
);

AOI22xp33_ASAP7_75t_L g922 ( 
.A1(n_770),
.A2(n_761),
.B1(n_684),
.B2(n_758),
.Y(n_922)
);

NOR2xp33_ASAP7_75t_L g923 ( 
.A(n_732),
.B(n_664),
.Y(n_923)
);

AND2x2_ASAP7_75t_L g924 ( 
.A(n_748),
.B(n_713),
.Y(n_924)
);

AOI21xp5_ASAP7_75t_L g925 ( 
.A1(n_716),
.A2(n_739),
.B(n_737),
.Y(n_925)
);

AOI21xp5_ASAP7_75t_L g926 ( 
.A1(n_752),
.A2(n_665),
.B(n_744),
.Y(n_926)
);

OAI21xp5_ASAP7_75t_L g927 ( 
.A1(n_677),
.A2(n_691),
.B(n_679),
.Y(n_927)
);

AND2x2_ASAP7_75t_L g928 ( 
.A(n_753),
.B(n_709),
.Y(n_928)
);

AO21x1_ASAP7_75t_L g929 ( 
.A1(n_736),
.A2(n_761),
.B(n_727),
.Y(n_929)
);

NOR2xp33_ASAP7_75t_L g930 ( 
.A(n_673),
.B(n_674),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_666),
.B(n_696),
.Y(n_931)
);

AND2x2_ASAP7_75t_L g932 ( 
.A(n_753),
.B(n_697),
.Y(n_932)
);

AOI21xp5_ASAP7_75t_L g933 ( 
.A1(n_665),
.A2(n_693),
.B(n_698),
.Y(n_933)
);

BUFx6f_ASAP7_75t_L g934 ( 
.A(n_731),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_707),
.B(n_719),
.Y(n_935)
);

A2O1A1Ixp33_ASAP7_75t_L g936 ( 
.A1(n_770),
.A2(n_652),
.B(n_724),
.C(n_725),
.Y(n_936)
);

AOI21xp5_ASAP7_75t_L g937 ( 
.A1(n_718),
.A2(n_735),
.B(n_723),
.Y(n_937)
);

AOI21xp33_ASAP7_75t_L g938 ( 
.A1(n_769),
.A2(n_784),
.B(n_718),
.Y(n_938)
);

BUFx6f_ASAP7_75t_L g939 ( 
.A(n_773),
.Y(n_939)
);

AOI21xp5_ASAP7_75t_L g940 ( 
.A1(n_718),
.A2(n_784),
.B(n_668),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_718),
.B(n_668),
.Y(n_941)
);

HB1xp67_ASAP7_75t_L g942 ( 
.A(n_718),
.Y(n_942)
);

AOI21xp5_ASAP7_75t_L g943 ( 
.A1(n_695),
.A2(n_722),
.B(n_728),
.Y(n_943)
);

BUFx6f_ASAP7_75t_L g944 ( 
.A(n_787),
.Y(n_944)
);

AOI21xp5_ASAP7_75t_L g945 ( 
.A1(n_695),
.A2(n_722),
.B(n_728),
.Y(n_945)
);

OAI21xp5_ASAP7_75t_L g946 ( 
.A1(n_695),
.A2(n_503),
.B(n_502),
.Y(n_946)
);

AOI21xp5_ASAP7_75t_L g947 ( 
.A1(n_695),
.A2(n_722),
.B(n_728),
.Y(n_947)
);

AO21x1_ASAP7_75t_L g948 ( 
.A1(n_662),
.A2(n_721),
.B(n_695),
.Y(n_948)
);

AOI21xp5_ASAP7_75t_L g949 ( 
.A1(n_695),
.A2(n_722),
.B(n_728),
.Y(n_949)
);

NAND3xp33_ASAP7_75t_L g950 ( 
.A(n_635),
.B(n_491),
.C(n_448),
.Y(n_950)
);

AOI21x1_ASAP7_75t_L g951 ( 
.A1(n_785),
.A2(n_762),
.B(n_722),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_690),
.B(n_650),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_690),
.B(n_633),
.Y(n_953)
);

A2O1A1Ixp33_ASAP7_75t_L g954 ( 
.A1(n_690),
.A2(n_468),
.B(n_749),
.C(n_741),
.Y(n_954)
);

O2A1O1Ixp33_ASAP7_75t_L g955 ( 
.A1(n_733),
.A2(n_670),
.B(n_644),
.C(n_515),
.Y(n_955)
);

NOR2xp33_ASAP7_75t_L g956 ( 
.A(n_635),
.B(n_334),
.Y(n_956)
);

NOR3xp33_ASAP7_75t_L g957 ( 
.A(n_757),
.B(n_578),
.C(n_513),
.Y(n_957)
);

OAI21xp5_ASAP7_75t_L g958 ( 
.A1(n_695),
.A2(n_503),
.B(n_502),
.Y(n_958)
);

NOR2xp33_ASAP7_75t_L g959 ( 
.A(n_635),
.B(n_334),
.Y(n_959)
);

BUFx6f_ASAP7_75t_L g960 ( 
.A(n_787),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_690),
.B(n_633),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_690),
.B(n_633),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_771),
.Y(n_963)
);

BUFx3_ASAP7_75t_L g964 ( 
.A(n_710),
.Y(n_964)
);

INVx2_ASAP7_75t_SL g965 ( 
.A(n_655),
.Y(n_965)
);

AND2x2_ASAP7_75t_L g966 ( 
.A(n_699),
.B(n_498),
.Y(n_966)
);

NOR2xp67_ASAP7_75t_L g967 ( 
.A(n_745),
.B(n_457),
.Y(n_967)
);

AOI21xp5_ASAP7_75t_L g968 ( 
.A1(n_695),
.A2(n_722),
.B(n_728),
.Y(n_968)
);

INVx2_ASAP7_75t_L g969 ( 
.A(n_701),
.Y(n_969)
);

AOI21xp5_ASAP7_75t_L g970 ( 
.A1(n_695),
.A2(n_722),
.B(n_728),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_SL g971 ( 
.A(n_690),
.B(n_533),
.Y(n_971)
);

AND2x2_ASAP7_75t_L g972 ( 
.A(n_699),
.B(n_498),
.Y(n_972)
);

O2A1O1Ixp33_ASAP7_75t_L g973 ( 
.A1(n_733),
.A2(n_670),
.B(n_644),
.C(n_515),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_953),
.B(n_961),
.Y(n_974)
);

AND2x4_ASAP7_75t_L g975 ( 
.A(n_840),
.B(n_837),
.Y(n_975)
);

AOI22xp5_ASAP7_75t_L g976 ( 
.A1(n_884),
.A2(n_959),
.B1(n_956),
.B2(n_841),
.Y(n_976)
);

AND2x2_ASAP7_75t_L g977 ( 
.A(n_966),
.B(n_972),
.Y(n_977)
);

AOI21xp33_ASAP7_75t_L g978 ( 
.A1(n_913),
.A2(n_919),
.B(n_915),
.Y(n_978)
);

OAI22xp5_ASAP7_75t_L g979 ( 
.A1(n_889),
.A2(n_908),
.B1(n_901),
.B2(n_963),
.Y(n_979)
);

BUFx2_ASAP7_75t_L g980 ( 
.A(n_812),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_864),
.Y(n_981)
);

INVx1_ASAP7_75t_SL g982 ( 
.A(n_855),
.Y(n_982)
);

OAI21x1_ASAP7_75t_SL g983 ( 
.A1(n_940),
.A2(n_941),
.B(n_890),
.Y(n_983)
);

HB1xp67_ASAP7_75t_L g984 ( 
.A(n_855),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_962),
.B(n_795),
.Y(n_985)
);

BUFx2_ASAP7_75t_L g986 ( 
.A(n_812),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_804),
.B(n_916),
.Y(n_987)
);

NOR2xp33_ASAP7_75t_L g988 ( 
.A(n_906),
.B(n_907),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_952),
.B(n_821),
.Y(n_989)
);

OR2x6_ASAP7_75t_L g990 ( 
.A(n_840),
.B(n_812),
.Y(n_990)
);

NOR2xp33_ASAP7_75t_R g991 ( 
.A(n_820),
.B(n_813),
.Y(n_991)
);

OAI21xp5_ASAP7_75t_L g992 ( 
.A1(n_946),
.A2(n_958),
.B(n_945),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_952),
.B(n_825),
.Y(n_993)
);

AOI22xp33_ASAP7_75t_L g994 ( 
.A1(n_884),
.A2(n_924),
.B1(n_890),
.B2(n_891),
.Y(n_994)
);

AOI21xp5_ASAP7_75t_L g995 ( 
.A1(n_946),
.A2(n_958),
.B(n_947),
.Y(n_995)
);

OR2x6_ASAP7_75t_L g996 ( 
.A(n_840),
.B(n_918),
.Y(n_996)
);

INVx2_ASAP7_75t_L g997 ( 
.A(n_811),
.Y(n_997)
);

AOI21xp5_ASAP7_75t_L g998 ( 
.A1(n_943),
.A2(n_968),
.B(n_949),
.Y(n_998)
);

OAI21x1_ASAP7_75t_L g999 ( 
.A1(n_970),
.A2(n_951),
.B(n_794),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_805),
.B(n_967),
.Y(n_1000)
);

OAI21x1_ASAP7_75t_L g1001 ( 
.A1(n_861),
.A2(n_859),
.B(n_808),
.Y(n_1001)
);

INVx2_ASAP7_75t_L g1002 ( 
.A(n_817),
.Y(n_1002)
);

INVx1_ASAP7_75t_SL g1003 ( 
.A(n_914),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_904),
.B(n_911),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_809),
.B(n_818),
.Y(n_1005)
);

AND2x2_ASAP7_75t_L g1006 ( 
.A(n_886),
.B(n_920),
.Y(n_1006)
);

NAND3xp33_ASAP7_75t_L g1007 ( 
.A(n_957),
.B(n_922),
.C(n_888),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_931),
.B(n_955),
.Y(n_1008)
);

OAI21x1_ASAP7_75t_L g1009 ( 
.A1(n_796),
.A2(n_831),
.B(n_824),
.Y(n_1009)
);

OAI21x1_ASAP7_75t_L g1010 ( 
.A1(n_836),
.A2(n_910),
.B(n_797),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_973),
.B(n_971),
.Y(n_1011)
);

OAI21x1_ASAP7_75t_SL g1012 ( 
.A1(n_948),
.A2(n_925),
.B(n_926),
.Y(n_1012)
);

INVx2_ASAP7_75t_L g1013 ( 
.A(n_876),
.Y(n_1013)
);

AND3x2_ASAP7_75t_L g1014 ( 
.A(n_921),
.B(n_928),
.C(n_932),
.Y(n_1014)
);

AO21x2_ASAP7_75t_L g1015 ( 
.A1(n_839),
.A2(n_806),
.B(n_929),
.Y(n_1015)
);

OAI22xp5_ASAP7_75t_L g1016 ( 
.A1(n_927),
.A2(n_829),
.B1(n_950),
.B2(n_930),
.Y(n_1016)
);

INVx2_ASAP7_75t_SL g1017 ( 
.A(n_964),
.Y(n_1017)
);

AOI21xp5_ASAP7_75t_L g1018 ( 
.A1(n_938),
.A2(n_849),
.B(n_798),
.Y(n_1018)
);

AOI21xp5_ASAP7_75t_SL g1019 ( 
.A1(n_896),
.A2(n_830),
.B(n_862),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_829),
.B(n_923),
.Y(n_1020)
);

A2O1A1Ixp33_ASAP7_75t_L g1021 ( 
.A1(n_927),
.A2(n_900),
.B(n_800),
.C(n_936),
.Y(n_1021)
);

O2A1O1Ixp33_ASAP7_75t_SL g1022 ( 
.A1(n_942),
.A2(n_878),
.B(n_816),
.C(n_843),
.Y(n_1022)
);

BUFx6f_ASAP7_75t_L g1023 ( 
.A(n_815),
.Y(n_1023)
);

A2O1A1Ixp33_ASAP7_75t_L g1024 ( 
.A1(n_860),
.A2(n_866),
.B(n_882),
.C(n_856),
.Y(n_1024)
);

AND2x4_ASAP7_75t_L g1025 ( 
.A(n_837),
.B(n_853),
.Y(n_1025)
);

INVx3_ASAP7_75t_L g1026 ( 
.A(n_815),
.Y(n_1026)
);

AND2x2_ASAP7_75t_L g1027 ( 
.A(n_846),
.B(n_965),
.Y(n_1027)
);

AOI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_828),
.A2(n_852),
.B(n_803),
.Y(n_1028)
);

OAI21x1_ASAP7_75t_L g1029 ( 
.A1(n_839),
.A2(n_842),
.B(n_814),
.Y(n_1029)
);

OAI21x1_ASAP7_75t_L g1030 ( 
.A1(n_806),
.A2(n_847),
.B(n_838),
.Y(n_1030)
);

O2A1O1Ixp5_ASAP7_75t_L g1031 ( 
.A1(n_883),
.A2(n_845),
.B(n_912),
.C(n_917),
.Y(n_1031)
);

AND2x2_ASAP7_75t_L g1032 ( 
.A(n_899),
.B(n_892),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_874),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_853),
.B(n_873),
.Y(n_1034)
);

OAI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_807),
.A2(n_801),
.B(n_802),
.Y(n_1035)
);

AOI21xp5_ASAP7_75t_L g1036 ( 
.A1(n_845),
.A2(n_933),
.B(n_848),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_873),
.B(n_879),
.Y(n_1037)
);

OR2x6_ASAP7_75t_L g1038 ( 
.A(n_830),
.B(n_896),
.Y(n_1038)
);

HB1xp67_ASAP7_75t_L g1039 ( 
.A(n_887),
.Y(n_1039)
);

OR2x2_ASAP7_75t_L g1040 ( 
.A(n_810),
.B(n_969),
.Y(n_1040)
);

AND2x4_ASAP7_75t_L g1041 ( 
.A(n_815),
.B(n_960),
.Y(n_1041)
);

AOI21xp5_ASAP7_75t_L g1042 ( 
.A1(n_863),
.A2(n_854),
.B(n_835),
.Y(n_1042)
);

INVx6_ASAP7_75t_L g1043 ( 
.A(n_960),
.Y(n_1043)
);

AOI221xp5_ASAP7_75t_L g1044 ( 
.A1(n_883),
.A2(n_885),
.B1(n_835),
.B2(n_856),
.C(n_854),
.Y(n_1044)
);

BUFx6f_ASAP7_75t_L g1045 ( 
.A(n_833),
.Y(n_1045)
);

AOI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_935),
.A2(n_871),
.B(n_822),
.Y(n_1046)
);

OAI21x1_ASAP7_75t_L g1047 ( 
.A1(n_893),
.A2(n_895),
.B(n_894),
.Y(n_1047)
);

A2O1A1Ixp33_ASAP7_75t_L g1048 ( 
.A1(n_832),
.A2(n_875),
.B(n_868),
.C(n_872),
.Y(n_1048)
);

OAI22xp5_ASAP7_75t_L g1049 ( 
.A1(n_867),
.A2(n_875),
.B1(n_823),
.B2(n_799),
.Y(n_1049)
);

BUFx8_ASAP7_75t_L g1050 ( 
.A(n_939),
.Y(n_1050)
);

OAI21x1_ASAP7_75t_L g1051 ( 
.A1(n_897),
.A2(n_902),
.B(n_898),
.Y(n_1051)
);

AOI22xp5_ASAP7_75t_L g1052 ( 
.A1(n_799),
.A2(n_887),
.B1(n_826),
.B2(n_865),
.Y(n_1052)
);

OAI21x1_ASAP7_75t_L g1053 ( 
.A1(n_834),
.A2(n_844),
.B(n_877),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_858),
.B(n_960),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_833),
.B(n_944),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_833),
.B(n_944),
.Y(n_1056)
);

OAI21xp5_ASAP7_75t_L g1057 ( 
.A1(n_827),
.A2(n_870),
.B(n_880),
.Y(n_1057)
);

BUFx8_ASAP7_75t_SL g1058 ( 
.A(n_939),
.Y(n_1058)
);

AND2x4_ASAP7_75t_L g1059 ( 
.A(n_850),
.B(n_944),
.Y(n_1059)
);

OAI22xp5_ASAP7_75t_L g1060 ( 
.A1(n_844),
.A2(n_850),
.B1(n_869),
.B2(n_881),
.Y(n_1060)
);

AOI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_903),
.A2(n_934),
.B(n_869),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_850),
.B(n_934),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_SL g1063 ( 
.A(n_869),
.B(n_881),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_934),
.Y(n_1064)
);

AOI21xp5_ASAP7_75t_L g1065 ( 
.A1(n_881),
.A2(n_909),
.B(n_851),
.Y(n_1065)
);

OAI21x1_ASAP7_75t_L g1066 ( 
.A1(n_909),
.A2(n_819),
.B(n_937),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_909),
.B(n_939),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_SL g1068 ( 
.A(n_841),
.B(n_533),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_953),
.B(n_961),
.Y(n_1069)
);

AOI221xp5_ASAP7_75t_L g1070 ( 
.A1(n_889),
.A2(n_733),
.B1(n_957),
.B2(n_915),
.C(n_919),
.Y(n_1070)
);

AND2x4_ASAP7_75t_SL g1071 ( 
.A(n_837),
.B(n_546),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_953),
.B(n_961),
.Y(n_1072)
);

INVx3_ASAP7_75t_L g1073 ( 
.A(n_815),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_SL g1074 ( 
.A(n_841),
.B(n_908),
.Y(n_1074)
);

OAI22xp5_ASAP7_75t_L g1075 ( 
.A1(n_889),
.A2(n_915),
.B1(n_841),
.B2(n_908),
.Y(n_1075)
);

AOI21xp5_ASAP7_75t_L g1076 ( 
.A1(n_889),
.A2(n_958),
.B(n_946),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_953),
.B(n_961),
.Y(n_1077)
);

INVx4_ASAP7_75t_L g1078 ( 
.A(n_815),
.Y(n_1078)
);

AND2x2_ASAP7_75t_L g1079 ( 
.A(n_966),
.B(n_972),
.Y(n_1079)
);

O2A1O1Ixp5_ASAP7_75t_L g1080 ( 
.A1(n_889),
.A2(n_948),
.B(n_662),
.C(n_721),
.Y(n_1080)
);

AOI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_889),
.A2(n_958),
.B(n_946),
.Y(n_1081)
);

INVx2_ASAP7_75t_L g1082 ( 
.A(n_811),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_SL g1083 ( 
.A(n_841),
.B(n_533),
.Y(n_1083)
);

AOI21x1_ASAP7_75t_SL g1084 ( 
.A1(n_915),
.A2(n_942),
.B(n_901),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_953),
.B(n_961),
.Y(n_1085)
);

AND2x4_ASAP7_75t_L g1086 ( 
.A(n_840),
.B(n_837),
.Y(n_1086)
);

AOI22xp33_ASAP7_75t_L g1087 ( 
.A1(n_884),
.A2(n_919),
.B1(n_916),
.B2(n_924),
.Y(n_1087)
);

A2O1A1Ixp33_ASAP7_75t_L g1088 ( 
.A1(n_841),
.A2(n_889),
.B(n_915),
.C(n_954),
.Y(n_1088)
);

AOI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_889),
.A2(n_958),
.B(n_946),
.Y(n_1089)
);

CKINVDCx20_ASAP7_75t_R g1090 ( 
.A(n_820),
.Y(n_1090)
);

A2O1A1Ixp33_ASAP7_75t_SL g1091 ( 
.A1(n_901),
.A2(n_776),
.B(n_781),
.C(n_767),
.Y(n_1091)
);

BUFx6f_ASAP7_75t_L g1092 ( 
.A(n_815),
.Y(n_1092)
);

BUFx6f_ASAP7_75t_L g1093 ( 
.A(n_815),
.Y(n_1093)
);

AOI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_889),
.A2(n_958),
.B(n_946),
.Y(n_1094)
);

BUFx6f_ASAP7_75t_L g1095 ( 
.A(n_815),
.Y(n_1095)
);

AOI22xp33_ASAP7_75t_L g1096 ( 
.A1(n_884),
.A2(n_919),
.B1(n_916),
.B2(n_924),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_953),
.B(n_961),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_953),
.B(n_961),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_953),
.B(n_961),
.Y(n_1099)
);

AND2x2_ASAP7_75t_L g1100 ( 
.A(n_966),
.B(n_972),
.Y(n_1100)
);

A2O1A1Ixp33_ASAP7_75t_L g1101 ( 
.A1(n_841),
.A2(n_889),
.B(n_915),
.C(n_954),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_864),
.Y(n_1102)
);

BUFx6f_ASAP7_75t_L g1103 ( 
.A(n_815),
.Y(n_1103)
);

AOI21x1_ASAP7_75t_L g1104 ( 
.A1(n_912),
.A2(n_905),
.B(n_796),
.Y(n_1104)
);

NOR2x1_ASAP7_75t_R g1105 ( 
.A(n_820),
.B(n_440),
.Y(n_1105)
);

NOR2x1_ASAP7_75t_L g1106 ( 
.A(n_964),
.B(n_533),
.Y(n_1106)
);

INVx1_ASAP7_75t_SL g1107 ( 
.A(n_982),
.Y(n_1107)
);

INVx2_ASAP7_75t_L g1108 ( 
.A(n_1002),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_981),
.Y(n_1109)
);

AND2x4_ASAP7_75t_L g1110 ( 
.A(n_990),
.B(n_975),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_1020),
.B(n_1074),
.Y(n_1111)
);

OAI22xp5_ASAP7_75t_L g1112 ( 
.A1(n_976),
.A2(n_994),
.B1(n_1075),
.B2(n_1088),
.Y(n_1112)
);

HB1xp67_ASAP7_75t_L g1113 ( 
.A(n_977),
.Y(n_1113)
);

AOI21xp5_ASAP7_75t_SL g1114 ( 
.A1(n_1021),
.A2(n_1008),
.B(n_979),
.Y(n_1114)
);

INVx2_ASAP7_75t_SL g1115 ( 
.A(n_1003),
.Y(n_1115)
);

INVx2_ASAP7_75t_SL g1116 ( 
.A(n_984),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_1102),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_1074),
.B(n_989),
.Y(n_1118)
);

CKINVDCx5p33_ASAP7_75t_R g1119 ( 
.A(n_1058),
.Y(n_1119)
);

CKINVDCx5p33_ASAP7_75t_R g1120 ( 
.A(n_991),
.Y(n_1120)
);

OAI21xp33_ASAP7_75t_SL g1121 ( 
.A1(n_1070),
.A2(n_978),
.B(n_994),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_SL g1122 ( 
.A(n_988),
.B(n_1070),
.Y(n_1122)
);

AOI222xp33_ASAP7_75t_L g1123 ( 
.A1(n_1087),
.A2(n_1096),
.B1(n_988),
.B2(n_1016),
.C1(n_1085),
.C2(n_1097),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_974),
.B(n_1069),
.Y(n_1124)
);

AOI22xp33_ASAP7_75t_L g1125 ( 
.A1(n_1087),
.A2(n_1096),
.B1(n_1007),
.B2(n_1006),
.Y(n_1125)
);

HB1xp67_ASAP7_75t_L g1126 ( 
.A(n_1079),
.Y(n_1126)
);

OAI22xp5_ASAP7_75t_L g1127 ( 
.A1(n_1072),
.A2(n_1077),
.B1(n_1098),
.B2(n_1099),
.Y(n_1127)
);

INVx2_ASAP7_75t_L g1128 ( 
.A(n_1013),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_1033),
.Y(n_1129)
);

A2O1A1Ixp33_ASAP7_75t_L g1130 ( 
.A1(n_1044),
.A2(n_1080),
.B(n_1083),
.C(n_1068),
.Y(n_1130)
);

AOI22xp33_ASAP7_75t_L g1131 ( 
.A1(n_1100),
.A2(n_1082),
.B1(n_1005),
.B2(n_985),
.Y(n_1131)
);

A2O1A1Ixp33_ASAP7_75t_L g1132 ( 
.A1(n_1044),
.A2(n_1080),
.B(n_1091),
.C(n_1011),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_993),
.B(n_1040),
.Y(n_1133)
);

AOI22xp5_ASAP7_75t_L g1134 ( 
.A1(n_1004),
.A2(n_1032),
.B1(n_984),
.B2(n_1027),
.Y(n_1134)
);

INVx5_ASAP7_75t_L g1135 ( 
.A(n_990),
.Y(n_1135)
);

O2A1O1Ixp33_ASAP7_75t_L g1136 ( 
.A1(n_1091),
.A2(n_1024),
.B(n_1022),
.C(n_1000),
.Y(n_1136)
);

AOI221x1_ASAP7_75t_L g1137 ( 
.A1(n_1076),
.A2(n_1094),
.B1(n_1089),
.B2(n_1081),
.C(n_998),
.Y(n_1137)
);

CKINVDCx5p33_ASAP7_75t_R g1138 ( 
.A(n_991),
.Y(n_1138)
);

AOI21xp5_ASAP7_75t_L g1139 ( 
.A1(n_1036),
.A2(n_1028),
.B(n_1019),
.Y(n_1139)
);

BUFx2_ASAP7_75t_L g1140 ( 
.A(n_1105),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_987),
.B(n_1076),
.Y(n_1141)
);

BUFx10_ASAP7_75t_L g1142 ( 
.A(n_1071),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_1081),
.B(n_1089),
.Y(n_1143)
);

AOI21xp5_ASAP7_75t_L g1144 ( 
.A1(n_1028),
.A2(n_1035),
.B(n_1018),
.Y(n_1144)
);

AO32x2_ASAP7_75t_L g1145 ( 
.A1(n_1049),
.A2(n_1094),
.A3(n_1084),
.B1(n_1015),
.B2(n_995),
.Y(n_1145)
);

AOI21xp5_ASAP7_75t_L g1146 ( 
.A1(n_1018),
.A2(n_995),
.B(n_992),
.Y(n_1146)
);

INVx2_ASAP7_75t_SL g1147 ( 
.A(n_1017),
.Y(n_1147)
);

AND2x2_ASAP7_75t_L g1148 ( 
.A(n_980),
.B(n_986),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_1037),
.Y(n_1149)
);

INVx1_ASAP7_75t_SL g1150 ( 
.A(n_1067),
.Y(n_1150)
);

BUFx6f_ASAP7_75t_L g1151 ( 
.A(n_975),
.Y(n_1151)
);

AOI222xp33_ASAP7_75t_L g1152 ( 
.A1(n_1050),
.A2(n_1086),
.B1(n_1054),
.B2(n_1025),
.C1(n_1106),
.C2(n_1090),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_1039),
.B(n_1086),
.Y(n_1153)
);

AND2x2_ASAP7_75t_L g1154 ( 
.A(n_996),
.B(n_1014),
.Y(n_1154)
);

AND2x2_ASAP7_75t_L g1155 ( 
.A(n_996),
.B(n_1014),
.Y(n_1155)
);

INVx4_ASAP7_75t_L g1156 ( 
.A(n_1023),
.Y(n_1156)
);

AND2x2_ASAP7_75t_L g1157 ( 
.A(n_996),
.B(n_1064),
.Y(n_1157)
);

AOI221xp5_ASAP7_75t_L g1158 ( 
.A1(n_1031),
.A2(n_1042),
.B1(n_983),
.B2(n_1048),
.C(n_1057),
.Y(n_1158)
);

INVx3_ASAP7_75t_L g1159 ( 
.A(n_1038),
.Y(n_1159)
);

BUFx2_ASAP7_75t_L g1160 ( 
.A(n_1050),
.Y(n_1160)
);

BUFx10_ASAP7_75t_L g1161 ( 
.A(n_1043),
.Y(n_1161)
);

INVx4_ASAP7_75t_L g1162 ( 
.A(n_1023),
.Y(n_1162)
);

AOI21xp33_ASAP7_75t_L g1163 ( 
.A1(n_1031),
.A2(n_1015),
.B(n_1012),
.Y(n_1163)
);

AO22x1_ASAP7_75t_L g1164 ( 
.A1(n_1041),
.A2(n_1059),
.B1(n_1062),
.B2(n_1073),
.Y(n_1164)
);

INVx4_ASAP7_75t_L g1165 ( 
.A(n_1023),
.Y(n_1165)
);

AND2x2_ASAP7_75t_L g1166 ( 
.A(n_1039),
.B(n_1052),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_SL g1167 ( 
.A(n_1034),
.B(n_1023),
.Y(n_1167)
);

INVx4_ASAP7_75t_L g1168 ( 
.A(n_1045),
.Y(n_1168)
);

BUFx6f_ASAP7_75t_L g1169 ( 
.A(n_1045),
.Y(n_1169)
);

BUFx3_ASAP7_75t_L g1170 ( 
.A(n_1043),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_1046),
.B(n_1065),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1043),
.Y(n_1172)
);

AND2x4_ASAP7_75t_L g1173 ( 
.A(n_1065),
.B(n_1078),
.Y(n_1173)
);

AND2x4_ASAP7_75t_L g1174 ( 
.A(n_1078),
.B(n_1026),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_1061),
.B(n_1073),
.Y(n_1175)
);

INVx3_ASAP7_75t_L g1176 ( 
.A(n_1045),
.Y(n_1176)
);

AND2x4_ASAP7_75t_L g1177 ( 
.A(n_1045),
.B(n_1103),
.Y(n_1177)
);

AOI22xp5_ASAP7_75t_L g1178 ( 
.A1(n_1063),
.A2(n_1056),
.B1(n_1055),
.B2(n_1060),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_1061),
.B(n_1093),
.Y(n_1179)
);

NAND2x1p5_ASAP7_75t_L g1180 ( 
.A(n_1092),
.B(n_1093),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_SL g1181 ( 
.A(n_1092),
.B(n_1103),
.Y(n_1181)
);

AND2x4_ASAP7_75t_L g1182 ( 
.A(n_1092),
.B(n_1103),
.Y(n_1182)
);

INVx5_ASAP7_75t_L g1183 ( 
.A(n_1093),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_1093),
.Y(n_1184)
);

NOR2xp33_ASAP7_75t_L g1185 ( 
.A(n_1095),
.B(n_1103),
.Y(n_1185)
);

AND2x2_ASAP7_75t_L g1186 ( 
.A(n_1095),
.B(n_1053),
.Y(n_1186)
);

AND2x4_ASAP7_75t_L g1187 ( 
.A(n_1095),
.B(n_1051),
.Y(n_1187)
);

AND2x2_ASAP7_75t_L g1188 ( 
.A(n_1095),
.B(n_1029),
.Y(n_1188)
);

AO21x1_ASAP7_75t_L g1189 ( 
.A1(n_1104),
.A2(n_1047),
.B(n_1030),
.Y(n_1189)
);

NAND3xp33_ASAP7_75t_L g1190 ( 
.A(n_1084),
.B(n_999),
.C(n_1010),
.Y(n_1190)
);

INVx1_ASAP7_75t_SL g1191 ( 
.A(n_1066),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_1001),
.B(n_1009),
.Y(n_1192)
);

INVx3_ASAP7_75t_L g1193 ( 
.A(n_1038),
.Y(n_1193)
);

OAI321xp33_ASAP7_75t_L g1194 ( 
.A1(n_1016),
.A2(n_994),
.A3(n_1070),
.B1(n_1075),
.B2(n_976),
.C(n_1020),
.Y(n_1194)
);

BUFx12f_ASAP7_75t_L g1195 ( 
.A(n_1050),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_1020),
.B(n_1074),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_981),
.Y(n_1197)
);

INVx5_ASAP7_75t_L g1198 ( 
.A(n_990),
.Y(n_1198)
);

CKINVDCx20_ASAP7_75t_R g1199 ( 
.A(n_1090),
.Y(n_1199)
);

BUFx2_ASAP7_75t_L g1200 ( 
.A(n_977),
.Y(n_1200)
);

INVx3_ASAP7_75t_SL g1201 ( 
.A(n_1090),
.Y(n_1201)
);

BUFx6f_ASAP7_75t_L g1202 ( 
.A(n_975),
.Y(n_1202)
);

OAI22xp5_ASAP7_75t_L g1203 ( 
.A1(n_976),
.A2(n_915),
.B1(n_889),
.B2(n_1020),
.Y(n_1203)
);

BUFx3_ASAP7_75t_L g1204 ( 
.A(n_1003),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_1020),
.B(n_1074),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_SL g1206 ( 
.A(n_988),
.B(n_841),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_1020),
.B(n_1074),
.Y(n_1207)
);

BUFx3_ASAP7_75t_L g1208 ( 
.A(n_1003),
.Y(n_1208)
);

NOR2xp33_ASAP7_75t_SL g1209 ( 
.A(n_1007),
.B(n_813),
.Y(n_1209)
);

INVx4_ASAP7_75t_L g1210 ( 
.A(n_1025),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_981),
.Y(n_1211)
);

INVx2_ASAP7_75t_SL g1212 ( 
.A(n_1003),
.Y(n_1212)
);

CKINVDCx6p67_ASAP7_75t_R g1213 ( 
.A(n_1090),
.Y(n_1213)
);

CKINVDCx5p33_ASAP7_75t_R g1214 ( 
.A(n_1058),
.Y(n_1214)
);

INVx2_ASAP7_75t_SL g1215 ( 
.A(n_1003),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_974),
.B(n_1069),
.Y(n_1216)
);

AOI21xp5_ASAP7_75t_L g1217 ( 
.A1(n_1021),
.A2(n_1075),
.B(n_857),
.Y(n_1217)
);

BUFx6f_ASAP7_75t_L g1218 ( 
.A(n_975),
.Y(n_1218)
);

INVx2_ASAP7_75t_L g1219 ( 
.A(n_997),
.Y(n_1219)
);

AOI22xp33_ASAP7_75t_L g1220 ( 
.A1(n_994),
.A2(n_414),
.B1(n_425),
.B2(n_884),
.Y(n_1220)
);

O2A1O1Ixp33_ASAP7_75t_L g1221 ( 
.A1(n_1075),
.A2(n_889),
.B(n_1101),
.C(n_1088),
.Y(n_1221)
);

BUFx3_ASAP7_75t_L g1222 ( 
.A(n_1003),
.Y(n_1222)
);

NOR2x1_ASAP7_75t_L g1223 ( 
.A(n_1054),
.B(n_964),
.Y(n_1223)
);

AND2x4_ASAP7_75t_L g1224 ( 
.A(n_990),
.B(n_975),
.Y(n_1224)
);

OR2x2_ASAP7_75t_L g1225 ( 
.A(n_977),
.B(n_1079),
.Y(n_1225)
);

NOR2xp67_ASAP7_75t_L g1226 ( 
.A(n_984),
.B(n_745),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_981),
.Y(n_1227)
);

AOI22xp5_ASAP7_75t_L g1228 ( 
.A1(n_976),
.A2(n_590),
.B1(n_884),
.B2(n_514),
.Y(n_1228)
);

AOI22xp33_ASAP7_75t_L g1229 ( 
.A1(n_994),
.A2(n_414),
.B1(n_425),
.B2(n_884),
.Y(n_1229)
);

INVx2_ASAP7_75t_L g1230 ( 
.A(n_997),
.Y(n_1230)
);

AND2x2_ASAP7_75t_L g1231 ( 
.A(n_977),
.B(n_1079),
.Y(n_1231)
);

BUFx2_ASAP7_75t_L g1232 ( 
.A(n_977),
.Y(n_1232)
);

INVxp67_ASAP7_75t_SL g1233 ( 
.A(n_984),
.Y(n_1233)
);

BUFx3_ASAP7_75t_L g1234 ( 
.A(n_1003),
.Y(n_1234)
);

OR2x6_ASAP7_75t_L g1235 ( 
.A(n_990),
.B(n_840),
.Y(n_1235)
);

OAI22xp5_ASAP7_75t_L g1236 ( 
.A1(n_976),
.A2(n_915),
.B1(n_889),
.B2(n_1020),
.Y(n_1236)
);

INVx2_ASAP7_75t_L g1237 ( 
.A(n_997),
.Y(n_1237)
);

HB1xp67_ASAP7_75t_L g1238 ( 
.A(n_977),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_1020),
.B(n_1074),
.Y(n_1239)
);

CKINVDCx20_ASAP7_75t_R g1240 ( 
.A(n_1090),
.Y(n_1240)
);

AOI21xp5_ASAP7_75t_L g1241 ( 
.A1(n_1021),
.A2(n_1075),
.B(n_857),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1143),
.Y(n_1242)
);

AND2x4_ASAP7_75t_L g1243 ( 
.A(n_1110),
.B(n_1224),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1141),
.Y(n_1244)
);

BUFx3_ASAP7_75t_L g1245 ( 
.A(n_1170),
.Y(n_1245)
);

AO21x1_ASAP7_75t_L g1246 ( 
.A1(n_1112),
.A2(n_1122),
.B(n_1203),
.Y(n_1246)
);

AND2x4_ASAP7_75t_L g1247 ( 
.A(n_1110),
.B(n_1224),
.Y(n_1247)
);

OAI22xp5_ASAP7_75t_L g1248 ( 
.A1(n_1228),
.A2(n_1206),
.B1(n_1112),
.B2(n_1236),
.Y(n_1248)
);

OAI21x1_ASAP7_75t_L g1249 ( 
.A1(n_1144),
.A2(n_1139),
.B(n_1146),
.Y(n_1249)
);

HB1xp67_ASAP7_75t_L g1250 ( 
.A(n_1113),
.Y(n_1250)
);

INVx1_ASAP7_75t_SL g1251 ( 
.A(n_1231),
.Y(n_1251)
);

CKINVDCx11_ASAP7_75t_R g1252 ( 
.A(n_1199),
.Y(n_1252)
);

INVx4_ASAP7_75t_L g1253 ( 
.A(n_1183),
.Y(n_1253)
);

AOI22xp33_ASAP7_75t_L g1254 ( 
.A1(n_1123),
.A2(n_1220),
.B1(n_1229),
.B2(n_1125),
.Y(n_1254)
);

OR2x2_ASAP7_75t_L g1255 ( 
.A(n_1233),
.B(n_1111),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1109),
.Y(n_1256)
);

AOI22xp33_ASAP7_75t_L g1257 ( 
.A1(n_1123),
.A2(n_1236),
.B1(n_1203),
.B2(n_1209),
.Y(n_1257)
);

BUFx2_ASAP7_75t_R g1258 ( 
.A(n_1119),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_1124),
.B(n_1127),
.Y(n_1259)
);

INVx1_ASAP7_75t_SL g1260 ( 
.A(n_1225),
.Y(n_1260)
);

AOI22xp33_ASAP7_75t_L g1261 ( 
.A1(n_1209),
.A2(n_1121),
.B1(n_1131),
.B2(n_1127),
.Y(n_1261)
);

AOI22xp33_ASAP7_75t_SL g1262 ( 
.A1(n_1154),
.A2(n_1155),
.B1(n_1194),
.B2(n_1239),
.Y(n_1262)
);

BUFx2_ASAP7_75t_R g1263 ( 
.A(n_1214),
.Y(n_1263)
);

HB1xp67_ASAP7_75t_L g1264 ( 
.A(n_1126),
.Y(n_1264)
);

BUFx3_ASAP7_75t_L g1265 ( 
.A(n_1151),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1171),
.Y(n_1266)
);

HB1xp67_ASAP7_75t_L g1267 ( 
.A(n_1238),
.Y(n_1267)
);

BUFx2_ASAP7_75t_SL g1268 ( 
.A(n_1183),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1145),
.Y(n_1269)
);

CKINVDCx16_ASAP7_75t_R g1270 ( 
.A(n_1240),
.Y(n_1270)
);

AO21x2_ASAP7_75t_L g1271 ( 
.A1(n_1163),
.A2(n_1132),
.B(n_1190),
.Y(n_1271)
);

BUFx3_ASAP7_75t_L g1272 ( 
.A(n_1202),
.Y(n_1272)
);

INVx1_ASAP7_75t_SL g1273 ( 
.A(n_1200),
.Y(n_1273)
);

AND2x4_ASAP7_75t_L g1274 ( 
.A(n_1235),
.B(n_1135),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1145),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1117),
.Y(n_1276)
);

AOI21xp33_ASAP7_75t_SL g1277 ( 
.A1(n_1201),
.A2(n_1138),
.B(n_1120),
.Y(n_1277)
);

AOI22xp33_ASAP7_75t_SL g1278 ( 
.A1(n_1194),
.A2(n_1239),
.B1(n_1196),
.B2(n_1111),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1129),
.Y(n_1279)
);

INVx1_ASAP7_75t_SL g1280 ( 
.A(n_1232),
.Y(n_1280)
);

AOI22xp33_ASAP7_75t_L g1281 ( 
.A1(n_1108),
.A2(n_1219),
.B1(n_1237),
.B2(n_1128),
.Y(n_1281)
);

AOI22xp33_ASAP7_75t_SL g1282 ( 
.A1(n_1196),
.A2(n_1205),
.B1(n_1207),
.B2(n_1217),
.Y(n_1282)
);

AOI21x1_ASAP7_75t_L g1283 ( 
.A1(n_1192),
.A2(n_1189),
.B(n_1241),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1197),
.Y(n_1284)
);

AOI22xp33_ASAP7_75t_L g1285 ( 
.A1(n_1230),
.A2(n_1124),
.B1(n_1216),
.B2(n_1134),
.Y(n_1285)
);

OAI22xp5_ASAP7_75t_L g1286 ( 
.A1(n_1221),
.A2(n_1114),
.B1(n_1118),
.B2(n_1205),
.Y(n_1286)
);

HB1xp67_ASAP7_75t_L g1287 ( 
.A(n_1116),
.Y(n_1287)
);

CKINVDCx16_ASAP7_75t_R g1288 ( 
.A(n_1195),
.Y(n_1288)
);

AOI22xp33_ASAP7_75t_L g1289 ( 
.A1(n_1166),
.A2(n_1207),
.B1(n_1133),
.B2(n_1150),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1211),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1227),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_L g1292 ( 
.A(n_1133),
.B(n_1118),
.Y(n_1292)
);

INVx2_ASAP7_75t_L g1293 ( 
.A(n_1188),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1149),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1145),
.Y(n_1295)
);

INVx1_ASAP7_75t_SL g1296 ( 
.A(n_1107),
.Y(n_1296)
);

INVx2_ASAP7_75t_SL g1297 ( 
.A(n_1183),
.Y(n_1297)
);

HB1xp67_ASAP7_75t_L g1298 ( 
.A(n_1153),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1153),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1157),
.Y(n_1300)
);

BUFx6f_ASAP7_75t_L g1301 ( 
.A(n_1202),
.Y(n_1301)
);

AND2x2_ASAP7_75t_L g1302 ( 
.A(n_1130),
.B(n_1186),
.Y(n_1302)
);

OAI21x1_ASAP7_75t_L g1303 ( 
.A1(n_1137),
.A2(n_1136),
.B(n_1179),
.Y(n_1303)
);

OA21x2_ASAP7_75t_L g1304 ( 
.A1(n_1163),
.A2(n_1158),
.B(n_1175),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1148),
.Y(n_1305)
);

AOI22xp33_ASAP7_75t_L g1306 ( 
.A1(n_1152),
.A2(n_1235),
.B1(n_1107),
.B2(n_1226),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1184),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_L g1308 ( 
.A(n_1210),
.B(n_1218),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1179),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1167),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1164),
.Y(n_1311)
);

BUFx12f_ASAP7_75t_L g1312 ( 
.A(n_1160),
.Y(n_1312)
);

AO21x2_ASAP7_75t_L g1313 ( 
.A1(n_1187),
.A2(n_1178),
.B(n_1181),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_L g1314 ( 
.A(n_1210),
.B(n_1218),
.Y(n_1314)
);

INVx3_ASAP7_75t_L g1315 ( 
.A(n_1169),
.Y(n_1315)
);

BUFx2_ASAP7_75t_L g1316 ( 
.A(n_1191),
.Y(n_1316)
);

INVx2_ASAP7_75t_L g1317 ( 
.A(n_1191),
.Y(n_1317)
);

OAI22xp5_ASAP7_75t_L g1318 ( 
.A1(n_1115),
.A2(n_1215),
.B1(n_1212),
.B2(n_1235),
.Y(n_1318)
);

AOI22xp5_ASAP7_75t_L g1319 ( 
.A1(n_1152),
.A2(n_1140),
.B1(n_1234),
.B2(n_1222),
.Y(n_1319)
);

HB1xp67_ASAP7_75t_L g1320 ( 
.A(n_1169),
.Y(n_1320)
);

BUFx3_ASAP7_75t_L g1321 ( 
.A(n_1202),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1159),
.Y(n_1322)
);

INVx3_ASAP7_75t_L g1323 ( 
.A(n_1169),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1193),
.Y(n_1324)
);

AOI22xp33_ASAP7_75t_L g1325 ( 
.A1(n_1198),
.A2(n_1204),
.B1(n_1208),
.B2(n_1173),
.Y(n_1325)
);

INVx2_ASAP7_75t_L g1326 ( 
.A(n_1173),
.Y(n_1326)
);

INVx4_ASAP7_75t_L g1327 ( 
.A(n_1177),
.Y(n_1327)
);

INVx1_ASAP7_75t_SL g1328 ( 
.A(n_1213),
.Y(n_1328)
);

OA21x2_ASAP7_75t_L g1329 ( 
.A1(n_1185),
.A2(n_1172),
.B(n_1177),
.Y(n_1329)
);

INVx1_ASAP7_75t_SL g1330 ( 
.A(n_1223),
.Y(n_1330)
);

OAI21xp5_ASAP7_75t_L g1331 ( 
.A1(n_1147),
.A2(n_1180),
.B(n_1176),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1182),
.Y(n_1332)
);

AOI22xp33_ASAP7_75t_L g1333 ( 
.A1(n_1174),
.A2(n_1142),
.B1(n_1156),
.B2(n_1162),
.Y(n_1333)
);

AND2x4_ASAP7_75t_L g1334 ( 
.A(n_1156),
.B(n_1162),
.Y(n_1334)
);

AND2x2_ASAP7_75t_L g1335 ( 
.A(n_1165),
.B(n_1168),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1165),
.Y(n_1336)
);

AOI21xp5_ASAP7_75t_SL g1337 ( 
.A1(n_1168),
.A2(n_1174),
.B(n_1142),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1161),
.Y(n_1338)
);

AOI22xp33_ASAP7_75t_L g1339 ( 
.A1(n_1161),
.A2(n_1123),
.B1(n_884),
.B2(n_414),
.Y(n_1339)
);

BUFx6f_ASAP7_75t_L g1340 ( 
.A(n_1151),
.Y(n_1340)
);

NOR2xp33_ASAP7_75t_L g1341 ( 
.A(n_1228),
.B(n_590),
.Y(n_1341)
);

AO21x1_ASAP7_75t_SL g1342 ( 
.A1(n_1143),
.A2(n_1163),
.B(n_1239),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1143),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1143),
.Y(n_1344)
);

OAI22xp5_ASAP7_75t_L g1345 ( 
.A1(n_1228),
.A2(n_976),
.B1(n_841),
.B2(n_915),
.Y(n_1345)
);

BUFx8_ASAP7_75t_L g1346 ( 
.A(n_1195),
.Y(n_1346)
);

AND2x2_ASAP7_75t_L g1347 ( 
.A(n_1112),
.B(n_1141),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1143),
.Y(n_1348)
);

CKINVDCx5p33_ASAP7_75t_R g1349 ( 
.A(n_1195),
.Y(n_1349)
);

OAI21xp5_ASAP7_75t_L g1350 ( 
.A1(n_1122),
.A2(n_889),
.B(n_976),
.Y(n_1350)
);

AND2x2_ASAP7_75t_L g1351 ( 
.A(n_1112),
.B(n_1141),
.Y(n_1351)
);

INVx4_ASAP7_75t_L g1352 ( 
.A(n_1183),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1143),
.Y(n_1353)
);

INVx3_ASAP7_75t_L g1354 ( 
.A(n_1187),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1143),
.Y(n_1355)
);

INVx2_ASAP7_75t_SL g1356 ( 
.A(n_1183),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1143),
.Y(n_1357)
);

HB1xp67_ASAP7_75t_L g1358 ( 
.A(n_1316),
.Y(n_1358)
);

OAI221xp5_ASAP7_75t_L g1359 ( 
.A1(n_1257),
.A2(n_1350),
.B1(n_1339),
.B2(n_1345),
.C(n_1248),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1309),
.Y(n_1360)
);

AND2x2_ASAP7_75t_L g1361 ( 
.A(n_1347),
.B(n_1351),
.Y(n_1361)
);

AND2x2_ASAP7_75t_L g1362 ( 
.A(n_1347),
.B(n_1351),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1266),
.Y(n_1363)
);

AND2x2_ASAP7_75t_L g1364 ( 
.A(n_1293),
.B(n_1242),
.Y(n_1364)
);

HB1xp67_ASAP7_75t_L g1365 ( 
.A(n_1316),
.Y(n_1365)
);

INVx3_ASAP7_75t_L g1366 ( 
.A(n_1249),
.Y(n_1366)
);

BUFx3_ASAP7_75t_L g1367 ( 
.A(n_1354),
.Y(n_1367)
);

OR2x2_ASAP7_75t_L g1368 ( 
.A(n_1269),
.B(n_1275),
.Y(n_1368)
);

AND2x2_ASAP7_75t_L g1369 ( 
.A(n_1343),
.B(n_1344),
.Y(n_1369)
);

BUFx2_ASAP7_75t_L g1370 ( 
.A(n_1249),
.Y(n_1370)
);

OR2x2_ASAP7_75t_L g1371 ( 
.A(n_1295),
.B(n_1348),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1353),
.Y(n_1372)
);

AND2x2_ASAP7_75t_L g1373 ( 
.A(n_1353),
.B(n_1355),
.Y(n_1373)
);

CKINVDCx20_ASAP7_75t_R g1374 ( 
.A(n_1252),
.Y(n_1374)
);

INVx2_ASAP7_75t_L g1375 ( 
.A(n_1357),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1244),
.Y(n_1376)
);

INVx3_ASAP7_75t_L g1377 ( 
.A(n_1303),
.Y(n_1377)
);

AO21x2_ASAP7_75t_L g1378 ( 
.A1(n_1271),
.A2(n_1246),
.B(n_1283),
.Y(n_1378)
);

AND2x2_ASAP7_75t_L g1379 ( 
.A(n_1342),
.B(n_1304),
.Y(n_1379)
);

INVx1_ASAP7_75t_SL g1380 ( 
.A(n_1296),
.Y(n_1380)
);

BUFx2_ASAP7_75t_L g1381 ( 
.A(n_1271),
.Y(n_1381)
);

AND2x2_ASAP7_75t_L g1382 ( 
.A(n_1342),
.B(n_1304),
.Y(n_1382)
);

BUFx2_ASAP7_75t_L g1383 ( 
.A(n_1271),
.Y(n_1383)
);

INVx2_ASAP7_75t_L g1384 ( 
.A(n_1304),
.Y(n_1384)
);

OAI22xp33_ASAP7_75t_L g1385 ( 
.A1(n_1259),
.A2(n_1341),
.B1(n_1251),
.B2(n_1286),
.Y(n_1385)
);

INVx1_ASAP7_75t_SL g1386 ( 
.A(n_1255),
.Y(n_1386)
);

OAI21xp5_ASAP7_75t_L g1387 ( 
.A1(n_1261),
.A2(n_1278),
.B(n_1254),
.Y(n_1387)
);

AND2x2_ASAP7_75t_L g1388 ( 
.A(n_1302),
.B(n_1317),
.Y(n_1388)
);

AND2x2_ASAP7_75t_L g1389 ( 
.A(n_1302),
.B(n_1282),
.Y(n_1389)
);

INVx5_ASAP7_75t_L g1390 ( 
.A(n_1253),
.Y(n_1390)
);

BUFx3_ASAP7_75t_L g1391 ( 
.A(n_1329),
.Y(n_1391)
);

AO21x2_ASAP7_75t_L g1392 ( 
.A1(n_1246),
.A2(n_1313),
.B(n_1310),
.Y(n_1392)
);

AND2x4_ASAP7_75t_L g1393 ( 
.A(n_1326),
.B(n_1274),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_L g1394 ( 
.A(n_1255),
.B(n_1292),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1256),
.Y(n_1395)
);

AND2x2_ASAP7_75t_L g1396 ( 
.A(n_1276),
.B(n_1279),
.Y(n_1396)
);

NAND2xp5_ASAP7_75t_L g1397 ( 
.A(n_1298),
.B(n_1299),
.Y(n_1397)
);

HB1xp67_ASAP7_75t_L g1398 ( 
.A(n_1250),
.Y(n_1398)
);

AO21x2_ASAP7_75t_L g1399 ( 
.A1(n_1284),
.A2(n_1290),
.B(n_1291),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1294),
.Y(n_1400)
);

BUFx12f_ASAP7_75t_L g1401 ( 
.A(n_1252),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1307),
.Y(n_1402)
);

OR2x2_ASAP7_75t_L g1403 ( 
.A(n_1264),
.B(n_1267),
.Y(n_1403)
);

HB1xp67_ASAP7_75t_L g1404 ( 
.A(n_1287),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_L g1405 ( 
.A(n_1289),
.B(n_1285),
.Y(n_1405)
);

AND2x2_ASAP7_75t_L g1406 ( 
.A(n_1305),
.B(n_1260),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1322),
.Y(n_1407)
);

BUFx3_ASAP7_75t_L g1408 ( 
.A(n_1274),
.Y(n_1408)
);

HB1xp67_ASAP7_75t_L g1409 ( 
.A(n_1324),
.Y(n_1409)
);

INVx2_ASAP7_75t_L g1410 ( 
.A(n_1311),
.Y(n_1410)
);

AO21x2_ASAP7_75t_L g1411 ( 
.A1(n_1331),
.A2(n_1332),
.B(n_1300),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1336),
.Y(n_1412)
);

NOR2xp33_ASAP7_75t_L g1413 ( 
.A(n_1273),
.B(n_1280),
.Y(n_1413)
);

INVx2_ASAP7_75t_L g1414 ( 
.A(n_1336),
.Y(n_1414)
);

INVx4_ASAP7_75t_SL g1415 ( 
.A(n_1274),
.Y(n_1415)
);

AND2x2_ASAP7_75t_L g1416 ( 
.A(n_1262),
.B(n_1327),
.Y(n_1416)
);

HB1xp67_ASAP7_75t_L g1417 ( 
.A(n_1320),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_L g1418 ( 
.A(n_1306),
.B(n_1325),
.Y(n_1418)
);

AND2x2_ASAP7_75t_L g1419 ( 
.A(n_1361),
.B(n_1323),
.Y(n_1419)
);

INVx2_ASAP7_75t_SL g1420 ( 
.A(n_1403),
.Y(n_1420)
);

OAI22xp5_ASAP7_75t_L g1421 ( 
.A1(n_1359),
.A2(n_1319),
.B1(n_1270),
.B2(n_1333),
.Y(n_1421)
);

INVx2_ASAP7_75t_SL g1422 ( 
.A(n_1403),
.Y(n_1422)
);

INVx5_ASAP7_75t_SL g1423 ( 
.A(n_1392),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1399),
.Y(n_1424)
);

AND2x2_ASAP7_75t_L g1425 ( 
.A(n_1361),
.B(n_1362),
.Y(n_1425)
);

AND2x2_ASAP7_75t_L g1426 ( 
.A(n_1361),
.B(n_1323),
.Y(n_1426)
);

BUFx3_ASAP7_75t_L g1427 ( 
.A(n_1401),
.Y(n_1427)
);

BUFx3_ASAP7_75t_L g1428 ( 
.A(n_1401),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1399),
.Y(n_1429)
);

NOR2x1_ASAP7_75t_L g1430 ( 
.A(n_1414),
.B(n_1337),
.Y(n_1430)
);

NAND2xp5_ASAP7_75t_L g1431 ( 
.A(n_1394),
.B(n_1245),
.Y(n_1431)
);

NAND3xp33_ASAP7_75t_L g1432 ( 
.A(n_1359),
.B(n_1338),
.C(n_1318),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1399),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1399),
.Y(n_1434)
);

AOI31xp33_ASAP7_75t_L g1435 ( 
.A1(n_1389),
.A2(n_1387),
.A3(n_1385),
.B(n_1362),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1399),
.Y(n_1436)
);

AND2x2_ASAP7_75t_L g1437 ( 
.A(n_1362),
.B(n_1315),
.Y(n_1437)
);

HB1xp67_ASAP7_75t_L g1438 ( 
.A(n_1358),
.Y(n_1438)
);

OAI221xp5_ASAP7_75t_L g1439 ( 
.A1(n_1387),
.A2(n_1330),
.B1(n_1338),
.B2(n_1308),
.C(n_1314),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_L g1440 ( 
.A(n_1394),
.B(n_1245),
.Y(n_1440)
);

NAND2xp5_ASAP7_75t_L g1441 ( 
.A(n_1380),
.B(n_1335),
.Y(n_1441)
);

HB1xp67_ASAP7_75t_L g1442 ( 
.A(n_1358),
.Y(n_1442)
);

AND2x2_ASAP7_75t_L g1443 ( 
.A(n_1388),
.B(n_1335),
.Y(n_1443)
);

AND2x2_ASAP7_75t_L g1444 ( 
.A(n_1388),
.B(n_1334),
.Y(n_1444)
);

AND2x2_ASAP7_75t_L g1445 ( 
.A(n_1388),
.B(n_1334),
.Y(n_1445)
);

OAI21xp33_ASAP7_75t_L g1446 ( 
.A1(n_1389),
.A2(n_1328),
.B(n_1337),
.Y(n_1446)
);

AND2x4_ASAP7_75t_L g1447 ( 
.A(n_1415),
.B(n_1352),
.Y(n_1447)
);

NOR2xp33_ASAP7_75t_L g1448 ( 
.A(n_1374),
.B(n_1277),
.Y(n_1448)
);

HB1xp67_ASAP7_75t_L g1449 ( 
.A(n_1365),
.Y(n_1449)
);

NAND2xp5_ASAP7_75t_L g1450 ( 
.A(n_1398),
.B(n_1356),
.Y(n_1450)
);

OR2x2_ASAP7_75t_L g1451 ( 
.A(n_1386),
.B(n_1288),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1375),
.Y(n_1452)
);

AND2x2_ASAP7_75t_L g1453 ( 
.A(n_1379),
.B(n_1243),
.Y(n_1453)
);

INVx2_ASAP7_75t_SL g1454 ( 
.A(n_1403),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_L g1455 ( 
.A(n_1398),
.B(n_1297),
.Y(n_1455)
);

AND2x2_ASAP7_75t_L g1456 ( 
.A(n_1379),
.B(n_1243),
.Y(n_1456)
);

INVx1_ASAP7_75t_SL g1457 ( 
.A(n_1374),
.Y(n_1457)
);

AND2x2_ASAP7_75t_L g1458 ( 
.A(n_1379),
.B(n_1247),
.Y(n_1458)
);

OR2x2_ASAP7_75t_L g1459 ( 
.A(n_1365),
.B(n_1368),
.Y(n_1459)
);

INVx2_ASAP7_75t_SL g1460 ( 
.A(n_1417),
.Y(n_1460)
);

OR2x2_ASAP7_75t_L g1461 ( 
.A(n_1368),
.B(n_1356),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1395),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_SL g1463 ( 
.A(n_1385),
.B(n_1301),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1395),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1364),
.Y(n_1465)
);

OR2x2_ASAP7_75t_L g1466 ( 
.A(n_1368),
.B(n_1268),
.Y(n_1466)
);

NAND3xp33_ASAP7_75t_L g1467 ( 
.A(n_1381),
.B(n_1301),
.C(n_1340),
.Y(n_1467)
);

INVx2_ASAP7_75t_SL g1468 ( 
.A(n_1417),
.Y(n_1468)
);

AOI211xp5_ASAP7_75t_L g1469 ( 
.A1(n_1389),
.A2(n_1349),
.B(n_1272),
.C(n_1321),
.Y(n_1469)
);

AOI22xp33_ASAP7_75t_L g1470 ( 
.A1(n_1418),
.A2(n_1281),
.B1(n_1265),
.B2(n_1272),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1364),
.Y(n_1471)
);

NAND2xp5_ASAP7_75t_L g1472 ( 
.A(n_1404),
.B(n_1301),
.Y(n_1472)
);

OR2x2_ASAP7_75t_L g1473 ( 
.A(n_1459),
.B(n_1371),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1420),
.B(n_1369),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_L g1475 ( 
.A(n_1422),
.B(n_1369),
.Y(n_1475)
);

AOI22xp5_ASAP7_75t_L g1476 ( 
.A1(n_1446),
.A2(n_1416),
.B1(n_1418),
.B2(n_1405),
.Y(n_1476)
);

OAI22xp33_ASAP7_75t_L g1477 ( 
.A1(n_1435),
.A2(n_1405),
.B1(n_1381),
.B2(n_1383),
.Y(n_1477)
);

NAND2xp33_ASAP7_75t_SL g1478 ( 
.A(n_1425),
.B(n_1382),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_SL g1479 ( 
.A(n_1446),
.B(n_1382),
.Y(n_1479)
);

AND2x2_ASAP7_75t_L g1480 ( 
.A(n_1425),
.B(n_1367),
.Y(n_1480)
);

OAI22xp33_ASAP7_75t_L g1481 ( 
.A1(n_1421),
.A2(n_1383),
.B1(n_1381),
.B2(n_1416),
.Y(n_1481)
);

NAND4xp25_ASAP7_75t_L g1482 ( 
.A(n_1432),
.B(n_1413),
.C(n_1412),
.D(n_1370),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1454),
.B(n_1431),
.Y(n_1483)
);

AND2x2_ASAP7_75t_L g1484 ( 
.A(n_1443),
.B(n_1367),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_L g1485 ( 
.A(n_1440),
.B(n_1373),
.Y(n_1485)
);

OA21x2_ASAP7_75t_L g1486 ( 
.A1(n_1424),
.A2(n_1384),
.B(n_1383),
.Y(n_1486)
);

AND2x2_ASAP7_75t_L g1487 ( 
.A(n_1443),
.B(n_1367),
.Y(n_1487)
);

AOI221xp5_ASAP7_75t_L g1488 ( 
.A1(n_1432),
.A2(n_1400),
.B1(n_1384),
.B2(n_1406),
.C(n_1396),
.Y(n_1488)
);

NAND2xp5_ASAP7_75t_L g1489 ( 
.A(n_1460),
.B(n_1396),
.Y(n_1489)
);

NOR2xp67_ASAP7_75t_L g1490 ( 
.A(n_1467),
.B(n_1384),
.Y(n_1490)
);

NOR3xp33_ASAP7_75t_L g1491 ( 
.A(n_1439),
.B(n_1463),
.C(n_1455),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_L g1492 ( 
.A(n_1468),
.B(n_1438),
.Y(n_1492)
);

AND2x2_ASAP7_75t_L g1493 ( 
.A(n_1419),
.B(n_1378),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_L g1494 ( 
.A(n_1468),
.B(n_1442),
.Y(n_1494)
);

AND2x2_ASAP7_75t_L g1495 ( 
.A(n_1426),
.B(n_1378),
.Y(n_1495)
);

NAND2xp5_ASAP7_75t_L g1496 ( 
.A(n_1449),
.B(n_1396),
.Y(n_1496)
);

OAI21xp5_ASAP7_75t_SL g1497 ( 
.A1(n_1457),
.A2(n_1416),
.B(n_1370),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_SL g1498 ( 
.A(n_1469),
.B(n_1390),
.Y(n_1498)
);

AND2x4_ASAP7_75t_L g1499 ( 
.A(n_1453),
.B(n_1408),
.Y(n_1499)
);

NAND3xp33_ASAP7_75t_L g1500 ( 
.A(n_1424),
.B(n_1412),
.C(n_1409),
.Y(n_1500)
);

OAI22xp5_ASAP7_75t_L g1501 ( 
.A1(n_1469),
.A2(n_1413),
.B1(n_1401),
.B2(n_1390),
.Y(n_1501)
);

NOR3xp33_ASAP7_75t_L g1502 ( 
.A(n_1450),
.B(n_1377),
.C(n_1366),
.Y(n_1502)
);

AND2x2_ASAP7_75t_L g1503 ( 
.A(n_1437),
.B(n_1378),
.Y(n_1503)
);

NAND4xp25_ASAP7_75t_L g1504 ( 
.A(n_1441),
.B(n_1370),
.C(n_1377),
.D(n_1414),
.Y(n_1504)
);

AND2x2_ASAP7_75t_L g1505 ( 
.A(n_1444),
.B(n_1378),
.Y(n_1505)
);

NAND2xp5_ASAP7_75t_L g1506 ( 
.A(n_1459),
.B(n_1406),
.Y(n_1506)
);

NAND3xp33_ASAP7_75t_L g1507 ( 
.A(n_1429),
.B(n_1409),
.C(n_1414),
.Y(n_1507)
);

NAND3xp33_ASAP7_75t_L g1508 ( 
.A(n_1429),
.B(n_1414),
.C(n_1360),
.Y(n_1508)
);

NOR3xp33_ASAP7_75t_L g1509 ( 
.A(n_1472),
.B(n_1377),
.C(n_1366),
.Y(n_1509)
);

OAI22xp5_ASAP7_75t_L g1510 ( 
.A1(n_1451),
.A2(n_1390),
.B1(n_1363),
.B2(n_1372),
.Y(n_1510)
);

AOI22xp33_ASAP7_75t_L g1511 ( 
.A1(n_1470),
.A2(n_1410),
.B1(n_1411),
.B2(n_1391),
.Y(n_1511)
);

AND2x2_ASAP7_75t_L g1512 ( 
.A(n_1444),
.B(n_1378),
.Y(n_1512)
);

NAND2xp5_ASAP7_75t_L g1513 ( 
.A(n_1465),
.B(n_1376),
.Y(n_1513)
);

NAND3xp33_ASAP7_75t_L g1514 ( 
.A(n_1433),
.B(n_1360),
.C(n_1407),
.Y(n_1514)
);

AND2x2_ASAP7_75t_L g1515 ( 
.A(n_1445),
.B(n_1377),
.Y(n_1515)
);

AND2x2_ASAP7_75t_SL g1516 ( 
.A(n_1447),
.B(n_1393),
.Y(n_1516)
);

OAI221xp5_ASAP7_75t_L g1517 ( 
.A1(n_1451),
.A2(n_1400),
.B1(n_1410),
.B2(n_1397),
.C(n_1402),
.Y(n_1517)
);

BUFx3_ASAP7_75t_L g1518 ( 
.A(n_1516),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1473),
.Y(n_1519)
);

OR2x2_ASAP7_75t_L g1520 ( 
.A(n_1473),
.B(n_1496),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1514),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1480),
.B(n_1493),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1508),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_L g1524 ( 
.A(n_1488),
.B(n_1485),
.Y(n_1524)
);

HB1xp67_ASAP7_75t_L g1525 ( 
.A(n_1492),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1513),
.Y(n_1526)
);

NOR2xp67_ASAP7_75t_L g1527 ( 
.A(n_1504),
.B(n_1467),
.Y(n_1527)
);

AND2x2_ASAP7_75t_L g1528 ( 
.A(n_1480),
.B(n_1493),
.Y(n_1528)
);

AND2x4_ASAP7_75t_L g1529 ( 
.A(n_1490),
.B(n_1447),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1474),
.Y(n_1530)
);

AND2x4_ASAP7_75t_L g1531 ( 
.A(n_1490),
.B(n_1447),
.Y(n_1531)
);

AND2x2_ASAP7_75t_L g1532 ( 
.A(n_1495),
.B(n_1503),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1475),
.Y(n_1533)
);

AOI21xp33_ASAP7_75t_L g1534 ( 
.A1(n_1477),
.A2(n_1434),
.B(n_1433),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_L g1535 ( 
.A(n_1505),
.B(n_1471),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_L g1536 ( 
.A(n_1505),
.B(n_1471),
.Y(n_1536)
);

INVx2_ASAP7_75t_L g1537 ( 
.A(n_1486),
.Y(n_1537)
);

AND2x2_ASAP7_75t_L g1538 ( 
.A(n_1495),
.B(n_1456),
.Y(n_1538)
);

INVx1_ASAP7_75t_SL g1539 ( 
.A(n_1483),
.Y(n_1539)
);

OR2x2_ASAP7_75t_L g1540 ( 
.A(n_1506),
.B(n_1461),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1489),
.Y(n_1541)
);

HB1xp67_ASAP7_75t_L g1542 ( 
.A(n_1494),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_L g1543 ( 
.A(n_1512),
.B(n_1461),
.Y(n_1543)
);

INVx2_ASAP7_75t_L g1544 ( 
.A(n_1486),
.Y(n_1544)
);

NOR2x1_ASAP7_75t_L g1545 ( 
.A(n_1498),
.B(n_1427),
.Y(n_1545)
);

AND2x2_ASAP7_75t_L g1546 ( 
.A(n_1503),
.B(n_1484),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1507),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_SL g1548 ( 
.A(n_1516),
.B(n_1427),
.Y(n_1548)
);

INVx2_ASAP7_75t_L g1549 ( 
.A(n_1486),
.Y(n_1549)
);

OR2x6_ASAP7_75t_L g1550 ( 
.A(n_1498),
.B(n_1430),
.Y(n_1550)
);

INVx2_ASAP7_75t_L g1551 ( 
.A(n_1512),
.Y(n_1551)
);

AND2x4_ASAP7_75t_L g1552 ( 
.A(n_1499),
.B(n_1447),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1500),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1517),
.Y(n_1554)
);

INVx4_ASAP7_75t_SL g1555 ( 
.A(n_1499),
.Y(n_1555)
);

INVxp67_ASAP7_75t_SL g1556 ( 
.A(n_1527),
.Y(n_1556)
);

OR2x2_ASAP7_75t_L g1557 ( 
.A(n_1554),
.B(n_1482),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1555),
.B(n_1484),
.Y(n_1558)
);

OR2x2_ASAP7_75t_L g1559 ( 
.A(n_1554),
.B(n_1497),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_L g1560 ( 
.A(n_1553),
.B(n_1491),
.Y(n_1560)
);

NAND2xp5_ASAP7_75t_L g1561 ( 
.A(n_1521),
.B(n_1462),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1553),
.B(n_1462),
.Y(n_1562)
);

OAI221xp5_ASAP7_75t_SL g1563 ( 
.A1(n_1524),
.A2(n_1476),
.B1(n_1481),
.B2(n_1511),
.C(n_1502),
.Y(n_1563)
);

OAI21xp5_ASAP7_75t_L g1564 ( 
.A1(n_1521),
.A2(n_1479),
.B(n_1501),
.Y(n_1564)
);

NAND2xp5_ASAP7_75t_L g1565 ( 
.A(n_1523),
.B(n_1547),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1519),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1555),
.B(n_1487),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1519),
.Y(n_1568)
);

AND2x2_ASAP7_75t_L g1569 ( 
.A(n_1555),
.B(n_1487),
.Y(n_1569)
);

OR2x2_ASAP7_75t_L g1570 ( 
.A(n_1523),
.B(n_1466),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1555),
.B(n_1499),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1526),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1526),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_L g1574 ( 
.A(n_1547),
.B(n_1464),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1520),
.Y(n_1575)
);

INVx2_ASAP7_75t_L g1576 ( 
.A(n_1544),
.Y(n_1576)
);

NAND2xp5_ASAP7_75t_L g1577 ( 
.A(n_1539),
.B(n_1464),
.Y(n_1577)
);

BUFx2_ASAP7_75t_L g1578 ( 
.A(n_1545),
.Y(n_1578)
);

AND2x4_ASAP7_75t_L g1579 ( 
.A(n_1555),
.B(n_1479),
.Y(n_1579)
);

AND2x2_ASAP7_75t_L g1580 ( 
.A(n_1522),
.B(n_1528),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1520),
.Y(n_1581)
);

INVx2_ASAP7_75t_SL g1582 ( 
.A(n_1518),
.Y(n_1582)
);

INVxp67_ASAP7_75t_SL g1583 ( 
.A(n_1527),
.Y(n_1583)
);

OR2x2_ASAP7_75t_L g1584 ( 
.A(n_1535),
.B(n_1478),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_L g1585 ( 
.A(n_1530),
.B(n_1452),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_L g1586 ( 
.A(n_1525),
.B(n_1515),
.Y(n_1586)
);

INVxp67_ASAP7_75t_SL g1587 ( 
.A(n_1545),
.Y(n_1587)
);

AND2x2_ASAP7_75t_L g1588 ( 
.A(n_1522),
.B(n_1515),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1530),
.Y(n_1589)
);

AND2x2_ASAP7_75t_L g1590 ( 
.A(n_1528),
.B(n_1458),
.Y(n_1590)
);

AND2x4_ASAP7_75t_L g1591 ( 
.A(n_1518),
.B(n_1550),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1533),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1533),
.Y(n_1593)
);

OAI32xp33_ASAP7_75t_L g1594 ( 
.A1(n_1518),
.A2(n_1478),
.A3(n_1428),
.B1(n_1509),
.B2(n_1510),
.Y(n_1594)
);

AND2x2_ASAP7_75t_L g1595 ( 
.A(n_1546),
.B(n_1458),
.Y(n_1595)
);

NAND2x1_ASAP7_75t_L g1596 ( 
.A(n_1578),
.B(n_1552),
.Y(n_1596)
);

INVx2_ASAP7_75t_L g1597 ( 
.A(n_1576),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1566),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1566),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1577),
.Y(n_1600)
);

XNOR2xp5_ASAP7_75t_L g1601 ( 
.A(n_1560),
.B(n_1349),
.Y(n_1601)
);

OR2x2_ASAP7_75t_L g1602 ( 
.A(n_1565),
.B(n_1540),
.Y(n_1602)
);

INVx2_ASAP7_75t_L g1603 ( 
.A(n_1576),
.Y(n_1603)
);

OAI22xp5_ASAP7_75t_L g1604 ( 
.A1(n_1556),
.A2(n_1550),
.B1(n_1548),
.B2(n_1529),
.Y(n_1604)
);

INVx2_ASAP7_75t_SL g1605 ( 
.A(n_1579),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_L g1606 ( 
.A(n_1583),
.B(n_1557),
.Y(n_1606)
);

OR2x2_ASAP7_75t_L g1607 ( 
.A(n_1557),
.B(n_1540),
.Y(n_1607)
);

NAND2x1p5_ASAP7_75t_L g1608 ( 
.A(n_1578),
.B(n_1430),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1561),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_L g1610 ( 
.A(n_1562),
.B(n_1561),
.Y(n_1610)
);

AOI22xp33_ASAP7_75t_L g1611 ( 
.A1(n_1559),
.A2(n_1534),
.B1(n_1423),
.B2(n_1544),
.Y(n_1611)
);

AOI21xp5_ASAP7_75t_L g1612 ( 
.A1(n_1563),
.A2(n_1550),
.B(n_1531),
.Y(n_1612)
);

NOR2xp33_ASAP7_75t_L g1613 ( 
.A(n_1559),
.B(n_1428),
.Y(n_1613)
);

AND2x2_ASAP7_75t_L g1614 ( 
.A(n_1571),
.B(n_1580),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1574),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1575),
.Y(n_1616)
);

INVx2_ASAP7_75t_L g1617 ( 
.A(n_1576),
.Y(n_1617)
);

HB1xp67_ASAP7_75t_L g1618 ( 
.A(n_1570),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1571),
.B(n_1580),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1575),
.Y(n_1620)
);

AND2x2_ASAP7_75t_L g1621 ( 
.A(n_1579),
.B(n_1552),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_L g1622 ( 
.A(n_1581),
.B(n_1542),
.Y(n_1622)
);

NOR2xp33_ASAP7_75t_L g1623 ( 
.A(n_1587),
.B(n_1258),
.Y(n_1623)
);

INVx2_ASAP7_75t_SL g1624 ( 
.A(n_1579),
.Y(n_1624)
);

OAI22xp5_ASAP7_75t_L g1625 ( 
.A1(n_1564),
.A2(n_1550),
.B1(n_1531),
.B2(n_1529),
.Y(n_1625)
);

AOI21xp33_ASAP7_75t_L g1626 ( 
.A1(n_1582),
.A2(n_1550),
.B(n_1436),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_L g1627 ( 
.A(n_1581),
.B(n_1541),
.Y(n_1627)
);

INVx3_ASAP7_75t_L g1628 ( 
.A(n_1579),
.Y(n_1628)
);

OR2x2_ASAP7_75t_L g1629 ( 
.A(n_1568),
.B(n_1570),
.Y(n_1629)
);

INVx2_ASAP7_75t_L g1630 ( 
.A(n_1589),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1558),
.B(n_1552),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1568),
.Y(n_1632)
);

OR2x2_ASAP7_75t_L g1633 ( 
.A(n_1589),
.B(n_1536),
.Y(n_1633)
);

AND2x4_ASAP7_75t_L g1634 ( 
.A(n_1591),
.B(n_1552),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1572),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_L g1636 ( 
.A(n_1592),
.B(n_1541),
.Y(n_1636)
);

INVx2_ASAP7_75t_L g1637 ( 
.A(n_1592),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1572),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1614),
.B(n_1582),
.Y(n_1639)
);

HB1xp67_ASAP7_75t_L g1640 ( 
.A(n_1630),
.Y(n_1640)
);

AND2x2_ASAP7_75t_L g1641 ( 
.A(n_1614),
.B(n_1558),
.Y(n_1641)
);

AND2x2_ASAP7_75t_L g1642 ( 
.A(n_1619),
.B(n_1567),
.Y(n_1642)
);

AND2x4_ASAP7_75t_SL g1643 ( 
.A(n_1634),
.B(n_1591),
.Y(n_1643)
);

AND2x2_ASAP7_75t_L g1644 ( 
.A(n_1619),
.B(n_1567),
.Y(n_1644)
);

AND2x2_ASAP7_75t_L g1645 ( 
.A(n_1621),
.B(n_1569),
.Y(n_1645)
);

OAI22xp5_ASAP7_75t_L g1646 ( 
.A1(n_1606),
.A2(n_1564),
.B1(n_1584),
.B2(n_1591),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1598),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1598),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_L g1649 ( 
.A(n_1618),
.B(n_1573),
.Y(n_1649)
);

HB1xp67_ASAP7_75t_L g1650 ( 
.A(n_1630),
.Y(n_1650)
);

AND2x2_ASAP7_75t_L g1651 ( 
.A(n_1621),
.B(n_1569),
.Y(n_1651)
);

INVx1_ASAP7_75t_SL g1652 ( 
.A(n_1601),
.Y(n_1652)
);

AND2x2_ASAP7_75t_L g1653 ( 
.A(n_1631),
.B(n_1588),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1599),
.Y(n_1654)
);

NAND2xp5_ASAP7_75t_L g1655 ( 
.A(n_1615),
.B(n_1573),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1631),
.B(n_1588),
.Y(n_1656)
);

INVx2_ASAP7_75t_L g1657 ( 
.A(n_1597),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1628),
.B(n_1590),
.Y(n_1658)
);

INVx2_ASAP7_75t_L g1659 ( 
.A(n_1597),
.Y(n_1659)
);

INVx2_ASAP7_75t_L g1660 ( 
.A(n_1603),
.Y(n_1660)
);

AND2x2_ASAP7_75t_L g1661 ( 
.A(n_1628),
.B(n_1590),
.Y(n_1661)
);

INVx2_ASAP7_75t_L g1662 ( 
.A(n_1603),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_L g1663 ( 
.A(n_1609),
.B(n_1593),
.Y(n_1663)
);

HB1xp67_ASAP7_75t_L g1664 ( 
.A(n_1637),
.Y(n_1664)
);

AND2x2_ASAP7_75t_L g1665 ( 
.A(n_1628),
.B(n_1595),
.Y(n_1665)
);

OAI21x1_ASAP7_75t_L g1666 ( 
.A1(n_1608),
.A2(n_1537),
.B(n_1544),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_L g1667 ( 
.A(n_1602),
.B(n_1593),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1599),
.Y(n_1668)
);

OAI21xp33_ASAP7_75t_L g1669 ( 
.A1(n_1607),
.A2(n_1594),
.B(n_1584),
.Y(n_1669)
);

OR2x2_ASAP7_75t_L g1670 ( 
.A(n_1610),
.B(n_1585),
.Y(n_1670)
);

CKINVDCx5p33_ASAP7_75t_R g1671 ( 
.A(n_1601),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1602),
.B(n_1585),
.Y(n_1672)
);

AND2x2_ASAP7_75t_L g1673 ( 
.A(n_1634),
.B(n_1595),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1638),
.Y(n_1674)
);

OAI31xp33_ASAP7_75t_L g1675 ( 
.A1(n_1646),
.A2(n_1612),
.A3(n_1611),
.B(n_1625),
.Y(n_1675)
);

OAI22xp33_ASAP7_75t_L g1676 ( 
.A1(n_1646),
.A2(n_1607),
.B1(n_1605),
.B2(n_1624),
.Y(n_1676)
);

NAND3xp33_ASAP7_75t_SL g1677 ( 
.A(n_1652),
.B(n_1608),
.C(n_1613),
.Y(n_1677)
);

OR2x2_ASAP7_75t_L g1678 ( 
.A(n_1667),
.B(n_1622),
.Y(n_1678)
);

OAI21xp5_ASAP7_75t_SL g1679 ( 
.A1(n_1669),
.A2(n_1624),
.B(n_1605),
.Y(n_1679)
);

AOI222xp33_ASAP7_75t_L g1680 ( 
.A1(n_1669),
.A2(n_1549),
.B1(n_1537),
.B2(n_1623),
.C1(n_1600),
.C2(n_1617),
.Y(n_1680)
);

INVxp67_ASAP7_75t_L g1681 ( 
.A(n_1652),
.Y(n_1681)
);

AO221x1_ASAP7_75t_L g1682 ( 
.A1(n_1643),
.A2(n_1604),
.B1(n_1620),
.B2(n_1616),
.C(n_1638),
.Y(n_1682)
);

NAND2x1_ASAP7_75t_L g1683 ( 
.A(n_1641),
.B(n_1634),
.Y(n_1683)
);

AOI211xp5_ASAP7_75t_L g1684 ( 
.A1(n_1640),
.A2(n_1594),
.B(n_1626),
.C(n_1629),
.Y(n_1684)
);

AOI22xp33_ASAP7_75t_SL g1685 ( 
.A1(n_1640),
.A2(n_1591),
.B1(n_1617),
.B2(n_1637),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1647),
.Y(n_1686)
);

AOI22xp5_ASAP7_75t_L g1687 ( 
.A1(n_1671),
.A2(n_1627),
.B1(n_1531),
.B2(n_1529),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1647),
.Y(n_1688)
);

NOR2xp33_ASAP7_75t_L g1689 ( 
.A(n_1643),
.B(n_1263),
.Y(n_1689)
);

AOI211xp5_ASAP7_75t_L g1690 ( 
.A1(n_1650),
.A2(n_1629),
.B(n_1635),
.C(n_1632),
.Y(n_1690)
);

OAI22xp5_ASAP7_75t_L g1691 ( 
.A1(n_1643),
.A2(n_1596),
.B1(n_1529),
.B2(n_1531),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1648),
.Y(n_1692)
);

AND2x2_ASAP7_75t_L g1693 ( 
.A(n_1673),
.B(n_1596),
.Y(n_1693)
);

AND2x2_ASAP7_75t_L g1694 ( 
.A(n_1673),
.B(n_1639),
.Y(n_1694)
);

NAND3xp33_ASAP7_75t_SL g1695 ( 
.A(n_1639),
.B(n_1608),
.C(n_1633),
.Y(n_1695)
);

NAND2xp5_ASAP7_75t_L g1696 ( 
.A(n_1639),
.B(n_1636),
.Y(n_1696)
);

AO22x1_ASAP7_75t_L g1697 ( 
.A1(n_1641),
.A2(n_1346),
.B1(n_1448),
.B2(n_1532),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1648),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_L g1699 ( 
.A(n_1658),
.B(n_1661),
.Y(n_1699)
);

AOI22xp33_ASAP7_75t_L g1700 ( 
.A1(n_1657),
.A2(n_1549),
.B1(n_1423),
.B2(n_1633),
.Y(n_1700)
);

AOI221x1_ASAP7_75t_SL g1701 ( 
.A1(n_1690),
.A2(n_1649),
.B1(n_1654),
.B2(n_1674),
.C(n_1668),
.Y(n_1701)
);

HB1xp67_ASAP7_75t_L g1702 ( 
.A(n_1681),
.Y(n_1702)
);

OAI21xp33_ASAP7_75t_L g1703 ( 
.A1(n_1679),
.A2(n_1643),
.B(n_1667),
.Y(n_1703)
);

NAND2xp5_ASAP7_75t_SL g1704 ( 
.A(n_1685),
.B(n_1650),
.Y(n_1704)
);

INVxp67_ASAP7_75t_L g1705 ( 
.A(n_1677),
.Y(n_1705)
);

AND2x2_ASAP7_75t_L g1706 ( 
.A(n_1694),
.B(n_1673),
.Y(n_1706)
);

INVx1_ASAP7_75t_SL g1707 ( 
.A(n_1699),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_L g1708 ( 
.A(n_1696),
.B(n_1658),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1686),
.Y(n_1709)
);

INVx8_ASAP7_75t_L g1710 ( 
.A(n_1693),
.Y(n_1710)
);

INVx3_ASAP7_75t_L g1711 ( 
.A(n_1683),
.Y(n_1711)
);

NAND2xp5_ASAP7_75t_L g1712 ( 
.A(n_1678),
.B(n_1658),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1688),
.Y(n_1713)
);

INVx2_ASAP7_75t_L g1714 ( 
.A(n_1692),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_1685),
.B(n_1661),
.Y(n_1715)
);

AOI22xp5_ASAP7_75t_L g1716 ( 
.A1(n_1680),
.A2(n_1660),
.B1(n_1657),
.B2(n_1659),
.Y(n_1716)
);

OAI22xp5_ASAP7_75t_L g1717 ( 
.A1(n_1684),
.A2(n_1644),
.B1(n_1641),
.B2(n_1642),
.Y(n_1717)
);

OR2x2_ASAP7_75t_L g1718 ( 
.A(n_1695),
.B(n_1672),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_L g1719 ( 
.A(n_1676),
.B(n_1661),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1698),
.Y(n_1720)
);

NAND3xp33_ASAP7_75t_L g1721 ( 
.A(n_1705),
.B(n_1675),
.C(n_1664),
.Y(n_1721)
);

AOI322xp5_ASAP7_75t_L g1722 ( 
.A1(n_1704),
.A2(n_1677),
.A3(n_1695),
.B1(n_1700),
.B2(n_1664),
.C1(n_1660),
.C2(n_1659),
.Y(n_1722)
);

AOI21xp5_ASAP7_75t_L g1723 ( 
.A1(n_1704),
.A2(n_1682),
.B(n_1689),
.Y(n_1723)
);

AOI221xp5_ASAP7_75t_L g1724 ( 
.A1(n_1701),
.A2(n_1668),
.B1(n_1674),
.B2(n_1654),
.C(n_1662),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_L g1725 ( 
.A(n_1702),
.B(n_1665),
.Y(n_1725)
);

NOR3xp33_ASAP7_75t_L g1726 ( 
.A(n_1705),
.B(n_1697),
.C(n_1691),
.Y(n_1726)
);

AOI221xp5_ASAP7_75t_L g1727 ( 
.A1(n_1717),
.A2(n_1662),
.B1(n_1657),
.B2(n_1659),
.C(n_1660),
.Y(n_1727)
);

AOI221xp5_ASAP7_75t_L g1728 ( 
.A1(n_1702),
.A2(n_1662),
.B1(n_1657),
.B2(n_1659),
.C(n_1660),
.Y(n_1728)
);

AOI221xp5_ASAP7_75t_L g1729 ( 
.A1(n_1715),
.A2(n_1662),
.B1(n_1649),
.B2(n_1663),
.C(n_1655),
.Y(n_1729)
);

AOI21xp5_ASAP7_75t_L g1730 ( 
.A1(n_1718),
.A2(n_1663),
.B(n_1655),
.Y(n_1730)
);

BUFx4f_ASAP7_75t_SL g1731 ( 
.A(n_1707),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1725),
.Y(n_1732)
);

NOR4xp25_ASAP7_75t_L g1733 ( 
.A(n_1721),
.B(n_1720),
.C(n_1713),
.D(n_1709),
.Y(n_1733)
);

NOR2xp33_ASAP7_75t_L g1734 ( 
.A(n_1731),
.B(n_1710),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1728),
.Y(n_1735)
);

NOR3xp33_ASAP7_75t_L g1736 ( 
.A(n_1723),
.B(n_1703),
.C(n_1719),
.Y(n_1736)
);

XNOR2x2_ASAP7_75t_L g1737 ( 
.A(n_1730),
.B(n_1716),
.Y(n_1737)
);

NOR2xp67_ASAP7_75t_L g1738 ( 
.A(n_1726),
.B(n_1711),
.Y(n_1738)
);

AOI21xp5_ASAP7_75t_L g1739 ( 
.A1(n_1724),
.A2(n_1710),
.B(n_1712),
.Y(n_1739)
);

NOR3xp33_ASAP7_75t_L g1740 ( 
.A(n_1727),
.B(n_1729),
.C(n_1714),
.Y(n_1740)
);

NAND2xp5_ASAP7_75t_SL g1741 ( 
.A(n_1738),
.B(n_1722),
.Y(n_1741)
);

OAI21xp33_ASAP7_75t_SL g1742 ( 
.A1(n_1733),
.A2(n_1711),
.B(n_1706),
.Y(n_1742)
);

NAND4xp25_ASAP7_75t_L g1743 ( 
.A(n_1734),
.B(n_1708),
.C(n_1687),
.D(n_1710),
.Y(n_1743)
);

AOI221xp5_ASAP7_75t_L g1744 ( 
.A1(n_1735),
.A2(n_1672),
.B1(n_1665),
.B2(n_1670),
.C(n_1549),
.Y(n_1744)
);

OAI211xp5_ASAP7_75t_L g1745 ( 
.A1(n_1736),
.A2(n_1642),
.B(n_1644),
.C(n_1665),
.Y(n_1745)
);

INVxp67_ASAP7_75t_SL g1746 ( 
.A(n_1741),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1745),
.Y(n_1747)
);

AOI22xp5_ASAP7_75t_L g1748 ( 
.A1(n_1744),
.A2(n_1740),
.B1(n_1742),
.B2(n_1732),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1743),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1745),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1745),
.Y(n_1751)
);

NOR2x1_ASAP7_75t_L g1752 ( 
.A(n_1749),
.B(n_1739),
.Y(n_1752)
);

AOI222xp33_ASAP7_75t_L g1753 ( 
.A1(n_1746),
.A2(n_1737),
.B1(n_1666),
.B2(n_1642),
.C1(n_1644),
.C2(n_1651),
.Y(n_1753)
);

AOI22xp5_ASAP7_75t_L g1754 ( 
.A1(n_1746),
.A2(n_1645),
.B1(n_1651),
.B2(n_1656),
.Y(n_1754)
);

NAND2x1_ASAP7_75t_L g1755 ( 
.A(n_1748),
.B(n_1645),
.Y(n_1755)
);

INVxp67_ASAP7_75t_SL g1756 ( 
.A(n_1747),
.Y(n_1756)
);

OA22x2_ASAP7_75t_L g1757 ( 
.A1(n_1754),
.A2(n_1751),
.B1(n_1750),
.B2(n_1645),
.Y(n_1757)
);

INVx3_ASAP7_75t_L g1758 ( 
.A(n_1755),
.Y(n_1758)
);

XNOR2x1_ASAP7_75t_L g1759 ( 
.A(n_1752),
.B(n_1346),
.Y(n_1759)
);

HB1xp67_ASAP7_75t_L g1760 ( 
.A(n_1759),
.Y(n_1760)
);

NAND3xp33_ASAP7_75t_SL g1761 ( 
.A(n_1760),
.B(n_1753),
.C(n_1756),
.Y(n_1761)
);

AO21x1_ASAP7_75t_L g1762 ( 
.A1(n_1761),
.A2(n_1757),
.B(n_1758),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1761),
.Y(n_1763)
);

OAI22xp33_ASAP7_75t_SL g1764 ( 
.A1(n_1763),
.A2(n_1346),
.B1(n_1670),
.B2(n_1312),
.Y(n_1764)
);

O2A1O1Ixp33_ASAP7_75t_L g1765 ( 
.A1(n_1762),
.A2(n_1670),
.B(n_1651),
.C(n_1656),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1765),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1764),
.Y(n_1767)
);

AOI221xp5_ASAP7_75t_L g1768 ( 
.A1(n_1766),
.A2(n_1767),
.B1(n_1656),
.B2(n_1653),
.C(n_1312),
.Y(n_1768)
);

AOI22xp5_ASAP7_75t_L g1769 ( 
.A1(n_1768),
.A2(n_1653),
.B1(n_1666),
.B2(n_1532),
.Y(n_1769)
);

AOI221xp5_ASAP7_75t_L g1770 ( 
.A1(n_1769),
.A2(n_1653),
.B1(n_1666),
.B2(n_1551),
.C(n_1586),
.Y(n_1770)
);

AOI211xp5_ASAP7_75t_L g1771 ( 
.A1(n_1770),
.A2(n_1546),
.B(n_1538),
.C(n_1543),
.Y(n_1771)
);


endmodule