module fake_jpeg_28344_n_323 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_323);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_323;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx4f_ASAP7_75t_SL g24 ( 
.A(n_1),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

CKINVDCx14_ASAP7_75t_R g29 ( 
.A(n_14),
.Y(n_29)
);

INVx6_ASAP7_75t_SL g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx10_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_9),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_16),
.Y(n_34)
);

CKINVDCx16_ASAP7_75t_R g35 ( 
.A(n_24),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_35),
.B(n_37),
.Y(n_53)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_17),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_38),
.B(n_39),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_29),
.B(n_8),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

INVx1_ASAP7_75t_SL g61 ( 
.A(n_44),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_36),
.A2(n_19),
.B1(n_28),
.B2(n_17),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_46),
.A2(n_49),
.B1(n_69),
.B2(n_43),
.Y(n_93)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g48 ( 
.A(n_35),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_48),
.B(n_35),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_36),
.A2(n_19),
.B1(n_28),
.B2(n_34),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_36),
.A2(n_28),
.B1(n_29),
.B2(n_23),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_50),
.A2(n_59),
.B1(n_64),
.B2(n_67),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_18),
.Y(n_52)
);

OR2x2_ASAP7_75t_L g87 ( 
.A(n_52),
.B(n_54),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_39),
.B(n_33),
.Y(n_54)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_55),
.Y(n_86)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_56),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_36),
.A2(n_30),
.B1(n_26),
.B2(n_25),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_39),
.B(n_31),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_60),
.B(n_62),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_37),
.B(n_31),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_37),
.A2(n_30),
.B1(n_20),
.B2(n_32),
.Y(n_64)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_66),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_37),
.A2(n_30),
.B1(n_20),
.B2(n_32),
.Y(n_67)
);

OA22x2_ASAP7_75t_L g68 ( 
.A1(n_43),
.A2(n_24),
.B1(n_31),
.B2(n_21),
.Y(n_68)
);

AO22x1_ASAP7_75t_L g79 ( 
.A1(n_68),
.A2(n_41),
.B1(n_44),
.B2(n_43),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_41),
.A2(n_34),
.B1(n_22),
.B2(n_25),
.Y(n_69)
);

INVx11_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_71),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_62),
.A2(n_44),
.B1(n_41),
.B2(n_43),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_72),
.A2(n_93),
.B1(n_38),
.B2(n_65),
.Y(n_113)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_53),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_73),
.B(n_74),
.Y(n_101)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_53),
.Y(n_74)
);

INVx11_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_76),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_77),
.Y(n_114)
);

INVx11_ASAP7_75t_L g78 ( 
.A(n_56),
.Y(n_78)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_78),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_79),
.Y(n_104)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_64),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_80),
.B(n_83),
.Y(n_107)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_67),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_58),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_84),
.B(n_51),
.Y(n_109)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_58),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_85),
.B(n_90),
.Y(n_108)
);

OR2x4_ASAP7_75t_L g88 ( 
.A(n_52),
.B(n_31),
.Y(n_88)
);

FAx1_ASAP7_75t_SL g116 ( 
.A(n_88),
.B(n_94),
.CI(n_68),
.CON(n_116),
.SN(n_116)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_52),
.B(n_41),
.C(n_38),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_89),
.B(n_38),
.C(n_42),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_66),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_56),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_91),
.Y(n_97)
);

INVx6_ASAP7_75t_SL g92 ( 
.A(n_48),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_92),
.Y(n_118)
);

AOI32xp33_ASAP7_75t_L g94 ( 
.A1(n_57),
.A2(n_44),
.A3(n_42),
.B1(n_22),
.B2(n_31),
.Y(n_94)
);

INVx11_ASAP7_75t_L g95 ( 
.A(n_55),
.Y(n_95)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_95),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g98 ( 
.A(n_81),
.B(n_60),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_98),
.B(n_117),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_81),
.B(n_57),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_99),
.B(n_102),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_73),
.B(n_54),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_74),
.B(n_54),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_106),
.B(n_110),
.Y(n_134)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_109),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_87),
.B(n_50),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_72),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_111),
.B(n_115),
.Y(n_131)
);

AO22x1_ASAP7_75t_SL g112 ( 
.A1(n_88),
.A2(n_45),
.B1(n_68),
.B2(n_59),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_112),
.A2(n_45),
.B1(n_61),
.B2(n_82),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_113),
.A2(n_45),
.B1(n_65),
.B2(n_68),
.Y(n_130)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_79),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_116),
.B(n_42),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_SL g119 ( 
.A(n_89),
.B(n_68),
.Y(n_119)
);

AOI32xp33_ASAP7_75t_L g153 ( 
.A1(n_119),
.A2(n_33),
.A3(n_42),
.B1(n_24),
.B2(n_21),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_87),
.B(n_63),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_120),
.B(n_124),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_80),
.B(n_23),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_121),
.B(n_122),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_83),
.B(n_61),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_96),
.B(n_63),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_110),
.A2(n_94),
.B(n_96),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_127),
.A2(n_136),
.B(n_141),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_111),
.A2(n_79),
.B1(n_51),
.B2(n_92),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_129),
.A2(n_140),
.B1(n_118),
.B2(n_71),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_130),
.A2(n_139),
.B1(n_148),
.B2(n_103),
.Y(n_173)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_109),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_133),
.B(n_146),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_101),
.B(n_84),
.Y(n_135)
);

CKINVDCx14_ASAP7_75t_R g161 ( 
.A(n_135),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_101),
.B(n_85),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_137),
.B(n_142),
.Y(n_162)
);

BUFx3_ASAP7_75t_L g138 ( 
.A(n_123),
.Y(n_138)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_138),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_107),
.A2(n_82),
.B1(n_75),
.B2(n_70),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_122),
.A2(n_61),
.B(n_1),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_108),
.Y(n_142)
);

OA21x2_ASAP7_75t_L g144 ( 
.A1(n_124),
.A2(n_24),
.B(n_21),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_144),
.A2(n_114),
.B(n_106),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_99),
.B(n_26),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_145),
.B(n_147),
.Y(n_180)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_107),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_113),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_104),
.A2(n_95),
.B1(n_70),
.B2(n_75),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_121),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_149),
.B(n_128),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_97),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_150),
.Y(n_164)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_100),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_151),
.B(n_152),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_120),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_153),
.B(n_117),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_97),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_154),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_125),
.B(n_98),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_155),
.B(n_165),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_150),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_156),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_147),
.A2(n_104),
.B1(n_115),
.B2(n_102),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_157),
.A2(n_173),
.B1(n_176),
.B2(n_182),
.Y(n_191)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_131),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_158),
.B(n_160),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_154),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_159),
.Y(n_212)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_140),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_163),
.A2(n_169),
.B1(n_133),
.B2(n_132),
.Y(n_189)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_139),
.B(n_148),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_167),
.A2(n_171),
.B(n_183),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_127),
.A2(n_112),
.B1(n_116),
.B2(n_119),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_174),
.B(n_175),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_141),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_146),
.A2(n_112),
.B1(n_116),
.B2(n_105),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_129),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_177),
.B(n_178),
.Y(n_187)
);

INVxp33_ASAP7_75t_L g178 ( 
.A(n_128),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_136),
.A2(n_152),
.B1(n_149),
.B2(n_142),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_179),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_136),
.Y(n_181)
);

INVx1_ASAP7_75t_SL g194 ( 
.A(n_181),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_132),
.A2(n_112),
.B1(n_103),
.B2(n_105),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_143),
.A2(n_123),
.B(n_33),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_143),
.B(n_90),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_185),
.Y(n_186)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_184),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_188),
.B(n_192),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_189),
.A2(n_193),
.B1(n_197),
.B2(n_201),
.Y(n_213)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_172),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_167),
.A2(n_144),
.B1(n_125),
.B2(n_134),
.Y(n_193)
);

OAI21xp33_ASAP7_75t_SL g195 ( 
.A1(n_158),
.A2(n_134),
.B(n_144),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_195),
.A2(n_204),
.B(n_210),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_155),
.B(n_126),
.C(n_100),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_196),
.B(n_208),
.C(n_211),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_167),
.A2(n_177),
.B1(n_169),
.B2(n_160),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_172),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_198),
.B(n_27),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_163),
.A2(n_180),
.B1(n_181),
.B2(n_173),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_182),
.A2(n_126),
.B1(n_151),
.B2(n_78),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_202),
.A2(n_209),
.B1(n_166),
.B2(n_91),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_168),
.A2(n_138),
.B(n_1),
.Y(n_204)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_162),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_206),
.B(n_188),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_165),
.B(n_42),
.C(n_91),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_175),
.A2(n_76),
.B1(n_65),
.B2(n_86),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_168),
.A2(n_0),
.B(n_1),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_179),
.B(n_185),
.C(n_183),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_191),
.A2(n_170),
.B1(n_164),
.B2(n_161),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_214),
.A2(n_218),
.B1(n_226),
.B2(n_236),
.Y(n_245)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_200),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_216),
.B(n_217),
.Y(n_240)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_200),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_205),
.A2(n_170),
.B1(n_164),
.B2(n_171),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_203),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_219),
.B(n_221),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_SL g220 ( 
.A(n_207),
.B(n_174),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_220),
.B(n_222),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_212),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_SL g222 ( 
.A(n_207),
.B(n_33),
.Y(n_222)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_224),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_196),
.B(n_42),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_225),
.B(n_229),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_205),
.A2(n_166),
.B1(n_86),
.B2(n_26),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_187),
.B(n_86),
.Y(n_227)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_227),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_SL g229 ( 
.A(n_211),
.B(n_33),
.Y(n_229)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_190),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_230),
.B(n_231),
.Y(n_246)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_209),
.Y(n_231)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_232),
.Y(n_253)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_201),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_233),
.B(n_218),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_198),
.B(n_42),
.Y(n_234)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_234),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_SL g235 ( 
.A(n_189),
.B(n_193),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_235),
.B(n_27),
.C(n_10),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_186),
.A2(n_197),
.B1(n_194),
.B2(n_199),
.Y(n_236)
);

INVx1_ASAP7_75t_SL g237 ( 
.A(n_194),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_237),
.B(n_227),
.Y(n_239)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_238),
.Y(n_255)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_239),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_228),
.A2(n_199),
.B(n_204),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_241),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_238),
.B(n_186),
.Y(n_243)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_243),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_223),
.B(n_208),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_247),
.B(n_258),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_213),
.A2(n_210),
.B1(n_27),
.B2(n_0),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_250),
.B(n_226),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_251),
.B(n_228),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_214),
.B(n_0),
.Y(n_256)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_256),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_236),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_257)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_257),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_215),
.B(n_10),
.C(n_4),
.Y(n_258)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_259),
.Y(n_275)
);

BUFx12_ASAP7_75t_L g262 ( 
.A(n_242),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_262),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_258),
.B(n_225),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_263),
.B(n_270),
.Y(n_279)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_265),
.Y(n_284)
);

OAI31xp33_ASAP7_75t_L g266 ( 
.A1(n_256),
.A2(n_241),
.A3(n_243),
.B(n_257),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_266),
.A2(n_267),
.B1(n_272),
.B2(n_264),
.Y(n_276)
);

A2O1A1O1Ixp25_ASAP7_75t_L g269 ( 
.A1(n_244),
.A2(n_220),
.B(n_235),
.C(n_215),
.D(n_229),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_269),
.B(n_248),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_246),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_248),
.B(n_222),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_273),
.B(n_274),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_253),
.B(n_237),
.Y(n_274)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_276),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_275),
.B(n_260),
.C(n_254),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_277),
.B(n_282),
.C(n_11),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_268),
.A2(n_245),
.B1(n_249),
.B2(n_261),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_278),
.B(n_285),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_269),
.B(n_244),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_280),
.B(n_283),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_271),
.B(n_245),
.C(n_239),
.Y(n_282)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_262),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_270),
.B(n_255),
.Y(n_286)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_286),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_268),
.B(n_240),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_288),
.B(n_289),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_262),
.B(n_251),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_287),
.B(n_250),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_290),
.B(n_294),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_284),
.A2(n_252),
.B1(n_234),
.B2(n_6),
.Y(n_293)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_293),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_282),
.B(n_10),
.C(n_5),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_295),
.B(n_297),
.C(n_278),
.Y(n_304)
);

OR2x6_ASAP7_75t_SL g296 ( 
.A(n_277),
.B(n_12),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_296),
.A2(n_14),
.B(n_5),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_289),
.A2(n_12),
.B1(n_5),
.B2(n_6),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_296),
.A2(n_279),
.B(n_281),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g313 ( 
.A1(n_302),
.A2(n_308),
.B(n_13),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_304),
.B(n_305),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_294),
.B(n_298),
.C(n_295),
.Y(n_305)
);

OAI21xp33_ASAP7_75t_L g314 ( 
.A1(n_306),
.A2(n_13),
.B(n_15),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_299),
.B(n_280),
.C(n_283),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_307),
.B(n_309),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_300),
.B(n_7),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_292),
.B(n_7),
.C(n_9),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_301),
.A2(n_291),
.B(n_9),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g316 ( 
.A1(n_310),
.A2(n_314),
.B(n_15),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_303),
.B(n_291),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_312),
.A2(n_308),
.B(n_15),
.Y(n_318)
);

INVxp67_ASAP7_75t_L g317 ( 
.A(n_313),
.Y(n_317)
);

OAI21x1_ASAP7_75t_SL g319 ( 
.A1(n_316),
.A2(n_318),
.B(n_16),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_319),
.B(n_315),
.C(n_317),
.Y(n_320)
);

AOI211xp5_ASAP7_75t_SL g321 ( 
.A1(n_320),
.A2(n_311),
.B(n_16),
.C(n_2),
.Y(n_321)
);

BUFx24_ASAP7_75t_SL g322 ( 
.A(n_321),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_322),
.B(n_2),
.Y(n_323)
);


endmodule