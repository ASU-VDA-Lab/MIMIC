module fake_jpeg_18047_n_269 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_269);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_269;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_14),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx6f_ASAP7_75t_SL g27 ( 
.A(n_5),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

INVxp67_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_27),
.Y(n_32)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_33),
.B(n_35),
.Y(n_42)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_36),
.B(n_37),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_38),
.B(n_40),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_18),
.B(n_0),
.Y(n_40)
);

BUFx10_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_41),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_40),
.B(n_16),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_43),
.B(n_17),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g44 ( 
.A(n_33),
.Y(n_44)
);

OR2x2_ASAP7_75t_L g70 ( 
.A(n_44),
.B(n_45),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_35),
.Y(n_45)
);

AND2x2_ASAP7_75t_SL g46 ( 
.A(n_38),
.B(n_20),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_46),
.B(n_20),
.C(n_37),
.Y(n_67)
);

CKINVDCx14_ASAP7_75t_SL g48 ( 
.A(n_32),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_39),
.B(n_31),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_49),
.B(n_50),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_39),
.B(n_31),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_34),
.B(n_18),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_51),
.B(n_55),
.Y(n_82)
);

OAI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_34),
.A2(n_26),
.B1(n_24),
.B2(n_23),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_54),
.A2(n_23),
.B1(n_26),
.B2(n_28),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_32),
.B(n_20),
.Y(n_55)
);

HB1xp67_ASAP7_75t_L g57 ( 
.A(n_32),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_57),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_59),
.B(n_64),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_56),
.B(n_17),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_60),
.B(n_63),
.Y(n_102)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_61),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_46),
.B(n_39),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_43),
.B(n_24),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_66),
.B(n_72),
.Y(n_107)
);

FAx1_ASAP7_75t_SL g94 ( 
.A(n_67),
.B(n_57),
.CI(n_21),
.CON(n_94),
.SN(n_94)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_53),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_68),
.B(n_71),
.Y(n_93)
);

NAND2xp33_ASAP7_75t_SL g86 ( 
.A(n_69),
.B(n_47),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_56),
.B(n_30),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_53),
.Y(n_72)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_41),
.Y(n_73)
);

BUFx4f_ASAP7_75t_SL g108 ( 
.A(n_73),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_44),
.B(n_21),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_75),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_49),
.A2(n_37),
.B1(n_36),
.B2(n_29),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_76),
.A2(n_55),
.B1(n_47),
.B2(n_45),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_46),
.B(n_30),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_77),
.B(n_79),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_51),
.A2(n_28),
.B1(n_25),
.B2(n_22),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_78),
.A2(n_15),
.B1(n_42),
.B2(n_55),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_50),
.B(n_25),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_51),
.B(n_22),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_80),
.B(n_81),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_51),
.B(n_16),
.Y(n_81)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_55),
.Y(n_84)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_84),
.Y(n_96)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_83),
.Y(n_85)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_85),
.Y(n_114)
);

AO21x1_ASAP7_75t_L g119 ( 
.A1(n_86),
.A2(n_81),
.B(n_80),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_74),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_87),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_88),
.B(n_92),
.Y(n_118)
);

INVx1_ASAP7_75t_SL g90 ( 
.A(n_70),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_90),
.B(n_98),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_91),
.A2(n_97),
.B1(n_101),
.B2(n_82),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_70),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_94),
.B(n_67),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_84),
.A2(n_47),
.B1(n_52),
.B2(n_36),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_70),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_79),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_100),
.B(n_71),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_63),
.A2(n_52),
.B1(n_15),
.B2(n_19),
.Y(n_101)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_62),
.Y(n_105)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_105),
.Y(n_112)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_62),
.Y(n_106)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_106),
.Y(n_120)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_74),
.Y(n_109)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_109),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_110),
.B(n_103),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_96),
.A2(n_82),
.B1(n_61),
.B2(n_68),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_113),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_116),
.A2(n_126),
.B1(n_91),
.B2(n_96),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_89),
.B(n_59),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_117),
.B(n_122),
.Y(n_151)
);

INVx1_ASAP7_75t_SL g161 ( 
.A(n_119),
.Y(n_161)
);

CKINVDCx14_ASAP7_75t_R g123 ( 
.A(n_93),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_123),
.B(n_127),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_85),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_124),
.B(n_129),
.Y(n_145)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_97),
.Y(n_125)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_125),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_105),
.A2(n_82),
.B1(n_62),
.B2(n_72),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_107),
.B(n_73),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_102),
.B(n_77),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_128),
.B(n_130),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_108),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_102),
.B(n_60),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_100),
.B(n_78),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_131),
.B(n_88),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_106),
.B(n_76),
.C(n_65),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_132),
.B(n_134),
.C(n_104),
.Y(n_153)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_109),
.Y(n_133)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_133),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_94),
.B(n_65),
.C(n_58),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_99),
.B(n_83),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_135),
.B(n_83),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_121),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_136),
.B(n_143),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_138),
.B(n_160),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_140),
.A2(n_141),
.B1(n_159),
.B2(n_1),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_125),
.A2(n_94),
.B1(n_95),
.B2(n_98),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_121),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_SL g182 ( 
.A(n_144),
.B(n_21),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_133),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_146),
.B(n_150),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_148),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_130),
.B(n_103),
.Y(n_149)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_149),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_129),
.B(n_101),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_128),
.B(n_115),
.Y(n_152)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_152),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_153),
.B(n_126),
.C(n_113),
.Y(n_168)
);

HB1xp67_ASAP7_75t_L g154 ( 
.A(n_124),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_154),
.B(n_156),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_116),
.B(n_104),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_114),
.Y(n_157)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_157),
.Y(n_174)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_114),
.Y(n_158)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_158),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_134),
.A2(n_95),
.B1(n_90),
.B2(n_92),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_131),
.B(n_21),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_132),
.B(n_21),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_162),
.B(n_112),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_157),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_164),
.B(n_170),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_139),
.A2(n_110),
.B(n_120),
.Y(n_165)
);

O2A1O1Ixp33_ASAP7_75t_L g198 ( 
.A1(n_165),
.A2(n_167),
.B(n_177),
.C(n_180),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_155),
.A2(n_161),
.B(n_139),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_168),
.B(n_179),
.C(n_182),
.Y(n_188)
);

INVx1_ASAP7_75t_SL g170 ( 
.A(n_136),
.Y(n_170)
);

NOR3xp33_ASAP7_75t_L g171 ( 
.A(n_151),
.B(n_138),
.C(n_160),
.Y(n_171)
);

NOR3xp33_ASAP7_75t_SL g203 ( 
.A(n_171),
.B(n_175),
.C(n_41),
.Y(n_203)
);

AOI322xp5_ASAP7_75t_L g175 ( 
.A1(n_153),
.A2(n_118),
.A3(n_120),
.B1(n_112),
.B2(n_119),
.C1(n_58),
.C2(n_108),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_178),
.B(n_74),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_144),
.B(n_108),
.C(n_111),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_137),
.B(n_111),
.Y(n_180)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_180),
.Y(n_189)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_147),
.Y(n_183)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_183),
.Y(n_190)
);

HB1xp67_ASAP7_75t_L g184 ( 
.A(n_147),
.Y(n_184)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_184),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_137),
.B(n_1),
.Y(n_185)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_185),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_186),
.A2(n_149),
.B1(n_145),
.B2(n_141),
.Y(n_193)
);

OAI21xp33_ASAP7_75t_L g187 ( 
.A1(n_161),
.A2(n_2),
.B(n_3),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_187),
.A2(n_155),
.B1(n_143),
.B2(n_146),
.Y(n_191)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_191),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_172),
.A2(n_142),
.B1(n_159),
.B2(n_152),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_192),
.A2(n_200),
.B1(n_5),
.B2(n_7),
.Y(n_217)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_193),
.Y(n_214)
);

NAND2x1_ASAP7_75t_L g194 ( 
.A(n_167),
.B(n_151),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_194),
.A2(n_174),
.B1(n_8),
.B2(n_9),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_165),
.A2(n_158),
.B1(n_58),
.B2(n_41),
.Y(n_195)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_195),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_198),
.A2(n_7),
.B(n_10),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_179),
.B(n_41),
.C(n_87),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_199),
.B(n_202),
.C(n_205),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_166),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_200)
);

AND2x2_ASAP7_75t_L g201 ( 
.A(n_186),
.B(n_4),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_201),
.A2(n_181),
.B(n_183),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_168),
.B(n_182),
.C(n_163),
.Y(n_202)
);

OA21x2_ASAP7_75t_SL g207 ( 
.A1(n_203),
.A2(n_173),
.B(n_166),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_169),
.B(n_4),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_206),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_207),
.A2(n_217),
.B1(n_219),
.B2(n_220),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_194),
.A2(n_163),
.B(n_164),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_209),
.A2(n_191),
.B1(n_195),
.B2(n_203),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_196),
.B(n_170),
.Y(n_210)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_210),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_202),
.B(n_185),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_211),
.B(n_221),
.C(n_199),
.Y(n_224)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_212),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_189),
.A2(n_181),
.B(n_176),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_213),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_204),
.B(n_176),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g233 ( 
.A(n_218),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_198),
.A2(n_174),
.B(n_8),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_222),
.B(n_10),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_224),
.B(n_234),
.C(n_228),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_215),
.A2(n_201),
.B1(n_190),
.B2(n_197),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_226),
.B(n_228),
.Y(n_241)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_227),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_215),
.A2(n_188),
.B1(n_200),
.B2(n_205),
.Y(n_228)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_229),
.Y(n_243)
);

AND2x2_ASAP7_75t_L g231 ( 
.A(n_210),
.B(n_208),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_231),
.A2(n_212),
.B(n_222),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_221),
.B(n_211),
.C(n_188),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_223),
.A2(n_216),
.B1(n_219),
.B2(n_209),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_236),
.A2(n_232),
.B1(n_233),
.B2(n_231),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_234),
.B(n_218),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_237),
.B(n_11),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_238),
.B(n_224),
.C(n_12),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g249 ( 
.A1(n_239),
.A2(n_11),
.B(n_12),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_230),
.A2(n_214),
.B(n_217),
.Y(n_240)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_240),
.Y(n_247)
);

AO22x1_ASAP7_75t_L g242 ( 
.A1(n_230),
.A2(n_213),
.B1(n_214),
.B2(n_12),
.Y(n_242)
);

OR2x2_ASAP7_75t_L g245 ( 
.A(n_242),
.B(n_226),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_225),
.B(n_10),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_244),
.B(n_243),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_245),
.B(n_249),
.Y(n_254)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_246),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_248),
.B(n_249),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_250),
.B(n_235),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_251),
.B(n_252),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_241),
.B(n_13),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_253),
.B(n_248),
.C(n_236),
.Y(n_260)
);

NAND2x1p5_ASAP7_75t_L g256 ( 
.A(n_245),
.B(n_242),
.Y(n_256)
);

NOR2x1_ASAP7_75t_L g262 ( 
.A(n_256),
.B(n_254),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_258),
.B(n_247),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_259),
.B(n_261),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_260),
.B(n_255),
.C(n_14),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_254),
.B(n_13),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_262),
.B(n_263),
.Y(n_266)
);

NOR2xp67_ASAP7_75t_L g263 ( 
.A(n_257),
.B(n_14),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_264),
.B(n_263),
.C(n_265),
.Y(n_268)
);

BUFx24_ASAP7_75t_SL g267 ( 
.A(n_266),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_267),
.B(n_268),
.Y(n_269)
);


endmodule