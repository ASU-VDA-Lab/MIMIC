module fake_jpeg_27610_n_55 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_55);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_55;

wire n_13;
wire n_21;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_47;
wire n_22;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

INVx1_ASAP7_75t_L g8 ( 
.A(n_0),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_2),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_1),
.Y(n_11)
);

INVxp67_ASAP7_75t_L g12 ( 
.A(n_7),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

INVx1_ASAP7_75t_SL g14 ( 
.A(n_3),
.Y(n_14)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx5_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_17),
.B(n_18),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_12),
.B(n_4),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_19),
.B(n_21),
.Y(n_25)
);

A2O1A1Ixp33_ASAP7_75t_L g20 ( 
.A1(n_12),
.A2(n_0),
.B(n_1),
.C(n_2),
.Y(n_20)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

OR2x4_ASAP7_75t_L g21 ( 
.A(n_14),
.B(n_1),
.Y(n_21)
);

OAI22xp33_ASAP7_75t_L g22 ( 
.A1(n_14),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_22),
.Y(n_29)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_23),
.B(n_15),
.Y(n_26)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_26),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_21),
.B(n_11),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_27),
.B(n_9),
.Y(n_31)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_32),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_28),
.B(n_13),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_33),
.A2(n_35),
.B1(n_32),
.B2(n_34),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_28),
.B(n_8),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_34),
.B(n_36),
.C(n_20),
.Y(n_41)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_25),
.B(n_18),
.Y(n_36)
);

OAI21x1_ASAP7_75t_L g45 ( 
.A1(n_38),
.A2(n_29),
.B(n_37),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_36),
.A2(n_29),
.B1(n_23),
.B2(n_17),
.Y(n_39)
);

XOR2xp5_ASAP7_75t_L g44 ( 
.A(n_39),
.B(n_41),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_40),
.B(n_30),
.C(n_41),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_42),
.B(n_43),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_39),
.B(n_36),
.C(n_35),
.Y(n_43)
);

OR2x2_ASAP7_75t_L g47 ( 
.A(n_45),
.B(n_16),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_44),
.B(n_8),
.Y(n_46)
);

AOI21xp5_ASAP7_75t_L g50 ( 
.A1(n_46),
.A2(n_47),
.B(n_10),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_48),
.B(n_10),
.C(n_16),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_49),
.B(n_50),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_49),
.B(n_47),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_51),
.B(n_46),
.Y(n_53)
);

MAJx2_ASAP7_75t_L g54 ( 
.A(n_53),
.B(n_52),
.C(n_6),
.Y(n_54)
);

XNOR2xp5_ASAP7_75t_L g55 ( 
.A(n_54),
.B(n_6),
.Y(n_55)
);


endmodule