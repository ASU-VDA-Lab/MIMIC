module fake_jpeg_31366_n_515 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_515);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_515;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_145;
wire n_20;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx16f_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx10_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_16),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_4),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_14),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

INVx1_ASAP7_75t_SL g32 ( 
.A(n_2),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_0),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_6),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_15),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_5),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_12),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_11),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_10),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_3),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_3),
.Y(n_48)
);

BUFx16f_ASAP7_75t_L g49 ( 
.A(n_6),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_0),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_3),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_6),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_30),
.Y(n_53)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_53),
.Y(n_134)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_17),
.Y(n_54)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_54),
.Y(n_119)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_27),
.Y(n_55)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_55),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_21),
.B(n_8),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_56),
.B(n_102),
.Y(n_116)
);

BUFx12_ASAP7_75t_L g57 ( 
.A(n_17),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_57),
.B(n_73),
.Y(n_110)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_26),
.Y(n_58)
);

INVx5_ASAP7_75t_L g162 ( 
.A(n_58),
.Y(n_162)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_27),
.Y(n_59)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_59),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_19),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_60),
.Y(n_111)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_27),
.Y(n_61)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_61),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_21),
.B(n_8),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_62),
.B(n_69),
.Y(n_126)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_29),
.Y(n_63)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_63),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_19),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_64),
.Y(n_124)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_29),
.Y(n_65)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_65),
.Y(n_117)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_30),
.Y(n_66)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_66),
.Y(n_145)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_30),
.Y(n_67)
);

INVx8_ASAP7_75t_L g163 ( 
.A(n_67),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_19),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_68),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_21),
.B(n_8),
.Y(n_69)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_31),
.Y(n_70)
);

BUFx2_ASAP7_75t_L g154 ( 
.A(n_70),
.Y(n_154)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_29),
.Y(n_71)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_71),
.Y(n_118)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_29),
.Y(n_72)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_72),
.Y(n_122)
);

OR2x2_ASAP7_75t_L g73 ( 
.A(n_23),
.B(n_9),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_42),
.Y(n_74)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_74),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_19),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_75),
.Y(n_155)
);

BUFx5_ASAP7_75t_L g76 ( 
.A(n_26),
.Y(n_76)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_76),
.Y(n_107)
);

BUFx4f_ASAP7_75t_L g77 ( 
.A(n_17),
.Y(n_77)
);

HB1xp67_ASAP7_75t_L g112 ( 
.A(n_77),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_23),
.B(n_9),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_78),
.B(n_90),
.Y(n_147)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_31),
.Y(n_79)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_79),
.Y(n_137)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_42),
.Y(n_80)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_80),
.Y(n_132)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_24),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_81),
.Y(n_158)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_24),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_82),
.Y(n_159)
);

INVx2_ASAP7_75t_SL g83 ( 
.A(n_17),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_83),
.B(n_101),
.Y(n_113)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_24),
.Y(n_84)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_84),
.Y(n_121)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_42),
.Y(n_85)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_85),
.Y(n_133)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_52),
.Y(n_86)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_86),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_24),
.Y(n_87)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_87),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_44),
.Y(n_88)
);

INVx6_ASAP7_75t_L g149 ( 
.A(n_88),
.Y(n_149)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_42),
.Y(n_89)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_89),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_23),
.B(n_9),
.Y(n_90)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_31),
.Y(n_91)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_91),
.Y(n_143)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_26),
.Y(n_92)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_92),
.Y(n_127)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_43),
.Y(n_93)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_93),
.Y(n_160)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_43),
.Y(n_94)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_94),
.Y(n_142)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_44),
.Y(n_95)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_95),
.Y(n_144)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_44),
.Y(n_96)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_96),
.Y(n_151)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_44),
.Y(n_97)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_97),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_26),
.Y(n_98)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_98),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_52),
.Y(n_99)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_99),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_52),
.Y(n_100)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_100),
.Y(n_136)
);

BUFx12f_ASAP7_75t_L g101 ( 
.A(n_17),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_49),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_49),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_103),
.B(n_48),
.Y(n_138)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_49),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_104),
.B(n_105),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_49),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g115 ( 
.A1(n_81),
.A2(n_32),
.B1(n_22),
.B2(n_37),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_115),
.A2(n_123),
.B1(n_135),
.B2(n_18),
.Y(n_167)
);

BUFx2_ASAP7_75t_R g120 ( 
.A(n_77),
.Y(n_120)
);

CKINVDCx14_ASAP7_75t_R g219 ( 
.A(n_120),
.Y(n_219)
);

OAI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_82),
.A2(n_32),
.B1(n_49),
.B2(n_50),
.Y(n_123)
);

OA22x2_ASAP7_75t_L g129 ( 
.A1(n_73),
.A2(n_32),
.B1(n_22),
.B2(n_37),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_129),
.B(n_46),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_60),
.A2(n_25),
.B1(n_28),
.B2(n_34),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_138),
.B(n_156),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_57),
.B(n_25),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_140),
.B(n_148),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_53),
.A2(n_25),
.B1(n_28),
.B2(n_34),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_141),
.A2(n_152),
.B1(n_33),
.B2(n_47),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_79),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_66),
.A2(n_28),
.B1(n_34),
.B2(n_36),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_101),
.B(n_40),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_101),
.B(n_83),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_157),
.B(n_164),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_54),
.B(n_40),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_94),
.B(n_40),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_165),
.B(n_166),
.Y(n_191)
);

NAND3xp33_ASAP7_75t_L g166 ( 
.A(n_84),
.B(n_39),
.C(n_36),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g239 ( 
.A(n_167),
.B(n_180),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_169),
.Y(n_228)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_109),
.Y(n_170)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_170),
.Y(n_222)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_117),
.Y(n_171)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_171),
.Y(n_226)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_118),
.Y(n_172)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_172),
.Y(n_234)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_119),
.Y(n_173)
);

INVx13_ASAP7_75t_L g244 ( 
.A(n_173),
.Y(n_244)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_127),
.Y(n_174)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_174),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_116),
.B(n_39),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_175),
.B(n_214),
.Y(n_221)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_122),
.Y(n_176)
);

INVx4_ASAP7_75t_SL g250 ( 
.A(n_176),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_126),
.B(n_39),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_177),
.B(n_182),
.Y(n_245)
);

BUFx2_ASAP7_75t_L g178 ( 
.A(n_137),
.Y(n_178)
);

INVx3_ASAP7_75t_L g249 ( 
.A(n_178),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_113),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_179),
.B(n_181),
.Y(n_233)
);

INVx6_ASAP7_75t_SL g180 ( 
.A(n_111),
.Y(n_180)
);

HB1xp67_ASAP7_75t_L g181 ( 
.A(n_145),
.Y(n_181)
);

INVx8_ASAP7_75t_L g183 ( 
.A(n_119),
.Y(n_183)
);

INVx6_ASAP7_75t_L g232 ( 
.A(n_183),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_131),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_184),
.B(n_190),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_123),
.A2(n_96),
.B1(n_64),
.B2(n_68),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_186),
.A2(n_198),
.B1(n_218),
.B2(n_33),
.Y(n_246)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_125),
.Y(n_187)
);

INVx4_ASAP7_75t_L g220 ( 
.A(n_187),
.Y(n_220)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_106),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_188),
.B(n_203),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_L g189 ( 
.A1(n_166),
.A2(n_88),
.B1(n_75),
.B2(n_87),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_L g254 ( 
.A1(n_189),
.A2(n_160),
.B1(n_107),
.B2(n_180),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_126),
.B(n_147),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_111),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_192),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g193 ( 
.A(n_110),
.B(n_48),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_SL g229 ( 
.A(n_193),
.B(n_194),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_129),
.B(n_147),
.Y(n_194)
);

INVx6_ASAP7_75t_L g195 ( 
.A(n_124),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_195),
.Y(n_227)
);

AND2x2_ASAP7_75t_SL g196 ( 
.A(n_132),
.B(n_105),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_196),
.B(n_160),
.C(n_137),
.Y(n_242)
);

BUFx12f_ASAP7_75t_L g197 ( 
.A(n_162),
.Y(n_197)
);

INVx3_ASAP7_75t_L g258 ( 
.A(n_197),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_121),
.A2(n_100),
.B1(n_99),
.B2(n_98),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_133),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_199),
.Y(n_230)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_139),
.Y(n_200)
);

INVx5_ASAP7_75t_L g240 ( 
.A(n_200),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_154),
.A2(n_91),
.B1(n_67),
.B2(n_36),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g256 ( 
.A1(n_201),
.A2(n_208),
.B1(n_211),
.B2(n_212),
.Y(n_256)
);

INVx6_ASAP7_75t_L g202 ( 
.A(n_124),
.Y(n_202)
);

INVx8_ASAP7_75t_L g231 ( 
.A(n_202),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_152),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_108),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_204),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_150),
.Y(n_206)
);

INVx8_ASAP7_75t_L g241 ( 
.A(n_206),
.Y(n_241)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_114),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_207),
.Y(n_243)
);

INVx5_ASAP7_75t_L g208 ( 
.A(n_107),
.Y(n_208)
);

OAI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_129),
.A2(n_22),
.B1(n_37),
.B2(n_46),
.Y(n_209)
);

OAI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_209),
.A2(n_128),
.B1(n_149),
.B2(n_158),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_154),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_210),
.B(n_213),
.Y(n_223)
);

INVx4_ASAP7_75t_L g211 ( 
.A(n_142),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_150),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_146),
.B(n_46),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_144),
.Y(n_214)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_143),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_215),
.B(n_217),
.Y(n_247)
);

NAND2xp33_ASAP7_75t_SL g216 ( 
.A(n_115),
.B(n_45),
.Y(n_216)
);

A2O1A1Ixp33_ASAP7_75t_L g235 ( 
.A1(n_216),
.A2(n_141),
.B(n_130),
.C(n_136),
.Y(n_235)
);

INVx4_ASAP7_75t_L g217 ( 
.A(n_143),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_121),
.A2(n_102),
.B1(n_18),
.B2(n_33),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_225),
.A2(n_251),
.B1(n_253),
.B2(n_259),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_235),
.B(n_260),
.Y(n_269)
);

CKINVDCx12_ASAP7_75t_R g237 ( 
.A(n_219),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_237),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_242),
.B(n_193),
.Y(n_266)
);

AOI22xp33_ASAP7_75t_L g284 ( 
.A1(n_246),
.A2(n_195),
.B1(n_212),
.B2(n_206),
.Y(n_284)
);

OAI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_216),
.A2(n_182),
.B1(n_191),
.B2(n_167),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_185),
.B(n_47),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_252),
.B(n_168),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_175),
.A2(n_128),
.B1(n_149),
.B2(n_158),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_254),
.A2(n_198),
.B1(n_218),
.B2(n_208),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_182),
.B(n_153),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_257),
.B(n_196),
.Y(n_272)
);

OAI22xp33_ASAP7_75t_L g259 ( 
.A1(n_186),
.A2(n_161),
.B1(n_155),
.B2(n_159),
.Y(n_259)
);

A2O1A1Ixp33_ASAP7_75t_L g260 ( 
.A1(n_194),
.A2(n_35),
.B(n_38),
.C(n_51),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_261),
.A2(n_293),
.B1(n_241),
.B2(n_231),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_247),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_263),
.Y(n_300)
);

INVx3_ASAP7_75t_L g264 ( 
.A(n_232),
.Y(n_264)
);

INVx4_ASAP7_75t_L g298 ( 
.A(n_264),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_SL g312 ( 
.A(n_265),
.B(n_238),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_266),
.B(n_275),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_252),
.B(n_205),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_267),
.B(n_272),
.Y(n_307)
);

AOI22xp33_ASAP7_75t_SL g268 ( 
.A1(n_228),
.A2(n_178),
.B1(n_197),
.B2(n_217),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g316 ( 
.A(n_268),
.Y(n_316)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_224),
.Y(n_270)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_270),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_228),
.A2(n_239),
.B1(n_221),
.B2(n_235),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_271),
.A2(n_278),
.B1(n_282),
.B2(n_289),
.Y(n_295)
);

A2O1A1Ixp33_ASAP7_75t_L g274 ( 
.A1(n_257),
.A2(n_194),
.B(n_193),
.C(n_196),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_SL g311 ( 
.A1(n_274),
.A2(n_277),
.B(n_287),
.Y(n_311)
);

AND2x2_ASAP7_75t_SL g275 ( 
.A(n_221),
.B(n_172),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_230),
.Y(n_276)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_276),
.Y(n_297)
);

AOI22xp33_ASAP7_75t_SL g277 ( 
.A1(n_256),
.A2(n_197),
.B1(n_215),
.B2(n_163),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_239),
.A2(n_248),
.B1(n_246),
.B2(n_245),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_223),
.B(n_171),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_279),
.B(n_280),
.Y(n_323)
);

CKINVDCx14_ASAP7_75t_R g280 ( 
.A(n_223),
.Y(n_280)
);

INVx3_ASAP7_75t_L g281 ( 
.A(n_232),
.Y(n_281)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_281),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_239),
.A2(n_155),
.B1(n_159),
.B2(n_202),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_242),
.B(n_176),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_283),
.B(n_290),
.Y(n_308)
);

AOI22xp33_ASAP7_75t_L g303 ( 
.A1(n_284),
.A2(n_285),
.B1(n_250),
.B2(n_243),
.Y(n_303)
);

AOI22xp33_ASAP7_75t_L g285 ( 
.A1(n_253),
.A2(n_151),
.B1(n_200),
.B2(n_199),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_247),
.Y(n_286)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_286),
.Y(n_324)
);

AOI22xp33_ASAP7_75t_SL g287 ( 
.A1(n_249),
.A2(n_163),
.B1(n_183),
.B2(n_173),
.Y(n_287)
);

OA22x2_ASAP7_75t_L g288 ( 
.A1(n_259),
.A2(n_211),
.B1(n_187),
.B2(n_50),
.Y(n_288)
);

CKINVDCx16_ASAP7_75t_R g306 ( 
.A(n_288),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_255),
.A2(n_192),
.B1(n_134),
.B2(n_112),
.Y(n_289)
);

HB1xp67_ASAP7_75t_L g290 ( 
.A(n_249),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_229),
.B(n_18),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_291),
.B(n_292),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_229),
.B(n_47),
.Y(n_292)
);

AOI22xp33_ASAP7_75t_SL g293 ( 
.A1(n_222),
.A2(n_112),
.B1(n_43),
.B2(n_48),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_L g294 ( 
.A1(n_260),
.A2(n_51),
.B(n_50),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_L g299 ( 
.A1(n_294),
.A2(n_233),
.B(n_35),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_L g329 ( 
.A1(n_296),
.A2(n_262),
.B1(n_264),
.B2(n_281),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_L g357 ( 
.A1(n_299),
.A2(n_20),
.B(n_7),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_266),
.B(n_222),
.C(n_236),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_301),
.B(n_315),
.C(n_320),
.Y(n_327)
);

AOI32xp33_ASAP7_75t_L g302 ( 
.A1(n_269),
.A2(n_271),
.A3(n_267),
.B1(n_263),
.B2(n_274),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_SL g328 ( 
.A1(n_302),
.A2(n_318),
.B(n_265),
.Y(n_328)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_303),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_278),
.A2(n_236),
.B1(n_243),
.B2(n_238),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_304),
.A2(n_319),
.B1(n_284),
.B2(n_285),
.Y(n_330)
);

NAND3xp33_ASAP7_75t_L g334 ( 
.A(n_312),
.B(n_289),
.C(n_262),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_280),
.A2(n_258),
.B1(n_231),
.B2(n_241),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g337 ( 
.A(n_314),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_283),
.B(n_274),
.C(n_292),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_275),
.B(n_226),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_317),
.B(n_288),
.Y(n_335)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_269),
.A2(n_294),
.B(n_282),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_261),
.A2(n_250),
.B1(n_227),
.B2(n_220),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_291),
.B(n_220),
.C(n_226),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_279),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_321),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_275),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_322),
.Y(n_351)
);

CKINVDCx16_ASAP7_75t_R g325 ( 
.A(n_286),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_325),
.B(n_275),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_L g326 ( 
.A1(n_272),
.A2(n_258),
.B(n_234),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_L g336 ( 
.A1(n_326),
.A2(n_240),
.B(n_234),
.Y(n_336)
);

AOI21xp5_ASAP7_75t_L g388 ( 
.A1(n_328),
.A2(n_333),
.B(n_298),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_329),
.A2(n_330),
.B1(n_321),
.B2(n_322),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_331),
.B(n_299),
.Y(n_376)
);

OAI21xp5_ASAP7_75t_SL g333 ( 
.A1(n_318),
.A2(n_290),
.B(n_273),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_334),
.B(n_355),
.Y(n_360)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_335),
.Y(n_369)
);

INVxp67_ASAP7_75t_L g368 ( 
.A(n_336),
.Y(n_368)
);

AO22x1_ASAP7_75t_L g338 ( 
.A1(n_300),
.A2(n_288),
.B1(n_250),
.B2(n_276),
.Y(n_338)
);

OA21x2_ASAP7_75t_L g384 ( 
.A1(n_338),
.A2(n_319),
.B(n_305),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_313),
.B(n_230),
.C(n_288),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_339),
.B(n_348),
.C(n_350),
.Y(n_366)
);

OAI32xp33_ASAP7_75t_L g341 ( 
.A1(n_323),
.A2(n_288),
.A3(n_51),
.B1(n_45),
.B2(n_35),
.Y(n_341)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_341),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_306),
.A2(n_227),
.B1(n_270),
.B2(n_224),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_L g386 ( 
.A1(n_342),
.A2(n_343),
.B1(n_354),
.B2(n_309),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_306),
.A2(n_270),
.B1(n_240),
.B2(n_244),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_323),
.B(n_45),
.Y(n_344)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_344),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_300),
.B(n_41),
.Y(n_345)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_345),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_312),
.B(n_244),
.Y(n_346)
);

CKINVDCx16_ASAP7_75t_R g358 ( 
.A(n_346),
.Y(n_358)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_317),
.Y(n_347)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_347),
.Y(n_379)
);

XOR2xp5_ASAP7_75t_L g348 ( 
.A(n_302),
.B(n_20),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_SL g349 ( 
.A(n_307),
.B(n_41),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_SL g359 ( 
.A(n_349),
.B(n_307),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_313),
.B(n_315),
.Y(n_350)
);

INVxp33_ASAP7_75t_SL g352 ( 
.A(n_314),
.Y(n_352)
);

INVxp67_ASAP7_75t_L g374 ( 
.A(n_352),
.Y(n_374)
);

AOI21xp5_ASAP7_75t_L g353 ( 
.A1(n_311),
.A2(n_10),
.B(n_16),
.Y(n_353)
);

OAI21xp5_ASAP7_75t_SL g362 ( 
.A1(n_353),
.A2(n_316),
.B(n_344),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_308),
.A2(n_41),
.B1(n_38),
.B2(n_2),
.Y(n_354)
);

AOI32xp33_ASAP7_75t_L g355 ( 
.A1(n_308),
.A2(n_20),
.A3(n_38),
.B1(n_9),
.B2(n_11),
.Y(n_355)
);

CKINVDCx16_ASAP7_75t_R g356 ( 
.A(n_324),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_356),
.B(n_304),
.Y(n_371)
);

INVxp67_ASAP7_75t_L g375 ( 
.A(n_357),
.Y(n_375)
);

CKINVDCx14_ASAP7_75t_R g401 ( 
.A(n_359),
.Y(n_401)
);

CKINVDCx16_ASAP7_75t_R g361 ( 
.A(n_345),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_SL g403 ( 
.A(n_361),
.B(n_370),
.Y(n_403)
);

AND2x2_ASAP7_75t_SL g406 ( 
.A(n_362),
.B(n_333),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_363),
.A2(n_365),
.B1(n_367),
.B2(n_372),
.Y(n_389)
);

XOR2xp5_ASAP7_75t_L g364 ( 
.A(n_350),
.B(n_315),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_L g391 ( 
.A(n_364),
.B(n_383),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_329),
.A2(n_324),
.B1(n_325),
.B2(n_295),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_337),
.A2(n_332),
.B1(n_338),
.B2(n_340),
.Y(n_367)
);

CKINVDCx16_ASAP7_75t_R g370 ( 
.A(n_347),
.Y(n_370)
);

CKINVDCx16_ASAP7_75t_R g395 ( 
.A(n_371),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_337),
.A2(n_295),
.B1(n_311),
.B2(n_296),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_376),
.B(n_386),
.Y(n_396)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_338),
.Y(n_380)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_380),
.Y(n_402)
);

AOI21xp5_ASAP7_75t_SL g381 ( 
.A1(n_335),
.A2(n_326),
.B(n_305),
.Y(n_381)
);

OAI21xp5_ASAP7_75t_L g399 ( 
.A1(n_381),
.A2(n_388),
.B(n_357),
.Y(n_399)
);

OAI21xp5_ASAP7_75t_SL g382 ( 
.A1(n_353),
.A2(n_301),
.B(n_303),
.Y(n_382)
);

AO21x1_ASAP7_75t_L g410 ( 
.A1(n_382),
.A2(n_355),
.B(n_341),
.Y(n_410)
);

XOR2xp5_ASAP7_75t_L g383 ( 
.A(n_327),
.B(n_320),
.Y(n_383)
);

AND2x2_ASAP7_75t_L g404 ( 
.A(n_384),
.B(n_343),
.Y(n_404)
);

XOR2xp5_ASAP7_75t_L g385 ( 
.A(n_327),
.B(n_310),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_L g407 ( 
.A(n_385),
.B(n_387),
.Y(n_407)
);

XOR2xp5_ASAP7_75t_L g387 ( 
.A(n_348),
.B(n_310),
.Y(n_387)
);

BUFx6f_ASAP7_75t_L g390 ( 
.A(n_380),
.Y(n_390)
);

HB1xp67_ASAP7_75t_L g423 ( 
.A(n_390),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_359),
.B(n_349),
.Y(n_392)
);

CKINVDCx16_ASAP7_75t_R g431 ( 
.A(n_392),
.Y(n_431)
);

A2O1A1O1Ixp25_ASAP7_75t_L g393 ( 
.A1(n_369),
.A2(n_328),
.B(n_340),
.C(n_351),
.D(n_336),
.Y(n_393)
);

XOR2xp5_ASAP7_75t_L g425 ( 
.A(n_393),
.B(n_388),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_363),
.A2(n_339),
.B1(n_332),
.B2(n_351),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_L g433 ( 
.A1(n_394),
.A2(n_368),
.B1(n_374),
.B2(n_369),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_378),
.B(n_356),
.Y(n_397)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_397),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_367),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_398),
.B(n_411),
.Y(n_430)
);

AOI21xp5_ASAP7_75t_L g426 ( 
.A1(n_399),
.A2(n_410),
.B(n_362),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_378),
.B(n_354),
.Y(n_400)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_400),
.Y(n_419)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_404),
.Y(n_424)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_379),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_405),
.B(n_408),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_406),
.B(n_382),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_377),
.B(n_342),
.Y(n_408)
);

AOI22xp33_ASAP7_75t_SL g409 ( 
.A1(n_373),
.A2(n_298),
.B1(n_309),
.B2(n_297),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_L g421 ( 
.A1(n_409),
.A2(n_374),
.B1(n_365),
.B2(n_372),
.Y(n_421)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_379),
.Y(n_411)
);

A2O1A1Ixp33_ASAP7_75t_SL g412 ( 
.A1(n_384),
.A2(n_330),
.B(n_298),
.C(n_297),
.Y(n_412)
);

OAI21xp5_ASAP7_75t_SL g418 ( 
.A1(n_412),
.A2(n_381),
.B(n_386),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_358),
.B(n_376),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_SL g437 ( 
.A(n_413),
.B(n_414),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_384),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_377),
.B(n_0),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_415),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_391),
.B(n_383),
.C(n_364),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_416),
.B(n_422),
.C(n_432),
.Y(n_445)
);

INVxp67_ASAP7_75t_L g443 ( 
.A(n_418),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_SL g420 ( 
.A(n_407),
.B(n_366),
.Y(n_420)
);

XOR2xp5_ASAP7_75t_L g449 ( 
.A(n_420),
.B(n_429),
.Y(n_449)
);

AOI22xp5_ASAP7_75t_L g447 ( 
.A1(n_421),
.A2(n_404),
.B1(n_389),
.B2(n_402),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_391),
.B(n_407),
.C(n_385),
.Y(n_422)
);

OR2x2_ASAP7_75t_L g448 ( 
.A(n_425),
.B(n_436),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_L g444 ( 
.A(n_426),
.B(n_406),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_394),
.B(n_366),
.C(n_387),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_433),
.A2(n_435),
.B1(n_402),
.B2(n_408),
.Y(n_439)
);

NAND3xp33_ASAP7_75t_L g434 ( 
.A(n_401),
.B(n_360),
.C(n_375),
.Y(n_434)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_434),
.Y(n_440)
);

AOI22xp5_ASAP7_75t_L g435 ( 
.A1(n_389),
.A2(n_373),
.B1(n_368),
.B2(n_375),
.Y(n_435)
);

FAx1_ASAP7_75t_SL g436 ( 
.A(n_406),
.B(n_20),
.CI(n_7),
.CON(n_436),
.SN(n_436)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_437),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_438),
.B(n_442),
.Y(n_464)
);

AOI22xp5_ASAP7_75t_L g459 ( 
.A1(n_439),
.A2(n_454),
.B1(n_404),
.B2(n_419),
.Y(n_459)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_423),
.Y(n_441)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_441),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_SL g442 ( 
.A(n_431),
.B(n_395),
.Y(n_442)
);

XOR2xp5_ASAP7_75t_L g458 ( 
.A(n_444),
.B(n_447),
.Y(n_458)
);

XNOR2xp5_ASAP7_75t_L g446 ( 
.A(n_432),
.B(n_396),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_446),
.B(n_422),
.C(n_416),
.Y(n_457)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_417),
.Y(n_450)
);

AOI22xp33_ASAP7_75t_SL g471 ( 
.A1(n_450),
.A2(n_451),
.B1(n_452),
.B2(n_418),
.Y(n_471)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_417),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_428),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_SL g453 ( 
.A(n_427),
.B(n_403),
.Y(n_453)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_453),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_SL g454 ( 
.A1(n_424),
.A2(n_390),
.B1(n_399),
.B2(n_396),
.Y(n_454)
);

BUFx24_ASAP7_75t_SL g455 ( 
.A(n_425),
.Y(n_455)
);

INVxp33_ASAP7_75t_SL g456 ( 
.A(n_455),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_457),
.B(n_20),
.Y(n_481)
);

XOR2xp5_ASAP7_75t_L g485 ( 
.A(n_459),
.B(n_0),
.Y(n_485)
);

AOI21xp5_ASAP7_75t_L g460 ( 
.A1(n_440),
.A2(n_429),
.B(n_426),
.Y(n_460)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_460),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_446),
.B(n_420),
.C(n_433),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_461),
.B(n_462),
.C(n_466),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_445),
.B(n_435),
.C(n_430),
.Y(n_462)
);

AOI22xp5_ASAP7_75t_L g465 ( 
.A1(n_439),
.A2(n_443),
.B1(n_454),
.B2(n_419),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_SL g482 ( 
.A1(n_465),
.A2(n_471),
.B1(n_7),
.B2(n_13),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_445),
.B(n_428),
.C(n_424),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_449),
.B(n_443),
.C(n_447),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_467),
.B(n_436),
.C(n_20),
.Y(n_480)
);

XOR2xp5_ASAP7_75t_SL g468 ( 
.A(n_444),
.B(n_393),
.Y(n_468)
);

AOI21xp33_ASAP7_75t_SL g478 ( 
.A1(n_468),
.A2(n_436),
.B(n_412),
.Y(n_478)
);

OAI21xp5_ASAP7_75t_SL g469 ( 
.A1(n_448),
.A2(n_411),
.B(n_405),
.Y(n_469)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_469),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_463),
.B(n_448),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_472),
.B(n_474),
.Y(n_491)
);

AOI22xp5_ASAP7_75t_L g473 ( 
.A1(n_458),
.A2(n_412),
.B1(n_410),
.B2(n_449),
.Y(n_473)
);

OAI22xp5_ASAP7_75t_L g496 ( 
.A1(n_473),
.A2(n_483),
.B1(n_11),
.B2(n_13),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_464),
.B(n_462),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_L g475 ( 
.A(n_461),
.B(n_397),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_475),
.B(n_476),
.Y(n_493)
);

OAI22xp5_ASAP7_75t_SL g476 ( 
.A1(n_459),
.A2(n_400),
.B1(n_412),
.B2(n_415),
.Y(n_476)
);

A2O1A1Ixp33_ASAP7_75t_SL g486 ( 
.A1(n_478),
.A2(n_468),
.B(n_467),
.C(n_465),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_SL g490 ( 
.A(n_480),
.B(n_481),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_482),
.B(n_485),
.Y(n_489)
);

AOI22xp5_ASAP7_75t_L g483 ( 
.A1(n_458),
.A2(n_7),
.B1(n_13),
.B2(n_12),
.Y(n_483)
);

XOR2xp5_ASAP7_75t_L g498 ( 
.A(n_486),
.B(n_496),
.Y(n_498)
);

A2O1A1Ixp33_ASAP7_75t_SL g487 ( 
.A1(n_479),
.A2(n_466),
.B(n_470),
.C(n_457),
.Y(n_487)
);

AOI21xp33_ASAP7_75t_L g502 ( 
.A1(n_487),
.A2(n_486),
.B(n_491),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_SL g488 ( 
.A(n_484),
.B(n_456),
.Y(n_488)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_488),
.Y(n_499)
);

AND2x2_ASAP7_75t_L g492 ( 
.A(n_477),
.B(n_10),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_492),
.B(n_495),
.Y(n_501)
);

AOI21xp5_ASAP7_75t_SL g494 ( 
.A1(n_475),
.A2(n_10),
.B(n_13),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_494),
.B(n_12),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_477),
.B(n_5),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_493),
.B(n_485),
.C(n_482),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_497),
.B(n_500),
.Y(n_506)
);

NOR2xp67_ASAP7_75t_SL g504 ( 
.A(n_502),
.B(n_487),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_489),
.B(n_473),
.Y(n_503)
);

XNOR2xp5_ASAP7_75t_L g507 ( 
.A(n_503),
.B(n_483),
.Y(n_507)
);

OAI21xp5_ASAP7_75t_L g508 ( 
.A1(n_504),
.A2(n_507),
.B(n_497),
.Y(n_508)
);

OAI21xp5_ASAP7_75t_SL g505 ( 
.A1(n_499),
.A2(n_490),
.B(n_480),
.Y(n_505)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_505),
.Y(n_509)
);

OAI21xp5_ASAP7_75t_SL g510 ( 
.A1(n_508),
.A2(n_506),
.B(n_498),
.Y(n_510)
);

AOI21xp5_ASAP7_75t_SL g511 ( 
.A1(n_510),
.A2(n_509),
.B(n_498),
.Y(n_511)
);

A2O1A1O1Ixp25_ASAP7_75t_L g512 ( 
.A1(n_511),
.A2(n_501),
.B(n_4),
.C(n_14),
.D(n_2),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_512),
.Y(n_513)
);

OAI22xp33_ASAP7_75t_SL g514 ( 
.A1(n_513),
.A2(n_4),
.B1(n_14),
.B2(n_3),
.Y(n_514)
);

OA21x2_ASAP7_75t_L g515 ( 
.A1(n_514),
.A2(n_1),
.B(n_2),
.Y(n_515)
);


endmodule