module fake_aes_2619_n_705 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_705);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_705;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_699;
wire n_693;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_420;
wire n_342;
wire n_423;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_78;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
BUFx3_ASAP7_75t_L g77 ( .A(n_47), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_19), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_21), .Y(n_79) );
CKINVDCx5p33_ASAP7_75t_R g80 ( .A(n_27), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_6), .Y(n_81) );
BUFx6f_ASAP7_75t_L g82 ( .A(n_11), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_20), .Y(n_83) );
CKINVDCx5p33_ASAP7_75t_R g84 ( .A(n_36), .Y(n_84) );
INVx2_ASAP7_75t_L g85 ( .A(n_12), .Y(n_85) );
CKINVDCx20_ASAP7_75t_R g86 ( .A(n_70), .Y(n_86) );
INVxp67_ASAP7_75t_SL g87 ( .A(n_72), .Y(n_87) );
INVxp33_ASAP7_75t_L g88 ( .A(n_12), .Y(n_88) );
CKINVDCx20_ASAP7_75t_R g89 ( .A(n_8), .Y(n_89) );
CKINVDCx20_ASAP7_75t_R g90 ( .A(n_29), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_48), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_2), .Y(n_92) );
INVx2_ASAP7_75t_L g93 ( .A(n_62), .Y(n_93) );
CKINVDCx20_ASAP7_75t_R g94 ( .A(n_43), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_42), .Y(n_95) );
CKINVDCx5p33_ASAP7_75t_R g96 ( .A(n_33), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_11), .Y(n_97) );
INVx2_ASAP7_75t_SL g98 ( .A(n_76), .Y(n_98) );
CKINVDCx16_ASAP7_75t_R g99 ( .A(n_66), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_75), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_28), .Y(n_101) );
CKINVDCx5p33_ASAP7_75t_R g102 ( .A(n_52), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_9), .Y(n_103) );
BUFx2_ASAP7_75t_L g104 ( .A(n_34), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_1), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_44), .Y(n_106) );
INVx2_ASAP7_75t_L g107 ( .A(n_38), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_4), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_14), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_57), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_23), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_16), .Y(n_112) );
INVxp67_ASAP7_75t_L g113 ( .A(n_31), .Y(n_113) );
CKINVDCx16_ASAP7_75t_R g114 ( .A(n_45), .Y(n_114) );
INVxp33_ASAP7_75t_L g115 ( .A(n_40), .Y(n_115) );
BUFx3_ASAP7_75t_L g116 ( .A(n_61), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_37), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_30), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_65), .Y(n_119) );
INVx2_ASAP7_75t_L g120 ( .A(n_64), .Y(n_120) );
INVxp67_ASAP7_75t_SL g121 ( .A(n_55), .Y(n_121) );
CKINVDCx5p33_ASAP7_75t_R g122 ( .A(n_15), .Y(n_122) );
CKINVDCx5p33_ASAP7_75t_R g123 ( .A(n_24), .Y(n_123) );
INVx2_ASAP7_75t_L g124 ( .A(n_56), .Y(n_124) );
CKINVDCx20_ASAP7_75t_R g125 ( .A(n_89), .Y(n_125) );
CKINVDCx5p33_ASAP7_75t_R g126 ( .A(n_86), .Y(n_126) );
INVx6_ASAP7_75t_L g127 ( .A(n_77), .Y(n_127) );
AND2x2_ASAP7_75t_L g128 ( .A(n_104), .B(n_0), .Y(n_128) );
INVx2_ASAP7_75t_L g129 ( .A(n_93), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_83), .Y(n_130) );
OAI22xp5_ASAP7_75t_SL g131 ( .A1(n_122), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_131) );
INVx2_ASAP7_75t_L g132 ( .A(n_93), .Y(n_132) );
BUFx8_ASAP7_75t_L g133 ( .A(n_104), .Y(n_133) );
OAI22xp5_ASAP7_75t_SL g134 ( .A1(n_122), .A2(n_88), .B1(n_92), .B2(n_112), .Y(n_134) );
BUFx6f_ASAP7_75t_L g135 ( .A(n_77), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g136 ( .A(n_98), .B(n_3), .Y(n_136) );
BUFx6f_ASAP7_75t_L g137 ( .A(n_116), .Y(n_137) );
BUFx2_ASAP7_75t_L g138 ( .A(n_99), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g139 ( .A(n_98), .B(n_3), .Y(n_139) );
INVx2_ASAP7_75t_L g140 ( .A(n_107), .Y(n_140) );
INVxp67_ASAP7_75t_L g141 ( .A(n_97), .Y(n_141) );
INVx2_ASAP7_75t_L g142 ( .A(n_107), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_83), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_91), .Y(n_144) );
INVx2_ASAP7_75t_L g145 ( .A(n_120), .Y(n_145) );
BUFx2_ASAP7_75t_L g146 ( .A(n_114), .Y(n_146) );
AND2x4_ASAP7_75t_L g147 ( .A(n_85), .B(n_4), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g148 ( .A(n_103), .B(n_5), .Y(n_148) );
CKINVDCx5p33_ASAP7_75t_R g149 ( .A(n_90), .Y(n_149) );
INVxp67_ASAP7_75t_L g150 ( .A(n_105), .Y(n_150) );
OR2x2_ASAP7_75t_L g151 ( .A(n_81), .B(n_5), .Y(n_151) );
BUFx3_ASAP7_75t_L g152 ( .A(n_116), .Y(n_152) );
BUFx6f_ASAP7_75t_L g153 ( .A(n_82), .Y(n_153) );
INVx3_ASAP7_75t_L g154 ( .A(n_82), .Y(n_154) );
INVx2_ASAP7_75t_L g155 ( .A(n_120), .Y(n_155) );
INVx2_ASAP7_75t_L g156 ( .A(n_124), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_91), .Y(n_157) );
INVx2_ASAP7_75t_L g158 ( .A(n_124), .Y(n_158) );
BUFx6f_ASAP7_75t_L g159 ( .A(n_82), .Y(n_159) );
CKINVDCx5p33_ASAP7_75t_R g160 ( .A(n_94), .Y(n_160) );
NOR2xp33_ASAP7_75t_L g161 ( .A(n_78), .B(n_6), .Y(n_161) );
AND2x2_ASAP7_75t_L g162 ( .A(n_115), .B(n_7), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_108), .B(n_7), .Y(n_163) );
AND2x4_ASAP7_75t_L g164 ( .A(n_85), .B(n_8), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_106), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_106), .Y(n_166) );
INVx2_ASAP7_75t_L g167 ( .A(n_110), .Y(n_167) );
AND2x2_ASAP7_75t_L g168 ( .A(n_128), .B(n_92), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_132), .Y(n_169) );
INVx2_ASAP7_75t_L g170 ( .A(n_135), .Y(n_170) );
INVx2_ASAP7_75t_L g171 ( .A(n_135), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_132), .Y(n_172) );
AND2x6_ASAP7_75t_L g173 ( .A(n_128), .B(n_111), .Y(n_173) );
INVx8_ASAP7_75t_L g174 ( .A(n_147), .Y(n_174) );
INVx2_ASAP7_75t_L g175 ( .A(n_135), .Y(n_175) );
AND2x4_ASAP7_75t_L g176 ( .A(n_147), .B(n_112), .Y(n_176) );
INVx2_ASAP7_75t_L g177 ( .A(n_135), .Y(n_177) );
NAND2xp5_ASAP7_75t_SL g178 ( .A(n_133), .B(n_80), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_132), .Y(n_179) );
INVxp67_ASAP7_75t_SL g180 ( .A(n_133), .Y(n_180) );
INVx1_ASAP7_75t_SL g181 ( .A(n_138), .Y(n_181) );
BUFx3_ASAP7_75t_L g182 ( .A(n_152), .Y(n_182) );
INVx2_ASAP7_75t_L g183 ( .A(n_135), .Y(n_183) );
INVx4_ASAP7_75t_L g184 ( .A(n_147), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_140), .Y(n_185) );
NOR2xp33_ASAP7_75t_L g186 ( .A(n_138), .B(n_113), .Y(n_186) );
NOR2x1p5_ASAP7_75t_L g187 ( .A(n_126), .B(n_123), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_140), .Y(n_188) );
NAND2xp5_ASAP7_75t_SL g189 ( .A(n_133), .B(n_146), .Y(n_189) );
BUFx2_ASAP7_75t_L g190 ( .A(n_133), .Y(n_190) );
INVx2_ASAP7_75t_L g191 ( .A(n_137), .Y(n_191) );
BUFx10_ASAP7_75t_L g192 ( .A(n_127), .Y(n_192) );
INVx2_ASAP7_75t_SL g193 ( .A(n_127), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_140), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_146), .B(n_123), .Y(n_195) );
AOI22xp33_ASAP7_75t_L g196 ( .A1(n_134), .A2(n_81), .B1(n_109), .B2(n_82), .Y(n_196) );
INVx2_ASAP7_75t_L g197 ( .A(n_137), .Y(n_197) );
INVx1_ASAP7_75t_L g198 ( .A(n_142), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_142), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_142), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_147), .Y(n_201) );
AND2x2_ASAP7_75t_L g202 ( .A(n_141), .B(n_102), .Y(n_202) );
INVx5_ASAP7_75t_L g203 ( .A(n_137), .Y(n_203) );
AND2x2_ASAP7_75t_L g204 ( .A(n_150), .B(n_102), .Y(n_204) );
AOI22xp33_ASAP7_75t_L g205 ( .A1(n_134), .A2(n_82), .B1(n_119), .B2(n_110), .Y(n_205) );
BUFx3_ASAP7_75t_L g206 ( .A(n_152), .Y(n_206) );
AND2x2_ASAP7_75t_L g207 ( .A(n_162), .B(n_118), .Y(n_207) );
INVx2_ASAP7_75t_L g208 ( .A(n_137), .Y(n_208) );
OAI22xp33_ASAP7_75t_L g209 ( .A1(n_151), .A2(n_80), .B1(n_118), .B2(n_84), .Y(n_209) );
OR2x2_ASAP7_75t_L g210 ( .A(n_151), .B(n_84), .Y(n_210) );
AND2x2_ASAP7_75t_L g211 ( .A(n_162), .B(n_96), .Y(n_211) );
BUFx3_ASAP7_75t_L g212 ( .A(n_152), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_164), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_130), .B(n_96), .Y(n_214) );
HB1xp67_ASAP7_75t_L g215 ( .A(n_149), .Y(n_215) );
INVx4_ASAP7_75t_L g216 ( .A(n_164), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_164), .Y(n_217) );
NAND2xp5_ASAP7_75t_SL g218 ( .A(n_130), .B(n_101), .Y(n_218) );
INVx3_ASAP7_75t_L g219 ( .A(n_164), .Y(n_219) );
NAND2xp5_ASAP7_75t_SL g220 ( .A(n_143), .B(n_100), .Y(n_220) );
BUFx6f_ASAP7_75t_L g221 ( .A(n_153), .Y(n_221) );
INVx1_ASAP7_75t_L g222 ( .A(n_154), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_154), .Y(n_223) );
INVx2_ASAP7_75t_SL g224 ( .A(n_127), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_154), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_154), .Y(n_226) );
INVx2_ASAP7_75t_L g227 ( .A(n_137), .Y(n_227) );
NOR2xp33_ASAP7_75t_L g228 ( .A(n_143), .B(n_95), .Y(n_228) );
AOI22xp5_ASAP7_75t_L g229 ( .A1(n_131), .A2(n_119), .B1(n_117), .B2(n_111), .Y(n_229) );
BUFx6f_ASAP7_75t_L g230 ( .A(n_153), .Y(n_230) );
NAND2xp5_ASAP7_75t_SL g231 ( .A(n_144), .B(n_79), .Y(n_231) );
HB1xp67_ASAP7_75t_L g232 ( .A(n_181), .Y(n_232) );
INVx2_ASAP7_75t_L g233 ( .A(n_170), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_174), .Y(n_234) );
INVx2_ASAP7_75t_L g235 ( .A(n_170), .Y(n_235) );
INVx3_ASAP7_75t_L g236 ( .A(n_184), .Y(n_236) );
AND2x2_ASAP7_75t_L g237 ( .A(n_202), .B(n_166), .Y(n_237) );
NOR2xp33_ASAP7_75t_L g238 ( .A(n_195), .B(n_139), .Y(n_238) );
BUFx2_ASAP7_75t_L g239 ( .A(n_190), .Y(n_239) );
AOI22xp33_ASAP7_75t_SL g240 ( .A1(n_190), .A2(n_131), .B1(n_160), .B2(n_125), .Y(n_240) );
A2O1A1Ixp33_ASAP7_75t_L g241 ( .A1(n_201), .A2(n_157), .B(n_166), .C(n_165), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_174), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_174), .Y(n_243) );
CKINVDCx5p33_ASAP7_75t_R g244 ( .A(n_180), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_214), .B(n_165), .Y(n_245) );
INVxp67_ASAP7_75t_L g246 ( .A(n_210), .Y(n_246) );
BUFx6f_ASAP7_75t_L g247 ( .A(n_174), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_202), .B(n_144), .Y(n_248) );
INVxp67_ASAP7_75t_L g249 ( .A(n_210), .Y(n_249) );
AND2x2_ASAP7_75t_L g250 ( .A(n_204), .B(n_157), .Y(n_250) );
NOR2xp33_ASAP7_75t_L g251 ( .A(n_186), .B(n_136), .Y(n_251) );
NOR2xp33_ASAP7_75t_L g252 ( .A(n_204), .B(n_148), .Y(n_252) );
BUFx3_ASAP7_75t_L g253 ( .A(n_174), .Y(n_253) );
INVx5_ASAP7_75t_L g254 ( .A(n_173), .Y(n_254) );
AOI22xp5_ASAP7_75t_L g255 ( .A1(n_173), .A2(n_161), .B1(n_163), .B2(n_167), .Y(n_255) );
NOR2x1p5_ASAP7_75t_L g256 ( .A(n_207), .B(n_87), .Y(n_256) );
NAND2xp5_ASAP7_75t_SL g257 ( .A(n_184), .B(n_117), .Y(n_257) );
BUFx3_ASAP7_75t_L g258 ( .A(n_182), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_176), .Y(n_259) );
HB1xp67_ASAP7_75t_L g260 ( .A(n_207), .Y(n_260) );
NAND2xp5_ASAP7_75t_SL g261 ( .A(n_184), .B(n_167), .Y(n_261) );
NAND2xp5_ASAP7_75t_SL g262 ( .A(n_184), .B(n_216), .Y(n_262) );
AND2x4_ASAP7_75t_L g263 ( .A(n_168), .B(n_129), .Y(n_263) );
NAND2x1p5_ASAP7_75t_L g264 ( .A(n_189), .B(n_129), .Y(n_264) );
BUFx6f_ASAP7_75t_L g265 ( .A(n_182), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_211), .B(n_168), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_211), .B(n_127), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_176), .Y(n_268) );
OAI22xp5_ASAP7_75t_SL g269 ( .A1(n_229), .A2(n_121), .B1(n_145), .B2(n_155), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_173), .B(n_158), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_176), .Y(n_271) );
BUFx4f_ASAP7_75t_SL g272 ( .A(n_178), .Y(n_272) );
INVx2_ASAP7_75t_SL g273 ( .A(n_176), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_201), .Y(n_274) );
INVx2_ASAP7_75t_L g275 ( .A(n_171), .Y(n_275) );
INVx2_ASAP7_75t_L g276 ( .A(n_171), .Y(n_276) );
AOI22xp33_ASAP7_75t_L g277 ( .A1(n_173), .A2(n_158), .B1(n_156), .B2(n_155), .Y(n_277) );
NOR2xp33_ASAP7_75t_L g278 ( .A(n_216), .B(n_145), .Y(n_278) );
INVxp67_ASAP7_75t_L g279 ( .A(n_215), .Y(n_279) );
INVx2_ASAP7_75t_L g280 ( .A(n_175), .Y(n_280) );
NOR2xp33_ASAP7_75t_L g281 ( .A(n_216), .B(n_156), .Y(n_281) );
NOR2xp33_ASAP7_75t_L g282 ( .A(n_216), .B(n_49), .Y(n_282) );
INVxp67_ASAP7_75t_SL g283 ( .A(n_213), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_213), .Y(n_284) );
INVx2_ASAP7_75t_L g285 ( .A(n_175), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_217), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_217), .Y(n_287) );
INVxp67_ASAP7_75t_L g288 ( .A(n_209), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_219), .Y(n_289) );
A2O1A1Ixp33_ASAP7_75t_L g290 ( .A1(n_219), .A2(n_228), .B(n_172), .C(n_198), .Y(n_290) );
NAND2xp5_ASAP7_75t_SL g291 ( .A(n_219), .B(n_159), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_219), .Y(n_292) );
OAI22xp5_ASAP7_75t_L g293 ( .A1(n_196), .A2(n_159), .B1(n_153), .B2(n_13), .Y(n_293) );
INVx2_ASAP7_75t_L g294 ( .A(n_177), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_169), .Y(n_295) );
INVx2_ASAP7_75t_SL g296 ( .A(n_173), .Y(n_296) );
AND2x2_ASAP7_75t_L g297 ( .A(n_173), .B(n_9), .Y(n_297) );
AOI22xp33_ASAP7_75t_L g298 ( .A1(n_173), .A2(n_153), .B1(n_159), .B2(n_14), .Y(n_298) );
HB1xp67_ASAP7_75t_L g299 ( .A(n_187), .Y(n_299) );
BUFx3_ASAP7_75t_L g300 ( .A(n_232), .Y(n_300) );
BUFx6f_ASAP7_75t_L g301 ( .A(n_247), .Y(n_301) );
AND2x2_ASAP7_75t_L g302 ( .A(n_246), .B(n_229), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_259), .Y(n_303) );
BUFx6f_ASAP7_75t_L g304 ( .A(n_247), .Y(n_304) );
OAI22xp5_ASAP7_75t_L g305 ( .A1(n_283), .A2(n_205), .B1(n_172), .B2(n_200), .Y(n_305) );
NOR2xp33_ASAP7_75t_SL g306 ( .A(n_254), .B(n_253), .Y(n_306) );
AOI22xp5_ASAP7_75t_L g307 ( .A1(n_252), .A2(n_231), .B1(n_220), .B2(n_218), .Y(n_307) );
INVx2_ASAP7_75t_L g308 ( .A(n_236), .Y(n_308) );
INVx2_ASAP7_75t_L g309 ( .A(n_236), .Y(n_309) );
O2A1O1Ixp5_ASAP7_75t_L g310 ( .A1(n_267), .A2(n_198), .B(n_185), .C(n_188), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_237), .B(n_187), .Y(n_311) );
OAI22xp5_ASAP7_75t_L g312 ( .A1(n_241), .A2(n_199), .B1(n_179), .B2(n_185), .Y(n_312) );
CKINVDCx5p33_ASAP7_75t_R g313 ( .A(n_244), .Y(n_313) );
AND2x2_ASAP7_75t_SL g314 ( .A(n_239), .B(n_199), .Y(n_314) );
A2O1A1Ixp33_ASAP7_75t_L g315 ( .A1(n_238), .A2(n_169), .B(n_188), .C(n_200), .Y(n_315) );
NOR2xp33_ASAP7_75t_L g316 ( .A(n_249), .B(n_212), .Y(n_316) );
BUFx6f_ASAP7_75t_L g317 ( .A(n_247), .Y(n_317) );
A2O1A1Ixp33_ASAP7_75t_L g318 ( .A1(n_290), .A2(n_179), .B(n_194), .C(n_182), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_268), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_271), .Y(n_320) );
AND2x4_ASAP7_75t_L g321 ( .A(n_239), .B(n_193), .Y(n_321) );
INVx2_ASAP7_75t_L g322 ( .A(n_236), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_237), .B(n_194), .Y(n_323) );
BUFx2_ASAP7_75t_L g324 ( .A(n_244), .Y(n_324) );
OAI22xp5_ASAP7_75t_L g325 ( .A1(n_273), .A2(n_212), .B1(n_206), .B2(n_224), .Y(n_325) );
OR2x6_ASAP7_75t_L g326 ( .A(n_253), .B(n_193), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_263), .Y(n_327) );
BUFx3_ASAP7_75t_L g328 ( .A(n_263), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_263), .Y(n_329) );
NAND2xp5_ASAP7_75t_SL g330 ( .A(n_247), .B(n_206), .Y(n_330) );
A2O1A1Ixp33_ASAP7_75t_SL g331 ( .A1(n_251), .A2(n_208), .B(n_227), .C(n_197), .Y(n_331) );
A2O1A1Ixp33_ASAP7_75t_L g332 ( .A1(n_290), .A2(n_224), .B(n_222), .C(n_226), .Y(n_332) );
INVx2_ASAP7_75t_L g333 ( .A(n_265), .Y(n_333) );
BUFx12f_ASAP7_75t_L g334 ( .A(n_256), .Y(n_334) );
INVx2_ASAP7_75t_L g335 ( .A(n_265), .Y(n_335) );
A2O1A1Ixp33_ASAP7_75t_L g336 ( .A1(n_241), .A2(n_222), .B(n_223), .C(n_226), .Y(n_336) );
O2A1O1Ixp5_ASAP7_75t_SL g337 ( .A1(n_291), .A2(n_225), .B(n_223), .C(n_153), .Y(n_337) );
BUFx6f_ASAP7_75t_L g338 ( .A(n_247), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_250), .B(n_192), .Y(n_339) );
INVx4_ASAP7_75t_L g340 ( .A(n_254), .Y(n_340) );
INVxp67_ASAP7_75t_L g341 ( .A(n_260), .Y(n_341) );
OAI21xp33_ASAP7_75t_L g342 ( .A1(n_248), .A2(n_250), .B(n_245), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_266), .B(n_192), .Y(n_343) );
INVx2_ASAP7_75t_L g344 ( .A(n_265), .Y(n_344) );
OR2x6_ASAP7_75t_L g345 ( .A(n_279), .B(n_208), .Y(n_345) );
NOR3xp33_ASAP7_75t_L g346 ( .A(n_240), .B(n_225), .C(n_177), .Y(n_346) );
AOI21xp5_ASAP7_75t_L g347 ( .A1(n_262), .A2(n_197), .B(n_227), .Y(n_347) );
NOR2xp33_ASAP7_75t_L g348 ( .A(n_288), .B(n_192), .Y(n_348) );
O2A1O1Ixp33_ASAP7_75t_L g349 ( .A1(n_274), .A2(n_191), .B(n_183), .C(n_192), .Y(n_349) );
CKINVDCx20_ASAP7_75t_R g350 ( .A(n_272), .Y(n_350) );
BUFx5_ASAP7_75t_L g351 ( .A(n_258), .Y(n_351) );
CKINVDCx16_ASAP7_75t_R g352 ( .A(n_300), .Y(n_352) );
HB1xp67_ASAP7_75t_L g353 ( .A(n_324), .Y(n_353) );
INVxp67_ASAP7_75t_SL g354 ( .A(n_314), .Y(n_354) );
OAI21x1_ASAP7_75t_L g355 ( .A1(n_337), .A2(n_264), .B(n_282), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_323), .Y(n_356) );
NOR2xp33_ASAP7_75t_L g357 ( .A(n_302), .B(n_299), .Y(n_357) );
OAI21xp5_ASAP7_75t_L g358 ( .A1(n_310), .A2(n_270), .B(n_292), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_342), .B(n_297), .Y(n_359) );
AND2x4_ASAP7_75t_L g360 ( .A(n_327), .B(n_254), .Y(n_360) );
AND2x6_ASAP7_75t_L g361 ( .A(n_301), .B(n_304), .Y(n_361) );
AOI22xp5_ASAP7_75t_L g362 ( .A1(n_313), .A2(n_269), .B1(n_297), .B2(n_273), .Y(n_362) );
AND2x4_ASAP7_75t_L g363 ( .A(n_329), .B(n_254), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_328), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_311), .Y(n_365) );
AOI221xp5_ASAP7_75t_L g366 ( .A1(n_341), .A2(n_284), .B1(n_286), .B2(n_287), .C(n_281), .Y(n_366) );
OAI21x1_ASAP7_75t_L g367 ( .A1(n_312), .A2(n_264), .B(n_291), .Y(n_367) );
AND2x2_ASAP7_75t_L g368 ( .A(n_342), .B(n_295), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_303), .B(n_255), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_319), .Y(n_370) );
INVxp67_ASAP7_75t_SL g371 ( .A(n_301), .Y(n_371) );
OAI21x1_ASAP7_75t_SL g372 ( .A1(n_312), .A2(n_296), .B(n_277), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_320), .Y(n_373) );
OA21x2_ASAP7_75t_L g374 ( .A1(n_318), .A2(n_332), .B(n_315), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_321), .Y(n_375) );
AOI21xp33_ASAP7_75t_L g376 ( .A1(n_348), .A2(n_296), .B(n_243), .Y(n_376) );
OAI21x1_ASAP7_75t_SL g377 ( .A1(n_340), .A2(n_298), .B(n_234), .Y(n_377) );
XNOR2xp5_ASAP7_75t_L g378 ( .A(n_350), .B(n_242), .Y(n_378) );
AOI21x1_ASAP7_75t_L g379 ( .A1(n_325), .A2(n_257), .B(n_191), .Y(n_379) );
NAND3xp33_ASAP7_75t_L g380 ( .A(n_316), .B(n_293), .C(n_278), .Y(n_380) );
A2O1A1Ixp33_ASAP7_75t_L g381 ( .A1(n_336), .A2(n_289), .B(n_257), .C(n_261), .Y(n_381) );
INVx2_ASAP7_75t_L g382 ( .A(n_308), .Y(n_382) );
AO21x1_ASAP7_75t_L g383 ( .A1(n_305), .A2(n_183), .B(n_261), .Y(n_383) );
AOI22xp33_ASAP7_75t_L g384 ( .A1(n_357), .A2(n_346), .B1(n_334), .B2(n_321), .Y(n_384) );
INVxp33_ASAP7_75t_SL g385 ( .A(n_378), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_356), .Y(n_386) );
AOI21xp5_ASAP7_75t_L g387 ( .A1(n_381), .A2(n_331), .B(n_349), .Y(n_387) );
AO21x2_ASAP7_75t_L g388 ( .A1(n_383), .A2(n_372), .B(n_355), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_357), .B(n_307), .Y(n_389) );
INVx2_ASAP7_75t_L g390 ( .A(n_382), .Y(n_390) );
AOI22xp5_ASAP7_75t_SL g391 ( .A1(n_378), .A2(n_301), .B1(n_304), .B2(n_317), .Y(n_391) );
INVx2_ASAP7_75t_L g392 ( .A(n_382), .Y(n_392) );
INVx2_ASAP7_75t_L g393 ( .A(n_370), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_373), .Y(n_394) );
AOI222xp33_ASAP7_75t_L g395 ( .A1(n_365), .A2(n_305), .B1(n_339), .B2(n_343), .C1(n_262), .C2(n_322), .Y(n_395) );
OAI221xp5_ASAP7_75t_L g396 ( .A1(n_362), .A2(n_307), .B1(n_345), .B2(n_326), .C(n_309), .Y(n_396) );
OAI22xp33_ASAP7_75t_L g397 ( .A1(n_352), .A2(n_345), .B1(n_306), .B2(n_254), .Y(n_397) );
AOI21xp33_ASAP7_75t_L g398 ( .A1(n_380), .A2(n_345), .B(n_326), .Y(n_398) );
INVx2_ASAP7_75t_L g399 ( .A(n_374), .Y(n_399) );
OAI21xp5_ASAP7_75t_L g400 ( .A1(n_381), .A2(n_330), .B(n_347), .Y(n_400) );
AND2x4_ASAP7_75t_L g401 ( .A(n_360), .B(n_340), .Y(n_401) );
AOI21xp5_ASAP7_75t_L g402 ( .A1(n_355), .A2(n_306), .B(n_344), .Y(n_402) );
OAI22xp5_ASAP7_75t_SL g403 ( .A1(n_354), .A2(n_326), .B1(n_304), .B2(n_317), .Y(n_403) );
OAI321xp33_ASAP7_75t_L g404 ( .A1(n_359), .A2(n_159), .A3(n_317), .B1(n_338), .B2(n_333), .C(n_335), .Y(n_404) );
OR2x6_ASAP7_75t_L g405 ( .A(n_375), .B(n_338), .Y(n_405) );
OAI211xp5_ASAP7_75t_L g406 ( .A1(n_353), .A2(n_203), .B(n_159), .C(n_338), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_368), .Y(n_407) );
AOI221xp5_ASAP7_75t_L g408 ( .A1(n_366), .A2(n_265), .B1(n_258), .B2(n_235), .C(n_233), .Y(n_408) );
AOI221xp5_ASAP7_75t_L g409 ( .A1(n_369), .A2(n_280), .B1(n_233), .B2(n_235), .C(n_275), .Y(n_409) );
OAI22xp5_ASAP7_75t_L g410 ( .A1(n_368), .A2(n_351), .B1(n_203), .B2(n_285), .Y(n_410) );
BUFx2_ASAP7_75t_L g411 ( .A(n_361), .Y(n_411) );
INVx4_ASAP7_75t_L g412 ( .A(n_411), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_407), .Y(n_413) );
AND2x2_ASAP7_75t_L g414 ( .A(n_407), .B(n_374), .Y(n_414) );
INVx2_ASAP7_75t_L g415 ( .A(n_399), .Y(n_415) );
INVx2_ASAP7_75t_L g416 ( .A(n_399), .Y(n_416) );
AND2x2_ASAP7_75t_L g417 ( .A(n_390), .B(n_374), .Y(n_417) );
INVx2_ASAP7_75t_SL g418 ( .A(n_411), .Y(n_418) );
INVx3_ASAP7_75t_L g419 ( .A(n_401), .Y(n_419) );
AND2x2_ASAP7_75t_L g420 ( .A(n_390), .B(n_383), .Y(n_420) );
AND2x2_ASAP7_75t_L g421 ( .A(n_392), .B(n_367), .Y(n_421) );
INVx2_ASAP7_75t_L g422 ( .A(n_392), .Y(n_422) );
INVx2_ASAP7_75t_L g423 ( .A(n_388), .Y(n_423) );
AND2x2_ASAP7_75t_L g424 ( .A(n_393), .B(n_367), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_393), .Y(n_425) );
AND2x2_ASAP7_75t_L g426 ( .A(n_386), .B(n_371), .Y(n_426) );
INVx2_ASAP7_75t_SL g427 ( .A(n_391), .Y(n_427) );
INVx2_ASAP7_75t_L g428 ( .A(n_388), .Y(n_428) );
AOI22xp5_ASAP7_75t_L g429 ( .A1(n_389), .A2(n_364), .B1(n_376), .B2(n_360), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_386), .Y(n_430) );
NAND2xp5_ASAP7_75t_SL g431 ( .A(n_404), .B(n_351), .Y(n_431) );
AO21x2_ASAP7_75t_L g432 ( .A1(n_387), .A2(n_377), .B(n_379), .Y(n_432) );
NAND2x1p5_ASAP7_75t_L g433 ( .A(n_401), .B(n_363), .Y(n_433) );
BUFx2_ASAP7_75t_L g434 ( .A(n_403), .Y(n_434) );
INVx2_ASAP7_75t_L g435 ( .A(n_388), .Y(n_435) );
OR2x2_ASAP7_75t_L g436 ( .A(n_394), .B(n_358), .Y(n_436) );
AND2x4_ASAP7_75t_L g437 ( .A(n_405), .B(n_401), .Y(n_437) );
HB1xp67_ASAP7_75t_L g438 ( .A(n_405), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_395), .B(n_361), .Y(n_439) );
BUFx3_ASAP7_75t_L g440 ( .A(n_405), .Y(n_440) );
AND2x2_ASAP7_75t_L g441 ( .A(n_400), .B(n_361), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_405), .B(n_361), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_384), .B(n_361), .Y(n_443) );
OAI22xp5_ASAP7_75t_L g444 ( .A1(n_396), .A2(n_363), .B1(n_360), .B2(n_361), .Y(n_444) );
CKINVDCx5p33_ASAP7_75t_R g445 ( .A(n_385), .Y(n_445) );
INVx4_ASAP7_75t_L g446 ( .A(n_397), .Y(n_446) );
AND2x2_ASAP7_75t_L g447 ( .A(n_398), .B(n_363), .Y(n_447) );
OR2x2_ASAP7_75t_L g448 ( .A(n_425), .B(n_410), .Y(n_448) );
INVx2_ASAP7_75t_L g449 ( .A(n_415), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_413), .B(n_402), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_413), .Y(n_451) );
AOI22xp33_ASAP7_75t_L g452 ( .A1(n_446), .A2(n_385), .B1(n_408), .B2(n_351), .Y(n_452) );
AND2x2_ASAP7_75t_L g453 ( .A(n_414), .B(n_10), .Y(n_453) );
AO21x2_ASAP7_75t_L g454 ( .A1(n_432), .A2(n_406), .B(n_280), .Y(n_454) );
OR2x2_ASAP7_75t_L g455 ( .A(n_425), .B(n_10), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_424), .Y(n_456) );
OR2x2_ASAP7_75t_L g457 ( .A(n_430), .B(n_13), .Y(n_457) );
CKINVDCx20_ASAP7_75t_R g458 ( .A(n_445), .Y(n_458) );
BUFx2_ASAP7_75t_SL g459 ( .A(n_427), .Y(n_459) );
AOI22xp33_ASAP7_75t_L g460 ( .A1(n_446), .A2(n_351), .B1(n_409), .B2(n_203), .Y(n_460) );
AND2x2_ASAP7_75t_L g461 ( .A(n_414), .B(n_15), .Y(n_461) );
INVx1_ASAP7_75t_SL g462 ( .A(n_426), .Y(n_462) );
AOI22xp33_ASAP7_75t_L g463 ( .A1(n_446), .A2(n_351), .B1(n_203), .B2(n_285), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_430), .B(n_16), .Y(n_464) );
NAND4xp25_ASAP7_75t_L g465 ( .A(n_429), .B(n_17), .C(n_294), .D(n_276), .Y(n_465) );
INVx1_ASAP7_75t_SL g466 ( .A(n_426), .Y(n_466) );
AND2x2_ASAP7_75t_L g467 ( .A(n_414), .B(n_17), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_424), .B(n_18), .Y(n_468) );
AND2x2_ASAP7_75t_L g469 ( .A(n_424), .B(n_22), .Y(n_469) );
INVx2_ASAP7_75t_L g470 ( .A(n_415), .Y(n_470) );
OR2x2_ASAP7_75t_L g471 ( .A(n_436), .B(n_203), .Y(n_471) );
INVx2_ASAP7_75t_SL g472 ( .A(n_437), .Y(n_472) );
HB1xp67_ASAP7_75t_L g473 ( .A(n_426), .Y(n_473) );
AND2x2_ASAP7_75t_L g474 ( .A(n_420), .B(n_25), .Y(n_474) );
AND2x2_ASAP7_75t_L g475 ( .A(n_420), .B(n_26), .Y(n_475) );
AND2x2_ASAP7_75t_L g476 ( .A(n_420), .B(n_32), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_415), .Y(n_477) );
OAI21xp33_ASAP7_75t_L g478 ( .A1(n_427), .A2(n_294), .B(n_276), .Y(n_478) );
NOR2x1_ASAP7_75t_L g479 ( .A(n_434), .B(n_275), .Y(n_479) );
AND2x2_ASAP7_75t_L g480 ( .A(n_422), .B(n_35), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_416), .Y(n_481) );
INVxp67_ASAP7_75t_SL g482 ( .A(n_422), .Y(n_482) );
INVxp67_ASAP7_75t_L g483 ( .A(n_434), .Y(n_483) );
AND2x2_ASAP7_75t_L g484 ( .A(n_422), .B(n_39), .Y(n_484) );
INVx2_ASAP7_75t_L g485 ( .A(n_416), .Y(n_485) );
INVxp67_ASAP7_75t_L g486 ( .A(n_438), .Y(n_486) );
INVx3_ASAP7_75t_L g487 ( .A(n_412), .Y(n_487) );
HB1xp67_ASAP7_75t_L g488 ( .A(n_419), .Y(n_488) );
AOI22xp33_ASAP7_75t_SL g489 ( .A1(n_446), .A2(n_203), .B1(n_221), .B2(n_230), .Y(n_489) );
HB1xp67_ASAP7_75t_L g490 ( .A(n_419), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_416), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_421), .Y(n_492) );
INVxp67_ASAP7_75t_L g493 ( .A(n_438), .Y(n_493) );
OAI31xp33_ASAP7_75t_L g494 ( .A1(n_444), .A2(n_41), .A3(n_46), .B(n_50), .Y(n_494) );
INVx2_ASAP7_75t_L g495 ( .A(n_421), .Y(n_495) );
INVx2_ASAP7_75t_L g496 ( .A(n_421), .Y(n_496) );
OR2x6_ASAP7_75t_SL g497 ( .A(n_444), .B(n_51), .Y(n_497) );
OR2x2_ASAP7_75t_L g498 ( .A(n_436), .B(n_53), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_473), .B(n_436), .Y(n_499) );
INVx2_ASAP7_75t_L g500 ( .A(n_449), .Y(n_500) );
AND2x2_ASAP7_75t_L g501 ( .A(n_456), .B(n_417), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_451), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_462), .B(n_429), .Y(n_503) );
OR2x2_ASAP7_75t_L g504 ( .A(n_462), .B(n_418), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_451), .Y(n_505) );
BUFx12f_ASAP7_75t_L g506 ( .A(n_457), .Y(n_506) );
OR2x2_ASAP7_75t_L g507 ( .A(n_466), .B(n_418), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_466), .B(n_447), .Y(n_508) );
AND2x4_ASAP7_75t_L g509 ( .A(n_472), .B(n_441), .Y(n_509) );
AND2x4_ASAP7_75t_L g510 ( .A(n_472), .B(n_441), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_455), .Y(n_511) );
AND2x2_ASAP7_75t_L g512 ( .A(n_456), .B(n_417), .Y(n_512) );
OR2x6_ASAP7_75t_L g513 ( .A(n_459), .B(n_427), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_453), .B(n_447), .Y(n_514) );
AOI21xp33_ASAP7_75t_L g515 ( .A1(n_479), .A2(n_443), .B(n_439), .Y(n_515) );
BUFx2_ASAP7_75t_L g516 ( .A(n_487), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_455), .Y(n_517) );
AND2x2_ASAP7_75t_L g518 ( .A(n_492), .B(n_417), .Y(n_518) );
AND2x2_ASAP7_75t_L g519 ( .A(n_453), .B(n_447), .Y(n_519) );
AND2x2_ASAP7_75t_L g520 ( .A(n_461), .B(n_419), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_461), .B(n_419), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_467), .Y(n_522) );
OR2x2_ASAP7_75t_L g523 ( .A(n_471), .B(n_418), .Y(n_523) );
OR2x2_ASAP7_75t_L g524 ( .A(n_471), .B(n_412), .Y(n_524) );
AND2x2_ASAP7_75t_L g525 ( .A(n_492), .B(n_435), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_467), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_457), .Y(n_527) );
OAI31xp33_ASAP7_75t_SL g528 ( .A1(n_465), .A2(n_437), .A3(n_442), .B(n_431), .Y(n_528) );
NAND2xp5_ASAP7_75t_SL g529 ( .A(n_478), .B(n_446), .Y(n_529) );
AND2x2_ASAP7_75t_L g530 ( .A(n_495), .B(n_435), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_483), .B(n_419), .Y(n_531) );
OR2x2_ASAP7_75t_L g532 ( .A(n_477), .B(n_412), .Y(n_532) );
INVx2_ASAP7_75t_L g533 ( .A(n_449), .Y(n_533) );
AND2x2_ASAP7_75t_L g534 ( .A(n_495), .B(n_423), .Y(n_534) );
AND2x2_ASAP7_75t_L g535 ( .A(n_495), .B(n_423), .Y(n_535) );
AND2x2_ASAP7_75t_L g536 ( .A(n_496), .B(n_423), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_496), .B(n_437), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_496), .B(n_437), .Y(n_538) );
AND2x2_ASAP7_75t_L g539 ( .A(n_477), .B(n_435), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_464), .B(n_437), .Y(n_540) );
AND2x2_ASAP7_75t_L g541 ( .A(n_481), .B(n_428), .Y(n_541) );
AND2x4_ASAP7_75t_L g542 ( .A(n_487), .B(n_441), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_481), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_491), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_491), .B(n_443), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_474), .B(n_440), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_474), .B(n_440), .Y(n_547) );
OAI21xp33_ASAP7_75t_L g548 ( .A1(n_465), .A2(n_439), .B(n_428), .Y(n_548) );
OR2x2_ASAP7_75t_L g549 ( .A(n_482), .B(n_412), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_486), .Y(n_550) );
AOI33xp33_ASAP7_75t_L g551 ( .A1(n_452), .A2(n_428), .A3(n_442), .B1(n_412), .B2(n_433), .B3(n_432), .Y(n_551) );
INVx1_ASAP7_75t_SL g552 ( .A(n_458), .Y(n_552) );
NOR2xp33_ASAP7_75t_L g553 ( .A(n_493), .B(n_440), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_475), .B(n_442), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_449), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_470), .Y(n_556) );
AND2x2_ASAP7_75t_L g557 ( .A(n_470), .B(n_432), .Y(n_557) );
BUFx3_ASAP7_75t_L g558 ( .A(n_552), .Y(n_558) );
OR2x2_ASAP7_75t_L g559 ( .A(n_508), .B(n_470), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_502), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_505), .Y(n_561) );
AOI21xp5_ASAP7_75t_L g562 ( .A1(n_528), .A2(n_431), .B(n_478), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_550), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_543), .Y(n_564) );
AND2x4_ASAP7_75t_L g565 ( .A(n_513), .B(n_487), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_501), .B(n_450), .Y(n_566) );
AND2x2_ASAP7_75t_L g567 ( .A(n_519), .B(n_487), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_544), .Y(n_568) );
NOR2xp33_ASAP7_75t_L g569 ( .A(n_506), .B(n_459), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_501), .B(n_450), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_527), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_512), .B(n_485), .Y(n_572) );
INVx2_ASAP7_75t_L g573 ( .A(n_500), .Y(n_573) );
NOR2xp33_ASAP7_75t_L g574 ( .A(n_506), .B(n_497), .Y(n_574) );
OR2x2_ASAP7_75t_L g575 ( .A(n_499), .B(n_485), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_511), .Y(n_576) );
NOR2xp33_ASAP7_75t_L g577 ( .A(n_531), .B(n_497), .Y(n_577) );
NOR2xp33_ASAP7_75t_SL g578 ( .A(n_513), .B(n_494), .Y(n_578) );
AND2x2_ASAP7_75t_L g579 ( .A(n_520), .B(n_490), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_512), .B(n_485), .Y(n_580) );
OR2x2_ASAP7_75t_L g581 ( .A(n_514), .B(n_488), .Y(n_581) );
AND2x2_ASAP7_75t_L g582 ( .A(n_518), .B(n_468), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_517), .Y(n_583) );
AND2x2_ASAP7_75t_L g584 ( .A(n_518), .B(n_468), .Y(n_584) );
INVx2_ASAP7_75t_L g585 ( .A(n_500), .Y(n_585) );
OR2x2_ASAP7_75t_L g586 ( .A(n_522), .B(n_448), .Y(n_586) );
OR2x2_ASAP7_75t_L g587 ( .A(n_526), .B(n_448), .Y(n_587) );
INVx1_ASAP7_75t_SL g588 ( .A(n_549), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_525), .B(n_479), .Y(n_589) );
HB1xp67_ASAP7_75t_L g590 ( .A(n_533), .Y(n_590) );
BUFx3_ASAP7_75t_L g591 ( .A(n_516), .Y(n_591) );
OR2x2_ASAP7_75t_L g592 ( .A(n_524), .B(n_469), .Y(n_592) );
NAND4xp25_ASAP7_75t_L g593 ( .A(n_551), .B(n_494), .C(n_475), .D(n_476), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_537), .Y(n_594) );
NOR2xp33_ASAP7_75t_L g595 ( .A(n_548), .B(n_498), .Y(n_595) );
INVx3_ASAP7_75t_SL g596 ( .A(n_513), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_525), .B(n_476), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_538), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_545), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_557), .B(n_432), .Y(n_600) );
AND2x2_ASAP7_75t_L g601 ( .A(n_509), .B(n_469), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_532), .Y(n_602) );
AND2x4_ASAP7_75t_SL g603 ( .A(n_542), .B(n_484), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_555), .Y(n_604) );
AND2x2_ASAP7_75t_L g605 ( .A(n_509), .B(n_454), .Y(n_605) );
INVx2_ASAP7_75t_L g606 ( .A(n_533), .Y(n_606) );
OR2x2_ASAP7_75t_L g607 ( .A(n_521), .B(n_498), .Y(n_607) );
OR2x2_ASAP7_75t_L g608 ( .A(n_504), .B(n_432), .Y(n_608) );
AND2x2_ASAP7_75t_SL g609 ( .A(n_551), .B(n_484), .Y(n_609) );
OAI21xp5_ASAP7_75t_SL g610 ( .A1(n_574), .A2(n_529), .B(n_503), .Y(n_610) );
AND2x4_ASAP7_75t_L g611 ( .A(n_591), .B(n_542), .Y(n_611) );
NAND2xp5_ASAP7_75t_SL g612 ( .A(n_578), .B(n_529), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_563), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_560), .Y(n_614) );
AOI22xp5_ASAP7_75t_L g615 ( .A1(n_577), .A2(n_553), .B1(n_509), .B2(n_510), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_594), .B(n_557), .Y(n_616) );
OR2x2_ASAP7_75t_L g617 ( .A(n_566), .B(n_507), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_598), .B(n_535), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_561), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_571), .Y(n_620) );
OAI22xp5_ASAP7_75t_L g621 ( .A1(n_574), .A2(n_554), .B1(n_546), .B2(n_547), .Y(n_621) );
AOI21xp5_ASAP7_75t_L g622 ( .A1(n_562), .A2(n_489), .B(n_454), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_576), .Y(n_623) );
NAND2xp33_ASAP7_75t_L g624 ( .A(n_596), .B(n_523), .Y(n_624) );
OAI22xp33_ASAP7_75t_L g625 ( .A1(n_593), .A2(n_540), .B1(n_542), .B2(n_553), .Y(n_625) );
INVxp67_ASAP7_75t_L g626 ( .A(n_558), .Y(n_626) );
A2O1A1Ixp33_ASAP7_75t_L g627 ( .A1(n_569), .A2(n_515), .B(n_510), .C(n_480), .Y(n_627) );
INVxp67_ASAP7_75t_L g628 ( .A(n_590), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_599), .B(n_530), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_583), .Y(n_630) );
AOI322xp5_ASAP7_75t_L g631 ( .A1(n_577), .A2(n_510), .A3(n_536), .B1(n_535), .B2(n_534), .C1(n_530), .C2(n_541), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_564), .Y(n_632) );
AOI22xp33_ASAP7_75t_L g633 ( .A1(n_609), .A2(n_536), .B1(n_534), .B2(n_433), .Y(n_633) );
INVx1_ASAP7_75t_L g634 ( .A(n_568), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_566), .B(n_541), .Y(n_635) );
OAI21xp5_ASAP7_75t_L g636 ( .A1(n_562), .A2(n_480), .B(n_460), .Y(n_636) );
NAND2xp5_ASAP7_75t_SL g637 ( .A(n_596), .B(n_556), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_575), .Y(n_638) );
OAI21xp5_ASAP7_75t_L g639 ( .A1(n_609), .A2(n_433), .B(n_463), .Y(n_639) );
INVx1_ASAP7_75t_SL g640 ( .A(n_588), .Y(n_640) );
O2A1O1Ixp33_ASAP7_75t_SL g641 ( .A1(n_595), .A2(n_433), .B(n_454), .C(n_539), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_572), .Y(n_642) );
AOI21xp33_ASAP7_75t_L g643 ( .A1(n_595), .A2(n_539), .B(n_58), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_572), .Y(n_644) );
OAI22xp5_ASAP7_75t_L g645 ( .A1(n_592), .A2(n_230), .B1(n_221), .B2(n_60), .Y(n_645) );
NOR2xp33_ASAP7_75t_L g646 ( .A(n_586), .B(n_54), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_614), .Y(n_647) );
INVxp67_ASAP7_75t_L g648 ( .A(n_640), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_619), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_632), .Y(n_650) );
AOI211xp5_ASAP7_75t_L g651 ( .A1(n_625), .A2(n_565), .B(n_605), .C(n_608), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_634), .Y(n_652) );
INVxp67_ASAP7_75t_SL g653 ( .A(n_628), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_631), .B(n_602), .Y(n_654) );
O2A1O1Ixp33_ASAP7_75t_L g655 ( .A1(n_612), .A2(n_600), .B(n_587), .C(n_570), .Y(n_655) );
AOI22xp5_ASAP7_75t_L g656 ( .A1(n_610), .A2(n_570), .B1(n_567), .B2(n_579), .Y(n_656) );
O2A1O1Ixp33_ASAP7_75t_L g657 ( .A1(n_626), .A2(n_600), .B(n_589), .C(n_581), .Y(n_657) );
NAND3x2_ASAP7_75t_L g658 ( .A(n_611), .B(n_565), .C(n_601), .Y(n_658) );
INVx1_ASAP7_75t_L g659 ( .A(n_617), .Y(n_659) );
AND2x2_ASAP7_75t_L g660 ( .A(n_638), .B(n_582), .Y(n_660) );
NOR2x1_ASAP7_75t_L g661 ( .A(n_624), .B(n_604), .Y(n_661) );
INVx1_ASAP7_75t_SL g662 ( .A(n_611), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_642), .B(n_580), .Y(n_663) );
INVx1_ASAP7_75t_L g664 ( .A(n_613), .Y(n_664) );
OAI22xp5_ASAP7_75t_L g665 ( .A1(n_633), .A2(n_597), .B1(n_603), .B2(n_580), .Y(n_665) );
INVxp67_ASAP7_75t_L g666 ( .A(n_620), .Y(n_666) );
NAND2xp33_ASAP7_75t_L g667 ( .A(n_639), .B(n_584), .Y(n_667) );
INVx1_ASAP7_75t_L g668 ( .A(n_623), .Y(n_668) );
AOI22xp33_ASAP7_75t_SL g669 ( .A1(n_621), .A2(n_597), .B1(n_589), .B2(n_607), .Y(n_669) );
XNOR2xp5_ASAP7_75t_L g670 ( .A(n_658), .B(n_651), .Y(n_670) );
INVx2_ASAP7_75t_L g671 ( .A(n_647), .Y(n_671) );
INVx1_ASAP7_75t_L g672 ( .A(n_649), .Y(n_672) );
OAI221xp5_ASAP7_75t_L g673 ( .A1(n_667), .A2(n_615), .B1(n_627), .B2(n_637), .C(n_636), .Y(n_673) );
OAI22xp5_ASAP7_75t_L g674 ( .A1(n_661), .A2(n_628), .B1(n_635), .B2(n_629), .Y(n_674) );
AOI21xp5_ASAP7_75t_L g675 ( .A1(n_667), .A2(n_641), .B(n_622), .Y(n_675) );
AOI22xp33_ASAP7_75t_L g676 ( .A1(n_654), .A2(n_644), .B1(n_643), .B2(n_646), .Y(n_676) );
O2A1O1Ixp33_ASAP7_75t_L g677 ( .A1(n_648), .A2(n_622), .B(n_630), .C(n_645), .Y(n_677) );
OAI21xp5_ASAP7_75t_L g678 ( .A1(n_655), .A2(n_618), .B(n_590), .Y(n_678) );
INVx1_ASAP7_75t_L g679 ( .A(n_650), .Y(n_679) );
AOI22xp5_ASAP7_75t_L g680 ( .A1(n_669), .A2(n_616), .B1(n_559), .B2(n_585), .Y(n_680) );
AOI22xp5_ASAP7_75t_L g681 ( .A1(n_656), .A2(n_606), .B1(n_573), .B2(n_230), .Y(n_681) );
AOI211xp5_ASAP7_75t_L g682 ( .A1(n_665), .A2(n_230), .B(n_221), .C(n_67), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_657), .B(n_59), .Y(n_683) );
HB1xp67_ASAP7_75t_L g684 ( .A(n_671), .Y(n_684) );
INVx1_ASAP7_75t_SL g685 ( .A(n_683), .Y(n_685) );
AOI21xp5_ASAP7_75t_L g686 ( .A1(n_670), .A2(n_653), .B(n_662), .Y(n_686) );
XNOR2x1_ASAP7_75t_L g687 ( .A(n_674), .B(n_659), .Y(n_687) );
AOI22xp33_ASAP7_75t_L g688 ( .A1(n_673), .A2(n_660), .B1(n_653), .B2(n_666), .Y(n_688) );
INVx1_ASAP7_75t_L g689 ( .A(n_672), .Y(n_689) );
AOI221xp5_ASAP7_75t_L g690 ( .A1(n_675), .A2(n_668), .B1(n_664), .B2(n_652), .C(n_663), .Y(n_690) );
INVx1_ASAP7_75t_L g691 ( .A(n_679), .Y(n_691) );
AOI22xp5_ASAP7_75t_L g692 ( .A1(n_688), .A2(n_676), .B1(n_680), .B2(n_681), .Y(n_692) );
NOR4xp25_ASAP7_75t_L g693 ( .A(n_690), .B(n_677), .C(n_678), .D(n_660), .Y(n_693) );
INVx1_ASAP7_75t_L g694 ( .A(n_689), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_686), .B(n_678), .Y(n_695) );
AND3x4_ASAP7_75t_L g696 ( .A(n_693), .B(n_687), .C(n_685), .Y(n_696) );
NAND2xp5_ASAP7_75t_SL g697 ( .A(n_695), .B(n_684), .Y(n_697) );
AND2x4_ASAP7_75t_L g698 ( .A(n_694), .B(n_691), .Y(n_698) );
AND2x4_ASAP7_75t_L g699 ( .A(n_698), .B(n_692), .Y(n_699) );
AOI21xp5_ASAP7_75t_L g700 ( .A1(n_696), .A2(n_684), .B(n_682), .Y(n_700) );
INVx2_ASAP7_75t_L g701 ( .A(n_699), .Y(n_701) );
INVx1_ASAP7_75t_L g702 ( .A(n_701), .Y(n_702) );
OAI222xp33_ASAP7_75t_L g703 ( .A1(n_702), .A2(n_700), .B1(n_697), .B2(n_69), .C1(n_71), .C2(n_73), .Y(n_703) );
AOI22x1_ASAP7_75t_L g704 ( .A1(n_703), .A2(n_221), .B1(n_230), .B2(n_74), .Y(n_704) );
AOI31xp33_ASAP7_75t_L g705 ( .A1(n_704), .A2(n_63), .A3(n_68), .B(n_221), .Y(n_705) );
endmodule