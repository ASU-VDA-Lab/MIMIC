module fake_jpeg_5233_n_108 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_108);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_108;

wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_106;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx12f_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

INVx5_ASAP7_75t_L g12 ( 
.A(n_9),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_7),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_6),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_23),
.B(n_24),
.Y(n_31)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_13),
.B(n_0),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_25),
.B(n_27),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

CKINVDCx16_ASAP7_75t_R g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_29),
.B(n_17),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_20),
.Y(n_30)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_30),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_24),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_34),
.B(n_37),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_27),
.B(n_22),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_39),
.Y(n_50)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_38),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_23),
.B(n_22),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_35),
.B(n_16),
.Y(n_42)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

A2O1A1Ixp33_ASAP7_75t_L g43 ( 
.A1(n_36),
.A2(n_13),
.B(n_19),
.C(n_14),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_43),
.B(n_48),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_39),
.B(n_11),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_44),
.B(n_51),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_19),
.Y(n_45)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_40),
.A2(n_29),
.B1(n_14),
.B2(n_21),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_46),
.A2(n_52),
.B1(n_15),
.B2(n_40),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_31),
.B(n_21),
.Y(n_49)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_36),
.B(n_11),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_40),
.A2(n_29),
.B1(n_18),
.B2(n_15),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_31),
.Y(n_53)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_53),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_57),
.B(n_28),
.Y(n_75)
);

NOR2x1_ASAP7_75t_L g58 ( 
.A(n_43),
.B(n_50),
.Y(n_58)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_58),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_50),
.B(n_37),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_59),
.B(n_44),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_48),
.A2(n_32),
.B1(n_33),
.B2(n_26),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_61),
.B(n_62),
.C(n_46),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_50),
.A2(n_33),
.B1(n_28),
.B2(n_26),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_41),
.A2(n_32),
.B1(n_33),
.B2(n_9),
.Y(n_64)
);

AOI21xp5_ASAP7_75t_L g71 ( 
.A1(n_64),
.A2(n_51),
.B(n_47),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_66),
.B(n_70),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_67),
.A2(n_71),
.B1(n_75),
.B2(n_63),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_SL g69 ( 
.A1(n_59),
.A2(n_41),
.B(n_53),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_SL g80 ( 
.A1(n_69),
.A2(n_56),
.B(n_63),
.Y(n_80)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_62),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_54),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_72),
.B(n_73),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_60),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_56),
.B(n_47),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_74),
.B(n_65),
.Y(n_84)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_74),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_76),
.B(n_78),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_70),
.A2(n_67),
.B1(n_68),
.B2(n_57),
.Y(n_77)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_77),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_80),
.A2(n_71),
.B(n_11),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_66),
.B(n_58),
.C(n_55),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_82),
.B(n_83),
.C(n_32),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_69),
.B(n_61),
.C(n_65),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_84),
.B(n_79),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_85),
.B(n_87),
.C(n_83),
.Y(n_92)
);

INVx1_ASAP7_75t_SL g89 ( 
.A(n_81),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_89),
.B(n_82),
.Y(n_94)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_90),
.Y(n_93)
);

HB1xp67_ASAP7_75t_L g91 ( 
.A(n_88),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_91),
.B(n_94),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_92),
.B(n_87),
.C(n_89),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_86),
.A2(n_77),
.B1(n_1),
.B2(n_2),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_95),
.B(n_0),
.C(n_2),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_96),
.A2(n_98),
.B(n_8),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_91),
.A2(n_93),
.B(n_2),
.Y(n_98)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_99),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_100),
.B(n_3),
.Y(n_104)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_97),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_102),
.B(n_10),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_103),
.B(n_104),
.C(n_101),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_105),
.A2(n_3),
.B(n_4),
.Y(n_106)
);

OAI21x1_ASAP7_75t_L g107 ( 
.A1(n_106),
.A2(n_3),
.B(n_4),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_107),
.B(n_4),
.Y(n_108)
);


endmodule