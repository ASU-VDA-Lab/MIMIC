module fake_jpeg_13680_n_193 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_193);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_193;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_26),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_5),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_22),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_15),
.Y(n_52)
);

INVx11_ASAP7_75t_SL g53 ( 
.A(n_38),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_18),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_8),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_6),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_9),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_13),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_39),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_3),
.Y(n_63)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

BUFx16f_ASAP7_75t_L g65 ( 
.A(n_7),
.Y(n_65)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_16),
.Y(n_66)
);

BUFx2_ASAP7_75t_L g67 ( 
.A(n_37),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_35),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_28),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_14),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_17),
.Y(n_72)
);

BUFx2_ASAP7_75t_L g73 ( 
.A(n_34),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_10),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_7),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_42),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_60),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_77),
.Y(n_94)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_56),
.Y(n_78)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_78),
.Y(n_90)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_47),
.Y(n_79)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_79),
.Y(n_95)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_55),
.Y(n_80)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_80),
.Y(n_88)
);

BUFx12f_ASAP7_75t_L g81 ( 
.A(n_63),
.Y(n_81)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_81),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_60),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_82),
.Y(n_100)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_65),
.Y(n_83)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_83),
.Y(n_93)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_70),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_84),
.B(n_85),
.Y(n_91)
);

BUFx8_ASAP7_75t_L g85 ( 
.A(n_53),
.Y(n_85)
);

INVx3_ASAP7_75t_SL g86 ( 
.A(n_57),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_86),
.B(n_76),
.Y(n_92)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_81),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_87),
.Y(n_115)
);

AO22x1_ASAP7_75t_SL g89 ( 
.A1(n_78),
.A2(n_53),
.B1(n_58),
.B2(n_65),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_89),
.A2(n_54),
.B1(n_48),
.B2(n_64),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_92),
.B(n_66),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_84),
.A2(n_67),
.B1(n_73),
.B2(n_47),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_96),
.A2(n_97),
.B(n_102),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_81),
.A2(n_73),
.B1(n_67),
.B2(n_76),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_78),
.B(n_68),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_98),
.B(n_72),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_80),
.B(n_75),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_101),
.B(n_62),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_81),
.A2(n_50),
.B1(n_59),
.B2(n_51),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_95),
.Y(n_103)
);

INVxp67_ASAP7_75t_SL g131 ( 
.A(n_103),
.Y(n_131)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_88),
.Y(n_104)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_104),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_91),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_105),
.B(n_124),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_98),
.B(n_74),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_106),
.B(n_108),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_107),
.B(n_119),
.Y(n_125)
);

BUFx2_ASAP7_75t_L g109 ( 
.A(n_99),
.Y(n_109)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_109),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_101),
.B(n_69),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_110),
.B(n_117),
.Y(n_145)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_90),
.Y(n_111)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_111),
.Y(n_141)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_93),
.Y(n_112)
);

HB1xp67_ASAP7_75t_L g127 ( 
.A(n_112),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_114),
.B(n_118),
.Y(n_134)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_91),
.Y(n_116)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_116),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_89),
.B(n_0),
.Y(n_117)
);

BUFx2_ASAP7_75t_L g119 ( 
.A(n_94),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_100),
.A2(n_71),
.B1(n_61),
.B2(n_2),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_120),
.A2(n_119),
.B1(n_113),
.B2(n_123),
.Y(n_135)
);

INVx1_ASAP7_75t_SL g121 ( 
.A(n_92),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_121),
.B(n_123),
.Y(n_130)
);

INVx8_ASAP7_75t_L g122 ( 
.A(n_87),
.Y(n_122)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_122),
.Y(n_146)
);

BUFx2_ASAP7_75t_L g123 ( 
.A(n_95),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_88),
.B(n_71),
.C(n_52),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_106),
.B(n_0),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_132),
.B(n_133),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_114),
.B(n_1),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_135),
.B(n_23),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_109),
.A2(n_49),
.B(n_2),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_136),
.B(n_4),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_115),
.Y(n_137)
);

BUFx2_ASAP7_75t_L g161 ( 
.A(n_137),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_108),
.B(n_1),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_138),
.B(n_24),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_121),
.B(n_3),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_139),
.B(n_144),
.Y(n_156)
);

AND2x2_ASAP7_75t_SL g142 ( 
.A(n_116),
.B(n_30),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_142),
.B(n_4),
.C(n_5),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_114),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_134),
.A2(n_29),
.B1(n_46),
.B2(n_45),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_147),
.A2(n_158),
.B1(n_125),
.B2(n_146),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_148),
.B(n_163),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_149),
.B(n_157),
.Y(n_171)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_126),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_150),
.B(n_152),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_128),
.B(n_6),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_151),
.B(n_153),
.Y(n_168)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_141),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_143),
.B(n_8),
.Y(n_153)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_127),
.Y(n_155)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_155),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_145),
.B(n_9),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_129),
.A2(n_11),
.B1(n_12),
.B2(n_19),
.Y(n_158)
);

AO21x1_ASAP7_75t_L g159 ( 
.A1(n_134),
.A2(n_20),
.B(n_21),
.Y(n_159)
);

OAI21xp33_ASAP7_75t_SL g164 ( 
.A1(n_159),
.A2(n_162),
.B(n_131),
.Y(n_164)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_140),
.Y(n_160)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_160),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_164),
.A2(n_161),
.B1(n_27),
.B2(n_31),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_156),
.B(n_130),
.Y(n_167)
);

CKINVDCx14_ASAP7_75t_R g175 ( 
.A(n_167),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_147),
.B(n_142),
.C(n_139),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_169),
.B(n_170),
.C(n_161),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_159),
.B(n_130),
.Y(n_170)
);

OR2x2_ASAP7_75t_L g176 ( 
.A(n_172),
.B(n_154),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_176),
.B(n_177),
.Y(n_183)
);

FAx1_ASAP7_75t_L g177 ( 
.A(n_167),
.B(n_149),
.CI(n_125),
.CON(n_177),
.SN(n_177)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_165),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_178),
.B(n_180),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_179),
.B(n_181),
.C(n_166),
.Y(n_182)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_173),
.Y(n_181)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_182),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_185),
.B(n_175),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_186),
.B(n_183),
.Y(n_187)
);

A2O1A1Ixp33_ASAP7_75t_SL g188 ( 
.A1(n_187),
.A2(n_177),
.B(n_175),
.C(n_184),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_188),
.B(n_171),
.Y(n_189)
);

FAx1_ASAP7_75t_SL g190 ( 
.A(n_189),
.B(n_168),
.CI(n_174),
.CON(n_190),
.SN(n_190)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_190),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_191),
.B(n_190),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_192),
.B(n_25),
.Y(n_193)
);


endmodule