module fake_netlist_6_3367_n_11214 (n_992, n_1671, n_1, n_801, n_1613, n_1234, n_1458, n_1199, n_1674, n_741, n_1027, n_1351, n_625, n_1189, n_223, n_1212, n_226, n_208, n_68, n_726, n_2157, n_212, n_700, n_50, n_1307, n_2003, n_1038, n_578, n_1581, n_1003, n_365, n_168, n_1237, n_1061, n_1357, n_1853, n_77, n_783, n_1738, n_2243, n_798, n_188, n_1575, n_1854, n_1923, n_509, n_1342, n_245, n_1209, n_1348, n_1387, n_2260, n_677, n_1708, n_805, n_1151, n_396, n_1739, n_350, n_78, n_2051, n_1380, n_442, n_480, n_142, n_1402, n_1688, n_1691, n_1975, n_1009, n_1743, n_62, n_1930, n_1160, n_883, n_1238, n_1991, n_2179, n_1724, n_1032, n_1247, n_1547, n_1553, n_893, n_1099, n_1264, n_1192, n_471, n_1844, n_424, n_1700, n_1555, n_1415, n_2211, n_1370, n_1786, n_369, n_287, n_415, n_830, n_65, n_230, n_461, n_873, n_141, n_383, n_1285, n_1371, n_200, n_1985, n_447, n_2184, n_1803, n_1172, n_852, n_71, n_229, n_1590, n_1532, n_1393, n_1517, n_1867, n_1704, n_1078, n_250, n_544, n_1711, n_2247, n_1140, n_1444, n_1670, n_1603, n_1579, n_35, n_1263, n_2019, n_836, n_375, n_2074, n_522, n_2129, n_1261, n_945, n_1649, n_2018, n_2094, n_1903, n_1511, n_1143, n_1422, n_1232, n_1772, n_1572, n_616, n_658, n_1874, n_1119, n_2013, n_428, n_1433, n_1902, n_1842, n_1620, n_2044, n_1954, n_1735, n_1541, n_1300, n_641, n_822, n_693, n_1313, n_1056, n_2212, n_758, n_516, n_1455, n_1163, n_1180, n_2256, n_943, n_1798, n_1550, n_491, n_1591, n_42, n_772, n_1344, n_666, n_371, n_940, n_770, n_567, n_1781, n_1971, n_2058, n_2090, n_405, n_213, n_538, n_2173, n_2004, n_1106, n_886, n_1471, n_343, n_953, n_1094, n_1345, n_1820, n_494, n_539, n_493, n_155, n_2108, n_45, n_454, n_1421, n_1936, n_638, n_1404, n_1211, n_2124, n_381, n_887, n_1660, n_1961, n_112, n_1280, n_713, n_1400, n_126, n_1467, n_58, n_976, n_2155, n_224, n_48, n_1445, n_1526, n_1560, n_734, n_1088, n_1894, n_196, n_1231, n_1978, n_2085, n_917, n_574, n_9, n_907, n_6, n_1446, n_14, n_659, n_1815, n_2214, n_407, n_913, n_1658, n_808, n_867, n_1230, n_473, n_1193, n_1967, n_1054, n_559, n_1333, n_44, n_1648, n_1911, n_1956, n_163, n_1644, n_2011, n_1558, n_1732, n_281, n_551, n_699, n_1986, n_564, n_451, n_824, n_279, n_686, n_757, n_594, n_1641, n_2113, n_1918, n_2190, n_577, n_166, n_1843, n_619, n_1367, n_1336, n_521, n_572, n_395, n_813, n_1909, n_2080, n_1481, n_323, n_606, n_1441, n_818, n_1123, n_1309, n_92, n_2104, n_513, n_645, n_1381, n_331, n_1699, n_916, n_2093, n_483, n_102, n_2207, n_1970, n_608, n_261, n_2101, n_630, n_2059, n_32, n_2198, n_541, n_512, n_2073, n_121, n_433, n_792, n_476, n_2, n_1328, n_1957, n_219, n_1907, n_264, n_263, n_1162, n_860, n_1530, n_788, n_939, n_1543, n_821, n_938, n_1302, n_1068, n_1599, n_329, n_982, n_549, n_1762, n_1910, n_1075, n_408, n_932, n_61, n_237, n_1876, n_1895, n_2123, n_1697, n_2143, n_243, n_979, n_1873, n_905, n_1866, n_1680, n_117, n_175, n_322, n_993, n_689, n_2031, n_354, n_2130, n_1330, n_1413, n_1605, n_2228, n_134, n_1988, n_1278, n_547, n_558, n_1064, n_1396, n_634, n_136, n_966, n_764, n_1663, n_2009, n_692, n_733, n_1793, n_1233, n_1289, n_2245, n_487, n_241, n_30, n_2068, n_1107, n_1014, n_1290, n_1703, n_882, n_2176, n_2072, n_1354, n_586, n_423, n_1865, n_1875, n_1701, n_318, n_1111, n_1713, n_715, n_1251, n_1265, n_88, n_1726, n_1950, n_530, n_1563, n_1912, n_277, n_1982, n_618, n_1297, n_1662, n_1312, n_199, n_1167, n_1359, n_674, n_871, n_922, n_268, n_1335, n_1760, n_1927, n_210, n_2028, n_1069, n_5, n_1664, n_1722, n_612, n_178, n_247, n_1165, n_355, n_702, n_347, n_2008, n_2192, n_2254, n_1926, n_1175, n_328, n_1386, n_1896, n_429, n_1747, n_1012, n_195, n_780, n_675, n_903, n_1540, n_1977, n_1802, n_1504, n_286, n_254, n_2193, n_1655, n_242, n_835, n_1214, n_928, n_47, n_690, n_850, n_1801, n_1886, n_2092, n_1654, n_816, n_1157, n_1750, n_1462, n_1188, n_1752, n_877, n_1813, n_2206, n_604, n_825, n_728, n_1063, n_1588, n_26, n_55, n_267, n_1124, n_1624, n_515, n_2096, n_1965, n_598, n_696, n_1515, n_961, n_437, n_1082, n_1317, n_593, n_514, n_687, n_697, n_890, n_637, n_295, n_701, n_2178, n_950, n_388, n_190, n_484, n_2036, n_2152, n_1709, n_1825, n_1757, n_1796, n_170, n_1792, n_891, n_2067, n_2136, n_2082, n_2252, n_1412, n_949, n_1630, n_678, n_283, n_2075, n_2194, n_91, n_1987, n_507, n_968, n_909, n_1369, n_881, n_1008, n_760, n_1546, n_590, n_63, n_362, n_148, n_161, n_22, n_462, n_1033, n_1052, n_1296, n_1990, n_304, n_694, n_2150, n_1294, n_1420, n_125, n_1634, n_2078, n_297, n_595, n_627, n_1767, n_1779, n_524, n_1465, n_342, n_1858, n_1044, n_2165, n_2133, n_1712, n_1391, n_449, n_131, n_1523, n_1208, n_1164, n_1295, n_1627, n_1072, n_1527, n_1495, n_1438, n_495, n_815, n_1100, n_585, n_1487, n_840, n_874, n_1756, n_1128, n_382, n_673, n_2230, n_1969, n_1071, n_1067, n_1565, n_1493, n_2145, n_1968, n_898, n_255, n_284, n_1952, n_865, n_925, n_1932, n_1101, n_15, n_1026, n_1880, n_38, n_289, n_1364, n_615, n_1249, n_59, n_1293, n_1127, n_1512, n_2151, n_1451, n_320, n_108, n_639, n_963, n_794, n_727, n_894, n_1839, n_685, n_1765, n_353, n_605, n_1514, n_1863, n_826, n_1646, n_872, n_1139, n_1714, n_86, n_104, n_718, n_1018, n_1521, n_1366, n_542, n_847, n_644, n_682, n_851, n_305, n_72, n_996, n_532, n_173, n_1308, n_2089, n_1376, n_1513, n_413, n_791, n_1913, n_510, n_837, n_2097, n_79, n_2170, n_1488, n_1808, n_948, n_704, n_2148, n_977, n_1005, n_1947, n_536, n_1788, n_1999, n_622, n_147, n_1469, n_2060, n_1838, n_1835, n_1766, n_1776, n_1959, n_2002, n_581, n_2138, n_765, n_432, n_987, n_1492, n_1340, n_1771, n_631, n_720, n_153, n_842, n_2262, n_1707, n_2239, n_1432, n_156, n_145, n_2208, n_843, n_656, n_989, n_1277, n_797, n_1473, n_2191, n_1723, n_1246, n_1878, n_899, n_189, n_738, n_2012, n_1304, n_1035, n_294, n_499, n_1426, n_705, n_11, n_1004, n_1176, n_2134, n_1529, n_1022, n_614, n_529, n_2069, n_425, n_684, n_1431, n_1615, n_1474, n_1571, n_1809, n_1577, n_1181, n_2119, n_1822, n_37, n_486, n_947, n_1117, n_1087, n_1448, n_1992, n_648, n_657, n_1049, n_2057, n_2103, n_1666, n_1505, n_803, n_290, n_118, n_1717, n_926, n_1817, n_927, n_1849, n_919, n_1698, n_478, n_2231, n_929, n_107, n_1228, n_417, n_446, n_89, n_1568, n_1490, n_777, n_1299, n_272, n_526, n_1183, n_1436, n_2251, n_1384, n_69, n_2238, n_293, n_53, n_458, n_1070, n_998, n_16, n_717, n_1665, n_18, n_154, n_1383, n_1178, n_98, n_2127, n_1424, n_1073, n_1000, n_796, n_252, n_1195, n_2137, n_1626, n_1507, n_184, n_552, n_1358, n_1811, n_1388, n_216, n_912, n_1857, n_1519, n_2144, n_745, n_1284, n_1604, n_1142, n_716, n_1475, n_623, n_1048, n_1201, n_1398, n_884, n_1774, n_1395, n_2110, n_2199, n_731, n_1502, n_1659, n_1955, n_755, n_931, n_1021, n_474, n_527, n_683, n_811, n_1207, n_312, n_1791, n_1368, n_66, n_1418, n_958, n_292, n_1250, n_100, n_1137, n_1897, n_2064, n_880, n_2053, n_2259, n_2121, n_889, n_150, n_1478, n_589, n_1310, n_819, n_1363, n_1334, n_1942, n_1966, n_767, n_1314, n_600, n_964, n_831, n_1837, n_2218, n_477, n_954, n_864, n_1110, n_2213, n_1410, n_399, n_1440, n_124, n_2132, n_2063, n_1382, n_1534, n_1564, n_1736, n_211, n_1483, n_1834, n_1372, n_231, n_40, n_1457, n_505, n_1719, n_319, n_1339, n_1787, n_537, n_1993, n_1427, n_311, n_1466, n_10, n_403, n_1919, n_1080, n_723, n_1877, n_596, n_123, n_546, n_562, n_1141, n_1268, n_386, n_1939, n_2030, n_1769, n_1220, n_1893, n_556, n_2209, n_162, n_1755, n_1602, n_1136, n_2025, n_128, n_1125, n_970, n_2224, n_1980, n_642, n_995, n_276, n_1159, n_1092, n_2237, n_441, n_221, n_1060, n_1951, n_2250, n_444, n_146, n_1252, n_1784, n_1223, n_303, n_511, n_193, n_1286, n_1773, n_1775, n_2115, n_1053, n_416, n_1681, n_520, n_418, n_1093, n_113, n_1783, n_1533, n_1597, n_4, n_266, n_296, n_775, n_651, n_1153, n_439, n_1618, n_217, n_518, n_1531, n_1185, n_453, n_215, n_1745, n_914, n_759, n_1831, n_426, n_317, n_1653, n_1679, n_1625, n_90, n_2160, n_54, n_1453, n_2146, n_2226, n_2131, n_488, n_497, n_773, n_1901, n_920, n_99, n_1374, n_1315, n_1647, n_13, n_1224, n_1614, n_1459, n_1892, n_1933, n_1135, n_1169, n_1179, n_401, n_324, n_1617, n_335, n_1470, n_463, n_1243, n_848, n_120, n_301, n_274, n_1096, n_2249, n_1091, n_1917, n_2000, n_1580, n_2227, n_1425, n_36, n_1881, n_1267, n_1281, n_1806, n_983, n_2023, n_427, n_2204, n_1520, n_496, n_2159, n_906, n_1390, n_688, n_1077, n_1733, n_1419, n_351, n_259, n_1731, n_177, n_2158, n_2087, n_1855, n_1636, n_1437, n_2135, n_1645, n_1832, n_385, n_1687, n_1439, n_1323, n_2202, n_858, n_2049, n_1331, n_613, n_736, n_501, n_956, n_960, n_663, n_856, n_2100, n_379, n_778, n_1668, n_1134, n_410, n_1129, n_554, n_602, n_1696, n_1995, n_1594, n_2181, n_664, n_1869, n_171, n_1764, n_169, n_1429, n_1610, n_1889, n_435, n_1905, n_2016, n_793, n_326, n_587, n_1593, n_580, n_762, n_1030, n_1202, n_1937, n_465, n_1790, n_1778, n_1635, n_1079, n_341, n_1744, n_828, n_2139, n_2142, n_607, n_316, n_419, n_28, n_1551, n_1103, n_144, n_2219, n_1203, n_820, n_951, n_106, n_2201, n_725, n_952, n_999, n_358, n_1254, n_160, n_186, n_0, n_368, n_575, n_994, n_2263, n_1508, n_732, n_974, n_2240, n_392, n_724, n_1934, n_1020, n_1042, n_628, n_1273, n_1434, n_1573, n_1728, n_557, n_1871, n_349, n_617, n_845, n_807, n_1036, n_140, n_1138, n_1661, n_1275, n_485, n_1549, n_67, n_443, n_1510, n_892, n_768, n_421, n_1468, n_1859, n_2102, n_238, n_1095, n_2024, n_1595, n_202, n_2156, n_1718, n_1749, n_1683, n_1916, n_597, n_280, n_1270, n_1187, n_610, n_1403, n_1669, n_1852, n_1024, n_1768, n_2153, n_198, n_1847, n_2052, n_179, n_248, n_517, n_1667, n_667, n_1206, n_621, n_1037, n_1397, n_1279, n_1115, n_750, n_901, n_1499, n_468, n_923, n_504, n_1409, n_1841, n_1639, n_1623, n_183, n_1015, n_1503, n_466, n_1057, n_603, n_991, n_1657, n_235, n_1126, n_1997, n_340, n_710, n_1108, n_1818, n_1182, n_1298, n_2177, n_39, n_2088, n_73, n_1611, n_785, n_746, n_609, n_1601, n_1960, n_2061, n_1686, n_101, n_167, n_1356, n_1589, n_127, n_1740, n_1497, n_1168, n_1216, n_1943, n_133, n_1320, n_96, n_1430, n_1316, n_1287, n_1452, n_1622, n_1586, n_302, n_1694, n_380, n_1535, n_137, n_1596, n_20, n_1190, n_1734, n_397, n_1983, n_1938, n_122, n_2220, n_34, n_1262, n_218, n_1891, n_2171, n_1213, n_70, n_2235, n_1350, n_1673, n_2232, n_1715, n_172, n_1443, n_1272, n_239, n_2037, n_97, n_782, n_1539, n_490, n_220, n_809, n_1043, n_1797, n_1608, n_986, n_2120, n_80, n_1472, n_2050, n_2164, n_2225, n_1081, n_402, n_1870, n_352, n_1692, n_800, n_1084, n_1171, n_460, n_2169, n_1827, n_1361, n_1864, n_2006, n_1491, n_2187, n_662, n_374, n_1152, n_1840, n_1705, n_450, n_2244, n_1684, n_921, n_1346, n_711, n_1642, n_579, n_1352, n_937, n_2257, n_1682, n_2017, n_370, n_1695, n_1828, n_2046, n_2200, n_650, n_1046, n_1940, n_1979, n_1145, n_330, n_1121, n_1102, n_1963, n_972, n_1405, n_258, n_1406, n_456, n_1332, n_260, n_313, n_624, n_962, n_1041, n_565, n_356, n_1569, n_936, n_1883, n_1288, n_1186, n_1062, n_885, n_896, n_83, n_2167, n_2084, n_654, n_411, n_152, n_1222, n_599, n_776, n_321, n_1823, n_105, n_227, n_1974, n_1720, n_204, n_482, n_934, n_1637, n_1407, n_1795, n_420, n_1341, n_394, n_1456, n_1845, n_1489, n_164, n_23, n_942, n_1524, n_543, n_2229, n_1964, n_1920, n_2099, n_1496, n_1271, n_1545, n_2007, n_2039, n_1946, n_1355, n_1225, n_1544, n_1485, n_2258, n_325, n_1640, n_804, n_464, n_1846, n_533, n_806, n_879, n_959, n_584, n_2141, n_244, n_1343, n_1522, n_76, n_548, n_1782, n_94, n_282, n_1676, n_833, n_1830, n_1567, n_523, n_1319, n_707, n_345, n_1900, n_799, n_1548, n_1155, n_139, n_2196, n_41, n_273, n_1633, n_2195, n_787, n_2172, n_1416, n_1528, n_1146, n_2021, n_2114, n_159, n_1086, n_1066, n_1948, n_157, n_2125, n_2026, n_1282, n_550, n_275, n_652, n_2154, n_560, n_1906, n_1484, n_1241, n_1321, n_1672, n_569, n_1758, n_1925, n_737, n_1318, n_1914, n_1235, n_1229, n_306, n_1292, n_1373, n_21, n_346, n_3, n_1029, n_1447, n_2056, n_790, n_138, n_1706, n_1498, n_1210, n_49, n_299, n_1248, n_1556, n_902, n_333, n_2189, n_2246, n_1047, n_1984, n_2236, n_1385, n_431, n_24, n_459, n_1269, n_1931, n_2083, n_502, n_672, n_1257, n_1751, n_285, n_1375, n_1941, n_85, n_2128, n_655, n_706, n_1045, n_1650, n_786, n_1794, n_1236, n_1962, n_1559, n_1725, n_1928, n_1872, n_834, n_19, n_29, n_75, n_743, n_766, n_430, n_1741, n_1325, n_1002, n_1746, n_1949, n_545, n_489, n_1804, n_1727, n_251, n_1019, n_636, n_2054, n_729, n_110, n_151, n_876, n_774, n_1337, n_660, n_2062, n_2041, n_438, n_1477, n_1360, n_1860, n_1904, n_1200, n_2070, n_479, n_1607, n_1353, n_1777, n_1908, n_1454, n_2126, n_869, n_1154, n_1113, n_1600, n_2253, n_646, n_528, n_391, n_1098, n_1329, n_2045, n_817, n_2261, n_2216, n_2210, n_262, n_187, n_897, n_846, n_2066, n_841, n_1476, n_1001, n_508, n_1800, n_2241, n_1050, n_1411, n_1463, n_1177, n_332, n_1150, n_1742, n_1562, n_1690, n_398, n_1191, n_1826, n_566, n_1023, n_1882, n_1076, n_1118, n_194, n_57, n_1007, n_1807, n_1929, n_1378, n_855, n_1592, n_1759, n_1814, n_1631, n_52, n_591, n_1377, n_1879, n_256, n_853, n_440, n_695, n_1542, n_875, n_209, n_367, n_680, n_1678, n_661, n_1716, n_278, n_1256, n_671, n_1953, n_7, n_933, n_740, n_703, n_978, n_384, n_1976, n_1291, n_1217, n_751, n_749, n_1824, n_310, n_1628, n_1324, n_1399, n_2122, n_2109, n_1435, n_969, n_988, n_2140, n_1065, n_84, n_1401, n_1255, n_568, n_1516, n_143, n_1536, n_180, n_2163, n_2186, n_2029, n_1204, n_823, n_1132, n_643, n_233, n_698, n_1074, n_1394, n_1327, n_1326, n_739, n_400, n_955, n_337, n_1379, n_214, n_246, n_1338, n_1097, n_935, n_781, n_789, n_1554, n_1130, n_181, n_1810, n_182, n_573, n_769, n_676, n_327, n_1120, n_832, n_1583, n_1730, n_555, n_389, n_814, n_1643, n_2020, n_1729, n_669, n_2048, n_176, n_114, n_300, n_222, n_2005, n_747, n_74, n_1389, n_1105, n_721, n_1461, n_742, n_535, n_691, n_372, n_2076, n_111, n_314, n_1408, n_378, n_1196, n_377, n_1598, n_863, n_2175, n_601, n_2182, n_338, n_1283, n_918, n_748, n_506, n_1114, n_1785, n_56, n_763, n_1147, n_1848, n_360, n_1754, n_2149, n_1506, n_119, n_1652, n_1812, n_957, n_1994, n_895, n_866, n_1227, n_191, n_387, n_452, n_744, n_971, n_946, n_344, n_761, n_1303, n_1205, n_1258, n_1392, n_174, n_1173, n_1924, n_525, n_1677, n_1116, n_611, n_1570, n_1702, n_1219, n_1780, n_1689, n_8, n_2180, n_1174, n_1944, n_1016, n_1347, n_795, n_1501, n_1221, n_1245, n_838, n_129, n_647, n_197, n_844, n_17, n_448, n_1017, n_2117, n_2234, n_1083, n_109, n_445, n_1561, n_930, n_888, n_1112, n_2081, n_2168, n_234, n_2022, n_1945, n_2203, n_910, n_1656, n_1721, n_1460, n_911, n_2112, n_2255, n_82, n_1464, n_27, n_236, n_653, n_1737, n_1414, n_752, n_908, n_944, n_2034, n_576, n_1028, n_2106, n_472, n_270, n_414, n_1922, n_563, n_2032, n_1011, n_1566, n_1215, n_25, n_93, n_839, n_708, n_1973, n_668, n_626, n_990, n_1500, n_779, n_1537, n_1821, n_2205, n_1104, n_854, n_1058, n_498, n_1122, n_870, n_904, n_1253, n_709, n_1266, n_366, n_2242, n_1509, n_103, n_1693, n_1109, n_185, n_2222, n_712, n_348, n_1276, n_376, n_2015, n_2118, n_2111, n_390, n_1148, n_31, n_2188, n_334, n_1989, n_1161, n_1085, n_232, n_2014, n_2042, n_46, n_1239, n_771, n_1584, n_470, n_475, n_924, n_298, n_1582, n_492, n_1149, n_265, n_1184, n_228, n_719, n_1972, n_1525, n_455, n_1585, n_1851, n_363, n_1799, n_1090, n_2147, n_592, n_1816, n_1518, n_829, n_1156, n_1362, n_393, n_984, n_1829, n_503, n_2035, n_1450, n_1638, n_132, n_868, n_570, n_859, n_2033, n_406, n_735, n_1789, n_1770, n_878, n_620, n_130, n_519, n_307, n_469, n_1218, n_500, n_1482, n_981, n_714, n_1349, n_291, n_1144, n_2071, n_357, n_985, n_2233, n_481, n_997, n_1710, n_2161, n_1301, n_802, n_561, n_33, n_980, n_1306, n_2010, n_1651, n_1198, n_2047, n_2095, n_1609, n_2174, n_436, n_116, n_409, n_1244, n_1685, n_1763, n_1998, n_1574, n_240, n_756, n_1619, n_1981, n_1606, n_810, n_1133, n_635, n_95, n_1194, n_1051, n_253, n_1552, n_583, n_1996, n_249, n_201, n_1039, n_1442, n_1034, n_2043, n_1480, n_1158, n_2248, n_754, n_941, n_975, n_1031, n_115, n_1305, n_553, n_43, n_849, n_753, n_1753, n_467, n_269, n_359, n_973, n_1921, n_1479, n_1055, n_1675, n_2197, n_2217, n_582, n_2065, n_861, n_857, n_967, n_571, n_2215, n_271, n_404, n_2001, n_158, n_2107, n_1884, n_206, n_2040, n_679, n_633, n_1170, n_665, n_1629, n_2221, n_588, n_225, n_1260, n_308, n_309, n_1819, n_2055, n_1010, n_149, n_1040, n_915, n_632, n_1166, n_2038, n_812, n_1131, n_1761, n_534, n_1578, n_1006, n_1861, n_373, n_87, n_1632, n_1890, n_1805, n_257, n_1557, n_1888, n_1833, n_730, n_1311, n_1494, n_670, n_203, n_1850, n_1898, n_2162, n_1868, n_207, n_2079, n_1089, n_1887, n_1587, n_1365, n_1417, n_205, n_1242, n_2086, n_2185, n_1836, n_681, n_1226, n_1274, n_1486, n_2166, n_412, n_640, n_1322, n_81, n_965, n_1899, n_1428, n_1616, n_1576, n_1856, n_1862, n_1958, n_2077, n_339, n_784, n_315, n_434, n_64, n_288, n_1059, n_1197, n_422, n_722, n_862, n_2105, n_135, n_165, n_2098, n_540, n_1423, n_1935, n_2027, n_457, n_2223, n_2091, n_364, n_1915, n_629, n_1621, n_1748, n_900, n_1449, n_531, n_827, n_60, n_361, n_1025, n_2116, n_336, n_12, n_1885, n_1013, n_1259, n_192, n_2183, n_1538, n_51, n_649, n_1612, n_1240, n_11214);

input n_992;
input n_1671;
input n_1;
input n_801;
input n_1613;
input n_1234;
input n_1458;
input n_1199;
input n_1674;
input n_741;
input n_1027;
input n_1351;
input n_625;
input n_1189;
input n_223;
input n_1212;
input n_226;
input n_208;
input n_68;
input n_726;
input n_2157;
input n_212;
input n_700;
input n_50;
input n_1307;
input n_2003;
input n_1038;
input n_578;
input n_1581;
input n_1003;
input n_365;
input n_168;
input n_1237;
input n_1061;
input n_1357;
input n_1853;
input n_77;
input n_783;
input n_1738;
input n_2243;
input n_798;
input n_188;
input n_1575;
input n_1854;
input n_1923;
input n_509;
input n_1342;
input n_245;
input n_1209;
input n_1348;
input n_1387;
input n_2260;
input n_677;
input n_1708;
input n_805;
input n_1151;
input n_396;
input n_1739;
input n_350;
input n_78;
input n_2051;
input n_1380;
input n_442;
input n_480;
input n_142;
input n_1402;
input n_1688;
input n_1691;
input n_1975;
input n_1009;
input n_1743;
input n_62;
input n_1930;
input n_1160;
input n_883;
input n_1238;
input n_1991;
input n_2179;
input n_1724;
input n_1032;
input n_1247;
input n_1547;
input n_1553;
input n_893;
input n_1099;
input n_1264;
input n_1192;
input n_471;
input n_1844;
input n_424;
input n_1700;
input n_1555;
input n_1415;
input n_2211;
input n_1370;
input n_1786;
input n_369;
input n_287;
input n_415;
input n_830;
input n_65;
input n_230;
input n_461;
input n_873;
input n_141;
input n_383;
input n_1285;
input n_1371;
input n_200;
input n_1985;
input n_447;
input n_2184;
input n_1803;
input n_1172;
input n_852;
input n_71;
input n_229;
input n_1590;
input n_1532;
input n_1393;
input n_1517;
input n_1867;
input n_1704;
input n_1078;
input n_250;
input n_544;
input n_1711;
input n_2247;
input n_1140;
input n_1444;
input n_1670;
input n_1603;
input n_1579;
input n_35;
input n_1263;
input n_2019;
input n_836;
input n_375;
input n_2074;
input n_522;
input n_2129;
input n_1261;
input n_945;
input n_1649;
input n_2018;
input n_2094;
input n_1903;
input n_1511;
input n_1143;
input n_1422;
input n_1232;
input n_1772;
input n_1572;
input n_616;
input n_658;
input n_1874;
input n_1119;
input n_2013;
input n_428;
input n_1433;
input n_1902;
input n_1842;
input n_1620;
input n_2044;
input n_1954;
input n_1735;
input n_1541;
input n_1300;
input n_641;
input n_822;
input n_693;
input n_1313;
input n_1056;
input n_2212;
input n_758;
input n_516;
input n_1455;
input n_1163;
input n_1180;
input n_2256;
input n_943;
input n_1798;
input n_1550;
input n_491;
input n_1591;
input n_42;
input n_772;
input n_1344;
input n_666;
input n_371;
input n_940;
input n_770;
input n_567;
input n_1781;
input n_1971;
input n_2058;
input n_2090;
input n_405;
input n_213;
input n_538;
input n_2173;
input n_2004;
input n_1106;
input n_886;
input n_1471;
input n_343;
input n_953;
input n_1094;
input n_1345;
input n_1820;
input n_494;
input n_539;
input n_493;
input n_155;
input n_2108;
input n_45;
input n_454;
input n_1421;
input n_1936;
input n_638;
input n_1404;
input n_1211;
input n_2124;
input n_381;
input n_887;
input n_1660;
input n_1961;
input n_112;
input n_1280;
input n_713;
input n_1400;
input n_126;
input n_1467;
input n_58;
input n_976;
input n_2155;
input n_224;
input n_48;
input n_1445;
input n_1526;
input n_1560;
input n_734;
input n_1088;
input n_1894;
input n_196;
input n_1231;
input n_1978;
input n_2085;
input n_917;
input n_574;
input n_9;
input n_907;
input n_6;
input n_1446;
input n_14;
input n_659;
input n_1815;
input n_2214;
input n_407;
input n_913;
input n_1658;
input n_808;
input n_867;
input n_1230;
input n_473;
input n_1193;
input n_1967;
input n_1054;
input n_559;
input n_1333;
input n_44;
input n_1648;
input n_1911;
input n_1956;
input n_163;
input n_1644;
input n_2011;
input n_1558;
input n_1732;
input n_281;
input n_551;
input n_699;
input n_1986;
input n_564;
input n_451;
input n_824;
input n_279;
input n_686;
input n_757;
input n_594;
input n_1641;
input n_2113;
input n_1918;
input n_2190;
input n_577;
input n_166;
input n_1843;
input n_619;
input n_1367;
input n_1336;
input n_521;
input n_572;
input n_395;
input n_813;
input n_1909;
input n_2080;
input n_1481;
input n_323;
input n_606;
input n_1441;
input n_818;
input n_1123;
input n_1309;
input n_92;
input n_2104;
input n_513;
input n_645;
input n_1381;
input n_331;
input n_1699;
input n_916;
input n_2093;
input n_483;
input n_102;
input n_2207;
input n_1970;
input n_608;
input n_261;
input n_2101;
input n_630;
input n_2059;
input n_32;
input n_2198;
input n_541;
input n_512;
input n_2073;
input n_121;
input n_433;
input n_792;
input n_476;
input n_2;
input n_1328;
input n_1957;
input n_219;
input n_1907;
input n_264;
input n_263;
input n_1162;
input n_860;
input n_1530;
input n_788;
input n_939;
input n_1543;
input n_821;
input n_938;
input n_1302;
input n_1068;
input n_1599;
input n_329;
input n_982;
input n_549;
input n_1762;
input n_1910;
input n_1075;
input n_408;
input n_932;
input n_61;
input n_237;
input n_1876;
input n_1895;
input n_2123;
input n_1697;
input n_2143;
input n_243;
input n_979;
input n_1873;
input n_905;
input n_1866;
input n_1680;
input n_117;
input n_175;
input n_322;
input n_993;
input n_689;
input n_2031;
input n_354;
input n_2130;
input n_1330;
input n_1413;
input n_1605;
input n_2228;
input n_134;
input n_1988;
input n_1278;
input n_547;
input n_558;
input n_1064;
input n_1396;
input n_634;
input n_136;
input n_966;
input n_764;
input n_1663;
input n_2009;
input n_692;
input n_733;
input n_1793;
input n_1233;
input n_1289;
input n_2245;
input n_487;
input n_241;
input n_30;
input n_2068;
input n_1107;
input n_1014;
input n_1290;
input n_1703;
input n_882;
input n_2176;
input n_2072;
input n_1354;
input n_586;
input n_423;
input n_1865;
input n_1875;
input n_1701;
input n_318;
input n_1111;
input n_1713;
input n_715;
input n_1251;
input n_1265;
input n_88;
input n_1726;
input n_1950;
input n_530;
input n_1563;
input n_1912;
input n_277;
input n_1982;
input n_618;
input n_1297;
input n_1662;
input n_1312;
input n_199;
input n_1167;
input n_1359;
input n_674;
input n_871;
input n_922;
input n_268;
input n_1335;
input n_1760;
input n_1927;
input n_210;
input n_2028;
input n_1069;
input n_5;
input n_1664;
input n_1722;
input n_612;
input n_178;
input n_247;
input n_1165;
input n_355;
input n_702;
input n_347;
input n_2008;
input n_2192;
input n_2254;
input n_1926;
input n_1175;
input n_328;
input n_1386;
input n_1896;
input n_429;
input n_1747;
input n_1012;
input n_195;
input n_780;
input n_675;
input n_903;
input n_1540;
input n_1977;
input n_1802;
input n_1504;
input n_286;
input n_254;
input n_2193;
input n_1655;
input n_242;
input n_835;
input n_1214;
input n_928;
input n_47;
input n_690;
input n_850;
input n_1801;
input n_1886;
input n_2092;
input n_1654;
input n_816;
input n_1157;
input n_1750;
input n_1462;
input n_1188;
input n_1752;
input n_877;
input n_1813;
input n_2206;
input n_604;
input n_825;
input n_728;
input n_1063;
input n_1588;
input n_26;
input n_55;
input n_267;
input n_1124;
input n_1624;
input n_515;
input n_2096;
input n_1965;
input n_598;
input n_696;
input n_1515;
input n_961;
input n_437;
input n_1082;
input n_1317;
input n_593;
input n_514;
input n_687;
input n_697;
input n_890;
input n_637;
input n_295;
input n_701;
input n_2178;
input n_950;
input n_388;
input n_190;
input n_484;
input n_2036;
input n_2152;
input n_1709;
input n_1825;
input n_1757;
input n_1796;
input n_170;
input n_1792;
input n_891;
input n_2067;
input n_2136;
input n_2082;
input n_2252;
input n_1412;
input n_949;
input n_1630;
input n_678;
input n_283;
input n_2075;
input n_2194;
input n_91;
input n_1987;
input n_507;
input n_968;
input n_909;
input n_1369;
input n_881;
input n_1008;
input n_760;
input n_1546;
input n_590;
input n_63;
input n_362;
input n_148;
input n_161;
input n_22;
input n_462;
input n_1033;
input n_1052;
input n_1296;
input n_1990;
input n_304;
input n_694;
input n_2150;
input n_1294;
input n_1420;
input n_125;
input n_1634;
input n_2078;
input n_297;
input n_595;
input n_627;
input n_1767;
input n_1779;
input n_524;
input n_1465;
input n_342;
input n_1858;
input n_1044;
input n_2165;
input n_2133;
input n_1712;
input n_1391;
input n_449;
input n_131;
input n_1523;
input n_1208;
input n_1164;
input n_1295;
input n_1627;
input n_1072;
input n_1527;
input n_1495;
input n_1438;
input n_495;
input n_815;
input n_1100;
input n_585;
input n_1487;
input n_840;
input n_874;
input n_1756;
input n_1128;
input n_382;
input n_673;
input n_2230;
input n_1969;
input n_1071;
input n_1067;
input n_1565;
input n_1493;
input n_2145;
input n_1968;
input n_898;
input n_255;
input n_284;
input n_1952;
input n_865;
input n_925;
input n_1932;
input n_1101;
input n_15;
input n_1026;
input n_1880;
input n_38;
input n_289;
input n_1364;
input n_615;
input n_1249;
input n_59;
input n_1293;
input n_1127;
input n_1512;
input n_2151;
input n_1451;
input n_320;
input n_108;
input n_639;
input n_963;
input n_794;
input n_727;
input n_894;
input n_1839;
input n_685;
input n_1765;
input n_353;
input n_605;
input n_1514;
input n_1863;
input n_826;
input n_1646;
input n_872;
input n_1139;
input n_1714;
input n_86;
input n_104;
input n_718;
input n_1018;
input n_1521;
input n_1366;
input n_542;
input n_847;
input n_644;
input n_682;
input n_851;
input n_305;
input n_72;
input n_996;
input n_532;
input n_173;
input n_1308;
input n_2089;
input n_1376;
input n_1513;
input n_413;
input n_791;
input n_1913;
input n_510;
input n_837;
input n_2097;
input n_79;
input n_2170;
input n_1488;
input n_1808;
input n_948;
input n_704;
input n_2148;
input n_977;
input n_1005;
input n_1947;
input n_536;
input n_1788;
input n_1999;
input n_622;
input n_147;
input n_1469;
input n_2060;
input n_1838;
input n_1835;
input n_1766;
input n_1776;
input n_1959;
input n_2002;
input n_581;
input n_2138;
input n_765;
input n_432;
input n_987;
input n_1492;
input n_1340;
input n_1771;
input n_631;
input n_720;
input n_153;
input n_842;
input n_2262;
input n_1707;
input n_2239;
input n_1432;
input n_156;
input n_145;
input n_2208;
input n_843;
input n_656;
input n_989;
input n_1277;
input n_797;
input n_1473;
input n_2191;
input n_1723;
input n_1246;
input n_1878;
input n_899;
input n_189;
input n_738;
input n_2012;
input n_1304;
input n_1035;
input n_294;
input n_499;
input n_1426;
input n_705;
input n_11;
input n_1004;
input n_1176;
input n_2134;
input n_1529;
input n_1022;
input n_614;
input n_529;
input n_2069;
input n_425;
input n_684;
input n_1431;
input n_1615;
input n_1474;
input n_1571;
input n_1809;
input n_1577;
input n_1181;
input n_2119;
input n_1822;
input n_37;
input n_486;
input n_947;
input n_1117;
input n_1087;
input n_1448;
input n_1992;
input n_648;
input n_657;
input n_1049;
input n_2057;
input n_2103;
input n_1666;
input n_1505;
input n_803;
input n_290;
input n_118;
input n_1717;
input n_926;
input n_1817;
input n_927;
input n_1849;
input n_919;
input n_1698;
input n_478;
input n_2231;
input n_929;
input n_107;
input n_1228;
input n_417;
input n_446;
input n_89;
input n_1568;
input n_1490;
input n_777;
input n_1299;
input n_272;
input n_526;
input n_1183;
input n_1436;
input n_2251;
input n_1384;
input n_69;
input n_2238;
input n_293;
input n_53;
input n_458;
input n_1070;
input n_998;
input n_16;
input n_717;
input n_1665;
input n_18;
input n_154;
input n_1383;
input n_1178;
input n_98;
input n_2127;
input n_1424;
input n_1073;
input n_1000;
input n_796;
input n_252;
input n_1195;
input n_2137;
input n_1626;
input n_1507;
input n_184;
input n_552;
input n_1358;
input n_1811;
input n_1388;
input n_216;
input n_912;
input n_1857;
input n_1519;
input n_2144;
input n_745;
input n_1284;
input n_1604;
input n_1142;
input n_716;
input n_1475;
input n_623;
input n_1048;
input n_1201;
input n_1398;
input n_884;
input n_1774;
input n_1395;
input n_2110;
input n_2199;
input n_731;
input n_1502;
input n_1659;
input n_1955;
input n_755;
input n_931;
input n_1021;
input n_474;
input n_527;
input n_683;
input n_811;
input n_1207;
input n_312;
input n_1791;
input n_1368;
input n_66;
input n_1418;
input n_958;
input n_292;
input n_1250;
input n_100;
input n_1137;
input n_1897;
input n_2064;
input n_880;
input n_2053;
input n_2259;
input n_2121;
input n_889;
input n_150;
input n_1478;
input n_589;
input n_1310;
input n_819;
input n_1363;
input n_1334;
input n_1942;
input n_1966;
input n_767;
input n_1314;
input n_600;
input n_964;
input n_831;
input n_1837;
input n_2218;
input n_477;
input n_954;
input n_864;
input n_1110;
input n_2213;
input n_1410;
input n_399;
input n_1440;
input n_124;
input n_2132;
input n_2063;
input n_1382;
input n_1534;
input n_1564;
input n_1736;
input n_211;
input n_1483;
input n_1834;
input n_1372;
input n_231;
input n_40;
input n_1457;
input n_505;
input n_1719;
input n_319;
input n_1339;
input n_1787;
input n_537;
input n_1993;
input n_1427;
input n_311;
input n_1466;
input n_10;
input n_403;
input n_1919;
input n_1080;
input n_723;
input n_1877;
input n_596;
input n_123;
input n_546;
input n_562;
input n_1141;
input n_1268;
input n_386;
input n_1939;
input n_2030;
input n_1769;
input n_1220;
input n_1893;
input n_556;
input n_2209;
input n_162;
input n_1755;
input n_1602;
input n_1136;
input n_2025;
input n_128;
input n_1125;
input n_970;
input n_2224;
input n_1980;
input n_642;
input n_995;
input n_276;
input n_1159;
input n_1092;
input n_2237;
input n_441;
input n_221;
input n_1060;
input n_1951;
input n_2250;
input n_444;
input n_146;
input n_1252;
input n_1784;
input n_1223;
input n_303;
input n_511;
input n_193;
input n_1286;
input n_1773;
input n_1775;
input n_2115;
input n_1053;
input n_416;
input n_1681;
input n_520;
input n_418;
input n_1093;
input n_113;
input n_1783;
input n_1533;
input n_1597;
input n_4;
input n_266;
input n_296;
input n_775;
input n_651;
input n_1153;
input n_439;
input n_1618;
input n_217;
input n_518;
input n_1531;
input n_1185;
input n_453;
input n_215;
input n_1745;
input n_914;
input n_759;
input n_1831;
input n_426;
input n_317;
input n_1653;
input n_1679;
input n_1625;
input n_90;
input n_2160;
input n_54;
input n_1453;
input n_2146;
input n_2226;
input n_2131;
input n_488;
input n_497;
input n_773;
input n_1901;
input n_920;
input n_99;
input n_1374;
input n_1315;
input n_1647;
input n_13;
input n_1224;
input n_1614;
input n_1459;
input n_1892;
input n_1933;
input n_1135;
input n_1169;
input n_1179;
input n_401;
input n_324;
input n_1617;
input n_335;
input n_1470;
input n_463;
input n_1243;
input n_848;
input n_120;
input n_301;
input n_274;
input n_1096;
input n_2249;
input n_1091;
input n_1917;
input n_2000;
input n_1580;
input n_2227;
input n_1425;
input n_36;
input n_1881;
input n_1267;
input n_1281;
input n_1806;
input n_983;
input n_2023;
input n_427;
input n_2204;
input n_1520;
input n_496;
input n_2159;
input n_906;
input n_1390;
input n_688;
input n_1077;
input n_1733;
input n_1419;
input n_351;
input n_259;
input n_1731;
input n_177;
input n_2158;
input n_2087;
input n_1855;
input n_1636;
input n_1437;
input n_2135;
input n_1645;
input n_1832;
input n_385;
input n_1687;
input n_1439;
input n_1323;
input n_2202;
input n_858;
input n_2049;
input n_1331;
input n_613;
input n_736;
input n_501;
input n_956;
input n_960;
input n_663;
input n_856;
input n_2100;
input n_379;
input n_778;
input n_1668;
input n_1134;
input n_410;
input n_1129;
input n_554;
input n_602;
input n_1696;
input n_1995;
input n_1594;
input n_2181;
input n_664;
input n_1869;
input n_171;
input n_1764;
input n_169;
input n_1429;
input n_1610;
input n_1889;
input n_435;
input n_1905;
input n_2016;
input n_793;
input n_326;
input n_587;
input n_1593;
input n_580;
input n_762;
input n_1030;
input n_1202;
input n_1937;
input n_465;
input n_1790;
input n_1778;
input n_1635;
input n_1079;
input n_341;
input n_1744;
input n_828;
input n_2139;
input n_2142;
input n_607;
input n_316;
input n_419;
input n_28;
input n_1551;
input n_1103;
input n_144;
input n_2219;
input n_1203;
input n_820;
input n_951;
input n_106;
input n_2201;
input n_725;
input n_952;
input n_999;
input n_358;
input n_1254;
input n_160;
input n_186;
input n_0;
input n_368;
input n_575;
input n_994;
input n_2263;
input n_1508;
input n_732;
input n_974;
input n_2240;
input n_392;
input n_724;
input n_1934;
input n_1020;
input n_1042;
input n_628;
input n_1273;
input n_1434;
input n_1573;
input n_1728;
input n_557;
input n_1871;
input n_349;
input n_617;
input n_845;
input n_807;
input n_1036;
input n_140;
input n_1138;
input n_1661;
input n_1275;
input n_485;
input n_1549;
input n_67;
input n_443;
input n_1510;
input n_892;
input n_768;
input n_421;
input n_1468;
input n_1859;
input n_2102;
input n_238;
input n_1095;
input n_2024;
input n_1595;
input n_202;
input n_2156;
input n_1718;
input n_1749;
input n_1683;
input n_1916;
input n_597;
input n_280;
input n_1270;
input n_1187;
input n_610;
input n_1403;
input n_1669;
input n_1852;
input n_1024;
input n_1768;
input n_2153;
input n_198;
input n_1847;
input n_2052;
input n_179;
input n_248;
input n_517;
input n_1667;
input n_667;
input n_1206;
input n_621;
input n_1037;
input n_1397;
input n_1279;
input n_1115;
input n_750;
input n_901;
input n_1499;
input n_468;
input n_923;
input n_504;
input n_1409;
input n_1841;
input n_1639;
input n_1623;
input n_183;
input n_1015;
input n_1503;
input n_466;
input n_1057;
input n_603;
input n_991;
input n_1657;
input n_235;
input n_1126;
input n_1997;
input n_340;
input n_710;
input n_1108;
input n_1818;
input n_1182;
input n_1298;
input n_2177;
input n_39;
input n_2088;
input n_73;
input n_1611;
input n_785;
input n_746;
input n_609;
input n_1601;
input n_1960;
input n_2061;
input n_1686;
input n_101;
input n_167;
input n_1356;
input n_1589;
input n_127;
input n_1740;
input n_1497;
input n_1168;
input n_1216;
input n_1943;
input n_133;
input n_1320;
input n_96;
input n_1430;
input n_1316;
input n_1287;
input n_1452;
input n_1622;
input n_1586;
input n_302;
input n_1694;
input n_380;
input n_1535;
input n_137;
input n_1596;
input n_20;
input n_1190;
input n_1734;
input n_397;
input n_1983;
input n_1938;
input n_122;
input n_2220;
input n_34;
input n_1262;
input n_218;
input n_1891;
input n_2171;
input n_1213;
input n_70;
input n_2235;
input n_1350;
input n_1673;
input n_2232;
input n_1715;
input n_172;
input n_1443;
input n_1272;
input n_239;
input n_2037;
input n_97;
input n_782;
input n_1539;
input n_490;
input n_220;
input n_809;
input n_1043;
input n_1797;
input n_1608;
input n_986;
input n_2120;
input n_80;
input n_1472;
input n_2050;
input n_2164;
input n_2225;
input n_1081;
input n_402;
input n_1870;
input n_352;
input n_1692;
input n_800;
input n_1084;
input n_1171;
input n_460;
input n_2169;
input n_1827;
input n_1361;
input n_1864;
input n_2006;
input n_1491;
input n_2187;
input n_662;
input n_374;
input n_1152;
input n_1840;
input n_1705;
input n_450;
input n_2244;
input n_1684;
input n_921;
input n_1346;
input n_711;
input n_1642;
input n_579;
input n_1352;
input n_937;
input n_2257;
input n_1682;
input n_2017;
input n_370;
input n_1695;
input n_1828;
input n_2046;
input n_2200;
input n_650;
input n_1046;
input n_1940;
input n_1979;
input n_1145;
input n_330;
input n_1121;
input n_1102;
input n_1963;
input n_972;
input n_1405;
input n_258;
input n_1406;
input n_456;
input n_1332;
input n_260;
input n_313;
input n_624;
input n_962;
input n_1041;
input n_565;
input n_356;
input n_1569;
input n_936;
input n_1883;
input n_1288;
input n_1186;
input n_1062;
input n_885;
input n_896;
input n_83;
input n_2167;
input n_2084;
input n_654;
input n_411;
input n_152;
input n_1222;
input n_599;
input n_776;
input n_321;
input n_1823;
input n_105;
input n_227;
input n_1974;
input n_1720;
input n_204;
input n_482;
input n_934;
input n_1637;
input n_1407;
input n_1795;
input n_420;
input n_1341;
input n_394;
input n_1456;
input n_1845;
input n_1489;
input n_164;
input n_23;
input n_942;
input n_1524;
input n_543;
input n_2229;
input n_1964;
input n_1920;
input n_2099;
input n_1496;
input n_1271;
input n_1545;
input n_2007;
input n_2039;
input n_1946;
input n_1355;
input n_1225;
input n_1544;
input n_1485;
input n_2258;
input n_325;
input n_1640;
input n_804;
input n_464;
input n_1846;
input n_533;
input n_806;
input n_879;
input n_959;
input n_584;
input n_2141;
input n_244;
input n_1343;
input n_1522;
input n_76;
input n_548;
input n_1782;
input n_94;
input n_282;
input n_1676;
input n_833;
input n_1830;
input n_1567;
input n_523;
input n_1319;
input n_707;
input n_345;
input n_1900;
input n_799;
input n_1548;
input n_1155;
input n_139;
input n_2196;
input n_41;
input n_273;
input n_1633;
input n_2195;
input n_787;
input n_2172;
input n_1416;
input n_1528;
input n_1146;
input n_2021;
input n_2114;
input n_159;
input n_1086;
input n_1066;
input n_1948;
input n_157;
input n_2125;
input n_2026;
input n_1282;
input n_550;
input n_275;
input n_652;
input n_2154;
input n_560;
input n_1906;
input n_1484;
input n_1241;
input n_1321;
input n_1672;
input n_569;
input n_1758;
input n_1925;
input n_737;
input n_1318;
input n_1914;
input n_1235;
input n_1229;
input n_306;
input n_1292;
input n_1373;
input n_21;
input n_346;
input n_3;
input n_1029;
input n_1447;
input n_2056;
input n_790;
input n_138;
input n_1706;
input n_1498;
input n_1210;
input n_49;
input n_299;
input n_1248;
input n_1556;
input n_902;
input n_333;
input n_2189;
input n_2246;
input n_1047;
input n_1984;
input n_2236;
input n_1385;
input n_431;
input n_24;
input n_459;
input n_1269;
input n_1931;
input n_2083;
input n_502;
input n_672;
input n_1257;
input n_1751;
input n_285;
input n_1375;
input n_1941;
input n_85;
input n_2128;
input n_655;
input n_706;
input n_1045;
input n_1650;
input n_786;
input n_1794;
input n_1236;
input n_1962;
input n_1559;
input n_1725;
input n_1928;
input n_1872;
input n_834;
input n_19;
input n_29;
input n_75;
input n_743;
input n_766;
input n_430;
input n_1741;
input n_1325;
input n_1002;
input n_1746;
input n_1949;
input n_545;
input n_489;
input n_1804;
input n_1727;
input n_251;
input n_1019;
input n_636;
input n_2054;
input n_729;
input n_110;
input n_151;
input n_876;
input n_774;
input n_1337;
input n_660;
input n_2062;
input n_2041;
input n_438;
input n_1477;
input n_1360;
input n_1860;
input n_1904;
input n_1200;
input n_2070;
input n_479;
input n_1607;
input n_1353;
input n_1777;
input n_1908;
input n_1454;
input n_2126;
input n_869;
input n_1154;
input n_1113;
input n_1600;
input n_2253;
input n_646;
input n_528;
input n_391;
input n_1098;
input n_1329;
input n_2045;
input n_817;
input n_2261;
input n_2216;
input n_2210;
input n_262;
input n_187;
input n_897;
input n_846;
input n_2066;
input n_841;
input n_1476;
input n_1001;
input n_508;
input n_1800;
input n_2241;
input n_1050;
input n_1411;
input n_1463;
input n_1177;
input n_332;
input n_1150;
input n_1742;
input n_1562;
input n_1690;
input n_398;
input n_1191;
input n_1826;
input n_566;
input n_1023;
input n_1882;
input n_1076;
input n_1118;
input n_194;
input n_57;
input n_1007;
input n_1807;
input n_1929;
input n_1378;
input n_855;
input n_1592;
input n_1759;
input n_1814;
input n_1631;
input n_52;
input n_591;
input n_1377;
input n_1879;
input n_256;
input n_853;
input n_440;
input n_695;
input n_1542;
input n_875;
input n_209;
input n_367;
input n_680;
input n_1678;
input n_661;
input n_1716;
input n_278;
input n_1256;
input n_671;
input n_1953;
input n_7;
input n_933;
input n_740;
input n_703;
input n_978;
input n_384;
input n_1976;
input n_1291;
input n_1217;
input n_751;
input n_749;
input n_1824;
input n_310;
input n_1628;
input n_1324;
input n_1399;
input n_2122;
input n_2109;
input n_1435;
input n_969;
input n_988;
input n_2140;
input n_1065;
input n_84;
input n_1401;
input n_1255;
input n_568;
input n_1516;
input n_143;
input n_1536;
input n_180;
input n_2163;
input n_2186;
input n_2029;
input n_1204;
input n_823;
input n_1132;
input n_643;
input n_233;
input n_698;
input n_1074;
input n_1394;
input n_1327;
input n_1326;
input n_739;
input n_400;
input n_955;
input n_337;
input n_1379;
input n_214;
input n_246;
input n_1338;
input n_1097;
input n_935;
input n_781;
input n_789;
input n_1554;
input n_1130;
input n_181;
input n_1810;
input n_182;
input n_573;
input n_769;
input n_676;
input n_327;
input n_1120;
input n_832;
input n_1583;
input n_1730;
input n_555;
input n_389;
input n_814;
input n_1643;
input n_2020;
input n_1729;
input n_669;
input n_2048;
input n_176;
input n_114;
input n_300;
input n_222;
input n_2005;
input n_747;
input n_74;
input n_1389;
input n_1105;
input n_721;
input n_1461;
input n_742;
input n_535;
input n_691;
input n_372;
input n_2076;
input n_111;
input n_314;
input n_1408;
input n_378;
input n_1196;
input n_377;
input n_1598;
input n_863;
input n_2175;
input n_601;
input n_2182;
input n_338;
input n_1283;
input n_918;
input n_748;
input n_506;
input n_1114;
input n_1785;
input n_56;
input n_763;
input n_1147;
input n_1848;
input n_360;
input n_1754;
input n_2149;
input n_1506;
input n_119;
input n_1652;
input n_1812;
input n_957;
input n_1994;
input n_895;
input n_866;
input n_1227;
input n_191;
input n_387;
input n_452;
input n_744;
input n_971;
input n_946;
input n_344;
input n_761;
input n_1303;
input n_1205;
input n_1258;
input n_1392;
input n_174;
input n_1173;
input n_1924;
input n_525;
input n_1677;
input n_1116;
input n_611;
input n_1570;
input n_1702;
input n_1219;
input n_1780;
input n_1689;
input n_8;
input n_2180;
input n_1174;
input n_1944;
input n_1016;
input n_1347;
input n_795;
input n_1501;
input n_1221;
input n_1245;
input n_838;
input n_129;
input n_647;
input n_197;
input n_844;
input n_17;
input n_448;
input n_1017;
input n_2117;
input n_2234;
input n_1083;
input n_109;
input n_445;
input n_1561;
input n_930;
input n_888;
input n_1112;
input n_2081;
input n_2168;
input n_234;
input n_2022;
input n_1945;
input n_2203;
input n_910;
input n_1656;
input n_1721;
input n_1460;
input n_911;
input n_2112;
input n_2255;
input n_82;
input n_1464;
input n_27;
input n_236;
input n_653;
input n_1737;
input n_1414;
input n_752;
input n_908;
input n_944;
input n_2034;
input n_576;
input n_1028;
input n_2106;
input n_472;
input n_270;
input n_414;
input n_1922;
input n_563;
input n_2032;
input n_1011;
input n_1566;
input n_1215;
input n_25;
input n_93;
input n_839;
input n_708;
input n_1973;
input n_668;
input n_626;
input n_990;
input n_1500;
input n_779;
input n_1537;
input n_1821;
input n_2205;
input n_1104;
input n_854;
input n_1058;
input n_498;
input n_1122;
input n_870;
input n_904;
input n_1253;
input n_709;
input n_1266;
input n_366;
input n_2242;
input n_1509;
input n_103;
input n_1693;
input n_1109;
input n_185;
input n_2222;
input n_712;
input n_348;
input n_1276;
input n_376;
input n_2015;
input n_2118;
input n_2111;
input n_390;
input n_1148;
input n_31;
input n_2188;
input n_334;
input n_1989;
input n_1161;
input n_1085;
input n_232;
input n_2014;
input n_2042;
input n_46;
input n_1239;
input n_771;
input n_1584;
input n_470;
input n_475;
input n_924;
input n_298;
input n_1582;
input n_492;
input n_1149;
input n_265;
input n_1184;
input n_228;
input n_719;
input n_1972;
input n_1525;
input n_455;
input n_1585;
input n_1851;
input n_363;
input n_1799;
input n_1090;
input n_2147;
input n_592;
input n_1816;
input n_1518;
input n_829;
input n_1156;
input n_1362;
input n_393;
input n_984;
input n_1829;
input n_503;
input n_2035;
input n_1450;
input n_1638;
input n_132;
input n_868;
input n_570;
input n_859;
input n_2033;
input n_406;
input n_735;
input n_1789;
input n_1770;
input n_878;
input n_620;
input n_130;
input n_519;
input n_307;
input n_469;
input n_1218;
input n_500;
input n_1482;
input n_981;
input n_714;
input n_1349;
input n_291;
input n_1144;
input n_2071;
input n_357;
input n_985;
input n_2233;
input n_481;
input n_997;
input n_1710;
input n_2161;
input n_1301;
input n_802;
input n_561;
input n_33;
input n_980;
input n_1306;
input n_2010;
input n_1651;
input n_1198;
input n_2047;
input n_2095;
input n_1609;
input n_2174;
input n_436;
input n_116;
input n_409;
input n_1244;
input n_1685;
input n_1763;
input n_1998;
input n_1574;
input n_240;
input n_756;
input n_1619;
input n_1981;
input n_1606;
input n_810;
input n_1133;
input n_635;
input n_95;
input n_1194;
input n_1051;
input n_253;
input n_1552;
input n_583;
input n_1996;
input n_249;
input n_201;
input n_1039;
input n_1442;
input n_1034;
input n_2043;
input n_1480;
input n_1158;
input n_2248;
input n_754;
input n_941;
input n_975;
input n_1031;
input n_115;
input n_1305;
input n_553;
input n_43;
input n_849;
input n_753;
input n_1753;
input n_467;
input n_269;
input n_359;
input n_973;
input n_1921;
input n_1479;
input n_1055;
input n_1675;
input n_2197;
input n_2217;
input n_582;
input n_2065;
input n_861;
input n_857;
input n_967;
input n_571;
input n_2215;
input n_271;
input n_404;
input n_2001;
input n_158;
input n_2107;
input n_1884;
input n_206;
input n_2040;
input n_679;
input n_633;
input n_1170;
input n_665;
input n_1629;
input n_2221;
input n_588;
input n_225;
input n_1260;
input n_308;
input n_309;
input n_1819;
input n_2055;
input n_1010;
input n_149;
input n_1040;
input n_915;
input n_632;
input n_1166;
input n_2038;
input n_812;
input n_1131;
input n_1761;
input n_534;
input n_1578;
input n_1006;
input n_1861;
input n_373;
input n_87;
input n_1632;
input n_1890;
input n_1805;
input n_257;
input n_1557;
input n_1888;
input n_1833;
input n_730;
input n_1311;
input n_1494;
input n_670;
input n_203;
input n_1850;
input n_1898;
input n_2162;
input n_1868;
input n_207;
input n_2079;
input n_1089;
input n_1887;
input n_1587;
input n_1365;
input n_1417;
input n_205;
input n_1242;
input n_2086;
input n_2185;
input n_1836;
input n_681;
input n_1226;
input n_1274;
input n_1486;
input n_2166;
input n_412;
input n_640;
input n_1322;
input n_81;
input n_965;
input n_1899;
input n_1428;
input n_1616;
input n_1576;
input n_1856;
input n_1862;
input n_1958;
input n_2077;
input n_339;
input n_784;
input n_315;
input n_434;
input n_64;
input n_288;
input n_1059;
input n_1197;
input n_422;
input n_722;
input n_862;
input n_2105;
input n_135;
input n_165;
input n_2098;
input n_540;
input n_1423;
input n_1935;
input n_2027;
input n_457;
input n_2223;
input n_2091;
input n_364;
input n_1915;
input n_629;
input n_1621;
input n_1748;
input n_900;
input n_1449;
input n_531;
input n_827;
input n_60;
input n_361;
input n_1025;
input n_2116;
input n_336;
input n_12;
input n_1885;
input n_1013;
input n_1259;
input n_192;
input n_2183;
input n_1538;
input n_51;
input n_649;
input n_1612;
input n_1240;

output n_11214;

wire n_5643;
wire n_2542;
wire n_2817;
wire n_4452;
wire n_6566;
wire n_2576;
wire n_5172;
wire n_11173;
wire n_4649;
wire n_5315;
wire n_10487;
wire n_6872;
wire n_5254;
wire n_6441;
wire n_8668;
wire n_6806;
wire n_5362;
wire n_4251;
wire n_10587;
wire n_5019;
wire n_2332;
wire n_8713;
wire n_7111;
wire n_6141;
wire n_10960;
wire n_3849;
wire n_11111;
wire n_7933;
wire n_7967;
wire n_5138;
wire n_10931;
wire n_4395;
wire n_4388;
wire n_6960;
wire n_3089;
wire n_8169;
wire n_9002;
wire n_9130;
wire n_7180;
wire n_5653;
wire n_4978;
wire n_8604;
wire n_5409;
wire n_5301;
wire n_7263;
wire n_3088;
wire n_8168;
wire n_3257;
wire n_4829;
wire n_5393;
wire n_3222;
wire n_7504;
wire n_7190;
wire n_6126;
wire n_6725;
wire n_4699;
wire n_4686;
wire n_8899;
wire n_2317;
wire n_5524;
wire n_10236;
wire n_5345;
wire n_11205;
wire n_8023;
wire n_10053;
wire n_3706;
wire n_5818;
wire n_8005;
wire n_8130;
wire n_8534;
wire n_5963;
wire n_5055;
wire n_9896;
wire n_3376;
wire n_4868;
wire n_10020;
wire n_3801;
wire n_7116;
wire n_5267;
wire n_10202;
wire n_4249;
wire n_5950;
wire n_3564;
wire n_9104;
wire n_6999;
wire n_11046;
wire n_11079;
wire n_5548;
wire n_10283;
wire n_5057;
wire n_11065;
wire n_8339;
wire n_8272;
wire n_7161;
wire n_3030;
wire n_7868;
wire n_5838;
wire n_5725;
wire n_6324;
wire n_2838;
wire n_5229;
wire n_5325;
wire n_11051;
wire n_3427;
wire n_5101;
wire n_2628;
wire n_3071;
wire n_7000;
wire n_8561;
wire n_7398;
wire n_2926;
wire n_10392;
wire n_5900;
wire n_4273;
wire n_5545;
wire n_8411;
wire n_2321;
wire n_8499;
wire n_8236;
wire n_5102;
wire n_3345;
wire n_6882;
wire n_2919;
wire n_4501;
wire n_9626;
wire n_10775;
wire n_11163;
wire n_9526;
wire n_6325;
wire n_4724;
wire n_9840;
wire n_5598;
wire n_7983;
wire n_10348;
wire n_10863;
wire n_9581;
wire n_7389;
wire n_4997;
wire n_2399;
wire n_10719;
wire n_9018;
wire n_4843;
wire n_8070;
wire n_4696;
wire n_6660;
wire n_9055;
wire n_4347;
wire n_5259;
wire n_6913;
wire n_8444;
wire n_10015;
wire n_10986;
wire n_7802;
wire n_6948;
wire n_5819;
wire n_2480;
wire n_7008;
wire n_3877;
wire n_3929;
wire n_8366;
wire n_3048;
wire n_8102;
wire n_9362;
wire n_7516;
wire n_7401;
wire n_7596;
wire n_6280;
wire n_6629;
wire n_5279;
wire n_2786;
wire n_5894;
wire n_10759;
wire n_8022;
wire n_5930;
wire n_9036;
wire n_9551;
wire n_10262;
wire n_8175;
wire n_8977;
wire n_9658;
wire n_5239;
wire n_8953;
wire n_5354;
wire n_8426;
wire n_10239;
wire n_5332;
wire n_9962;
wire n_4814;
wire n_3979;
wire n_5908;
wire n_10373;
wire n_3077;
wire n_2873;
wire n_11104;
wire n_3452;
wire n_8913;
wire n_9525;
wire n_3107;
wire n_10816;
wire n_9725;
wire n_4956;
wire n_7686;
wire n_3664;
wire n_6914;
wire n_5337;
wire n_10335;
wire n_5129;
wire n_5420;
wire n_5070;
wire n_10381;
wire n_6243;
wire n_3047;
wire n_4414;
wire n_6585;
wire n_2625;
wire n_6374;
wire n_4646;
wire n_7651;
wire n_2843;
wire n_10947;
wire n_6628;
wire n_8125;
wire n_3760;
wire n_6015;
wire n_10226;
wire n_4262;
wire n_6526;
wire n_7956;
wire n_7369;
wire n_6570;
wire n_8556;
wire n_7196;
wire n_3347;
wire n_10767;
wire n_5136;
wire n_8040;
wire n_5638;
wire n_9100;
wire n_4110;
wire n_6784;
wire n_10755;
wire n_4950;
wire n_10868;
wire n_9067;
wire n_10161;
wire n_9842;
wire n_4729;
wire n_4268;
wire n_6323;
wire n_9614;
wire n_10682;
wire n_6110;
wire n_3999;
wire n_3928;
wire n_6371;
wire n_8079;
wire n_10699;
wire n_2613;
wire n_3535;
wire n_4751;
wire n_7846;
wire n_8595;
wire n_2708;
wire n_9400;
wire n_5151;
wire n_8142;
wire n_5684;
wire n_8598;
wire n_10022;
wire n_5729;
wire n_7256;
wire n_6404;
wire n_7331;
wire n_7774;
wire n_7856;
wire n_5680;
wire n_6674;
wire n_9680;
wire n_6148;
wire n_6951;
wire n_7625;
wire n_4102;
wire n_3871;
wire n_9106;
wire n_2735;
wire n_4662;
wire n_8869;
wire n_6989;
wire n_4671;
wire n_7863;
wire n_3959;
wire n_2268;
wire n_8381;
wire n_5504;
wire n_5522;
wire n_5828;
wire n_7342;
wire n_4314;
wire n_9520;
wire n_8958;
wire n_5099;
wire n_6896;
wire n_7770;
wire n_10606;
wire n_8421;
wire n_11164;
wire n_7623;
wire n_6968;
wire n_7217;
wire n_4296;
wire n_10114;
wire n_10357;
wire n_7147;
wire n_2770;
wire n_8115;
wire n_4507;
wire n_8389;
wire n_9398;
wire n_5902;
wire n_3484;
wire n_4677;
wire n_5063;
wire n_6196;
wire n_9037;
wire n_2917;
wire n_2616;
wire n_5275;
wire n_5306;
wire n_3923;
wire n_9042;
wire n_3900;
wire n_8412;
wire n_9267;
wire n_3488;
wire n_3732;
wire n_2811;
wire n_6485;
wire n_8987;
wire n_10177;
wire n_6107;
wire n_9652;
wire n_2832;
wire n_4226;
wire n_5493;
wire n_8849;
wire n_9059;
wire n_3980;
wire n_2998;
wire n_5346;
wire n_4366;
wire n_3446;
wire n_5252;
wire n_5309;
wire n_7796;
wire n_6282;
wire n_6863;
wire n_6994;
wire n_10012;
wire n_4294;
wire n_4698;
wire n_4445;
wire n_4810;
wire n_7564;
wire n_3859;
wire n_2692;
wire n_9446;
wire n_11129;
wire n_10204;
wire n_6768;
wire n_9453;
wire n_6383;
wire n_7234;
wire n_3914;
wire n_4456;
wire n_8119;
wire n_10296;
wire n_3397;
wire n_8641;
wire n_3575;
wire n_8151;
wire n_8118;
wire n_9718;
wire n_9128;
wire n_2469;
wire n_10281;
wire n_9038;
wire n_9872;
wire n_10310;
wire n_11139;
wire n_8748;
wire n_3927;
wire n_8436;
wire n_5452;
wire n_6794;
wire n_3888;
wire n_6151;
wire n_8718;
wire n_7110;
wire n_5476;
wire n_2764;
wire n_9935;
wire n_2895;
wire n_6431;
wire n_6990;
wire n_8659;
wire n_2922;
wire n_8223;
wire n_3882;
wire n_4856;
wire n_10097;
wire n_3492;
wire n_4369;
wire n_9135;
wire n_7849;
wire n_8915;
wire n_4331;
wire n_7297;
wire n_9866;
wire n_10018;
wire n_4972;
wire n_4993;
wire n_7298;
wire n_5536;
wire n_9129;
wire n_9858;
wire n_10141;
wire n_7533;
wire n_7221;
wire n_4375;
wire n_10656;
wire n_6575;
wire n_6055;
wire n_8727;
wire n_8224;
wire n_2678;
wire n_3935;
wire n_5130;
wire n_4291;
wire n_5532;
wire n_5897;
wire n_8246;
wire n_8952;
wire n_4613;
wire n_2434;
wire n_9070;
wire n_2878;
wire n_3875;
wire n_3012;
wire n_10266;
wire n_5609;
wire n_2428;
wire n_4717;
wire n_10827;
wire n_10897;
wire n_4877;
wire n_3247;
wire n_5922;
wire n_10449;
wire n_7861;
wire n_2641;
wire n_7734;
wire n_7062;
wire n_7569;
wire n_7823;
wire n_8955;
wire n_5658;
wire n_4731;
wire n_9477;
wire n_3052;
wire n_7039;
wire n_8577;
wire n_8594;
wire n_5046;
wire n_8428;
wire n_9829;
wire n_2749;
wire n_3298;
wire n_8848;
wire n_5058;
wire n_10685;
wire n_3273;
wire n_4467;
wire n_7077;
wire n_5667;
wire n_8259;
wire n_10607;
wire n_2624;
wire n_5865;
wire n_8349;
wire n_6836;
wire n_2350;
wire n_5042;
wire n_5305;
wire n_4681;
wire n_8164;
wire n_4072;
wire n_10628;
wire n_4752;
wire n_4220;
wire n_7905;
wire n_5281;
wire n_8776;
wire n_9143;
wire n_8287;
wire n_10256;
wire n_7753;
wire n_10368;
wire n_6771;
wire n_10769;
wire n_7950;
wire n_9947;
wire n_9088;
wire n_8607;
wire n_2514;
wire n_10138;
wire n_6248;
wire n_10183;
wire n_10375;
wire n_6952;
wire n_6795;
wire n_5314;
wire n_10452;
wire n_7806;
wire n_3942;
wire n_3997;
wire n_2468;
wire n_4381;
wire n_11143;
wire n_7595;
wire n_5144;
wire n_7648;
wire n_3968;
wire n_10383;
wire n_4466;
wire n_4418;
wire n_8066;
wire n_6831;
wire n_11074;
wire n_3434;
wire n_4510;
wire n_6776;
wire n_5795;
wire n_4473;
wire n_6043;
wire n_5552;
wire n_7452;
wire n_5226;
wire n_9269;
wire n_10320;
wire n_6715;
wire n_6714;
wire n_7677;
wire n_10903;
wire n_5457;
wire n_8416;
wire n_10396;
wire n_2812;
wire n_4518;
wire n_10724;
wire n_8404;
wire n_8997;
wire n_6584;
wire n_11084;
wire n_9988;
wire n_7009;
wire n_8453;
wire n_10693;
wire n_2393;
wire n_2657;
wire n_9113;
wire n_7149;
wire n_5291;
wire n_2921;
wire n_10363;
wire n_2409;
wire n_3237;
wire n_8949;
wire n_10831;
wire n_3500;
wire n_3834;
wire n_9131;
wire n_10517;
wire n_4589;
wire n_10323;
wire n_2972;
wire n_10842;
wire n_3542;
wire n_7519;
wire n_7400;
wire n_10876;
wire n_2763;
wire n_2762;
wire n_9137;
wire n_11180;
wire n_9724;
wire n_11146;
wire n_9281;
wire n_3192;
wire n_8995;
wire n_10883;
wire n_10101;
wire n_9393;
wire n_4394;
wire n_6581;
wire n_2279;
wire n_6010;
wire n_3352;
wire n_8711;
wire n_3073;
wire n_7013;
wire n_5343;
wire n_3696;
wire n_4082;
wire n_7290;
wire n_10820;
wire n_4921;
wire n_9687;
wire n_4329;
wire n_5135;
wire n_7303;
wire n_3021;
wire n_6616;
wire n_8306;
wire n_10123;
wire n_10781;
wire n_7488;
wire n_2558;
wire n_7315;
wire n_9886;
wire n_10651;
wire n_8887;
wire n_9426;
wire n_4697;
wire n_4289;
wire n_4288;
wire n_3763;
wire n_6185;
wire n_2712;
wire n_5529;
wire n_3733;
wire n_7889;
wire n_10943;
wire n_6042;
wire n_9102;
wire n_9578;
wire n_3614;
wire n_5183;
wire n_8500;
wire n_7438;
wire n_7337;
wire n_7268;
wire n_4964;
wire n_9489;
wire n_5957;
wire n_6965;
wire n_10728;
wire n_4228;
wire n_3423;
wire n_6357;
wire n_10094;
wire n_9144;
wire n_6800;
wire n_10084;
wire n_4636;
wire n_10468;
wire n_7461;
wire n_8285;
wire n_4322;
wire n_10655;
wire n_3644;
wire n_9797;
wire n_6955;
wire n_8483;
wire n_4946;
wire n_2706;
wire n_4767;
wire n_4287;
wire n_2693;
wire n_4137;
wire n_9521;
wire n_8332;
wire n_9478;
wire n_9932;
wire n_2767;
wire n_7278;
wire n_6509;
wire n_4576;
wire n_7454;
wire n_10670;
wire n_5929;
wire n_9020;
wire n_4615;
wire n_5787;
wire n_3179;
wire n_3400;
wire n_9895;
wire n_8741;
wire n_4000;
wire n_9351;
wire n_5445;
wire n_2897;
wire n_4389;
wire n_3970;
wire n_5342;
wire n_5501;
wire n_6839;
wire n_7232;
wire n_4345;
wire n_7377;
wire n_6646;
wire n_8648;
wire n_9189;
wire n_4664;
wire n_4156;
wire n_7098;
wire n_7069;
wire n_7904;
wire n_6033;
wire n_3158;
wire n_8851;
wire n_8921;
wire n_4873;
wire n_9410;
wire n_9801;
wire n_2643;
wire n_5748;
wire n_3782;
wire n_9356;
wire n_8773;
wire n_6097;
wire n_6369;
wire n_10712;
wire n_8394;
wire n_3470;
wire n_11155;
wire n_5076;
wire n_5870;
wire n_4713;
wire n_9175;
wire n_7093;
wire n_4098;
wire n_6508;
wire n_5026;
wire n_4476;
wire n_7168;
wire n_3700;
wire n_4995;
wire n_7542;
wire n_7970;
wire n_7091;
wire n_3166;
wire n_10959;
wire n_3104;
wire n_6809;
wire n_3435;
wire n_5636;
wire n_7840;
wire n_10972;
wire n_4310;
wire n_6359;
wire n_7782;
wire n_5212;
wire n_10024;
wire n_10945;
wire n_8800;
wire n_10845;
wire n_7080;
wire n_2689;
wire n_6636;
wire n_5286;
wire n_8229;
wire n_4528;
wire n_8410;
wire n_5811;
wire n_10711;
wire n_7739;
wire n_6766;
wire n_7624;
wire n_4914;
wire n_4939;
wire n_7629;
wire n_3418;
wire n_9735;
wire n_9186;
wire n_10818;
wire n_5530;
wire n_2473;
wire n_5397;
wire n_10624;
wire n_4634;
wire n_11069;
wire n_2362;
wire n_4096;
wire n_2539;
wire n_4123;
wire n_2698;
wire n_5595;
wire n_9941;
wire n_7003;
wire n_3119;
wire n_5427;
wire n_10788;
wire n_3735;
wire n_2297;
wire n_4379;
wire n_10563;
wire n_8810;
wire n_5388;
wire n_4718;
wire n_9802;
wire n_5901;
wire n_6538;
wire n_5962;
wire n_3631;
wire n_5599;
wire n_7010;
wire n_8107;
wire n_11108;
wire n_9728;
wire n_11004;
wire n_2445;
wire n_5324;
wire n_6519;
wire n_8983;
wire n_10422;
wire n_3770;
wire n_9818;
wire n_2772;
wire n_6530;
wire n_7219;
wire n_9662;
wire n_4440;
wire n_8774;
wire n_4402;
wire n_10566;
wire n_10178;
wire n_5052;
wire n_7299;
wire n_4541;
wire n_5009;
wire n_4872;
wire n_6402;
wire n_9936;
wire n_4551;
wire n_2857;
wire n_6195;
wire n_7326;
wire n_6609;
wire n_7243;
wire n_9530;
wire n_10115;
wire n_5326;
wire n_7471;
wire n_7067;
wire n_10455;
wire n_4627;
wire n_4079;
wire n_2494;
wire n_5300;
wire n_9909;
wire n_8691;
wire n_8620;
wire n_3342;
wire n_6748;
wire n_7741;
wire n_5035;
wire n_9466;
wire n_7790;
wire n_6149;
wire n_10052;
wire n_10109;
wire n_7484;
wire n_3390;
wire n_3656;
wire n_7002;
wire n_10448;
wire n_6414;
wire n_11196;
wire n_8424;
wire n_9571;
wire n_3025;
wire n_2482;
wire n_7528;
wire n_8026;
wire n_9470;
wire n_3810;
wire n_4798;
wire n_9638;
wire n_2532;
wire n_3006;
wire n_10265;
wire n_8174;
wire n_7941;
wire n_11175;
wire n_5010;
wire n_2296;
wire n_3633;
wire n_5352;
wire n_5089;
wire n_2849;
wire n_10040;
wire n_5394;
wire n_4592;
wire n_9405;
wire n_6264;
wire n_2661;
wire n_8861;
wire n_5359;
wire n_8644;
wire n_8907;
wire n_11080;
wire n_10984;
wire n_5137;
wire n_6902;
wire n_5104;
wire n_3331;
wire n_10100;
wire n_7117;
wire n_9894;
wire n_5741;
wire n_8324;
wire n_2773;
wire n_6205;
wire n_9441;
wire n_6380;
wire n_10906;
wire n_7478;
wire n_7913;
wire n_5405;
wire n_7136;
wire n_6754;
wire n_7883;
wire n_5288;
wire n_7456;
wire n_3606;
wire n_3591;
wire n_7939;
wire n_2788;
wire n_8503;
wire n_9612;
wire n_4756;
wire n_8196;
wire n_10380;
wire n_10790;
wire n_6449;
wire n_2797;
wire n_6723;
wire n_7458;
wire n_9108;
wire n_9787;
wire n_6440;
wire n_7436;
wire n_10846;
wire n_4746;
wire n_6461;
wire n_3892;
wire n_4970;
wire n_4069;
wire n_2748;
wire n_8446;
wire n_5194;
wire n_9376;
wire n_9786;
wire n_9033;
wire n_2331;
wire n_2292;
wire n_7435;
wire n_3441;
wire n_9537;
wire n_3534;
wire n_6997;
wire n_10509;
wire n_5952;
wire n_3964;
wire n_2416;
wire n_5947;
wire n_8923;
wire n_3944;
wire n_6124;
wire n_6736;
wire n_7685;
wire n_7363;
wire n_8192;
wire n_5985;
wire n_8197;
wire n_3605;
wire n_6622;
wire n_9443;
wire n_9996;
wire n_4633;
wire n_6891;
wire n_7800;
wire n_10031;
wire n_3306;
wire n_9115;
wire n_3026;
wire n_4584;
wire n_3090;
wire n_5232;
wire n_3724;
wire n_7663;
wire n_4276;
wire n_10898;
wire n_5116;
wire n_2990;
wire n_3847;
wire n_5001;
wire n_2552;
wire n_5176;
wire n_7443;
wire n_7747;
wire n_9779;
wire n_9938;
wire n_8082;
wire n_4428;
wire n_8730;
wire n_3323;
wire n_7917;
wire n_7261;
wire n_9023;
wire n_6528;
wire n_2274;
wire n_9203;
wire n_9977;
wire n_7532;
wire n_8051;
wire n_9613;
wire n_5761;
wire n_9242;
wire n_6773;
wire n_4618;
wire n_7375;
wire n_4679;
wire n_3479;
wire n_4496;
wire n_7968;
wire n_6382;
wire n_7455;
wire n_4805;
wire n_8651;
wire n_3454;
wire n_9141;
wire n_5760;
wire n_6885;
wire n_9201;
wire n_10732;
wire n_6531;
wire n_10952;
wire n_10851;
wire n_11027;
wire n_10660;
wire n_7430;
wire n_5472;
wire n_3547;
wire n_10221;
wire n_9559;
wire n_8377;
wire n_9299;
wire n_9937;
wire n_5679;
wire n_11162;
wire n_7912;
wire n_9913;
wire n_5100;
wire n_2575;
wire n_9286;
wire n_8015;
wire n_5973;
wire n_7921;
wire n_10044;
wire n_7728;
wire n_4410;
wire n_8281;
wire n_10819;
wire n_3816;
wire n_4807;
wire n_8842;
wire n_4411;
wire n_9184;
wire n_3214;
wire n_9704;
wire n_2928;
wire n_5166;
wire n_9046;
wire n_6339;
wire n_8024;
wire n_7730;
wire n_8814;
wire n_8530;
wire n_2822;
wire n_4180;
wire n_9193;
wire n_8467;
wire n_7281;
wire n_3109;
wire n_9717;
wire n_3354;
wire n_2572;
wire n_7711;
wire n_3126;
wire n_11090;
wire n_8984;
wire n_3663;
wire n_2863;
wire n_3299;
wire n_5688;
wire n_6417;
wire n_9290;
wire n_5740;
wire n_5820;
wire n_5648;
wire n_5745;
wire n_4707;
wire n_4676;
wire n_9403;
wire n_10996;
wire n_9875;
wire n_5180;
wire n_6763;
wire n_8956;
wire n_5182;
wire n_7858;
wire n_8676;
wire n_5534;
wire n_8003;
wire n_4880;
wire n_8785;
wire n_9853;
wire n_3566;
wire n_7448;
wire n_6542;
wire n_4126;
wire n_2781;
wire n_2829;
wire n_3845;
wire n_6556;
wire n_8692;
wire n_6889;
wire n_7230;
wire n_9183;
wire n_3804;
wire n_7989;
wire n_4207;
wire n_9778;
wire n_5196;
wire n_6199;
wire n_9823;
wire n_5171;
wire n_10698;
wire n_10852;
wire n_4470;
wire n_6726;
wire n_9529;
wire n_4813;
wire n_5542;
wire n_3901;
wire n_7011;
wire n_8998;
wire n_10538;
wire n_5261;
wire n_10870;
wire n_4014;
wire n_4704;
wire n_11066;
wire n_10315;
wire n_4252;
wire n_9123;
wire n_4028;
wire n_6576;
wire n_6471;
wire n_2448;
wire n_8906;
wire n_5949;
wire n_4048;
wire n_4596;
wire n_4444;
wire n_5255;
wire n_3756;
wire n_8482;
wire n_6478;
wire n_7952;
wire n_3406;
wire n_6100;
wire n_6516;
wire n_3919;
wire n_8462;
wire n_6977;
wire n_9380;
wire n_10062;
wire n_7660;
wire n_6915;
wire n_7834;
wire n_5185;
wire n_6911;
wire n_8409;
wire n_6599;
wire n_6522;
wire n_8979;
wire n_4952;
wire n_2656;
wire n_5023;
wire n_2375;
wire n_5906;
wire n_8429;
wire n_8930;
wire n_10514;
wire n_5660;
wire n_3981;
wire n_7890;
wire n_3973;
wire n_2756;
wire n_7245;
wire n_5334;
wire n_6024;
wire n_9347;
wire n_4761;
wire n_6675;
wire n_6270;
wire n_6808;
wire n_2884;
wire n_7620;
wire n_7265;
wire n_7986;
wire n_5783;
wire n_6207;
wire n_7006;
wire n_6931;
wire n_3120;
wire n_5821;
wire n_6245;
wire n_6079;
wire n_7948;
wire n_3797;
wire n_9082;
wire n_10925;
wire n_4770;
wire n_9879;
wire n_11158;
wire n_3474;
wire n_9861;
wire n_6963;
wire n_8685;
wire n_2549;
wire n_4690;
wire n_3864;
wire n_8264;
wire n_5556;
wire n_4932;
wire n_8250;
wire n_8492;
wire n_7381;
wire n_10601;
wire n_5456;
wire n_9158;
wire n_2302;
wire n_8135;
wire n_10618;
wire n_9594;
wire n_7837;
wire n_9832;
wire n_7717;
wire n_8445;
wire n_9518;
wire n_6427;
wire n_6580;
wire n_5143;
wire n_9898;
wire n_3592;
wire n_5500;
wire n_6412;
wire n_4230;
wire n_10497;
wire n_9445;
wire n_2637;
wire n_7627;
wire n_9803;
wire n_3967;
wire n_7601;
wire n_6437;
wire n_8298;
wire n_3195;
wire n_6346;
wire n_2526;
wire n_4274;
wire n_5215;
wire n_7860;
wire n_8408;
wire n_3277;
wire n_2548;
wire n_5386;
wire n_10661;
wire n_7335;
wire n_4189;
wire n_9815;
wire n_8895;
wire n_9495;
wire n_3817;
wire n_10028;
wire n_7811;
wire n_11044;
wire n_3659;
wire n_2559;
wire n_2595;
wire n_5003;
wire n_10512;
wire n_4827;
wire n_2694;
wire n_8450;
wire n_3648;
wire n_8273;
wire n_9867;
wire n_6059;
wire n_7499;
wire n_3042;
wire n_6065;
wire n_9688;
wire n_9761;
wire n_7292;
wire n_5094;
wire n_4610;
wire n_10967;
wire n_9087;
wire n_4472;
wire n_5433;
wire n_7870;
wire n_9043;
wire n_6075;
wire n_3228;
wire n_3657;
wire n_7397;
wire n_3081;
wire n_10789;
wire n_11134;
wire n_6117;
wire n_7977;
wire n_8886;
wire n_10434;
wire n_7211;
wire n_10933;
wire n_5618;
wire n_6861;
wire n_8312;
wire n_6781;
wire n_7847;
wire n_8506;
wire n_2264;
wire n_3464;
wire n_6494;
wire n_6133;
wire n_3723;
wire n_8963;
wire n_7822;
wire n_4380;
wire n_6453;
wire n_5978;
wire n_9307;
wire n_5247;
wire n_4996;
wire n_4990;
wire n_6127;
wire n_10762;
wire n_4398;
wire n_2498;
wire n_8078;
wire n_7785;
wire n_6217;
wire n_4515;
wire n_5031;
wire n_6006;
wire n_10797;
wire n_7289;
wire n_4193;
wire n_3570;
wire n_7926;
wire n_5082;
wire n_6598;
wire n_7399;
wire n_5338;
wire n_3828;
wire n_7354;
wire n_8352;
wire n_2392;
wire n_3424;
wire n_4131;
wire n_10360;
wire n_7960;
wire n_9450;
wire n_2298;
wire n_2326;
wire n_3594;
wire n_5689;
wire n_7482;
wire n_10312;
wire n_4090;
wire n_6115;
wire n_4165;
wire n_8143;
wire n_2305;
wire n_4626;
wire n_9223;
wire n_10480;
wire n_6048;
wire n_4144;
wire n_6416;
wire n_2964;
wire n_10131;
wire n_6838;
wire n_10068;
wire n_6867;
wire n_9693;
wire n_6139;
wire n_4077;
wire n_5931;
wire n_2371;
wire n_3485;
wire n_10633;
wire n_6256;
wire n_7965;
wire n_3262;
wire n_6613;
wire n_4008;
wire n_3356;
wire n_5221;
wire n_10273;
wire n_5641;
wire n_10209;
wire n_3210;
wire n_6361;
wire n_9880;
wire n_4689;
wire n_8183;
wire n_4547;
wire n_9685;
wire n_6085;
wire n_7474;
wire n_11169;
wire n_5731;
wire n_6329;
wire n_8650;
wire n_6678;
wire n_3329;
wire n_8662;
wire n_10503;
wire n_9694;
wire n_3826;
wire n_4905;
wire n_7158;
wire n_4601;
wire n_9905;
wire n_9948;
wire n_10465;
wire n_10590;
wire n_3647;
wire n_3681;
wire n_4300;
wire n_8526;
wire n_4623;
wire n_7325;
wire n_10887;
wire n_9456;
wire n_5007;
wire n_7044;
wire n_3320;
wire n_9710;
wire n_6370;
wire n_8623;
wire n_11113;
wire n_9923;
wire n_2518;
wire n_5883;
wire n_7166;
wire n_6554;
wire n_7356;
wire n_5754;
wire n_6759;
wire n_10786;
wire n_3988;
wire n_6560;
wire n_3476;
wire n_7028;
wire n_4842;
wire n_7838;
wire n_9890;
wire n_5629;
wire n_3439;
wire n_4135;
wire n_7873;
wire n_2688;
wire n_6535;
wire n_7518;
wire n_2798;
wire n_7414;
wire n_9744;
wire n_9817;
wire n_6147;
wire n_2852;
wire n_9199;
wire n_10063;
wire n_9548;
wire n_8973;
wire n_11160;
wire n_6448;
wire n_7791;
wire n_8419;
wire n_9782;
wire n_2753;
wire n_3292;
wire n_9862;
wire n_5434;
wire n_5934;
wire n_7431;
wire n_10805;
wire n_3437;
wire n_4111;
wire n_6643;
wire n_7146;
wire n_9471;
wire n_3712;
wire n_4608;
wire n_2310;
wire n_2506;
wire n_10091;
wire n_6157;
wire n_4859;
wire n_9363;
wire n_2626;
wire n_5880;
wire n_4037;
wire n_8351;
wire n_8430;
wire n_10747;
wire n_9069;
wire n_3562;
wire n_5852;
wire n_2973;
wire n_8603;
wire n_9422;
wire n_5218;
wire n_8249;
wire n_7052;
wire n_3665;
wire n_10496;
wire n_3007;
wire n_3528;
wire n_5960;
wire n_4571;
wire n_10843;
wire n_3698;
wire n_7888;
wire n_5358;
wire n_6397;
wire n_3355;
wire n_2454;
wire n_8234;
wire n_3174;
wire n_5321;
wire n_9960;
wire n_10997;
wire n_4215;
wire n_9010;
wire n_10998;
wire n_9003;
wire n_9280;
wire n_6073;
wire n_7502;
wire n_6331;
wire n_5290;
wire n_4185;
wire n_3752;
wire n_7312;
wire n_7919;
wire n_2283;
wire n_5145;
wire n_4219;
wire n_10800;
wire n_7085;
wire n_3958;
wire n_9341;
wire n_6939;
wire n_7848;
wire n_3985;
wire n_2427;
wire n_4196;
wire n_4774;
wire n_5210;
wire n_6689;
wire n_10993;
wire n_7632;
wire n_4242;
wire n_5109;
wire n_3389;
wire n_9172;
wire n_4232;
wire n_4190;
wire n_4902;
wire n_3000;
wire n_6405;
wire n_7580;
wire n_5149;
wire n_8980;
wire n_5571;
wire n_2680;
wire n_10112;
wire n_10765;
wire n_3375;
wire n_3899;
wire n_6698;
wire n_7304;
wire n_3713;
wire n_9734;
wire n_2668;
wire n_7288;
wire n_8558;
wire n_10489;
wire n_7707;
wire n_3197;
wire n_7223;
wire n_7833;
wire n_4987;
wire n_5512;
wire n_7274;
wire n_9297;
wire n_10159;
wire n_10495;
wire n_9004;
wire n_4736;
wire n_2398;
wire n_3743;
wire n_6206;
wire n_9068;
wire n_8136;
wire n_5033;
wire n_9808;
wire n_2695;
wire n_4035;
wire n_3818;
wire n_6610;
wire n_7445;
wire n_3124;
wire n_10612;
wire n_11086;
wire n_7466;
wire n_6529;
wire n_10260;
wire n_3759;
wire n_2671;
wire n_4516;
wire n_6363;
wire n_6750;
wire n_2715;
wire n_8619;
wire n_2508;
wire n_3511;
wire n_6290;
wire n_10253;
wire n_7429;
wire n_6025;
wire n_11038;
wire n_9150;
wire n_10134;
wire n_7277;
wire n_6455;
wire n_2614;
wire n_8146;
wire n_4492;
wire n_2833;
wire n_2758;
wire n_8813;
wire n_5607;
wire n_3694;
wire n_7695;
wire n_2937;
wire n_10194;
wire n_7179;
wire n_10356;
wire n_7122;
wire n_10173;
wire n_7165;
wire n_7869;
wire n_4789;
wire n_5999;
wire n_8910;
wire n_4376;
wire n_6203;
wire n_6408;
wire n_6555;
wire n_9448;
wire n_7683;
wire n_10739;
wire n_6150;
wire n_7630;
wire n_10077;
wire n_4708;
wire n_8470;
wire n_4657;
wire n_9587;
wire n_5341;
wire n_8643;
wire n_4512;
wire n_9278;
wire n_10671;
wire n_10889;
wire n_10010;
wire n_10193;
wire n_8565;
wire n_10821;
wire n_11170;
wire n_8550;
wire n_4081;
wire n_9396;
wire n_4542;
wire n_6892;
wire n_11094;
wire n_4462;
wire n_7061;
wire n_10599;
wire n_9667;
wire n_6401;
wire n_7322;
wire n_9053;
wire n_6685;
wire n_4931;
wire n_9739;
wire n_10573;
wire n_4536;
wire n_9480;
wire n_5562;
wire n_3303;
wire n_4324;
wire n_7051;
wire n_10850;
wire n_8477;
wire n_9185;
wire n_7880;
wire n_9793;
wire n_4382;
wire n_2905;
wire n_8230;
wire n_6679;
wire n_8092;
wire n_3954;
wire n_5911;
wire n_10546;
wire n_5622;
wire n_3503;
wire n_9919;
wire n_3160;
wire n_6574;
wire n_11116;
wire n_6571;
wire n_5577;
wire n_9541;
wire n_8876;
wire n_5124;
wire n_9151;
wire n_3951;
wire n_8829;
wire n_7824;
wire n_9359;
wire n_3569;
wire n_7094;
wire n_3874;
wire n_2528;
wire n_5123;
wire n_7097;
wire n_4639;
wire n_5413;
wire n_8140;
wire n_8971;
wire n_8060;
wire n_10558;
wire n_3027;
wire n_7036;
wire n_4083;
wire n_9579;
wire n_9475;
wire n_11124;
wire n_6392;
wire n_5915;
wire n_8527;
wire n_9049;
wire n_7351;
wire n_4480;
wire n_9352;
wire n_2295;
wire n_2746;
wire n_7608;
wire n_5779;
wire n_6260;
wire n_6832;
wire n_7394;
wire n_11045;
wire n_7909;
wire n_7413;
wire n_4171;
wire n_6303;
wire n_3652;
wire n_8935;
wire n_10734;
wire n_6286;
wire n_7675;
wire n_8267;
wire n_4023;
wire n_7027;
wire n_7992;
wire n_6912;
wire n_10330;
wire n_7175;
wire n_8276;
wire n_3617;
wire n_10395;
wire n_6019;
wire n_10174;
wire n_3567;
wire n_7524;
wire n_4344;
wire n_2935;
wire n_8027;
wire n_4705;
wire n_4046;
wire n_3807;
wire n_8925;
wire n_6214;
wire n_9978;
wire n_9370;
wire n_11125;
wire n_9670;
wire n_4027;
wire n_3154;
wire n_9334;
wire n_7783;
wire n_6692;
wire n_2485;
wire n_3898;
wire n_10276;
wire n_3520;
wire n_8978;
wire n_10594;
wire n_8093;
wire n_8245;
wire n_6036;
wire n_8471;
wire n_4391;
wire n_9956;
wire n_9800;
wire n_8454;
wire n_6552;
wire n_4095;
wire n_8327;
wire n_9413;
wire n_10991;
wire n_2881;
wire n_10098;
wire n_8891;
wire n_4947;
wire n_3551;
wire n_3064;
wire n_9487;
wire n_3897;
wire n_5591;
wire n_3372;
wire n_7697;
wire n_6403;
wire n_7306;
wire n_7947;
wire n_10118;
wire n_7470;
wire n_7547;
wire n_6013;
wire n_7733;
wire n_7693;
wire n_9557;
wire n_3215;
wire n_6491;
wire n_3853;
wire n_4740;
wire n_4631;
wire n_6348;
wire n_6744;
wire n_8582;
wire n_10441;
wire n_5518;
wire n_6982;
wire n_10002;
wire n_5068;
wire n_6293;
wire n_6661;
wire n_9124;
wire n_5847;
wire n_7345;
wire n_6049;
wire n_9762;
wire n_8847;
wire n_8957;
wire n_7385;
wire n_10923;
wire n_5159;
wire n_2862;
wire n_2615;
wire n_4068;
wire n_6558;
wire n_4625;
wire n_11149;
wire n_10841;
wire n_2474;
wire n_3703;
wire n_2437;
wire n_2444;
wire n_3962;
wire n_2743;
wire n_4766;
wire n_8488;
wire n_9271;
wire n_4863;
wire n_2267;
wire n_9543;
wire n_3035;
wire n_4166;
wire n_8356;
wire n_6136;
wire n_9660;
wire n_9483;
wire n_3378;
wire n_6855;
wire n_3745;
wire n_3362;
wire n_10665;
wire n_4744;
wire n_8888;
wire n_4188;
wire n_5357;
wire n_2934;
wire n_3667;
wire n_6091;
wire n_3523;
wire n_9328;
wire n_7857;
wire n_3176;
wire n_7481;
wire n_6551;
wire n_7691;
wire n_7907;
wire n_5541;
wire n_5568;
wire n_10576;
wire n_6312;
wire n_8747;
wire n_2505;
wire n_9539;
wire n_4817;
wire n_6668;
wire n_9415;
wire n_4115;
wire n_2999;
wire n_9385;
wire n_3697;
wire n_9147;
wire n_11209;
wire n_7653;
wire n_3680;
wire n_5381;
wire n_8354;
wire n_2408;
wire n_9785;
wire n_5723;
wire n_6859;
wire n_5918;
wire n_3468;
wire n_6959;
wire n_8353;
wire n_8922;
wire n_6388;
wire n_5045;
wire n_10237;
wire n_11053;
wire n_9027;
wire n_9434;
wire n_4383;
wire n_6995;
wire n_10902;
wire n_4491;
wire n_5696;
wire n_8348;
wire n_7032;
wire n_8211;
wire n_4486;
wire n_9515;
wire n_10420;
wire n_6971;
wire n_9642;
wire n_9233;
wire n_6131;
wire n_9681;
wire n_5848;
wire n_3024;
wire n_7475;
wire n_10485;
wire n_4612;
wire n_6435;
wire n_10536;
wire n_5673;
wire n_5443;
wire n_2531;
wire n_6351;
wire n_9079;
wire n_9382;
wire n_10282;
wire n_5163;
wire n_6212;
wire n_7668;
wire n_9775;
wire n_10444;
wire n_4529;
wire n_3361;
wire n_3478;
wire n_8018;
wire n_8653;
wire n_3936;
wire n_8920;
wire n_10913;
wire n_7937;
wire n_9176;
wire n_6829;
wire n_2723;
wire n_10950;
wire n_5485;
wire n_7819;
wire n_10631;
wire n_5823;
wire n_7305;
wire n_2800;
wire n_3496;
wire n_11071;
wire n_5473;
wire n_10072;
wire n_6682;
wire n_6334;
wire n_6823;
wire n_10708;
wire n_10703;
wire n_9089;
wire n_9666;
wire n_4390;
wire n_3096;
wire n_8678;
wire n_10565;
wire n_10011;
wire n_2651;
wire n_8884;
wire n_8803;
wire n_3239;
wire n_8942;
wire n_7993;
wire n_7181;
wire n_9865;
wire n_3161;
wire n_2799;
wire n_5537;
wire n_10978;
wire n_8222;
wire n_6822;
wire n_3902;
wire n_4062;
wire n_3295;
wire n_4396;
wire n_8553;
wire n_7071;
wire n_9706;
wire n_3101;
wire n_10642;
wire n_4233;
wire n_10187;
wire n_3374;
wire n_10387;
wire n_11014;
wire n_2640;
wire n_3288;
wire n_2918;
wire n_8751;
wire n_4307;
wire n_3992;
wire n_3876;
wire n_11007;
wire n_11006;
wire n_9564;
wire n_3125;
wire n_7391;
wire n_8790;
wire n_9230;
wire n_6617;
wire n_4293;
wire n_10219;
wire n_3552;
wire n_7511;
wire n_6533;
wire n_10768;
wire n_10316;
wire n_9795;
wire n_4684;
wire n_3116;
wire n_9591;
wire n_6429;
wire n_6407;
wire n_4091;
wire n_6389;
wire n_5027;
wire n_3095;
wire n_6137;
wire n_10364;
wire n_2471;
wire n_10479;
wire n_8338;
wire n_6983;
wire n_10494;
wire n_8398;
wire n_4412;
wire n_2807;
wire n_8178;
wire n_6801;
wire n_8491;
wire n_3618;
wire n_4580;
wire n_5630;
wire n_4758;
wire n_4781;
wire n_10065;
wire n_10212;
wire n_9283;
wire n_8700;
wire n_4148;
wire n_2461;
wire n_4057;
wire n_5379;
wire n_5335;
wire n_10268;
wire n_3444;
wire n_3059;
wire n_6113;
wire n_9468;
wire n_10070;
wire n_9425;
wire n_2634;
wire n_11172;
wire n_10089;
wire n_5424;
wire n_8750;
wire n_3017;
wire n_2477;
wire n_5505;
wire n_5868;
wire n_10305;
wire n_8560;
wire n_10559;
wire n_2308;
wire n_2333;
wire n_8439;
wire n_3001;
wire n_9641;
wire n_10004;
wire n_3795;
wire n_7321;
wire n_3852;
wire n_5289;
wire n_4138;
wire n_8200;
wire n_11110;
wire n_7154;
wire n_5018;
wire n_6129;
wire n_6518;
wire n_8304;
wire n_3815;
wire n_3896;
wire n_6655;
wire n_8674;
wire n_5274;
wire n_9138;
wire n_3274;
wire n_5401;
wire n_7584;
wire n_9958;
wire n_4457;
wire n_7537;
wire n_10516;
wire n_4093;
wire n_8675;
wire n_6254;
wire n_5989;
wire n_10892;
wire n_10493;
wire n_9367;
wire n_7320;
wire n_4928;
wire n_5769;
wire n_10405;
wire n_4794;
wire n_5613;
wire n_8212;
wire n_5612;
wire n_4197;
wire n_7964;
wire n_4482;
wire n_9016;
wire n_2547;
wire n_2415;
wire n_6278;
wire n_6786;
wire n_7022;
wire n_10026;
wire n_9729;
wire n_5073;
wire n_8846;
wire n_8315;
wire n_11033;
wire n_4834;
wire n_11040;
wire n_9194;
wire n_8760;
wire n_9756;
wire n_4762;
wire n_5581;
wire n_9029;
wire n_9411;
wire n_3113;
wire n_6837;
wire n_10353;
wire n_3813;
wire n_3660;
wire n_10847;
wire n_3766;
wire n_10451;
wire n_11043;
wire n_5303;
wire n_7486;
wire n_6756;
wire n_9414;
wire n_3266;
wire n_7023;
wire n_3574;
wire n_9615;
wire n_7496;
wire n_4154;
wire n_4907;
wire n_5077;
wire n_5034;
wire n_10866;
wire n_7410;
wire n_9940;
wire n_10779;
wire n_8563;
wire n_6200;
wire n_4504;
wire n_3844;
wire n_8777;
wire n_4975;
wire n_2534;
wire n_11061;
wire n_8465;
wire n_6670;
wire n_3741;
wire n_8535;
wire n_10653;
wire n_6373;
wire n_5375;
wire n_9221;
wire n_2451;
wire n_5370;
wire n_4898;
wire n_4815;
wire n_5601;
wire n_5784;
wire n_9811;
wire n_3443;
wire n_7899;
wire n_8631;
wire n_4819;
wire n_7906;
wire n_5248;
wire n_9951;
wire n_7131;
wire n_6411;
wire n_9424;
wire n_9586;
wire n_10285;
wire n_4370;
wire n_8909;
wire n_11032;
wire n_2359;
wire n_5112;
wire n_3332;
wire n_4134;
wire n_10507;
wire n_10520;
wire n_7302;
wire n_2570;
wire n_4092;
wire n_10045;
wire n_11174;
wire n_4645;
wire n_7797;
wire n_3668;
wire n_6381;
wire n_7030;
wire n_6656;
wire n_9730;
wire n_7687;
wire n_2491;
wire n_9554;
wire n_10294;
wire n_4755;
wire n_4359;
wire n_4960;
wire n_10106;
wire n_4087;
wire n_5635;
wire n_7582;
wire n_9934;
wire n_4933;
wire n_10541;
wire n_5091;
wire n_3487;
wire n_4591;
wire n_6546;
wire n_5528;
wire n_4302;
wire n_9234;
wire n_10674;
wire n_5111;
wire n_8959;
wire n_6534;
wire n_3340;
wire n_10614;
wire n_5227;
wire n_7809;
wire n_10417;
wire n_3946;
wire n_6265;
wire n_2989;
wire n_5778;
wire n_8425;
wire n_8087;
wire n_9910;
wire n_3395;
wire n_7060;
wire n_7607;
wire n_10217;
wire n_8938;
wire n_4474;
wire n_5665;
wire n_2509;
wire n_2513;
wire n_6898;
wire n_6596;
wire n_3757;
wire n_5363;
wire n_4178;
wire n_10743;
wire n_5165;
wire n_4884;
wire n_10853;
wire n_7867;
wire n_9651;
wire n_3275;
wire n_10249;
wire n_8361;
wire n_6135;
wire n_7761;
wire n_10705;
wire n_8007;
wire n_9246;
wire n_10338;
wire n_10270;
wire n_3678;
wire n_6814;
wire n_10557;
wire n_3440;
wire n_11115;
wire n_8669;
wire n_8001;
wire n_7525;
wire n_2356;
wire n_7257;
wire n_9372;
wire n_7553;
wire n_7529;
wire n_4692;
wire n_6791;
wire n_8496;
wire n_3165;
wire n_6824;
wire n_5788;
wire n_11016;
wire n_9326;
wire n_2739;
wire n_3890;
wire n_3750;
wire n_3607;
wire n_7650;
wire n_3316;
wire n_8568;
wire n_6903;
wire n_2418;
wire n_2864;
wire n_8852;
wire n_4311;
wire n_8637;
wire n_2703;
wire n_6168;
wire n_6881;
wire n_3371;
wire n_4722;
wire n_4606;
wire n_10339;
wire n_9908;
wire n_10908;
wire n_9486;
wire n_6450;
wire n_9544;
wire n_3261;
wire n_7520;
wire n_9831;
wire n_4187;
wire n_6309;
wire n_7903;
wire n_9697;
wire n_2660;
wire n_6733;
wire n_8864;
wire n_7384;
wire n_8456;
wire n_5317;
wire n_5430;
wire n_5942;
wire n_8610;
wire n_7894;
wire n_4962;
wire n_4563;
wire n_7137;
wire n_9902;
wire n_5056;
wire n_8362;
wire n_4820;
wire n_2394;
wire n_5540;
wire n_9900;
wire n_6300;
wire n_8256;
wire n_3532;
wire n_9920;
wire n_7055;
wire n_7202;
wire n_5716;
wire n_8520;
wire n_9310;
wire n_10132;
wire n_3948;
wire n_9039;
wire n_8573;
wire n_8265;
wire n_4619;
wire n_7639;
wire n_8704;
wire n_5762;
wire n_6132;
wire n_4327;
wire n_5211;
wire n_5336;
wire n_3765;
wire n_5447;
wire n_4125;
wire n_7743;
wire n_9294;
wire n_5036;
wire n_4221;
wire n_3297;
wire n_6179;
wire n_6395;
wire n_10327;
wire n_7054;
wire n_7605;
wire n_3067;
wire n_11001;
wire n_9512;
wire n_10437;
wire n_2686;
wire n_5327;
wire n_10021;
wire n_9146;
wire n_2364;
wire n_9125;
wire n_4392;
wire n_9170;
wire n_9139;
wire n_2996;
wire n_7433;
wire n_9616;
wire n_8131;
wire n_3803;
wire n_8941;
wire n_5014;
wire n_5747;
wire n_3639;
wire n_9073;
wire n_10075;
wire n_10423;
wire n_5192;
wire n_4334;
wire n_3351;
wire n_6171;
wire n_8775;
wire n_9302;
wire n_5519;
wire n_9062;
wire n_4047;
wire n_6269;
wire n_5753;
wire n_3413;
wire n_7092;
wire n_6980;
wire n_11213;
wire n_9171;
wire n_10886;
wire n_5233;
wire n_3412;
wire n_8279;
wire n_6654;
wire n_9358;
wire n_9580;
wire n_8019;
wire n_9972;
wire n_3791;
wire n_6083;
wire n_3164;
wire n_4575;
wire n_6434;
wire n_6387;
wire n_4320;
wire n_9565;
wire n_9157;
wire n_8257;
wire n_10192;
wire n_7832;
wire n_3884;
wire n_9465;
wire n_9540;
wire n_9324;
wire n_5808;
wire n_8390;
wire n_11137;
wire n_8898;
wire n_7726;
wire n_8807;
wire n_5436;
wire n_5139;
wire n_5231;
wire n_6120;
wire n_8613;
wire n_6068;
wire n_6933;
wire n_8521;
wire n_4141;
wire n_3438;
wire n_10436;
wire n_8464;
wire n_6547;
wire n_8799;
wire n_5193;
wire n_6423;
wire n_9442;
wire n_2850;
wire n_6342;
wire n_6641;
wire n_6984;
wire n_3373;
wire n_5789;
wire n_10763;
wire n_7441;
wire n_9957;
wire n_10124;
wire n_7106;
wire n_7213;
wire n_3883;
wire n_10245;
wire n_5961;
wire n_10905;
wire n_9449;
wire n_5866;
wire n_9050;
wire n_3728;
wire n_6507;
wire n_2925;
wire n_4499;
wire n_6399;
wire n_6687;
wire n_9313;
wire n_5822;
wire n_9173;
wire n_5195;
wire n_6690;
wire n_6121;
wire n_7412;
wire n_9959;
wire n_3949;
wire n_5726;
wire n_9563;
wire n_11015;
wire n_2792;
wire n_9160;
wire n_5364;
wire n_9974;
wire n_11166;
wire n_3315;
wire n_7031;
wire n_9285;
wire n_5533;
wire n_7763;
wire n_3798;
wire n_9631;
wire n_8033;
wire n_4257;
wire n_4458;
wire n_6194;
wire n_2674;
wire n_5103;
wire n_4641;
wire n_8393;
wire n_7133;
wire n_4720;
wire n_10784;
wire n_4893;
wire n_3857;
wire n_4107;
wire n_8463;
wire n_8153;
wire n_3630;
wire n_6524;
wire n_3518;
wire n_10944;
wire n_10211;
wire n_10129;
wire n_10431;
wire n_9945;
wire n_8661;
wire n_7424;
wire n_3714;
wire n_7523;
wire n_8654;
wire n_5039;
wire n_2455;
wire n_2876;
wire n_4772;
wire n_6790;
wire n_8746;
wire n_5953;
wire n_11183;
wire n_10019;
wire n_3099;
wire n_11156;
wire n_8531;
wire n_10611;
wire n_7141;
wire n_5198;
wire n_10715;
wire n_4468;
wire n_5718;
wire n_4161;
wire n_6505;
wire n_6459;
wire n_8379;
wire n_8609;
wire n_4172;
wire n_3403;
wire n_7626;
wire n_2714;
wire n_4961;
wire n_7310;
wire n_4454;
wire n_3294;
wire n_2457;
wire n_6686;
wire n_4119;
wire n_6001;
wire n_7311;
wire n_9209;
wire n_3686;
wire n_7669;
wire n_4502;
wire n_5958;
wire n_8793;
wire n_8103;
wire n_9838;
wire n_2971;
wire n_9767;
wire n_10195;
wire n_4277;
wire n_4526;
wire n_9300;
wire n_3490;
wire n_4849;
wire n_4319;
wire n_7327;
wire n_3369;
wire n_8873;
wire n_8367;
wire n_7367;
wire n_5792;
wire n_11021;
wire n_3581;
wire n_8543;
wire n_3069;
wire n_6183;
wire n_6023;
wire n_7323;
wire n_7189;
wire n_7301;
wire n_10730;
wire n_6258;
wire n_3715;
wire n_6905;
wire n_10243;
wire n_9700;
wire n_10564;
wire n_8682;
wire n_3725;
wire n_8089;
wire n_9218;
wire n_6704;
wire n_3933;
wire n_8533;
wire n_9118;
wire n_11122;
wire n_6657;
wire n_7655;
wire n_5554;
wire n_7244;
wire n_10745;
wire n_7368;
wire n_2311;
wire n_3691;
wire n_10596;
wire n_5553;
wire n_4485;
wire n_8011;
wire n_4066;
wire n_7633;
wire n_4146;
wire n_5711;
wire n_9437;
wire n_10263;
wire n_4340;
wire n_5790;
wire n_8640;
wire n_8063;
wire n_3961;
wire n_4855;
wire n_2347;
wire n_3917;
wire n_6186;
wire n_7878;
wire n_6803;
wire n_9514;
wire n_6210;
wire n_8437;
wire n_6500;
wire n_8427;
wire n_8032;
wire n_10280;
wire n_7427;
wire n_10605;
wire n_4004;
wire n_11029;
wire n_2967;
wire n_5404;
wire n_9933;
wire n_2916;
wire n_11190;
wire n_5739;
wire n_10951;
wire n_4292;
wire n_9892;
wire n_8570;
wire n_6163;
wire n_7628;
wire n_9462;
wire n_9074;
wire n_5972;
wire n_10519;
wire n_2467;
wire n_5549;
wire n_9408;
wire n_3145;
wire n_6785;
wire n_6553;
wire n_10163;
wire n_10454;
wire n_3983;
wire n_4940;
wire n_5444;
wire n_3538;
wire n_3280;
wire n_8039;
wire n_5757;
wire n_8902;
wire n_8916;
wire n_7557;
wire n_10087;
wire n_4356;
wire n_3510;
wire n_2824;
wire n_8843;
wire n_9891;
wire n_10146;
wire n_7128;
wire n_9946;
wire n_2377;
wire n_6849;
wire n_9885;
wire n_7594;
wire n_8129;
wire n_8162;
wire n_7457;
wire n_10643;
wire n_8744;
wire n_3009;
wire n_10504;
wire n_5824;
wire n_3719;
wire n_2525;
wire n_7788;
wire n_4361;
wire n_10872;
wire n_5488;
wire n_6760;
wire n_10701;
wire n_3827;
wire n_5154;
wire n_10658;
wire n_7752;
wire n_3889;
wire n_2687;
wire n_2887;
wire n_9509;
wire n_4245;
wire n_4136;
wire n_8286;
wire n_3526;
wire n_2619;
wire n_5329;
wire n_9015;
wire n_4367;
wire n_9757;
wire n_5637;
wire n_9925;
wire n_10874;
wire n_6825;
wire n_7586;
wire n_10008;
wire n_6452;
wire n_9628;
wire n_7767;
wire n_8294;
wire n_2271;
wire n_9419;
wire n_6611;
wire n_8562;
wire n_2583;
wire n_4560;
wire n_2606;
wire n_4899;
wire n_10250;
wire n_5728;
wire n_5471;
wire n_2794;
wire n_10032;
wire n_10592;
wire n_5164;
wire n_9277;
wire n_9257;
wire n_2391;
wire n_2431;
wire n_7207;
wire n_8218;
wire n_9806;
wire n_5843;
wire n_8170;
wire n_9159;
wire n_7744;
wire n_7021;
wire n_2932;
wire n_3431;
wire n_10595;
wire n_7748;
wire n_8537;
wire n_3450;
wire n_6827;
wire n_10126;
wire n_4663;
wire n_2893;
wire n_11073;
wire n_5484;
wire n_6355;
wire n_2954;
wire n_2728;
wire n_6227;
wire n_7215;
wire n_7485;
wire n_3421;
wire n_9066;
wire n_3183;
wire n_4802;
wire n_2493;
wire n_5523;
wire n_2705;
wire n_10302;
wire n_3405;
wire n_8016;
wire n_8671;
wire n_5423;
wire n_10645;
wire n_10604;
wire n_5074;
wire n_11096;
wire n_4044;
wire n_6564;
wire n_3436;
wire n_11161;
wire n_9671;
wire n_8709;
wire n_8782;
wire n_3442;
wire n_3366;
wire n_2631;
wire n_6468;
wire n_3937;
wire n_10080;
wire n_10570;
wire n_9857;
wire n_3159;
wire n_4701;
wire n_10966;
wire n_10057;
wire n_10882;
wire n_9338;
wire n_6857;
wire n_3240;
wire n_8144;
wire n_3576;
wire n_10435;
wire n_9542;
wire n_3385;
wire n_10795;
wire n_10921;
wire n_7171;
wire n_4851;
wire n_6442;
wire n_3293;
wire n_3922;
wire n_11085;
wire n_8049;
wire n_5204;
wire n_7762;
wire n_5333;
wire n_9467;
wire n_7068;
wire n_7925;
wire n_7186;
wire n_10609;
wire n_11157;
wire n_4991;
wire n_5594;
wire n_2554;
wire n_9097;
wire n_5422;
wire n_6871;
wire n_9783;
wire n_9510;
wire n_9389;
wire n_4934;
wire n_9404;
wire n_8357;
wire n_6904;
wire n_10912;
wire n_5087;
wire n_9916;
wire n_5526;
wire n_5292;
wire n_2517;
wire n_2713;
wire n_9314;
wire n_7017;
wire n_7777;
wire n_9752;
wire n_5000;
wire n_2765;
wire n_5403;
wire n_2590;
wire n_5551;
wire n_7652;
wire n_3150;
wire n_10220;
wire n_8701;
wire n_10341;
wire n_4479;
wire n_2608;
wire n_6499;
wire n_10550;
wire n_7830;
wire n_4011;
wire n_5131;
wire n_3133;
wire n_7138;
wire n_5257;
wire n_8097;
wire n_9679;
wire n_8084;
wire n_9306;
wire n_8645;
wire n_4753;
wire n_4688;
wire n_8712;
wire n_10232;
wire n_4058;
wire n_10461;
wire n_8289;
wire n_11178;
wire n_3611;
wire n_3082;
wire n_4848;
wire n_7966;
wire n_8591;
wire n_5059;
wire n_8837;
wire n_5887;
wire n_8811;
wire n_8824;
wire n_2604;
wire n_2407;
wire n_2816;
wire n_7191;
wire n_3799;
wire n_7712;
wire n_2574;
wire n_4475;
wire n_10412;
wire n_5242;
wire n_10326;
wire n_5219;
wire n_8417;
wire n_2675;
wire n_6276;
wire n_9721;
wire n_5631;
wire n_3537;
wire n_10499;
wire n_8340;
wire n_4443;
wire n_3887;
wire n_6008;
wire n_9197;
wire n_7997;
wire n_6420;
wire n_5854;
wire n_2667;
wire n_5460;
wire n_4587;
wire n_4114;
wire n_2948;
wire n_8455;
wire n_7208;
wire n_9210;
wire n_7961;
wire n_9770;
wire n_6893;
wire n_5899;
wire n_5686;
wire n_7406;
wire n_8681;
wire n_8905;
wire n_3223;
wire n_10617;
wire n_3140;
wire n_7807;
wire n_3185;
wire n_4749;
wire n_9592;
wire n_2605;
wire n_5155;
wire n_7680;
wire n_9180;
wire n_10922;
wire n_10544;
wire n_3654;
wire n_2848;
wire n_8172;
wire n_9917;
wire n_10718;
wire n_8106;
wire n_9502;
wire n_4100;
wire n_6447;
wire n_4264;
wire n_5981;
wire n_3788;
wire n_9625;
wire n_4891;
wire n_5937;
wire n_6422;
wire n_6751;
wire n_5339;
wire n_3837;
wire n_2718;
wire n_11087;
wire n_3325;
wire n_9873;
wire n_6040;
wire n_8375;
wire n_4085;
wire n_4464;
wire n_8612;
wire n_4624;
wire n_4818;
wire n_6851;
wire n_6460;
wire n_8345;
wire n_10095;
wire n_4659;
wire n_10309;
wire n_3600;
wire n_6741;
wire n_8459;
wire n_5217;
wire n_5465;
wire n_11099;
wire n_5015;
wire n_8974;
wire n_4339;
wire n_8268;
wire n_2338;
wire n_3324;
wire n_6160;
wire n_9871;
wire n_6650;
wire n_8221;
wire n_10050;
wire n_7066;
wire n_9164;
wire n_8255;
wire n_7183;
wire n_7789;
wire n_10306;
wire n_10878;
wire n_7606;
wire n_8461;
wire n_6192;
wire n_6368;
wire n_10056;
wire n_7140;
wire n_7193;
wire n_3987;
wire n_6039;
wire n_4487;
wire n_6583;
wire n_4866;
wire n_4889;
wire n_10450;
wire n_5721;
wire n_3638;
wire n_9114;
wire n_4816;
wire n_8515;
wire n_10529;
wire n_5719;
wire n_5773;
wire n_5482;
wire n_3393;
wire n_8812;
wire n_6012;
wire n_3451;
wire n_9392;
wire n_10429;
wire n_4937;
wire n_10904;
wire n_5277;
wire n_8792;
wire n_3615;
wire n_7344;
wire n_9888;
wire n_3072;
wire n_3087;
wire n_10037;
wire n_4222;
wire n_6707;
wire n_9698;
wire n_4874;
wire n_4401;
wire n_2710;
wire n_6064;
wire n_11136;
wire n_9903;
wire n_3142;
wire n_4015;
wire n_5793;
wire n_9644;
wire n_6787;
wire n_11102;
wire n_8523;
wire n_4709;
wire n_9228;
wire n_10179;
wire n_4976;
wire n_7710;
wire n_2389;
wire n_9499;
wire n_7892;
wire n_2892;
wire n_6647;
wire n_4120;
wire n_6275;
wire n_9522;
wire n_5578;
wire n_4658;
wire n_2860;
wire n_2330;
wire n_5296;
wire n_11076;
wire n_9366;
wire n_3718;
wire n_7915;
wire n_5893;
wire n_7750;
wire n_9077;
wire n_6769;
wire n_9148;
wire n_2281;
wire n_11054;
wire n_8406;
wire n_6277;
wire n_2617;
wire n_2776;
wire n_10754;
wire n_5742;
wire n_5207;
wire n_11050;
wire n_3705;
wire n_3211;
wire n_6463;
wire n_3909;
wire n_5676;
wire n_8554;
wire n_10920;
wire n_9275;
wire n_10223;
wire n_6051;
wire n_8896;
wire n_2301;
wire n_4665;
wire n_3582;
wire n_7206;
wire n_4223;
wire n_11126;
wire n_7538;
wire n_2387;
wire n_5674;
wire n_3270;
wire n_5539;
wire n_6895;
wire n_2846;
wire n_5282;
wire n_10295;
wire n_2488;
wire n_9409;
wire n_5464;
wire n_6799;
wire n_10336;
wire n_10228;
wire n_4362;
wire n_3311;
wire n_3913;
wire n_7716;
wire n_6487;
wire n_5121;
wire n_8758;
wire n_9768;
wire n_6026;
wire n_6070;
wire n_8818;
wire n_4430;
wire n_3302;
wire n_8617;
wire n_4348;
wire n_9881;
wire n_5013;
wire n_6807;
wire n_8954;
wire n_9463;
wire n_7251;
wire n_4489;
wire n_4839;
wire n_7254;
wire n_10466;
wire n_2596;
wire n_3163;
wire n_7540;
wire n_4404;
wire n_5589;
wire n_6563;
wire n_10776;
wire n_7882;
wire n_2828;
wire n_8552;
wire n_10425;
wire n_7554;
wire n_2384;
wire n_8069;
wire n_7558;
wire n_4261;
wire n_4204;
wire n_8373;
wire n_10848;
wire n_2724;
wire n_6481;
wire n_2585;
wire n_5628;
wire n_4825;
wire n_2352;
wire n_7765;
wire n_3986;
wire n_5006;
wire n_4513;
wire n_7816;
wire n_4006;
wire n_11089;
wire n_2801;
wire n_9997;
wire n_6341;
wire n_10164;
wire n_6384;
wire n_3869;
wire n_7421;
wire n_2556;
wire n_10166;
wire n_7489;
wire n_4747;
wire n_6906;
wire n_7541;
wire n_5251;
wire n_3753;
wire n_2306;
wire n_3742;
wire n_9844;
wire n_3683;
wire n_8318;
wire n_4801;
wire n_3260;
wire n_10366;
wire n_2550;
wire n_8341;
wire n_9970;
wire n_11193;
wire n_3175;
wire n_9595;
wire n_7188;
wire n_3736;
wire n_5475;
wire n_7334;
wire n_6923;
wire n_5807;
wire n_4448;
wire n_9287;
wire n_7991;
wire n_6233;
wire n_10877;
wire n_6377;
wire n_9265;
wire n_5216;
wire n_3284;
wire n_10225;
wire n_4869;
wire n_8239;
wire n_8926;
wire n_6257;
wire n_2315;
wire n_4132;
wire n_4386;
wire n_10361;
wire n_2995;
wire n_5273;
wire n_7898;
wire n_10766;
wire n_4438;
wire n_4844;
wire n_8383;
wire n_10086;
wire n_4836;
wire n_5439;
wire n_7143;
wire n_9789;
wire n_10424;
wire n_4955;
wire n_8965;
wire n_4149;
wire n_5936;
wire n_9608;
wire n_4355;
wire n_7646;
wire n_3234;
wire n_2276;
wire n_9052;
wire n_2803;
wire n_8817;
wire n_8190;
wire n_2777;
wire n_3202;
wire n_2830;
wire n_3220;
wire n_6587;
wire n_6987;
wire n_7781;
wire n_7360;
wire n_11037;
wire n_6069;
wire n_2911;
wire n_7497;
wire n_4655;
wire n_5706;
wire n_2826;
wire n_7665;
wire n_9354;
wire n_3429;
wire n_10501;
wire n_10817;
wire n_2379;
wire n_7793;
wire n_8355;
wire n_3554;
wire n_6991;
wire n_10556;
wire n_7101;
wire n_7671;
wire n_9436;
wire n_7530;
wire n_8489;
wire n_5431;
wire n_7248;
wire n_4067;
wire n_4357;
wire n_10350;
wire n_7204;
wire n_9860;
wire n_8649;
wire n_6887;
wire n_10567;
wire n_7578;
wire n_3462;
wire n_7654;
wire n_2851;
wire n_8303;
wire n_6153;
wire n_4374;
wire n_5132;
wire n_6637;
wire n_8369;
wire n_9022;
wire n_9238;
wire n_8059;
wire n_6633;
wire n_10230;
wire n_2420;
wire n_5627;
wire n_9103;
wire n_11031;
wire n_5774;
wire n_6579;
wire n_3722;
wire n_4400;
wire n_4846;
wire n_5798;
wire n_2984;
wire n_11138;
wire n_5187;
wire n_5875;
wire n_9839;
wire n_4024;
wire n_8831;
wire n_5621;
wire n_5608;
wire n_7900;
wire n_6569;
wire n_2983;
wire n_6335;
wire n_7120;
wire n_8728;
wire n_10807;
wire n_2538;
wire n_3250;
wire n_6789;
wire n_8386;
wire n_8853;
wire n_4582;
wire n_6252;
wire n_4860;
wire n_6211;
wire n_10511;
wire n_5844;
wire n_8862;
wire n_3414;
wire n_10580;
wire n_4870;
wire n_6164;
wire n_7576;
wire n_6173;
wire n_8081;
wire n_9675;
wire n_7786;
wire n_11023;
wire n_3651;
wire n_7313;
wire n_10058;
wire n_2563;
wire n_10873;
wire n_4989;
wire n_7676;
wire n_7609;
wire n_7757;
wire n_3449;
wire n_2598;
wire n_8900;
wire n_6630;
wire n_6934;
wire n_9017;
wire n_10484;
wire n_4304;
wire n_4558;
wire n_6737;
wire n_4488;
wire n_3767;
wire n_8396;
wire n_6612;
wire n_8478;
wire n_6606;
wire n_2544;
wire n_6695;
wire n_3550;
wire n_8865;
wire n_10288;
wire n_10337;
wire n_4211;
wire n_7779;
wire n_8999;
wire n_6189;
wire n_10388;
wire n_4016;
wire n_11072;
wire n_5867;
wire n_5508;
wire n_4656;
wire n_6479;
wire n_10791;
wire n_10506;
wire n_3839;
wire n_8497;
wire n_2823;
wire n_10770;
wire n_8820;
wire n_6410;
wire n_9318;
wire n_6158;
wire n_5597;
wire n_9028;
wire n_4915;
wire n_4328;
wire n_9492;
wire n_6413;
wire n_6090;
wire n_8020;
wire n_9374;
wire n_7419;
wire n_6506;
wire n_2785;
wire n_5515;
wire n_5662;
wire n_2636;
wire n_3131;
wire n_3730;
wire n_6935;
wire n_9727;
wire n_10413;
wire n_10593;
wire n_5862;
wire n_4397;
wire n_3399;
wire n_5050;
wire n_10636;
wire n_2740;
wire n_4808;
wire n_7667;
wire n_5697;
wire n_3416;
wire n_10203;
wire n_3498;
wire n_10980;
wire n_9174;
wire n_5767;
wire n_2401;
wire n_8992;
wire n_4712;
wire n_8880;
wire n_10369;
wire n_8690;
wire n_2309;
wire n_2900;
wire n_6234;
wire n_2957;
wire n_2737;
wire n_6821;
wire n_3994;
wire n_5462;
wire n_9983;
wire n_9375;
wire n_10082;
wire n_6688;
wire n_5980;
wire n_8580;
wire n_7818;
wire n_9993;
wire n_8770;
wire n_3672;
wire n_7182;
wire n_5318;
wire n_7365;
wire n_6608;
wire n_10467;
wire n_3533;
wire n_9109;
wire n_9849;
wire n_6105;
wire n_4725;
wire n_6022;
wire n_11207;
wire n_9856;
wire n_10964;
wire n_4406;
wire n_3382;
wire n_3132;
wire n_5498;
wire n_2571;
wire n_3138;
wire n_8075;
wire n_6798;
wire n_10838;
wire n_10530;
wire n_5053;
wire n_7896;
wire n_7841;
wire n_9458;
wire n_9237;
wire n_7885;
wire n_6860;
wire n_6557;
wire n_8466;
wire n_6753;
wire n_6527;
wire n_7341;
wire n_2988;
wire n_9349;
wire n_4908;
wire n_3136;
wire n_11200;
wire n_11091;
wire n_8094;
wire n_4192;
wire n_4109;
wire n_10940;
wire n_6639;
wire n_4824;
wire n_2808;
wire n_4567;
wire n_6430;
wire n_5150;
wire n_8832;
wire n_10987;
wire n_3819;
wire n_4778;
wire n_5477;
wire n_5175;
wire n_8839;
wire n_7996;
wire n_4595;
wire n_4174;
wire n_11098;
wire n_10533;
wire n_11059;
wire n_5987;
wire n_5179;
wire n_7957;
wire n_4904;
wire n_10938;
wire n_10176;
wire n_7517;
wire n_6627;
wire n_8080;
wire n_3544;
wire n_4150;
wire n_2904;
wire n_5988;
wire n_5585;
wire n_6058;
wire n_7745;
wire n_3105;
wire n_2872;
wire n_6666;
wire n_3692;
wire n_10927;
wire n_4616;
wire n_8321;
wire n_8772;
wire n_8735;
wire n_9954;
wire n_4982;
wire n_2272;
wire n_8592;
wire n_8786;
wire n_11204;
wire n_8684;
wire n_6190;
wire n_2760;
wire n_4643;
wire n_6249;
wire n_2738;
wire n_8083;
wire n_5348;
wire n_11060;
wire n_10578;
wire n_6594;
wire n_9805;
wire n_5480;
wire n_10155;
wire n_4323;
wire n_8157;
wire n_2346;
wire n_4831;
wire n_7095;
wire n_3045;
wire n_3821;
wire n_10714;
wire n_6969;
wire n_6615;
wire n_6161;
wire n_7459;
wire n_2970;
wire n_2342;
wire n_7294;
wire n_3676;
wire n_4896;
wire n_8206;
wire n_2882;
wire n_3666;
wire n_3675;
wire n_4017;
wire n_4260;
wire n_4916;
wire n_9110;
wire n_10569;
wire n_2541;
wire n_8622;
wire n_2940;
wire n_5904;
wire n_4739;
wire n_7184;
wire n_9617;
wire n_6607;
wire n_9335;
wire n_6062;
wire n_7908;
wire n_9452;
wire n_4122;
wire n_7974;
wire n_7551;
wire n_10051;
wire n_4209;
wire n_8104;
wire n_10414;
wire n_8344;
wire n_2768;
wire n_3858;
wire n_5284;
wire n_4298;
wire n_2314;
wire n_8120;
wire n_3502;
wire n_8513;
wire n_10120;
wire n_9474;
wire n_5461;
wire n_3003;
wire n_9075;
wire n_6482;
wire n_9427;
wire n_4128;
wire n_10746;
wire n_9188;
wire n_6294;
wire n_5147;
wire n_9611;
wire n_4271;
wire n_4644;
wire n_9021;
wire n_8779;
wire n_9810;
wire n_8621;
wire n_5503;
wire n_5845;
wire n_9250;
wire n_5945;
wire n_9550;
wire n_11212;
wire n_10697;
wire n_10641;
wire n_2390;
wire n_6246;
wire n_8868;
wire n_2562;
wire n_8134;
wire n_4716;
wire n_4312;
wire n_9975;
wire n_2734;
wire n_7250;
wire n_5600;
wire n_5755;
wire n_8762;
wire n_8043;
wire n_8694;
wire n_5048;
wire n_6053;
wire n_7252;
wire n_3246;
wire n_3381;
wire n_9207;
wire n_4944;
wire n_3208;
wire n_10103;
wire n_5245;
wire n_4343;
wire n_6843;
wire n_10926;
wire n_4715;
wire n_6123;
wire n_8897;
wire n_11000;
wire n_10626;
wire n_6901;
wire n_4935;
wire n_4694;
wire n_8191;
wire n_10325;
wire n_6841;
wire n_4672;
wire n_10153;
wire n_8101;
wire n_5054;
wire n_10298;
wire n_2962;
wire n_8171;
wire n_8376;
wire n_5448;
wire n_6922;
wire n_9006;
wire n_2939;
wire n_7698;
wire n_5749;
wire n_6774;
wire n_6271;
wire n_6489;
wire n_8600;
wire n_4407;
wire n_7402;
wire n_8431;
wire n_8710;
wire n_3517;
wire n_4045;
wire n_3893;
wire n_3061;
wire n_4598;
wire n_2945;
wire n_3932;
wire n_3469;
wire n_8599;
wire n_2960;
wire n_8549;
wire n_10172;
wire n_5993;
wire n_8054;
wire n_10400;
wire n_6716;
wire n_9637;
wire n_3258;
wire n_9418;
wire n_8616;
wire n_4524;
wire n_3143;
wire n_6020;
wire n_9177;
wire n_9060;
wire n_9096;
wire n_9081;
wire n_4084;
wire n_3149;
wire n_6844;
wire n_9236;
wire n_7914;
wire n_8628;
wire n_3365;
wire n_6521;
wire n_7891;
wire n_3379;
wire n_8857;
wire n_8517;
wire n_4850;
wire n_8547;
wire n_10156;
wire n_4424;
wire n_9040;
wire n_7113;
wire n_9607;
wire n_3008;
wire n_6162;
wire n_10433;
wire n_2840;
wire n_6779;
wire n_8010;
wire n_3939;
wire n_4776;
wire n_6432;
wire n_9116;
wire n_10774;
wire n_3972;
wire n_4153;
wire n_10901;
wire n_11034;
wire n_10549;
wire n_10839;
wire n_3506;
wire n_7216;
wire n_3855;
wire n_10825;
wire n_3091;
wire n_4317;
wire n_8275;
wire n_4723;
wire n_6198;
wire n_4269;
wire n_5418;
wire n_6543;
wire n_9830;
wire n_6762;
wire n_6178;
wire n_9621;
wire n_4088;
wire n_3398;
wire n_5685;
wire n_10761;
wire n_2761;
wire n_2793;
wire n_3776;
wire n_3711;
wire n_4235;
wire n_5459;
wire n_9035;
wire n_10398;
wire n_8291;
wire n_4170;
wire n_4143;
wire n_3642;
wire n_2845;
wire n_4650;
wire n_7706;
wire n_4719;
wire n_5173;
wire n_7477;
wire n_5016;
wire n_2874;
wire n_2588;
wire n_6458;
wire n_4967;
wire n_7642;
wire n_9678;
wire n_8247;
wire n_6577;
wire n_6740;
wire n_3308;
wire n_6315;
wire n_2366;
wire n_10581;
wire n_4912;
wire n_4799;
wire n_9284;
wire n_4423;
wire n_5086;
wire n_5283;
wire n_9111;
wire n_7156;
wire n_4735;
wire n_9163;
wire n_3602;
wire n_3300;
wire n_2978;
wire n_2516;
wire n_5170;
wire n_6910;
wire n_6262;
wire n_7604;
wire n_2827;
wire n_7703;
wire n_3515;
wire n_9606;
wire n_6319;
wire n_2951;
wire n_10470;
wire n_2949;
wire n_10297;
wire n_5028;
wire n_5839;
wire n_6536;
wire n_6175;
wire n_3806;
wire n_7040;
wire n_8827;
wire n_10625;
wire n_8280;
wire n_5514;
wire n_2931;
wire n_8388;
wire n_2569;
wire n_10235;
wire n_3866;
wire n_6978;
wire n_9589;
wire n_5351;
wire n_5909;
wire n_9344;
wire n_10865;
wire n_9549;
wire n_6093;
wire n_4543;
wire n_10445;
wire n_7378;
wire n_10738;
wire n_4157;
wire n_8988;
wire n_6845;
wire n_9798;
wire n_9190;
wire n_6947;
wire n_4229;
wire n_9482;
wire n_5293;
wire n_8203;
wire n_6099;
wire n_3865;
wire n_4073;
wire n_8569;
wire n_3629;
wire n_5400;
wire n_3920;
wire n_4892;
wire n_3255;
wire n_6140;
wire n_8877;
wire n_9412;
wire n_7498;
wire n_10679;
wire n_10799;
wire n_3846;
wire n_6321;
wire n_3512;
wire n_6819;
wire n_7501;
wire n_5201;
wire n_9506;
wire n_10136;
wire n_10421;
wire n_5890;
wire n_6415;
wire n_10976;
wire n_6465;
wire n_9447;
wire n_4439;
wire n_10585;
wire n_4783;
wire n_7931;
wire n_8688;
wire n_10828;
wire n_9092;
wire n_10034;
wire n_9451;
wire n_4910;
wire n_11148;
wire n_3083;
wire n_6899;
wire n_7549;
wire n_10692;
wire n_7373;
wire n_7895;
wire n_6592;
wire n_3049;
wire n_8686;
wire n_8871;
wire n_9712;
wire n_6626;
wire n_8585;
wire n_8951;
wire n_5389;
wire n_5142;
wire n_11114;
wire n_9011;
wire n_8418;
wire n_3830;
wire n_7740;
wire n_8403;
wire n_3679;
wire n_5891;
wire n_7613;
wire n_3541;
wire n_6101;
wire n_9220;
wire n_3117;
wire n_5935;
wire n_7556;
wire n_10528;
wire n_10860;
wire n_4930;
wire n_8588;
wire n_5623;
wire n_8564;
wire n_6944;
wire n_9121;
wire n_10471;
wire n_2385;
wire n_4112;
wire n_9012;
wire n_2396;
wire n_4557;
wire n_4917;
wire n_8698;
wire n_8924;
wire n_3739;
wire n_4432;
wire n_2450;
wire n_2284;
wire n_10376;
wire n_4352;
wire n_7515;
wire n_6928;
wire n_4416;
wire n_10880;
wire n_4593;
wire n_7238;
wire n_9994;
wire n_2769;
wire n_4465;
wire n_3622;
wire n_8780;
wire n_7309;
wire n_5114;
wire n_7958;
wire n_4980;
wire n_8047;
wire n_8559;
wire n_5693;
wire n_4495;
wire n_6273;
wire n_5117;
wire n_5663;
wire n_7572;
wire n_2463;
wire n_3363;
wire n_8214;
wire n_10224;
wire n_5990;
wire n_7043;
wire n_10777;
wire n_3721;
wire n_3062;
wire n_2679;
wire n_5024;
wire n_9391;
wire n_7760;
wire n_4559;
wire n_8514;
wire n_9134;
wire n_9753;
wire n_8722;
wire n_10214;
wire n_8241;
wire n_8589;
wire n_3969;
wire n_3336;
wire n_7573;
wire n_4160;
wire n_8442;
wire n_4231;
wire n_6281;
wire n_10649;
wire n_7364;
wire n_2952;
wire n_5647;
wire n_4256;
wire n_2779;
wire n_4938;
wire n_5396;
wire n_9572;
wire n_8608;
wire n_5203;
wire n_6846;
wire n_6311;
wire n_10469;
wire n_9229;
wire n_11194;
wire n_7590;
wire n_9342;
wire n_2620;
wire n_5162;
wire n_6134;
wire n_9329;
wire n_5426;
wire n_10175;
wire n_5803;
wire n_2430;
wire n_9868;
wire n_5285;
wire n_9602;
wire n_7048;
wire n_6886;
wire n_2721;
wire n_9311;
wire n_4335;
wire n_6593;
wire n_8630;
wire n_2683;
wire n_9884;
wire n_5365;
wire n_9876;
wire n_8583;
wire n_2744;
wire n_4521;
wire n_8145;
wire n_8405;
wire n_10447;
wire n_9260;
wire n_7176;
wire n_8928;
wire n_7682;
wire n_9353;
wire n_6231;
wire n_8948;
wire n_8672;
wire n_10406;
wire n_3204;
wire n_5715;
wire n_4920;
wire n_8295;
wire n_6932;
wire n_6746;
wire n_8447;
wire n_7901;
wire n_5395;
wire n_10522;
wire n_6443;
wire n_5709;
wire n_7658;
wire n_6446;
wire n_10278;
wire n_10055;
wire n_10979;
wire n_7980;
wire n_3802;
wire n_3256;
wire n_6996;
wire n_7218;
wire n_8828;
wire n_9430;
wire n_9750;
wire n_9749;
wire n_2915;
wire n_6749;
wire n_9263;
wire n_11082;
wire n_8440;
wire n_7005;
wire n_10408;
wire n_2802;
wire n_8572;
wire n_10798;
wire n_10965;
wire n_7732;
wire n_6337;
wire n_3643;
wire n_6181;
wire n_7447;
wire n_2425;
wire n_9776;
wire n_6777;
wire n_4265;
wire n_8227;
wire n_2950;
wire n_5634;
wire n_5672;
wire n_8475;
wire n_3060;
wire n_10482;
wire n_3098;
wire n_6924;
wire n_8029;
wire n_9804;
wire n_4105;
wire n_4861;
wire n_9304;
wire n_5799;
wire n_8859;
wire n_8380;
wire n_4064;
wire n_7405;
wire n_4926;
wire n_3123;
wire n_8314;
wire n_3380;
wire n_9386;
wire n_10154;
wire n_5617;
wire n_7922;
wire n_10377;
wire n_5580;
wire n_5266;
wire n_4828;
wire n_10033;
wire n_9926;
wire n_3038;
wire n_11121;
wire n_6310;
wire n_10003;
wire n_8311;
wire n_2523;
wire n_10858;
wire n_10321;
wire n_5450;
wire n_2413;
wire n_3769;
wire n_11147;
wire n_5310;
wire n_9661;
wire n_9843;
wire n_9877;
wire n_8764;
wire n_3863;
wire n_3669;
wire n_6953;
wire n_3130;
wire n_4316;
wire n_5722;
wire n_4640;
wire n_5122;
wire n_5390;
wire n_9901;
wire n_5593;
wire n_2805;
wire n_6683;
wire n_4769;
wire n_10683;
wire n_5764;
wire n_9834;
wire n_8934;
wire n_2282;
wire n_6365;
wire n_4628;
wire n_6920;
wire n_9921;
wire n_8407;
wire n_6229;
wire n_5385;
wire n_8567;
wire n_8729;
wire n_10359;
wire n_5237;
wire n_3344;
wire n_2334;
wire n_5133;
wire n_11042;
wire n_5322;
wire n_6907;
wire n_10726;
wire n_3989;
wire n_7089;
wire n_2490;
wire n_7144;
wire n_7286;
wire n_4460;
wire n_4108;
wire n_8048;
wire n_3786;
wire n_3841;
wire n_7072;
wire n_4254;
wire n_8253;
wire n_6177;
wire n_6332;
wire n_2867;
wire n_2726;
wire n_4303;
wire n_5853;
wire n_8283;
wire n_5982;
wire n_10930;
wire n_8749;
wire n_8088;
wire n_7403;
wire n_10722;
wire n_5011;
wire n_10666;
wire n_7338;
wire n_5917;
wire n_7129;
wire n_3147;
wire n_2662;
wire n_4909;
wire n_6696;
wire n_3925;
wire n_9882;
wire n_9527;
wire n_3180;
wire n_8566;
wire n_7343;
wire n_2795;
wire n_3472;
wire n_8516;
wire n_8302;
wire n_10637;
wire n_8317;
wire n_5376;
wire n_5106;
wire n_6116;
wire n_9205;
wire n_9511;
wire n_8167;
wire n_7859;
wire n_6730;
wire n_7492;
wire n_7872;
wire n_7972;
wire n_4768;
wire n_9071;
wire n_7916;
wire n_3717;
wire n_9368;
wire n_7480;
wire n_7694;
wire n_5561;
wire n_10415;
wire n_5410;
wire n_8944;
wire n_6167;
wire n_8008;
wire n_10023;
wire n_10999;
wire n_6170;
wire n_8109;
wire n_9459;
wire n_5156;
wire n_2553;
wire n_6307;
wire n_10410;
wire n_6094;
wire n_9098;
wire n_7987;
wire n_7483;
wire n_4447;
wire n_9133;
wire n_7434;
wire n_4826;
wire n_3445;
wire n_9009;
wire n_6155;
wire n_7269;
wire n_9777;
wire n_9504;
wire n_8975;
wire n_6267;
wire n_9063;
wire n_7787;
wire n_3903;
wire n_5998;
wire n_2325;
wire n_9268;
wire n_5304;
wire n_3854;
wire n_3235;
wire n_6568;
wire n_8673;
wire n_7507;
wire n_7159;
wire n_5378;
wire n_6028;
wire n_9101;
wire n_10456;
wire n_6261;
wire n_3673;
wire n_4281;
wire n_5916;
wire n_4648;
wire n_10096;
wire n_3094;
wire n_10025;
wire n_10627;
wire n_10475;
wire n_10189;
wire n_8697;
wire n_6299;
wire n_6813;
wire n_8825;
wire n_7425;
wire n_6669;
wire n_8581;
wire n_8266;
wire n_5691;
wire n_4951;
wire n_8981;
wire n_8420;
wire n_4957;
wire n_8297;
wire n_11150;
wire n_3079;
wire n_4360;
wire n_8771;
wire n_10881;
wire n_4039;
wire n_3070;
wire n_3800;
wire n_4566;
wire n_3263;
wire n_6316;
wire n_6292;
wire n_4853;
wire n_9726;
wire n_10404;
wire n_8639;
wire n_8058;
wire n_8138;
wire n_9308;
wire n_3504;
wire n_6638;
wire n_10508;
wire n_7719;
wire n_4272;
wire n_10811;
wire n_8333;
wire n_5615;
wire n_2930;
wire n_6220;
wire n_7562;
wire n_3111;
wire n_7619;
wire n_6985;
wire n_7170;
wire n_9211;
wire n_8176;
wire n_8124;
wire n_8823;
wire n_7366;
wire n_9395;
wire n_5269;
wire n_10891;
wire n_9026;
wire n_3054;
wire n_10803;
wire n_8147;
wire n_5468;
wire n_6188;
wire n_4730;
wire n_5399;
wire n_8127;
wire n_9402;
wire n_5262;
wire n_10700;
wire n_3254;
wire n_3684;
wire n_7938;
wire n_4670;
wire n_10968;
wire n_4882;
wire n_4620;
wire n_3152;
wire n_7935;
wire n_4738;
wire n_5421;
wire n_3579;
wire n_8458;
wire n_6772;
wire n_8113;
wire n_3335;
wire n_9716;
wire n_4177;
wire n_3783;
wire n_3178;
wire n_4127;
wire n_5206;
wire n_6077;
wire n_5713;
wire n_5256;
wire n_6318;
wire n_2353;
wire n_4099;
wire n_7918;
wire n_4517;
wire n_4168;
wire n_5188;
wire n_6916;
wire n_4490;
wire n_6651;
wire n_10290;
wire n_10783;
wire n_10147;
wire n_10725;
wire n_3952;
wire n_7845;
wire n_5550;
wire n_3911;
wire n_8290;
wire n_7536;
wire n_7472;
wire n_9433;
wire n_9737;
wire n_9298;
wire n_4285;
wire n_3465;
wire n_10812;
wire n_6366;
wire n_6230;
wire n_2997;
wire n_6604;
wire n_2386;
wire n_5161;
wire n_5373;
wire n_10001;
wire n_3708;
wire n_11107;
wire n_4078;
wire n_9301;
wire n_3046;
wire n_11088;
wire n_5573;
wire n_2956;
wire n_5939;
wire n_5509;
wire n_5382;
wire n_6391;
wire n_8160;
wire n_10284;
wire n_5659;
wire n_8099;
wire n_8840;
wire n_3619;
wire n_5881;
wire n_8522;
wire n_7222;
wire n_7942;
wire n_6473;
wire n_8578;
wire n_4198;
wire n_2382;
wire n_3754;
wire n_10046;
wire n_2291;
wire n_9083;
wire n_7725;
wire n_2886;
wire n_2974;
wire n_4213;
wire n_10977;
wire n_10397;
wire n_2982;
wire n_6483;
wire n_10615;
wire n_10994;
wire n_4065;
wire n_5863;
wire n_7647;
wire n_8626;
wire n_10385;
wire n_10936;
wire n_2645;
wire n_3904;
wire n_8611;
wire n_8036;
wire n_8819;
wire n_2630;
wire n_9835;
wire n_7300;
wire n_6697;
wire n_9054;
wire n_7875;
wire n_6975;
wire n_2470;
wire n_4446;
wire n_10532;
wire n_4417;
wire n_5466;
wire n_7643;
wire n_11048;
wire n_4733;
wire n_6728;
wire n_6729;
wire n_4764;
wire n_3879;
wire n_2286;
wire n_4743;
wire n_10207;
wire n_3080;
wire n_10401;
wire n_5955;
wire n_7242;
wire n_10013;
wire n_10771;
wire n_2865;
wire n_2825;
wire n_8441;
wire n_6076;
wire n_8933;
wire n_3023;
wire n_3232;
wire n_7778;
wire n_5851;
wire n_7073;
wire n_9755;
wire n_4060;
wire n_5110;
wire n_9774;
wire n_8397;
wire n_4879;
wire n_6390;
wire n_10139;
wire n_5796;
wire n_10104;
wire n_8726;
wire n_2806;
wire n_6665;
wire n_8797;
wire n_10723;
wire n_7224;
wire n_9117;
wire n_9720;
wire n_3028;
wire n_7746;
wire n_3662;
wire n_9381;
wire n_2981;
wire n_6958;
wire n_3076;
wire n_10169;
wire n_7563;
wire n_3624;
wire n_4556;
wire n_6549;
wire n_8414;
wire n_6297;
wire n_6523;
wire n_6653;
wire n_8434;
wire n_10477;
wire n_6096;
wire n_4117;
wire n_7853;
wire n_4687;
wire n_2836;
wire n_7531;
wire n_8890;
wire n_5492;
wire n_5995;
wire n_9965;
wire n_8615;
wire n_11062;
wire n_2378;
wire n_7721;
wire n_7192;
wire n_5905;
wire n_11206;
wire n_9887;
wire n_9149;
wire n_2655;
wire n_4600;
wire n_7035;
wire n_6193;
wire n_6501;
wire n_8316;
wire n_4250;
wire n_9990;
wire n_5829;
wire n_3906;
wire n_10005;
wire n_8057;
wire n_4954;
wire n_5191;
wire n_2599;
wire n_8505;
wire n_9273;
wire n_3963;
wire n_3368;
wire n_7884;
wire n_9345;
wire n_2370;
wire n_2612;
wire n_8970;
wire n_7527;
wire n_7417;
wire n_9682;
wire n_2591;
wire n_4881;
wire n_4253;
wire n_10640;
wire n_6582;
wire n_5734;
wire n_2593;
wire n_4255;
wire n_4071;
wire n_10729;
wire n_7388;
wire n_3568;
wire n_3850;
wire n_9924;
wire n_8717;
wire n_5770;
wire n_2496;
wire n_5705;
wire n_3313;
wire n_4605;
wire n_9064;
wire n_3189;
wire n_7635;
wire n_5525;
wire n_2725;
wire n_2277;
wire n_4691;
wire n_7090;
wire n_9254;
wire n_3943;
wire n_2300;
wire n_8571;
wire n_4305;
wire n_7227;
wire n_10492;
wire n_7415;
wire n_11211;
wire n_6745;
wire n_6972;
wire n_10048;
wire n_4297;
wire n_8030;
wire n_9247;
wire n_6052;
wire n_8378;
wire n_8687;
wire n_2907;
wire n_5374;
wire n_10526;
wire n_5575;
wire n_8725;
wire n_9570;
wire n_5675;
wire n_9738;
wire n_4227;
wire n_2778;
wire n_6240;
wire n_11077;
wire n_8243;
wire n_6347;
wire n_8633;
wire n_5020;
wire n_9593;
wire n_7689;
wire n_9846;
wire n_6511;
wire n_5297;
wire n_7121;
wire n_9469;
wire n_10764;
wire n_9677;
wire n_2961;
wire n_3934;
wire n_4033;
wire n_4415;
wire n_6515;
wire n_7099;
wire n_6804;
wire n_8449;
wire n_6358;
wire n_2669;
wire n_4094;
wire n_6603;
wire n_4765;
wire n_2546;
wire n_3193;
wire n_2522;
wire n_4364;
wire n_7534;
wire n_9406;
wire n_8201;
wire n_8967;
wire n_4354;
wire n_6986;
wire n_4732;
wire n_3912;
wire n_8801;
wire n_9322;
wire n_3118;
wire n_10438;
wire n_5959;
wire n_11201;
wire n_3720;
wire n_10531;
wire n_2529;
wire n_8031;
wire n_8918;
wire n_9348;
wire n_8219;
wire n_8696;
wire n_4745;
wire n_6396;
wire n_8932;
wire n_5642;
wire n_9232;
wire n_10575;
wire n_4581;
wire n_6890;
wire n_11028;
wire n_4377;
wire n_9249;
wire n_7827;
wire n_8180;
wire n_10741;
wire n_6109;
wire n_10760;
wire n_4792;
wire n_9444;
wire n_7731;
wire n_3842;
wire n_10772;
wire n_7114;
wire n_4878;
wire n_3514;
wire n_10915;
wire n_4979;
wire n_9535;
wire n_6770;
wire n_2654;
wire n_3036;
wire n_7943;
wire n_8892;
wire n_5302;
wire n_4511;
wire n_2908;
wire n_9707;
wire n_3357;
wire n_5639;
wire n_5781;
wire n_3895;
wire n_8943;
wire n_8486;
wire n_10279;
wire n_4520;
wire n_5299;
wire n_3455;
wire n_4118;
wire n_4503;
wire n_10680;
wire n_2459;
wire n_10127;
wire n_3599;
wire n_5543;
wire n_5361;
wire n_7081;
wire n_2711;
wire n_7132;
wire n_4199;
wire n_5885;
wire n_6663;
wire n_9723;
wire n_5356;
wire n_4441;
wire n_7319;
wire n_3872;
wire n_3772;
wire n_5458;
wire n_7644;
wire n_11176;
wire n_9883;
wire n_11135;
wire n_8155;
wire n_5668;
wire n_5038;
wire n_5330;
wire n_4585;
wire n_7199;
wire n_2664;
wire n_10039;
wire n_10854;
wire n_5463;
wire n_3022;
wire n_8098;
wire n_8833;
wire n_9191;
wire n_5489;
wire n_5892;
wire n_7828;
wire n_10142;
wire n_4773;
wire n_7940;
wire n_9918;
wire n_7910;
wire n_5654;
wire n_6782;
wire n_6009;
wire n_3281;
wire n_2345;
wire n_9034;
wire n_6503;
wire n_6376;
wire n_4427;
wire n_7084;
wire n_5923;
wire n_9390;
wire n_5113;
wire n_10069;
wire n_5479;
wire n_3549;
wire n_5714;
wire n_8541;
wire n_2804;
wire n_2453;
wire n_8074;
wire n_8485;
wire n_8860;
wire n_5510;
wire n_2676;
wire n_3940;
wire n_6621;
wire n_7001;
wire n_9650;
wire n_4822;
wire n_8271;
wire n_5692;
wire n_8473;
wire n_4800;
wire n_9266;
wire n_3453;
wire n_5555;
wire n_3410;
wire n_10027;
wire n_3768;
wire n_4958;
wire n_2810;
wire n_4043;
wire n_2319;
wire n_5441;
wire n_6783;
wire n_9664;
wire n_6066;
wire n_8699;
wire n_3785;
wire n_6897;
wire n_2963;
wire n_10616;
wire n_8587;
wire n_9619;
wire n_11171;
wire n_5366;
wire n_2602;
wire n_6925;
wire n_6878;
wire n_3873;
wire n_8225;
wire n_9078;
wire n_9536;
wire n_2980;
wire n_4886;
wire n_9931;
wire n_3227;
wire n_2733;
wire n_3289;
wire n_6296;
wire n_9187;
wire n_7708;
wire n_4055;
wire n_10328;
wire n_5968;
wire n_11063;
wire n_2644;
wire n_3326;
wire n_10753;
wire n_6497;
wire n_8319;
wire n_9989;
wire n_4200;
wire n_3460;
wire n_2411;
wire n_7108;
wire n_6470;
wire n_8368;
wire n_9259;
wire n_8322;
wire n_7333;
wire n_6187;
wire n_3519;
wire n_7876;
wire n_8546;
wire n_10963;
wire n_8300;
wire n_7371;
wire n_9378;
wire n_8152;
wire n_10826;
wire n_7463;
wire n_8525;
wire n_6573;
wire n_9656;
wire n_7634;
wire n_5078;
wire n_3707;
wire n_8148;
wire n_8150;
wire n_3578;
wire n_6693;
wire n_10483;
wire n_4737;
wire n_4925;
wire n_9620;
wire n_4116;
wire n_5415;
wire n_8986;
wire n_7285;
wire n_5419;
wire n_3805;
wire n_8929;
wire n_9360;
wire n_7260;
wire n_2943;
wire n_5205;
wire n_6409;
wire n_3252;
wire n_3253;
wire n_7954;
wire n_9824;
wire n_11119;
wire n_2622;
wire n_7951;
wire n_2658;
wire n_7552;
wire n_8096;
wire n_2665;
wire n_8233;
wire n_6130;
wire n_4603;
wire n_7273;
wire n_9683;
wire n_10646;
wire n_7231;
wire n_5080;
wire n_5976;
wire n_3128;
wire n_5732;
wire n_5372;
wire n_2691;
wire n_2913;
wire n_4471;
wire n_7449;
wire n_7772;
wire n_8763;
wire n_2690;
wire n_5208;
wire n_8679;
wire n_7239;
wire n_9848;
wire n_5690;
wire n_9227;
wire n_8187;
wire n_10751;
wire n_7050;
wire n_10240;
wire n_9399;
wire n_8996;
wire n_10691;
wire n_2573;
wire n_2646;
wire n_2535;
wire n_6623;
wire n_9561;
wire n_10378;
wire n_9714;
wire n_9740;
wire n_3078;
wire n_9773;
wire n_2436;
wire n_10313;
wire n_3838;
wire n_5371;
wire n_4651;
wire n_9745;
wire n_3941;
wire n_3793;
wire n_10216;
wire n_8139;
wire n_9764;
wire n_4854;
wire n_5071;
wire n_3789;
wire n_7597;
wire n_5801;
wire n_10150;
wire n_6047;
wire n_8292;
wire n_3037;
wire n_10133;
wire n_3729;
wire n_8601;
wire n_10773;
wire n_4994;
wire n_6652;
wire n_9377;
wire n_2537;
wire n_10971;
wire n_8830;
wire n_4483;
wire n_5347;
wire n_6921;
wire n_6970;
wire n_5168;
wire n_4661;
wire n_4988;
wire n_7674;
wire n_9826;
wire n_3171;
wire n_7568;
wire n_6354;
wire n_7272;
wire n_3608;
wire n_4540;
wire n_6344;
wire n_3459;
wire n_9772;
wire n_2853;
wire n_3053;
wire n_3358;
wire n_6021;
wire n_7949;
wire n_7724;
wire n_3499;
wire n_6624;
wire n_9630;
wire n_6956;
wire n_4284;
wire n_6305;
wire n_9255;
wire n_6209;
wire n_8310;
wire n_10231;
wire n_9758;
wire n_3426;
wire n_4971;
wire n_8936;
wire n_5656;
wire n_7126;
wire n_5125;
wire n_5857;
wire n_7329;
wire n_8646;
wire n_7408;
wire n_9691;
wire n_10259;
wire n_2650;
wire n_7107;
wire n_5652;
wire n_6457;
wire n_8597;
wire n_10488;
wire n_7690;
wire n_8969;
wire n_7123;
wire n_10752;
wire n_5499;
wire n_8117;
wire n_10067;
wire n_3229;
wire n_3348;
wire n_10399;
wire n_10213;
wire n_6950;
wire n_8208;
wire n_10038;
wire n_9048;
wire n_5228;
wire n_11010;
wire n_2933;
wire n_10274;
wire n_9590;
wire n_2717;
wire n_6694;
wire n_3497;
wire n_6880;
wire n_5066;
wire n_7418;
wire n_9168;
wire n_3580;
wire n_2842;
wire n_2335;
wire n_9497;
wire n_8536;
wire n_9435;
wire n_7229;
wire n_8350;
wire n_2307;
wire n_3704;
wire n_9219;
wire n_5507;
wire n_5569;
wire n_8028;
wire n_4280;
wire n_8328;
wire n_8914;
wire n_7258;
wire n_5190;
wire n_8391;
wire n_10579;
wire n_10832;
wire n_3173;
wire n_3677;
wire n_8336;
wire n_6856;
wire n_3996;
wire n_6466;
wire n_7864;
wire n_6727;
wire n_4097;
wire n_10584;
wire n_4218;
wire n_5392;
wire n_2449;
wire n_3880;
wire n_3685;
wire n_8216;
wire n_2868;
wire n_10332;
wire n_7709;
wire n_3609;
wire n_9982;
wire n_10171;
wire n_5455;
wire n_5442;
wire n_6386;
wire n_5948;
wire n_7804;
wire n_4459;
wire n_4545;
wire n_9852;
wire n_6820;
wire n_2896;
wire n_8313;
wire n_3019;
wire n_2639;
wire n_3471;
wire n_5511;
wire n_2898;
wire n_7656;
wire n_6208;
wire n_5295;
wire n_6739;
wire n_2368;
wire n_8041;
wire n_10676;
wire n_8202;
wire n_8263;
wire n_4175;
wire n_10299;
wire n_6438;
wire n_5490;
wire n_10540;
wire n_10374;
wire n_3200;
wire n_4771;
wire n_10200;
wire n_7332;
wire n_3259;
wire n_2524;
wire n_10382;
wire n_3167;
wire n_2460;
wire n_5836;
wire n_7185;
wire n_6291;
wire n_3867;
wire n_10269;
wire n_3593;
wire n_4455;
wire n_8374;
wire n_9169;
wire n_4514;
wire n_5834;
wire n_3191;
wire n_10229;
wire n_5584;
wire n_7512;
wire n_4140;
wire n_2481;
wire n_3561;
wire n_4806;
wire n_7386;
wire n_9939;
wire n_7766;
wire n_10981;
wire n_8738;
wire n_11018;
wire n_9126;
wire n_6469;
wire n_6700;
wire n_2682;
wire n_3032;
wire n_6223;
wire n_6758;
wire n_9438;
wire n_5160;
wire n_7808;
wire n_6544;
wire n_8798;
wire n_9481;
wire n_9600;
wire n_2877;
wire n_9122;
wire n_8085;
wire n_5098;
wire n_8123;
wire n_10344;
wire n_7955;
wire n_5707;
wire n_5140;
wire n_4992;
wire n_5197;
wire n_7287;
wire n_9927;
wire n_5497;
wire n_10076;
wire n_8721;
wire n_6464;
wire n_9912;
wire n_6356;
wire n_3505;
wire n_3540;
wire n_3577;
wire n_7637;
wire n_2432;
wire n_10148;
wire n_10318;
wire n_4796;
wire n_3598;
wire n_4442;
wire n_2581;
wire n_3777;
wire n_3641;
wire n_4203;
wire n_7127;
wire n_4533;
wire n_9635;
wire n_5481;
wire n_3590;
wire n_8666;
wire n_2435;
wire n_5344;
wire n_9264;
wire n_4419;
wire n_8326;
wire n_8670;
wire n_5308;
wire n_5184;
wire n_5794;
wire n_7638;
wire n_5408;
wire n_7801;
wire n_9155;
wire n_4053;
wire n_10234;
wire n_8460;
wire n_3848;
wire n_10416;
wire n_3327;
wire n_8836;
wire n_7959;
wire n_7019;
wire n_8181;
wire n_2701;
wire n_2511;
wire n_8254;
wire n_4167;
wire n_8071;
wire n_2745;
wire n_7735;
wire n_8004;
wire n_6667;
wire n_7409;
wire n_5271;
wire n_10731;
wire n_10583;
wire n_10735;
wire n_9878;
wire n_5964;
wire n_6004;
wire n_10806;
wire n_2323;
wire n_9825;
wire n_2784;
wire n_5494;
wire n_7444;
wire n_5234;
wire n_4431;
wire n_7546;
wire n_2421;
wire n_6272;
wire n_4387;
wire n_2618;
wire n_6588;
wire n_3265;
wire n_2464;
wire n_3755;
wire n_4042;
wire n_5128;
wire n_9001;
wire n_10393;
wire n_2329;
wire n_10513;
wire n_5467;
wire n_10439;
wire n_7296;
wire n_8013;
wire n_4299;
wire n_4890;
wire n_7575;
wire n_3571;
wire n_9045;
wire n_7083;
wire n_2410;
wire n_7720;
wire n_6222;
wire n_9373;
wire n_6268;
wire n_5827;
wire n_4176;
wire n_2929;
wire n_5199;
wire n_6456;
wire n_11103;
wire n_11181;
wire n_9967;
wire n_7521;
wire n_3407;
wire n_5992;
wire n_5313;
wire n_10663;
wire n_3856;
wire n_4236;
wire n_7187;
wire n_9971;
wire n_3425;
wire n_10894;
wire n_3894;
wire n_9524;
wire n_3127;
wire n_2621;
wire n_5312;
wire n_3623;
wire n_6467;
wire n_9182;
wire n_9243;
wire n_9282;
wire n_5079;
wire n_9365;
wire n_6540;
wire n_6625;
wire n_10909;
wire n_6336;
wire n_10083;
wire n_6796;
wire n_2502;
wire n_3646;
wire n_9224;
wire n_10347;
wire n_5513;
wire n_5614;
wire n_6541;
wire n_4830;
wire n_4706;
wire n_5225;
wire n_4570;
wire n_2754;
wire n_2783;
wire n_10208;
wire n_7722;
wire n_3188;
wire n_2462;
wire n_3243;
wire n_2889;
wire n_8487;
wire n_4034;
wire n_4056;
wire n_9240;
wire n_10804;
wire n_8293;
wire n_6486;
wire n_4622;
wire n_3960;
wire n_8141;
wire n_7603;
wire n_10667;
wire n_4887;
wire n_8438;
wire n_10548;
wire n_11020;
wire n_2732;
wire n_4693;
wire n_4206;
wire n_8791;
wire n_10793;
wire n_8288;
wire n_3862;
wire n_4267;
wire n_5835;
wire n_10481;
wire n_6732;
wire n_7979;
wire n_6876;
wire n_2270;
wire n_5049;
wire n_10678;
wire n_6757;
wire n_9573;
wire n_5846;
wire n_2289;
wire n_8323;
wire n_8006;
wire n_8296;
wire n_8657;
wire n_7636;
wire n_9695;
wire n_9799;
wire n_10391;
wire n_2955;
wire n_11083;
wire n_5592;
wire n_6954;
wire n_6938;
wire n_4609;
wire n_7866;
wire n_3051;
wire n_9784;
wire n_11198;
wire n_3367;
wire n_7205;
wire n_8757;
wire n_2328;
wire n_7990;
wire n_7020;
wire n_2859;
wire n_10036;
wire n_5278;
wire n_8596;
wire n_3525;
wire n_5157;
wire n_3314;
wire n_2993;
wire n_3016;
wire n_4754;
wire n_4647;
wire n_9556;
wire n_3688;
wire n_8590;
wire n_8720;
wire n_10261;
wire n_4003;
wire n_5708;
wire n_3751;
wire n_5223;
wire n_6298;
wire n_4894;
wire n_5474;
wire n_4113;
wire n_10813;
wire n_10757;
wire n_4760;
wire n_5649;
wire n_6421;
wire n_7407;
wire n_9827;
wire n_3466;
wire n_10907;
wire n_5704;
wire n_4983;
wire n_7148;
wire n_6328;
wire n_5956;
wire n_5287;
wire n_6236;
wire n_9417;
wire n_5083;
wire n_7214;
wire n_4509;
wire n_6007;
wire n_2875;
wire n_3907;
wire n_6144;
wire n_10135;
wire n_3338;
wire n_4217;
wire n_6197;
wire n_6658;
wire n_4906;
wire n_6835;
wire n_8834;
wire n_3636;
wire n_2327;
wire n_8826;
wire n_5516;
wire n_2841;
wire n_6247;
wire n_7075;
wire n_4897;
wire n_10822;
wire n_10919;
wire n_7104;
wire n_9152;
wire n_7124;
wire n_3539;
wire n_3291;
wire n_7467;
wire n_4399;
wire n_2304;
wire n_7799;
wire n_8364;
wire n_2487;
wire n_5698;
wire n_11092;
wire n_3276;
wire n_2597;
wire n_9534;
wire n_3194;
wire n_5084;
wire n_5771;
wire n_7544;
wire n_9792;
wire n_7513;
wire n_10720;
wire n_9336;
wire n_10535;
wire n_3572;
wire n_6602;
wire n_10924;
wire n_3886;
wire n_6708;
wire n_8854;
wire n_11186;
wire n_8917;
wire n_9647;
wire n_6645;
wire n_9742;
wire n_10727;
wire n_10885;
wire n_6484;
wire n_4710;
wire n_4420;
wire n_3637;
wire n_6242;
wire n_4574;
wire n_2855;
wire n_9312;
wire n_9019;
wire n_8985;
wire n_7692;
wire n_9214;
wire n_5174;
wire n_4234;
wire n_7469;
wire n_5538;
wire n_4101;
wire n_3548;
wire n_7776;
wire n_5017;
wire n_10418;
wire n_10895;
wire n_3974;
wire n_3634;
wire n_10875;
wire n_7560;
wire n_9864;
wire n_8548;
wire n_10672;
wire n_7645;
wire n_3236;
wire n_5096;
wire n_3141;
wire n_2755;
wire n_4660;
wire n_9533;
wire n_9494;
wire n_5241;
wire n_10308;
wire n_9145;
wire n_7082;
wire n_3112;
wire n_10623;
wire n_9754;
wire n_4797;
wire n_3108;
wire n_6285;
wire n_9315;
wire n_4270;
wire n_5428;
wire n_4151;
wire n_7451;
wire n_4945;
wire n_8260;
wire n_3417;
wire n_9000;
wire n_5677;
wire n_9454;
wire n_4124;
wire n_6734;
wire n_7476;
wire n_10864;
wire n_10586;
wire n_5570;
wire n_6418;
wire n_8742;
wire n_8307;
wire n_5153;
wire n_9383;
wire n_9253;
wire n_10571;
wire n_4611;
wire n_8874;
wire n_5927;
wire n_7495;
wire n_7392;
wire n_9566;
wire n_5435;
wire n_2337;
wire n_9765;
wire n_3213;
wire n_9807;
wire n_4333;
wire n_3820;
wire n_5200;
wire n_8706;
wire n_9057;
wire n_6400;
wire n_2607;
wire n_7666;
wire n_7945;
wire n_8894;
wire n_2890;
wire n_5115;
wire n_6941;
wire n_5566;
wire n_7829;
wire n_3249;
wire n_7543;
wire n_8680;
wire n_2722;
wire n_2854;
wire n_7877;
wire n_7963;
wire n_9672;
wire n_2499;
wire n_4152;
wire n_5487;
wire n_8855;
wire n_6398;
wire n_8885;
wire n_10394;
wire n_8329;
wire n_5486;
wire n_9503;
wire n_5092;
wire n_5244;
wire n_3172;
wire n_8270;
wire n_4832;
wire n_2902;
wire n_5889;
wire n_3217;
wire n_7284;
wire n_7264;
wire n_5391;
wire n_9763;
wire n_7737;
wire n_6537;
wire n_8614;
wire n_2472;
wire n_7328;
wire n_10702;
wire n_11070;
wire n_10958;
wire n_9479;
wire n_3394;
wire n_9162;
wire n_9568;
wire n_3536;
wire n_8816;
wire n_3957;
wire n_2894;
wire n_3710;
wire n_9119;
wire n_4195;
wire n_10319;
wire n_5849;
wire n_9654;
wire n_9181;
wire n_4554;
wire n_10322;
wire n_7135;
wire n_6578;
wire n_6224;
wire n_3040;
wire n_8802;
wire n_9859;
wire n_3279;
wire n_8555;
wire n_5240;
wire n_10695;
wire n_8636;
wire n_7024;
wire n_2402;
wire n_6092;
wire n_10879;
wire n_5951;
wire n_6241;
wire n_6589;
wire n_8508;
wire n_6614;
wire n_5912;
wire n_8667;
wire n_3402;
wire n_10639;
wire n_3475;
wire n_3501;
wire n_8121;
wire n_3905;
wire n_8207;
wire n_9645;
wire n_9276;
wire n_8035;
wire n_6735;
wire n_7754;
wire n_4680;
wire n_3013;
wire n_10491;
wire n_2789;
wire n_5152;
wire n_5265;
wire n_9943;
wire n_4927;
wire n_5574;
wire n_9821;
wire n_11112;
wire n_4258;
wire n_2699;
wire n_7152;
wire n_9575;
wire n_6165;
wire n_8320;
wire n_9796;
wire n_10409;
wire n_4548;
wire n_4862;
wire n_10521;
wire n_9610;
wire n_2376;
wire n_5469;
wire n_8766;
wire n_3878;
wire n_6567;
wire n_9165;
wire n_2670;
wire n_2700;
wire n_5910;
wire n_5895;
wire n_5804;
wire n_9508;
wire n_10527;
wire n_3134;
wire n_5965;
wire n_9596;
wire n_3115;
wire n_7240;
wire n_7570;
wire n_4553;
wire n_3278;
wire n_7033;
wire n_4875;
wire n_10476;
wire n_9966;
wire n_7817;
wire n_5682;
wire n_10710;
wire n_5387;
wire n_5557;
wire n_2458;
wire n_8850;
wire n_3050;
wire n_9928;
wire n_2673;
wire n_2456;
wire n_8002;
wire n_9741;
wire n_2527;
wire n_2635;
wire n_3307;
wire n_2871;
wire n_4321;
wire n_10180;
wire n_4183;
wire n_8370;
wire n_7237;
wire n_5681;
wire n_10650;
wire n_9090;
wire n_10157;
wire n_6877;
wire n_7423;
wire n_10402;
wire n_6949;
wire n_7566;
wire n_6119;
wire n_4145;
wire n_4821;
wire n_3121;
wire n_4901;
wire n_9217;
wire n_9261;
wire n_9166;
wire n_4040;
wire n_10518;
wire n_8301;
wire n_2406;
wire n_7617;
wire n_9771;
wire n_5316;
wire n_7718;
wire n_6940;
wire n_9893;
wire n_7396;
wire n_10942;
wire n_5703;
wire n_7835;
wire n_6320;
wire n_8126;
wire n_7998;
wire n_10362;
wire n_9239;
wire n_3930;
wire n_4943;
wire n_10953;
wire n_4757;
wire n_3044;
wire n_7561;
wire n_6810;
wire n_7842;
wire n_2629;
wire n_2809;
wire n_6202;
wire n_9969;
wire n_10099;
wire n_4682;
wire n_9961;
wire n_5564;
wire n_5620;
wire n_7163;
wire n_4530;
wire n_10343;
wire n_10836;
wire n_4942;
wire n_9899;
wire n_9258;
wire n_10181;
wire n_10286;
wire n_5406;
wire n_8072;
wire n_10371;
wire n_2561;
wire n_8277;
wire n_7236;
wire n_4604;
wire n_10257;
wire n_3305;
wire n_7130;
wire n_2992;
wire n_5724;
wire n_7201;
wire n_4841;
wire n_3157;
wire n_10047;
wire n_3221;
wire n_3267;
wire n_2422;
wire n_5806;
wire n_10949;
wire n_4338;
wire n_3457;
wire n_10486;
wire n_3762;
wire n_8724;
wire n_5738;
wire n_3005;
wire n_3151;
wire n_3411;
wire n_4840;
wire n_4519;
wire n_3779;
wire n_2388;
wire n_5355;
wire n_3984;
wire n_5320;
wire n_7491;
wire n_5353;
wire n_9995;
wire n_5186;
wire n_5710;
wire n_9076;
wire n_2417;
wire n_9105;
wire n_6792;
wire n_5093;
wire n_4052;
wire n_9316;
wire n_5979;
wire n_9636;
wire n_9668;
wire n_3558;
wire n_10372;
wire n_7559;
wire n_5438;
wire n_6044;
wire n_8867;
wire n_9491;
wire n_4326;
wire n_2834;
wire n_5517;
wire n_3207;
wire n_5605;
wire n_2441;
wire n_3401;
wire n_10744;
wire n_3242;
wire n_11008;
wire n_9870;
wire n_9833;
wire n_3613;
wire n_6125;
wire n_7314;
wire n_9095;
wire n_4726;
wire n_7678;
wire n_5907;
wire n_6045;
wire n_9914;
wire n_8132;
wire n_6731;
wire n_9178;
wire n_7526;
wire n_5040;
wire n_6063;
wire n_10736;
wire n_10917;
wire n_6504;
wire n_3761;
wire n_4315;
wire n_2888;
wire n_2923;
wire n_7004;
wire n_7821;
wire n_8308;
wire n_6154;
wire n_6943;
wire n_4301;
wire n_10597;
wire n_3744;
wire n_8165;
wire n_4788;
wire n_8400;
wire n_10458;
wire n_8210;
wire n_5977;
wire n_10446;
wire n_7879;
wire n_10271;
wire n_3814;
wire n_3781;
wire n_10888;
wire n_2484;
wire n_10116;
wire n_7696;
wire n_6003;
wire n_6684;
wire n_3843;
wire n_5746;
wire n_6600;
wire n_5451;
wire n_9323;
wire n_3687;
wire n_5402;
wire n_6673;
wire n_10696;
wire n_7355;
wire n_6961;
wire n_3543;
wire n_9331;
wire n_3621;
wire n_6031;
wire n_9922;
wire n_10170;
wire n_8331;
wire n_8217;
wire n_10603;
wire n_6962;
wire n_2903;
wire n_3216;
wire n_3808;
wire n_8858;
wire n_7887;
wire n_7246;
wire n_4365;
wire n_6060;
wire n_7929;
wire n_10255;
wire n_10572;
wire n_3726;
wire n_2369;
wire n_2719;
wire n_7270;
wire n_3758;
wire n_8689;
wire n_10648;
wire n_5417;
wire n_6967;
wire n_2587;
wire n_10113;
wire n_7550;
wire n_3199;
wire n_9760;
wire n_10690;
wire n_3339;
wire n_6742;
wire n_6853;
wire n_10188;
wire n_4923;
wire n_2400;
wire n_5864;
wire n_10686;
wire n_9841;
wire n_6691;
wire n_8743;
wire n_7087;
wire n_8753;
wire n_6191;
wire n_4741;
wire n_10689;
wire n_6172;
wire n_3343;
wire n_10974;
wire n_11067;
wire n_2752;
wire n_8627;
wire n_9513;
wire n_9863;
wire n_4885;
wire n_10233;
wire n_10500;
wire n_10555;
wire n_5432;
wire n_10314;
wire n_4550;
wire n_6988;
wire n_4652;
wire n_10810;
wire n_11075;
wire n_7851;
wire n_6894;
wire n_9791;
wire n_10311;
wire n_9179;
wire n_2358;
wire n_5453;
wire n_3658;
wire n_9140;
wire n_8752;
wire n_6834;
wire n_4900;
wire n_2815;
wire n_3034;
wire n_11177;
wire n_4408;
wire n_4577;
wire n_4748;
wire n_6817;
wire n_5842;
wire n_10937;
wire n_6927;
wire n_5814;
wire n_2814;
wire n_7798;
wire n_5253;
wire n_5209;
wire n_10857;
wire n_6215;
wire n_3231;
wire n_11165;
wire n_4212;
wire n_9736;
wire n_2979;
wire n_5699;
wire n_5531;
wire n_5765;
wire n_2953;
wire n_6517;
wire n_6284;
wire n_4295;
wire n_5943;
wire n_10167;
wire n_7862;
wire n_9225;
wire n_2946;
wire n_2500;
wire n_3430;
wire n_2269;
wire n_10630;
wire n_8105;
wire n_6088;
wire n_9031;
wire n_5777;
wire n_4225;
wire n_6883;
wire n_8808;
wire n_10061;
wire n_10428;
wire n_8528;
wire n_8204;
wire n_11068;
wire n_11035;
wire n_2565;
wire n_5495;
wire n_10694;
wire n_10602;
wire n_7100;
wire n_3583;
wire n_3860;
wire n_11041;
wire n_9420;
wire n_3851;
wire n_5655;
wire n_6393;
wire n_9708;
wire n_5064;
wire n_7825;
wire n_10079;
wire n_7119;
wire n_5610;
wire n_7212;
wire n_8154;
wire n_6966;
wire n_8889;
wire n_3015;
wire n_9790;
wire n_10502;
wire n_11131;
wire n_4009;
wire n_5002;
wire n_5759;
wire n_10778;
wire n_6722;
wire n_6035;
wire n_3473;
wire n_7874;
wire n_8490;
wire n_7622;
wire n_9014;
wire n_10329;
wire n_9979;
wire n_8509;
wire n_8767;
wire n_11123;
wire n_8512;
wire n_9505;
wire n_8634;
wire n_9531;
wire n_2566;
wire n_6364;
wire n_8635;
wire n_2702;
wire n_3241;
wire n_7102;
wire n_7420;
wire n_2906;
wire n_4342;
wire n_10855;
wire n_7995;
wire n_6114;
wire n_4568;
wire n_11003;
wire n_6061;
wire n_10662;
wire n_5559;
wire n_2438;
wire n_6253;
wire n_7831;
wire n_2914;
wire n_10258;
wire n_5786;
wire n_8532;
wire n_10227;
wire n_10588;
wire n_8624;
wire n_8991;
wire n_11022;
wire n_10574;
wire n_8065;
wire n_10247;
wire n_3100;
wire n_11140;
wire n_2858;
wire n_5377;
wire n_3573;
wire n_6201;
wire n_8796;
wire n_4106;
wire n_5737;
wire n_3604;
wire n_10733;
wire n_4373;
wire n_8518;
wire n_8919;
wire n_10472;
wire n_4711;
wire n_3068;
wire n_10066;
wire n_2685;
wire n_6419;
wire n_7784;
wire n_8372;
wire n_9272;
wire n_5768;
wire n_3553;
wire n_10088;
wire n_2465;
wire n_2275;
wire n_7225;
wire n_8077;
wire n_2568;
wire n_3811;
wire n_3494;
wire n_6244;
wire n_9812;
wire n_6900;
wire n_9337;
wire n_3486;
wire n_4086;
wire n_6755;
wire n_7361;
wire n_6565;
wire n_9432;
wire n_9949;
wire n_10289;
wire n_6942;
wire n_7705;
wire n_2265;
wire n_7228;
wire n_5350;
wire n_5470;
wire n_4812;
wire n_7932;
wire n_4409;
wire n_9576;
wire n_7509;
wire n_10145;
wire n_5872;
wire n_6862;
wire n_7058;
wire n_11005;
wire n_5858;
wire n_4629;
wire n_6255;
wire n_4638;
wire n_6840;
wire n_3181;
wire n_6338;
wire n_8262;
wire n_8423;
wire n_5700;
wire n_6037;
wire n_7981;
wire n_9577;
wire n_9874;
wire n_3699;
wire n_4913;
wire n_2312;
wire n_5874;
wire n_6266;
wire n_6488;
wire n_8337;
wire n_7164;
wire n_9231;
wire n_3328;
wire n_6635;
wire n_7973;
wire n_6815;
wire n_3868;
wire n_9569;
wire n_4266;
wire n_8632;
wire n_2466;
wire n_2530;
wire n_7018;
wire n_5873;
wire n_7975;
wire n_9719;
wire n_8358;
wire n_10009;
wire n_9552;
wire n_11100;
wire n_9279;
wire n_6317;
wire n_8199;
wire n_5588;
wire n_2318;
wire n_3286;
wire n_4012;
wire n_3170;
wire n_10443;
wire n_8656;
wire n_7167;
wire n_10756;
wire n_6480;
wire n_3645;
wire n_10918;
wire n_5075;
wire n_3682;
wire n_3304;
wire n_2592;
wire n_4968;
wire n_3771;
wire n_7865;
wire n_2666;
wire n_10384;
wire n_9289;
wire n_2564;
wire n_5085;
wire n_5736;
wire n_4259;
wire n_2433;
wire n_6561;
wire n_7978;
wire n_7820;
wire n_11127;
wire n_10293;
wire n_8881;
wire n_7844;
wire n_7134;
wire n_9633;
wire n_11153;
wire n_3422;
wire n_10074;
wire n_4572;
wire n_4845;
wire n_4104;
wire n_3086;
wire n_9547;
wire n_6875;
wire n_10934;
wire n_10197;
wire n_8346;
wire n_5120;
wire n_3285;
wire n_4208;
wire n_8761;
wire n_9085;
wire n_9632;
wire n_10042;
wire n_8226;
wire n_8402;
wire n_10478;
wire n_7079;
wire n_9690;
wire n_9084;
wire n_5928;
wire n_4089;
wire n_5478;
wire n_6016;
wire n_3219;
wire n_9371;
wire n_3702;
wire n_9711;
wire n_8754;
wire n_9431;
wire n_9847;
wire n_4779;
wire n_7267;
wire n_10367;
wire n_3233;
wire n_4599;
wire n_4437;
wire n_5222;
wire n_9889;
wire n_7316;
wire n_7850;
wire n_10867;
wire n_3310;
wire n_3264;
wire n_7812;
wire n_7103;
wire n_9080;
wire n_4061;
wire n_8133;
wire n_10168;
wire n_7460;
wire n_6176;
wire n_9519;
wire n_6367;
wire n_3881;
wire n_4508;
wire n_4727;
wire n_4594;
wire n_2426;
wire n_10621;
wire n_2478;
wire n_7056;
wire n_9731;
wire n_8193;
wire n_6572;
wire n_8714;
wire n_4429;
wire n_9604;
wire n_7962;
wire n_4642;
wire n_4051;
wire n_7813;
wire n_10085;
wire n_7755;
wire n_7514;
wire n_7649;
wire n_11151;
wire n_6080;
wire n_4865;
wire n_8182;
wire n_8387;
wire n_6078;
wire n_10613;
wire n_10716;
wire n_6056;
wire n_6717;
wire n_5832;
wire n_10664;
wire n_7473;
wire n_7200;
wire n_3206;
wire n_2363;
wire n_2578;
wire n_7688;
wire n_4562;
wire n_3383;
wire n_8707;
wire n_4903;
wire n_3709;
wire n_10561;
wire n_3738;
wire n_9208;
wire n_7611;
wire n_6873;
wire n_4186;
wire n_8494;
wire n_5812;
wire n_2540;
wire n_5743;
wire n_9429;
wire n_8544;
wire n_3610;
wire n_11152;
wire n_4998;
wire n_10749;
wire n_3330;
wire n_7795;
wire n_2879;
wire n_8788;
wire n_4522;
wire n_10122;
wire n_10935;
wire n_7038;
wire n_10992;
wire n_7723;
wire n_4341;
wire n_10160;
wire n_9327;
wire n_10560;
wire n_7404;
wire n_5368;
wire n_4263;
wire n_8177;
wire n_3555;
wire n_9854;
wire n_7059;
wire n_7450;
wire n_8962;
wire n_9538;
wire n_5971;
wire n_6327;
wire n_7362;
wire n_6145;
wire n_3155;
wire n_6539;
wire n_6926;
wire n_3110;
wire n_7271;
wire n_7826;
wire n_9713;
wire n_5933;
wire n_8993;
wire n_6204;
wire n_7076;
wire n_4780;
wire n_10300;
wire n_9588;
wire n_2697;
wire n_3908;
wire n_4973;
wire n_6842;
wire n_3467;
wire n_6866;
wire n_9044;
wire n_3916;
wire n_3527;
wire n_4803;
wire n_2512;
wire n_3950;
wire n_9423;
wire n_9387;
wire n_6030;
wire n_2927;
wire n_4750;
wire n_6451;
wire n_9813;
wire n_3039;
wire n_9127;
wire n_6514;
wire n_3740;
wire n_9794;
wire n_5996;
wire n_2899;
wire n_3186;
wire n_7105;
wire n_10140;
wire n_9244;
wire n_9869;
wire n_11142;
wire n_7049;
wire n_5903;
wire n_5986;
wire n_3065;
wire n_2632;
wire n_6710;
wire n_4984;
wire n_8278;
wire n_2579;
wire n_6345;
wire n_9715;
wire n_8618;
wire n_3387;
wire n_9094;
wire n_5782;
wire n_7535;
wire n_5041;
wire n_3420;
wire n_4275;
wire n_10862;
wire n_4283;
wire n_4959;
wire n_8248;
wire n_8911;
wire n_9056;
wire n_4426;
wire n_9407;
wire n_2912;
wire n_2659;
wire n_4425;
wire n_3409;
wire n_9985;
wire n_4449;
wire n_2320;
wire n_7057;
wire n_3002;
wire n_6957;
wire n_9361;
wire n_4809;
wire n_8495;
wire n_8783;
wire n_3392;
wire n_8529;
wire n_8733;
wire n_8990;
wire n_6050;
wire n_7976;
wire n_6444;
wire n_10254;
wire n_7944;
wire n_11208;
wire n_7262;
wire n_3773;
wire n_8647;
wire n_8574;
wire n_7016;
wire n_10782;
wire n_3301;
wire n_4241;
wire n_10386;
wire n_6379;
wire n_2324;
wire n_5563;
wire n_11026;
wire n_8044;
wire n_2977;
wire n_5840;
wire n_6719;
wire n_7178;
wire n_9439;
wire n_9553;
wire n_2847;
wire n_7506;
wire n_2557;
wire n_8551;
wire n_8330;
wire n_2405;
wire n_4050;
wire n_2647;
wire n_6232;
wire n_9132;
wire n_2336;
wire n_5717;
wire n_6017;
wire n_9696;
wire n_10861;
wire n_2521;
wire n_9120;
wire n_8879;
wire n_11203;
wire n_11159;
wire n_8052;
wire n_4578;
wire n_6362;
wire n_4777;
wire n_5720;
wire n_9332;
wire n_8903;
wire n_11030;
wire n_2672;
wire n_4702;
wire n_2299;
wire n_4179;
wire n_4895;
wire n_5871;
wire n_7142;
wire n_10182;
wire n_6326;
wire n_5898;
wire n_7125;
wire n_6858;
wire n_9252;
wire n_9464;
wire n_6649;
wire n_6283;
wire n_4026;
wire n_10073;
wire n_4531;
wire n_3282;
wire n_3626;
wire n_5072;
wire n_2313;
wire n_11017;
wire n_7241;
wire n_7247;
wire n_10419;
wire n_7172;
wire n_3106;
wire n_10333;
wire n_2344;
wire n_10317;
wire n_2365;
wire n_4666;
wire n_7893;
wire n_6213;
wire n_4029;
wire n_3031;
wire n_7235;
wire n_8540;
wire n_2447;
wire n_6239;
wire n_9915;
wire n_4617;
wire n_2340;
wire n_9325;
wire n_9196;
wire n_4010;
wire n_5896;
wire n_4555;
wire n_5882;
wire n_5940;
wire n_6089;
wire n_5650;
wire n_7588;
wire n_9384;
wire n_4969;
wire n_6057;
wire n_6216;
wire n_10017;
wire n_7340;
wire n_6974;
wire n_11141;
wire n_5105;
wire n_10893;
wire n_4308;
wire n_11093;
wire n_5021;
wire n_9251;
wire n_3463;
wire n_8939;
wire n_9973;
wire n_5263;
wire n_11117;
wire n_2510;
wire n_6713;
wire n_8064;
wire n_9030;
wire n_7657;
wire n_8468;
wire n_2791;
wire n_4325;
wire n_3251;
wire n_4602;
wire n_5044;
wire n_9665;
wire n_10201;
wire n_5134;
wire n_7096;
wire n_3063;
wire n_2729;
wire n_2582;
wire n_8778;
wire n_11197;
wire n_3998;
wire n_7442;
wire n_3632;
wire n_10093;
wire n_3122;
wire n_5567;
wire n_8343;
wire n_6174;
wire n_2730;
wire n_2495;
wire n_7999;
wire n_10128;
wire n_10675;
wire n_6087;
wire n_7593;
wire n_5249;
wire n_2603;
wire n_8068;
wire n_9955;
wire n_3829;
wire n_10539;
wire n_4164;
wire n_5625;
wire n_9007;
wire n_10143;
wire n_7764;
wire n_4919;
wire n_3737;
wire n_10107;
wire n_5969;
wire n_3655;
wire n_10121;
wire n_10196;
wire n_8198;
wire n_3825;
wire n_3225;
wire n_2880;
wire n_7780;
wire n_6828;
wire n_5158;
wire n_7255;
wire n_8693;
wire n_6454;
wire n_5022;
wire n_9270;
wire n_8452;
wire n_7041;
wire n_7307;
wire n_10742;
wire n_5670;
wire n_10829;
wire n_8557;
wire n_6041;
wire n_6918;
wire n_9099;
wire n_9309;
wire n_3296;
wire n_7350;
wire n_10620;
wire n_10303;
wire n_10814;
wire n_5276;
wire n_9627;
wire n_8012;
wire n_7672;
wire n_2551;
wire n_6664;
wire n_5047;
wire n_7318;
wire n_2985;
wire n_6472;
wire n_10218;
wire n_8114;
wire n_3792;
wire n_4202;
wire n_3938;
wire n_4791;
wire n_11154;
wire n_3507;
wire n_5879;
wire n_8062;
wire n_4403;
wire n_5238;
wire n_6166;
wire n_5855;
wire n_3269;
wire n_3531;
wire n_9136;
wire n_6375;
wire n_10975;
wire n_6352;
wire n_9460;
wire n_8542;
wire n_10859;
wire n_7063;
wire n_7047;
wire n_4139;
wire n_6632;
wire n_4549;
wire n_11056;
wire n_8576;
wire n_6238;
wire n_10542;
wire n_8038;
wire n_2397;
wire n_3931;
wire n_4349;
wire n_10681;
wire n_6081;
wire n_9732;
wire n_10459;
wire n_5141;
wire n_3603;
wire n_10222;
wire n_6724;
wire n_10524;
wire n_5429;
wire n_6545;
wire n_8716;
wire n_6705;
wire n_3822;
wire n_9766;
wire n_8629;
wire n_4163;
wire n_9517;
wire n_10463;
wire n_5535;
wire n_7074;
wire n_3910;
wire n_3812;
wire n_8734;
wire n_9204;
wire n_9476;
wire n_9689;
wire n_2633;
wire n_10659;
wire n_6591;
wire n_7585;
wire n_4948;
wire n_5268;
wire n_9780;
wire n_6946;
wire n_2696;
wire n_3482;
wire n_4080;
wire n_6002;
wire n_3319;
wire n_10403;
wire n_2273;
wire n_6289;
wire n_7037;
wire n_3748;
wire n_3272;
wire n_6424;
wire n_4941;
wire n_5506;
wire n_5298;
wire n_9025;
wire n_8524;
wire n_3396;
wire n_11210;
wire n_7599;
wire n_7928;
wire n_8768;
wire n_4393;
wire n_10884;
wire n_6532;
wire n_4372;
wire n_7293;
wire n_5640;
wire n_11191;
wire n_7600;
wire n_10547;
wire n_2831;
wire n_4318;
wire n_6778;
wire n_4158;
wire n_3978;
wire n_3317;
wire n_6721;
wire n_5560;
wire n_6644;
wire n_6512;
wire n_5544;
wire n_4074;
wire n_3716;
wire n_4795;
wire n_6108;
wire n_8258;
wire n_10370;
wire n_4918;
wire n_3824;
wire n_9597;
wire n_5067;
wire n_5744;
wire n_4013;
wire n_6703;
wire n_5384;
wire n_4544;
wire n_3248;
wire n_5841;
wire n_7614;
wire n_9343;
wire n_2941;
wire n_7839;
wire n_5108;
wire n_8299;
wire n_7347;
wire n_4032;
wire n_6086;
wire n_9837;
wire n_11057;
wire n_2355;
wire n_4147;
wire n_10896;
wire n_10969;
wire n_4477;
wire n_3168;
wire n_7383;
wire n_2751;
wire n_6805;
wire n_4337;
wire n_8863;
wire n_4130;
wire n_10562;
wire n_5941;
wire n_7759;
wire n_10210;
wire n_5611;
wire n_3601;
wire n_6340;
wire n_10054;
wire n_3092;
wire n_6219;
wire n_3055;
wire n_6706;
wire n_7479;
wire n_3966;
wire n_10355;
wire n_9692;
wire n_2866;
wire n_7395;
wire n_10598;
wire n_8947;
wire n_4742;
wire n_3734;
wire n_9609;
wire n_10717;
wire n_11118;
wire n_10029;
wire n_7078;
wire n_8188;
wire n_2580;
wire n_6761;
wire n_8972;
wire n_10007;
wire n_3649;
wire n_2821;
wire n_5701;
wire n_3746;
wire n_6067;
wire n_10801;
wire n_9206;
wire n_8510;
wire n_3384;
wire n_9567;
wire n_6811;
wire n_9061;
wire n_3419;
wire n_9942;
wire n_9703;
wire n_4478;
wire n_7372;
wire n_2818;
wire n_5367;
wire n_3794;
wire n_3921;
wire n_6868;
wire n_8664;
wire n_10704;
wire n_4838;
wire n_5970;
wire n_7174;
wire n_9421;
wire n_5202;
wire n_10740;
wire n_10457;
wire n_4965;
wire n_8021;
wire n_3346;
wire n_9705;
wire n_7803;
wire n_11012;
wire n_2965;
wire n_6111;
wire n_3058;
wire n_9624;
wire n_3861;
wire n_9701;
wire n_10389;
wire n_3891;
wire n_6659;
wire n_4523;
wire n_9709;
wire n_6011;
wire n_9295;
wire n_9416;
wire n_4371;
wire n_6225;
wire n_10990;
wire n_2994;
wire n_5502;
wire n_3428;
wire n_3153;
wire n_4552;
wire n_6218;
wire n_3689;
wire n_8982;
wire n_9929;
wire n_10264;
wire n_5850;
wire n_4673;
wire n_2519;
wire n_9953;
wire n_7086;
wire n_3415;
wire n_6648;
wire n_4607;
wire n_10955;
wire n_7226;
wire n_6182;
wire n_7927;
wire n_9013;
wire n_4041;
wire n_2947;
wire n_6520;
wire n_3918;
wire n_9634;
wire n_9532;
wire n_11011;
wire n_5876;
wire n_9998;
wire n_5521;
wire n_4837;
wire n_2476;
wire n_9850;
wire n_6601;
wire n_10916;
wire n_8584;
wire n_9346;
wire n_7920;
wire n_7810;
wire n_8501;
wire n_4169;
wire n_8480;
wire n_10301;
wire n_3271;
wire n_5088;
wire n_4248;
wire n_8034;
wire n_7025;
wire n_9364;
wire n_8228;
wire n_2976;
wire n_2652;
wire n_8076;
wire n_10440;
wire n_6826;
wire n_5856;
wire n_8484;
wire n_9472;
wire n_9836;
wire n_2497;
wire n_10929;
wire n_9107;
wire n_3809;
wire n_3139;
wire n_8100;
wire n_4070;
wire n_10837;
wire n_3545;
wire n_3885;
wire n_10554;
wire n_8014;
wire n_3993;
wire n_8994;
wire n_8091;
wire n_8413;
wire n_4685;
wire n_4031;
wire n_5837;
wire n_4675;
wire n_10149;
wire n_10970;
wire n_7768;
wire n_2663;
wire n_8638;
wire n_5825;
wire n_4018;
wire n_5491;
wire n_2987;
wire n_2938;
wire n_3780;
wire n_5496;
wire n_5802;
wire n_7982;
wire n_8804;
wire n_3337;
wire n_4002;
wire n_3209;
wire n_5178;
wire n_9317;
wire n_9769;
wire n_5547;
wire n_8158;
wire n_2750;
wire n_11167;
wire n_2775;
wire n_6879;
wire n_8469;
wire n_7567;
wire n_10238;
wire n_8765;
wire n_3477;
wire n_8433;
wire n_10102;
wire n_2349;
wire n_8931;
wire n_5596;
wire n_6074;
wire n_2684;
wire n_5983;
wire n_8213;
wire n_3146;
wire n_3953;
wire n_4588;
wire n_10534;
wire n_4653;
wire n_4435;
wire n_10932;
wire n_10619;
wire n_7684;
wire n_11049;
wire n_5604;
wire n_8451;
wire n_5411;
wire n_8334;
wire n_4019;
wire n_8731;
wire n_10589;
wire n_8385;
wire n_10890;
wire n_9156;
wire n_11202;
wire n_4728;
wire n_4999;
wire n_4385;
wire n_6642;
wire n_6847;
wire n_10707;
wire n_4922;
wire n_10552;
wire n_10248;
wire n_5815;
wire n_3616;
wire n_7370;
wire n_9748;
wire n_6595;
wire n_4191;
wire n_7771;
wire n_9350;
wire n_5695;
wire n_6027;
wire n_2870;
wire n_8539;
wire n_10205;
wire n_7026;
wire n_7701;
wire n_7053;
wire n_2341;
wire n_9226;
wire n_3727;
wire n_5235;
wire n_10110;
wire n_2707;
wire n_6306;
wire n_6720;
wire n_10608;
wire n_6888;
wire n_7173;
wire n_4350;
wire n_3747;
wire n_7042;
wire n_8122;
wire n_6095;
wire n_8432;
wire n_5331;
wire n_4330;
wire n_7592;
wire n_5311;
wire n_9528;
wire n_6590;
wire n_10638;
wire n_7583;
wire n_3522;
wire n_6559;
wire n_2747;
wire n_3924;
wire n_9112;
wire n_4621;
wire n_4216;
wire n_5797;
wire n_9235;
wire n_10610;
wire n_11187;
wire n_4240;
wire n_5572;
wire n_3491;
wire n_9333;
wire n_7151;
wire n_4162;
wire n_5565;
wire n_8950;
wire n_2339;
wire n_10758;
wire n_2861;
wire n_10190;
wire n_5520;
wire n_2731;
wire n_3353;
wire n_3975;
wire n_3018;
wire n_5800;
wire n_6562;
wire n_5984;
wire n_6287;
wire n_2638;
wire n_4785;
wire n_8347;
wire n_4683;
wire n_7353;
wire n_9330;
wire n_7758;
wire n_4021;
wire n_2414;
wire n_9490;
wire n_3014;
wire n_2316;
wire n_4103;
wire n_9355;
wire n_11052;
wire n_5060;
wire n_9523;
wire n_3148;
wire n_4022;
wire n_4986;
wire n_5888;
wire n_5669;
wire n_9024;
wire n_9574;
wire n_5772;
wire n_7571;
wire n_9582;
wire n_4775;
wire n_5884;
wire n_10060;
wire n_6671;
wire n_11009;
wire n_6812;
wire n_4864;
wire n_9288;
wire n_9686;
wire n_9488;
wire n_5758;
wire n_10748;
wire n_4674;
wire n_4481;
wire n_6308;
wire n_7897;
wire n_10910;
wire n_10162;
wire n_8242;
wire n_3775;
wire n_4669;
wire n_7118;
wire n_8284;
wire n_9964;
wire n_7792;
wire n_8161;
wire n_9702;
wire n_7510;
wire n_9819;
wire n_6662;
wire n_8184;
wire n_5603;
wire n_9154;
wire n_6525;
wire n_7422;
wire n_3312;
wire n_3835;
wire n_6738;
wire n_4286;
wire n_5763;
wire n_2958;
wire n_8703;
wire n_10014;
wire n_7109;
wire n_3731;
wire n_2936;
wire n_3224;
wire n_6128;
wire n_2489;
wire n_6029;
wire n_8822;
wire n_10677;
wire n_5751;
wire n_2771;
wire n_3020;
wire n_5264;
wire n_4525;
wire n_5924;
wire n_9992;
wire n_7253;
wire n_8384;
wire n_5712;
wire n_6445;
wire n_3557;
wire n_2610;
wire n_3129;
wire n_8476;
wire n_6702;
wire n_3620;
wire n_11179;
wire n_6701;
wire n_7339;
wire n_3832;
wire n_2520;
wire n_8359;
wire n_7380;
wire n_4484;
wire n_3693;
wire n_8736;
wire n_8545;
wire n_9051;
wire n_4497;
wire n_7749;
wire n_10078;
wire n_2372;
wire n_10105;
wire n_9500;
wire n_8705;
wire n_10215;
wire n_7508;
wire n_3674;
wire n_2959;
wire n_2501;
wire n_5694;
wire n_3203;
wire n_9455;
wire n_10251;
wire n_4871;
wire n_8708;
wire n_10834;
wire n_7574;
wire n_2403;
wire n_2837;
wire n_4700;
wire n_4883;
wire n_9980;
wire n_4306;
wire n_4224;
wire n_10706;
wire n_3341;
wire n_6005;
wire n_8872;
wire n_4453;
wire n_9555;
wire n_11133;
wire n_5449;
wire n_3559;
wire n_4005;
wire n_6169;
wire n_8238;
wire n_3546;
wire n_3661;
wire n_7713;
wire n_4564;
wire n_9200;
wire n_5146;
wire n_10709;
wire n_3056;
wire n_2424;
wire n_3201;
wire n_10871;
wire n_3447;
wire n_7352;
wire n_3971;
wire n_5926;
wire n_3103;
wire n_2354;
wire n_4573;
wire n_5398;
wire n_5860;
wire n_10304;
wire n_6936;
wire n_2589;
wire n_4535;
wire n_10244;
wire n_7704;
wire n_7487;
wire n_9986;
wire n_8844;
wire n_6302;
wire n_2442;
wire n_7641;
wire n_3627;
wire n_6106;
wire n_3480;
wire n_7203;
wire n_9397;
wire n_7169;
wire n_10407;
wire n_7670;
wire n_3612;
wire n_9673;
wire n_4695;
wire n_6848;
wire n_2545;
wire n_8642;
wire n_3509;
wire n_10043;
wire n_9855;
wire n_10568;
wire n_5919;
wire n_4368;
wire n_8159;
wire n_8912;
wire n_2966;
wire n_2294;
wire n_7439;
wire n_9496;
wire n_3196;
wire n_8110;
wire n_5319;
wire n_2504;
wire n_10796;
wire n_2623;
wire n_10016;
wire n_9008;
wire n_6343;
wire n_5270;
wire n_10030;
wire n_8805;
wire n_6850;
wire n_5005;
wire n_9653;
wire n_10272;
wire n_8989;
wire n_9640;
wire n_6098;
wire n_6014;
wire n_7209;
wire n_7112;
wire n_2475;
wire n_5181;
wire n_6979;
wire n_7815;
wire n_7934;
wire n_9545;
wire n_3144;
wire n_8111;
wire n_3244;
wire n_9629;
wire n_9603;
wire n_6865;
wire n_10432;
wire n_7276;
wire n_10342;
wire n_8056;
wire n_3287;
wire n_3322;
wire n_5043;
wire n_8739;
wire n_6747;
wire n_9674;
wire n_2357;
wire n_5583;
wire n_4654;
wire n_6433;
wire n_10462;
wire n_3640;
wire n_3481;
wire n_6640;
wire n_8856;
wire n_3033;
wire n_6142;
wire n_9930;
wire n_5775;
wire n_6462;
wire n_7769;
wire n_2374;
wire n_6034;
wire n_9781;
wire n_10291;
wire n_4597;
wire n_9659;
wire n_3364;
wire n_3226;
wire n_4020;
wire n_2780;
wire n_7233;
wire n_8732;
wire n_7602;
wire n_9296;
wire n_7034;
wire n_9897;
wire n_5220;
wire n_9241;
wire n_7390;
wire n_10787;
wire n_4867;
wire n_10669;
wire n_6870;
wire n_6221;
wire n_8231;
wire n_8185;
wire n_6279;
wire n_5061;
wire n_6775;
wire n_9291;
wire n_7881;
wire n_4063;
wire n_9906;
wire n_9369;
wire n_4237;
wire n_2601;
wire n_5029;
wire n_5127;
wire n_6071;
wire n_2920;
wire n_7598;
wire n_9583;
wire n_8908;
wire n_10185;
wire n_11182;
wire n_2648;
wire n_3212;
wire n_10092;
wire n_8220;
wire n_6833;
wire n_6793;
wire n_6767;
wire n_6295;
wire n_3370;
wire n_3386;
wire n_4721;
wire n_3093;
wire n_8090;
wire n_8053;
wire n_10184;
wire n_10111;
wire n_6385;
wire n_9262;
wire n_7426;
wire n_4247;
wire n_8137;
wire n_7045;
wire n_9851;
wire n_3169;
wire n_8740;
wire n_8009;
wire n_7852;
wire n_3205;
wire n_9987;
wire n_10983;
wire n_7984;
wire n_6788;
wire n_7014;
wire n_2720;
wire n_10430;
wire n_8305;
wire n_4614;
wire n_3360;
wire n_10277;
wire n_3956;
wire n_8163;
wire n_4001;
wire n_7220;
wire n_6709;
wire n_2627;
wire n_4422;
wire n_10948;
wire n_6550;
wire n_6712;
wire n_10525;
wire n_9507;
wire n_7416;
wire n_6143;
wire n_3004;
wire n_8841;
wire n_3870;
wire n_5177;
wire n_9657;
wire n_5483;
wire n_3625;
wire n_6743;
wire n_4632;
wire n_10354;
wire n_3084;
wire n_5785;
wire n_2343;
wire n_7465;
wire n_5967;
wire n_4546;
wire n_10049;
wire n_4583;
wire n_4963;
wire n_3749;
wire n_6672;
wire n_9457;
wire n_2942;
wire n_4966;
wire n_9485;
wire n_5780;
wire n_4714;
wire n_7679;
wire n_5037;
wire n_2515;
wire n_7936;
wire n_8966;
wire n_6084;
wire n_4847;
wire n_10287;
wire n_4054;
wire n_8538;
wire n_11039;
wire n_7738;
wire n_2555;
wire n_10119;
wire n_11145;
wire n_3586;
wire n_3653;
wire n_8395;
wire n_10900;
wire n_5966;
wire n_10349;
wire n_6634;
wire n_4668;
wire n_3349;
wire n_5213;
wire n_8961;
wire n_10849;
wire n_7462;
wire n_4635;
wire n_5735;
wire n_7490;
wire n_2278;
wire n_7545;
wire n_10792;
wire n_8625;
wire n_7160;
wire n_7464;
wire n_8937;
wire n_4214;
wire n_9809;
wire n_6919;
wire n_10750;
wire n_3448;
wire n_7805;
wire n_10995;
wire n_7115;
wire n_7295;
wire n_2924;
wire n_9192;
wire n_3595;
wire n_7348;
wire n_5752;
wire n_5360;
wire n_10673;
wire n_6681;
wire n_6104;
wire n_8179;
wire n_10537;
wire n_3991;
wire n_6548;
wire n_3516;
wire n_3926;
wire n_6082;
wire n_6993;
wire n_8511;
wire n_6973;
wire n_10426;
wire n_4405;
wire n_4413;
wire n_9558;
wire n_7453;
wire n_9167;
wire n_8715;
wire n_9655;
wire n_10241;
wire n_4036;
wire n_10684;
wire n_4759;
wire n_7162;
wire n_3670;
wire n_2381;
wire n_4667;
wire n_5081;
wire n_4182;
wire n_3230;
wire n_8371;
wire n_8702;
wire n_8116;
wire n_7946;
wire n_8195;
wire n_8806;
wire n_5877;
wire n_9991;
wire n_7681;
wire n_8845;
wire n_6018;
wire n_6619;
wire n_5189;
wire n_7702;
wire n_6676;
wire n_2819;
wire n_8149;
wire n_10823;
wire n_3041;
wire n_4637;
wire n_9976;
wire n_2423;
wire n_8042;
wire n_10390;
wire n_11106;
wire n_2412;
wire n_8392;
wire n_9560;
wire n_8095;
wire n_7210;
wire n_5869;
wire n_10830;
wire n_2439;
wire n_11132;
wire n_2404;
wire n_6718;
wire n_3635;
wire n_5118;
wire n_7503;
wire n_10824;
wire n_4155;
wire n_6854;
wire n_4238;
wire n_3011;
wire n_2757;
wire n_4977;
wire n_5632;
wire n_8519;
wire n_5582;
wire n_5425;
wire n_5886;
wire n_8269;
wire n_2716;
wire n_6032;
wire n_9047;
wire n_2452;
wire n_3650;
wire n_8968;
wire n_9319;
wire n_9215;
wire n_5446;
wire n_3010;
wire n_7855;
wire n_3043;
wire n_11047;
wire n_8050;
wire n_5224;
wire n_4590;
wire n_8399;
wire n_2543;
wire n_5090;
wire n_3137;
wire n_9599;
wire n_2486;
wire n_3560;
wire n_10985;
wire n_9072;
wire n_3177;
wire n_4929;
wire n_9401;
wire n_5678;
wire n_9428;
wire n_10340;
wire n_10946;
wire n_6981;
wire n_7065;
wire n_2577;
wire n_9216;
wire n_3238;
wire n_3529;
wire n_4835;
wire n_11109;
wire n_11195;
wire n_4038;
wire n_6122;
wire n_2790;
wire n_7911;
wire n_6765;
wire n_9747;
wire n_4565;
wire n_5414;
wire n_4159;
wire n_3784;
wire n_7330;
wire n_5437;
wire n_8883;
wire n_10634;
wire n_8586;
wire n_9202;
wire n_4586;
wire n_11058;
wire n_9058;
wire n_7336;
wire n_2373;
wire n_7446;
wire n_3628;
wire n_8401;
wire n_7854;
wire n_10351;
wire n_5454;
wire n_8186;
wire n_10577;
wire n_4734;
wire n_7493;
wire n_10961;
wire n_10460;
wire n_10780;
wire n_7357;
wire n_8756;
wire n_8737;
wire n_10334;
wire n_4434;
wire n_5307;
wire n_7923;
wire n_10379;
wire n_10151;
wire n_6439;
wire n_4290;
wire n_8602;
wire n_2586;
wire n_2446;
wire n_8240;
wire n_7714;
wire n_5407;
wire n_10411;
wire n_9484;
wire n_10989;
wire n_8422;
wire n_3029;
wire n_10939;
wire n_3597;
wire n_5913;
wire n_7088;
wire n_2560;
wire n_9305;
wire n_9394;
wire n_9999;
wire n_2704;
wire n_8878;
wire n_11144;
wire n_10090;
wire n_6406;
wire n_7440;
wire n_6945;
wire n_8112;
wire n_3790;
wire n_10962;
wire n_7029;
wire n_2766;
wire n_11128;
wire n_9292;
wire n_9622;
wire n_10721;
wire n_8593;
wire n_10186;
wire n_3318;
wire n_4833;
wire n_11025;
wire n_5062;
wire n_6618;
wire n_6474;
wire n_10191;
wire n_5230;
wire n_5944;
wire n_6226;
wire n_4888;
wire n_7317;
wire n_10856;
wire n_6000;
wire n_2479;
wire n_3350;
wire n_2782;
wire n_9584;
wire n_3977;
wire n_8194;
wire n_9461;
wire n_8055;
wire n_11168;
wire n_8579;
wire n_6816;
wire n_10914;
wire n_10911;
wire n_10928;
wire n_8360;
wire n_3588;
wire n_4279;
wire n_5008;
wire n_6425;
wire n_5004;
wire n_5294;
wire n_6493;
wire n_9845;
wire n_6502;
wire n_6250;
wire n_7374;
wire n_6288;
wire n_5974;
wire n_7522;
wire n_6492;
wire n_10071;
wire n_8755;
wire n_4133;
wire n_4527;
wire n_2288;
wire n_6046;
wire n_8251;
wire n_5323;
wire n_3388;
wire n_4790;
wire n_4181;
wire n_3184;
wire n_9618;
wire n_6118;
wire n_5810;
wire n_4561;
wire n_4461;
wire n_3245;
wire n_3075;
wire n_7046;
wire n_11192;
wire n_4007;
wire n_10956;
wire n_4949;
wire n_6852;
wire n_2642;
wire n_4239;
wire n_8677;
wire n_7468;
wire n_9091;
wire n_11013;
wire n_2383;
wire n_5991;
wire n_4184;
wire n_2351;
wire n_5069;
wire n_2986;
wire n_5702;
wire n_10035;
wire n_6251;
wire n_9828;
wire n_3915;
wire n_2536;
wire n_9699;
wire n_3489;
wire n_8108;
wire n_2835;
wire n_5243;
wire n_5914;
wire n_2820;
wire n_2293;
wire n_10252;
wire n_5250;
wire n_3074;
wire n_6869;
wire n_3102;
wire n_10041;
wire n_9321;
wire n_5590;
wire n_10345;
wire n_10059;
wire n_5260;
wire n_8325;
wire n_9751;
wire n_7621;
wire n_7359;
wire n_8498;
wire n_3321;
wire n_2567;
wire n_5809;
wire n_2322;
wire n_10543;
wire n_2727;
wire n_3377;
wire n_7924;
wire n_4782;
wire n_7659;
wire n_2533;
wire n_9005;
wire n_3530;
wire n_9161;
wire n_2869;
wire n_8875;
wire n_4378;
wire n_5349;
wire n_8274;
wire n_9585;
wire n_7153;
wire n_11101;
wire n_2759;
wire n_7836;
wire n_2361;
wire n_10737;
wire n_2266;
wire n_4876;
wire n_6146;
wire n_8504;
wire n_10464;
wire n_7280;
wire n_10644;
wire n_5813;
wire n_9293;
wire n_10365;
wire n_5833;
wire n_2611;
wire n_2901;
wire n_11055;
wire n_7886;
wire n_4358;
wire n_10982;
wire n_5616;
wire n_5805;
wire n_9648;
wire n_2653;
wire n_6884;
wire n_7664;
wire n_7012;
wire n_10591;
wire n_6631;
wire n_4469;
wire n_9498;
wire n_7376;
wire n_7577;
wire n_7308;
wire n_5169;
wire n_5816;
wire n_3156;
wire n_10809;
wire n_8927;
wire n_10899;
wire n_9639;
wire n_10137;
wire n_6228;
wire n_6711;
wire n_3483;
wire n_5416;
wire n_8946;
wire n_4493;
wire n_4924;
wire n_7279;
wire n_7971;
wire n_9646;
wire n_8017;
wire n_8474;
wire n_9984;
wire n_3524;
wire n_7275;
wire n_8232;
wire n_2885;
wire n_8795;
wire n_7195;
wire n_10600;
wire n_10794;
wire n_6102;
wire n_9649;
wire n_8904;
wire n_11199;
wire n_6274;
wire n_10833;
wire n_8838;
wire n_10629;
wire n_9562;
wire n_3097;
wire n_7007;
wire n_7070;
wire n_4539;
wire n_2975;
wire n_8382;
wire n_4421;
wire n_6072;
wire n_7610;
wire n_2839;
wire n_9501;
wire n_2856;
wire n_4793;
wire n_4498;
wire n_10006;
wire n_7259;
wire n_9759;
wire n_6353;
wire n_4953;
wire n_6992;
wire n_11185;
wire n_2348;
wire n_2944;
wire n_8128;
wire n_6818;
wire n_3831;
wire n_10206;
wire n_6322;
wire n_5167;
wire n_5661;
wire n_5932;
wire n_5830;
wire n_3589;
wire n_7539;
wire n_3391;
wire n_8794;
wire n_7616;
wire n_9733;
wire n_8189;
wire n_6498;
wire n_8481;
wire n_10275;
wire n_11081;
wire n_3458;
wire n_7775;
wire n_4505;
wire n_9981;
wire n_3190;
wire n_7930;
wire n_5558;
wire n_8787;
wire n_5687;
wire n_7661;
wire n_6378;
wire n_5383;
wire n_5126;
wire n_8205;
wire n_5051;
wire n_9907;
wire n_5587;
wire n_6976;
wire n_10941;
wire n_11024;
wire n_6304;
wire n_5236;
wire n_7640;
wire n_9816;
wire n_10498;
wire n_5012;
wire n_10292;
wire n_7969;
wire n_6864;
wire n_8605;
wire n_10358;
wire n_3787;
wire n_7548;
wire n_3585;
wire n_10635;
wire n_3565;
wire n_9944;
wire n_4450;
wire n_5954;
wire n_6156;
wire n_5025;
wire n_6998;
wire n_8067;
wire n_7587;
wire n_7064;
wire n_4173;
wire n_3135;
wire n_9643;
wire n_7615;
wire n_5651;
wire n_6930;
wire n_4630;
wire n_9605;
wire n_8000;
wire n_10064;
wire n_7197;
wire n_5645;
wire n_9676;
wire n_3990;
wire n_7393;
wire n_6917;
wire n_6937;
wire n_7591;
wire n_9963;
wire n_5766;
wire n_7727;
wire n_7358;
wire n_2796;
wire n_7324;
wire n_2507;
wire n_9950;
wire n_5878;
wire n_5671;
wire n_10152;
wire n_4534;
wire n_6301;
wire n_9788;
wire n_6929;
wire n_8719;
wire n_8045;
wire n_10785;
wire n_7729;
wire n_2787;
wire n_2969;
wire n_2395;
wire n_4494;
wire n_6436;
wire n_5412;
wire n_8209;
wire n_10802;
wire n_2380;
wire n_4786;
wire n_10815;
wire n_7565;
wire n_6699;
wire n_9213;
wire n_4579;
wire n_7291;
wire n_7631;
wire n_8784;
wire n_2290;
wire n_7382;
wire n_4811;
wire n_6874;
wire n_7387;
wire n_6259;
wire n_9212;
wire n_9340;
wire n_9473;
wire n_4857;
wire n_10490;
wire n_7437;
wire n_6677;
wire n_3432;
wire n_2736;
wire n_2883;
wire n_7618;
wire n_4282;
wire n_10647;
wire n_3493;
wire n_9320;
wire n_10523;
wire n_8769;
wire n_6764;
wire n_8575;
wire n_10081;
wire n_3774;
wire n_5733;
wire n_10324;
wire n_6780;
wire n_11189;
wire n_8815;
wire n_2910;
wire n_6620;
wire n_6597;
wire n_9303;
wire n_3268;
wire n_11105;
wire n_3057;
wire n_3701;
wire n_5148;
wire n_8261;
wire n_2584;
wire n_7673;
wire n_6830;
wire n_8655;
wire n_7282;
wire n_2287;
wire n_6586;
wire n_9968;
wire n_10808;
wire n_6333;
wire n_10474;
wire n_7139;
wire n_8745;
wire n_5791;
wire n_5727;
wire n_10657;
wire n_8086;
wire n_5946;
wire n_8789;
wire n_5997;
wire n_2492;
wire n_7953;
wire n_3778;
wire n_6428;
wire n_5328;
wire n_7379;
wire n_10687;
wire n_9722;
wire n_5657;
wire n_8901;
wire n_11078;
wire n_11130;
wire n_8695;
wire n_4974;
wire n_5975;
wire n_4911;
wire n_8173;
wire n_4436;
wire n_8363;
wire n_5119;
wire n_10652;
wire n_4569;
wire n_10545;
wire n_9669;
wire n_8665;
wire n_6510;
wire n_8282;
wire n_3334;
wire n_9388;
wire n_5938;
wire n_6237;
wire n_5602;
wire n_9379;
wire n_5097;
wire n_4985;
wire n_7751;
wire n_10869;
wire n_3823;
wire n_4384;
wire n_3114;
wire n_2741;
wire n_7581;
wire n_6360;
wire n_5246;
wire n_3584;
wire n_10453;
wire n_4858;
wire n_4678;
wire n_9952;
wire n_2649;
wire n_3556;
wire n_9911;
wire n_3836;
wire n_5579;
wire n_8835;
wire n_9256;
wire n_10668;
wire n_10346;
wire n_5750;
wire n_10688;
wire n_4823;
wire n_5831;
wire n_4309;
wire n_4363;
wire n_7742;
wire n_9274;
wire n_10473;
wire n_5107;
wire n_5095;
wire n_3456;
wire n_8493;
wire n_7346;
wire n_10331;
wire n_10957;
wire n_4243;
wire n_7579;
wire n_10352;
wire n_4025;
wire n_11188;
wire n_7428;
wire n_3404;
wire n_5666;
wire n_4059;
wire n_9195;
wire n_10442;
wire n_4121;
wire n_3290;
wire n_8870;
wire n_7150;
wire n_7155;
wire n_8252;
wire n_4313;
wire n_3309;
wire n_3671;
wire n_4142;
wire n_6475;
wire n_7015;
wire n_3982;
wire n_7283;
wire n_7699;
wire n_8507;
wire n_6314;
wire n_8415;
wire n_10632;
wire n_9623;
wire n_6103;
wire n_2609;
wire n_5546;
wire n_7249;
wire n_10713;
wire n_3796;
wire n_6394;
wire n_8781;
wire n_6964;
wire n_3840;
wire n_3461;
wire n_6680;
wire n_3408;
wire n_7985;
wire n_10954;
wire n_4246;
wire n_7432;
wire n_8365;
wire n_3513;
wire n_3690;
wire n_2483;
wire n_4532;
wire n_8893;
wire n_6372;
wire n_3995;
wire n_4076;
wire n_2594;
wire n_5994;
wire n_6495;
wire n_7194;
wire n_9516;
wire n_4244;
wire n_2503;
wire n_4049;
wire n_6752;
wire n_8976;
wire n_6426;
wire n_2600;
wire n_7505;
wire n_5626;
wire n_3508;
wire n_8025;
wire n_8502;
wire n_10165;
wire n_8244;
wire n_10130;
wire n_7612;
wire n_8156;
wire n_7494;
wire n_4353;
wire n_11120;
wire n_9222;
wire n_8435;
wire n_6350;
wire n_8882;
wire n_4787;
wire n_7736;
wire n_10622;
wire n_5633;
wire n_9546;
wire n_5664;
wire n_7589;
wire n_5921;
wire n_6797;
wire n_3596;
wire n_4537;
wire n_4346;
wire n_8759;
wire n_4351;
wire n_6159;
wire n_7177;
wire n_7814;
wire n_8660;
wire n_2429;
wire n_8479;
wire n_2440;
wire n_6054;
wire n_11095;
wire n_3521;
wire n_8723;
wire n_11019;
wire n_8606;
wire n_9663;
wire n_2681;
wire n_6235;
wire n_7843;
wire n_8235;
wire n_2360;
wire n_3764;
wire n_7662;
wire n_4784;
wire n_6152;
wire n_4075;
wire n_9820;
wire n_7773;
wire n_7902;
wire n_5340;
wire n_3947;
wire n_9743;
wire n_6496;
wire n_3066;
wire n_7756;
wire n_2844;
wire n_8342;
wire n_8940;
wire n_2303;
wire n_2285;
wire n_5280;
wire n_8448;
wire n_8472;
wire n_7700;
wire n_4451;
wire n_4332;
wire n_7555;
wire n_10000;
wire n_4538;
wire n_4506;
wire n_10158;
wire n_2742;
wire n_10582;
wire n_3695;
wire n_10427;
wire n_3976;
wire n_10199;
wire n_7988;
wire n_8658;
wire n_3563;
wire n_6513;
wire n_7500;
wire n_2367;
wire n_10246;
wire n_3198;
wire n_3495;
wire n_5925;
wire n_2909;
wire n_9248;
wire n_6138;
wire n_5369;
wire n_8061;
wire n_8866;
wire n_9822;
wire n_10835;
wire n_5730;
wire n_5576;
wire n_11184;
wire n_3359;
wire n_5272;
wire n_10125;
wire n_6330;
wire n_10117;
wire n_9065;
wire n_3187;
wire n_10844;
wire n_3218;
wire n_8457;
wire n_6802;
wire n_10654;
wire n_9153;
wire n_9086;
wire n_10505;
wire n_9339;
wire n_10198;
wire n_6909;
wire n_7157;
wire n_11064;
wire n_6908;
wire n_8237;
wire n_7411;
wire n_9601;
wire n_9093;
wire n_4201;
wire n_4336;
wire n_2968;
wire n_7266;
wire n_8046;
wire n_7871;
wire n_5646;
wire n_11097;
wire n_5624;
wire n_4852;
wire n_4210;
wire n_4981;
wire n_10840;
wire n_6477;
wire n_9746;
wire n_6263;
wire n_10515;
wire n_8073;
wire n_5440;
wire n_2891;
wire n_6490;
wire n_2709;
wire n_8652;
wire n_9198;
wire n_8821;
wire n_7198;
wire n_8335;
wire n_9904;
wire n_10242;
wire n_9142;
wire n_9440;
wire n_10144;
wire n_3955;
wire n_9684;
wire n_2280;
wire n_3945;
wire n_6184;
wire n_5817;
wire n_5214;
wire n_10973;
wire n_2443;
wire n_4936;
wire n_4205;
wire n_9493;
wire n_4763;
wire n_3587;
wire n_4278;
wire n_5586;
wire n_11036;
wire n_8663;
wire n_3433;
wire n_4463;
wire n_7794;
wire n_10267;
wire n_6038;
wire n_10551;
wire n_5861;
wire n_3833;
wire n_10553;
wire n_2774;
wire n_3162;
wire n_8309;
wire n_3333;
wire n_4129;
wire n_5258;
wire n_8945;
wire n_11002;
wire n_6605;
wire n_5032;
wire n_8964;
wire n_10988;
wire n_9032;
wire n_9814;
wire n_6313;
wire n_4804;
wire n_5619;
wire n_6112;
wire n_3965;
wire n_7145;
wire n_9041;
wire n_5859;
wire n_5380;
wire n_4500;
wire n_9245;
wire n_5065;
wire n_5776;
wire n_8166;
wire n_4433;
wire n_3085;
wire n_5606;
wire n_9357;
wire n_5644;
wire n_2813;
wire n_5826;
wire n_10108;
wire n_8960;
wire n_5920;
wire n_2991;
wire n_10307;
wire n_5030;
wire n_4194;
wire n_7994;
wire n_4703;
wire n_8443;
wire n_7349;
wire n_9598;
wire n_8215;
wire n_7715;
wire n_2419;
wire n_6180;
wire n_8683;
wire n_8809;
wire n_5683;
wire n_6349;
wire n_10510;
wire n_2677;
wire n_3182;
wire n_5756;
wire n_5527;
wire n_3283;
wire n_6476;
wire n_8037;
wire n_4030;

CKINVDCx5p33_ASAP7_75t_R g2264 ( 
.A(n_2022),
.Y(n_2264)
);

CKINVDCx5p33_ASAP7_75t_R g2265 ( 
.A(n_1570),
.Y(n_2265)
);

INVx1_ASAP7_75t_L g2266 ( 
.A(n_1835),
.Y(n_2266)
);

INVx1_ASAP7_75t_L g2267 ( 
.A(n_2113),
.Y(n_2267)
);

CKINVDCx5p33_ASAP7_75t_R g2268 ( 
.A(n_56),
.Y(n_2268)
);

CKINVDCx5p33_ASAP7_75t_R g2269 ( 
.A(n_1822),
.Y(n_2269)
);

CKINVDCx5p33_ASAP7_75t_R g2270 ( 
.A(n_1088),
.Y(n_2270)
);

CKINVDCx5p33_ASAP7_75t_R g2271 ( 
.A(n_1391),
.Y(n_2271)
);

INVx1_ASAP7_75t_L g2272 ( 
.A(n_158),
.Y(n_2272)
);

INVxp67_ASAP7_75t_L g2273 ( 
.A(n_787),
.Y(n_2273)
);

CKINVDCx5p33_ASAP7_75t_R g2274 ( 
.A(n_1764),
.Y(n_2274)
);

INVx1_ASAP7_75t_L g2275 ( 
.A(n_2157),
.Y(n_2275)
);

CKINVDCx20_ASAP7_75t_R g2276 ( 
.A(n_2121),
.Y(n_2276)
);

INVx1_ASAP7_75t_L g2277 ( 
.A(n_716),
.Y(n_2277)
);

INVx1_ASAP7_75t_L g2278 ( 
.A(n_713),
.Y(n_2278)
);

INVx1_ASAP7_75t_L g2279 ( 
.A(n_1351),
.Y(n_2279)
);

CKINVDCx20_ASAP7_75t_R g2280 ( 
.A(n_2226),
.Y(n_2280)
);

INVx2_ASAP7_75t_L g2281 ( 
.A(n_1680),
.Y(n_2281)
);

CKINVDCx20_ASAP7_75t_R g2282 ( 
.A(n_1012),
.Y(n_2282)
);

CKINVDCx5p33_ASAP7_75t_R g2283 ( 
.A(n_1825),
.Y(n_2283)
);

CKINVDCx5p33_ASAP7_75t_R g2284 ( 
.A(n_1961),
.Y(n_2284)
);

CKINVDCx5p33_ASAP7_75t_R g2285 ( 
.A(n_2094),
.Y(n_2285)
);

CKINVDCx5p33_ASAP7_75t_R g2286 ( 
.A(n_1734),
.Y(n_2286)
);

CKINVDCx5p33_ASAP7_75t_R g2287 ( 
.A(n_234),
.Y(n_2287)
);

CKINVDCx5p33_ASAP7_75t_R g2288 ( 
.A(n_141),
.Y(n_2288)
);

CKINVDCx5p33_ASAP7_75t_R g2289 ( 
.A(n_178),
.Y(n_2289)
);

CKINVDCx5p33_ASAP7_75t_R g2290 ( 
.A(n_436),
.Y(n_2290)
);

CKINVDCx5p33_ASAP7_75t_R g2291 ( 
.A(n_1871),
.Y(n_2291)
);

CKINVDCx5p33_ASAP7_75t_R g2292 ( 
.A(n_1395),
.Y(n_2292)
);

CKINVDCx5p33_ASAP7_75t_R g2293 ( 
.A(n_762),
.Y(n_2293)
);

HB1xp67_ASAP7_75t_L g2294 ( 
.A(n_349),
.Y(n_2294)
);

INVx1_ASAP7_75t_SL g2295 ( 
.A(n_893),
.Y(n_2295)
);

INVx1_ASAP7_75t_L g2296 ( 
.A(n_2104),
.Y(n_2296)
);

INVx1_ASAP7_75t_L g2297 ( 
.A(n_299),
.Y(n_2297)
);

CKINVDCx5p33_ASAP7_75t_R g2298 ( 
.A(n_754),
.Y(n_2298)
);

CKINVDCx5p33_ASAP7_75t_R g2299 ( 
.A(n_1287),
.Y(n_2299)
);

INVx1_ASAP7_75t_SL g2300 ( 
.A(n_1885),
.Y(n_2300)
);

CKINVDCx5p33_ASAP7_75t_R g2301 ( 
.A(n_31),
.Y(n_2301)
);

CKINVDCx5p33_ASAP7_75t_R g2302 ( 
.A(n_2131),
.Y(n_2302)
);

CKINVDCx5p33_ASAP7_75t_R g2303 ( 
.A(n_1385),
.Y(n_2303)
);

CKINVDCx5p33_ASAP7_75t_R g2304 ( 
.A(n_2147),
.Y(n_2304)
);

CKINVDCx5p33_ASAP7_75t_R g2305 ( 
.A(n_590),
.Y(n_2305)
);

INVx1_ASAP7_75t_SL g2306 ( 
.A(n_600),
.Y(n_2306)
);

CKINVDCx5p33_ASAP7_75t_R g2307 ( 
.A(n_160),
.Y(n_2307)
);

BUFx6f_ASAP7_75t_L g2308 ( 
.A(n_845),
.Y(n_2308)
);

CKINVDCx5p33_ASAP7_75t_R g2309 ( 
.A(n_1733),
.Y(n_2309)
);

CKINVDCx5p33_ASAP7_75t_R g2310 ( 
.A(n_2118),
.Y(n_2310)
);

BUFx3_ASAP7_75t_L g2311 ( 
.A(n_751),
.Y(n_2311)
);

INVxp67_ASAP7_75t_L g2312 ( 
.A(n_1909),
.Y(n_2312)
);

CKINVDCx5p33_ASAP7_75t_R g2313 ( 
.A(n_2154),
.Y(n_2313)
);

INVx1_ASAP7_75t_L g2314 ( 
.A(n_5),
.Y(n_2314)
);

CKINVDCx5p33_ASAP7_75t_R g2315 ( 
.A(n_677),
.Y(n_2315)
);

CKINVDCx5p33_ASAP7_75t_R g2316 ( 
.A(n_259),
.Y(n_2316)
);

INVx2_ASAP7_75t_L g2317 ( 
.A(n_1878),
.Y(n_2317)
);

CKINVDCx5p33_ASAP7_75t_R g2318 ( 
.A(n_1680),
.Y(n_2318)
);

CKINVDCx5p33_ASAP7_75t_R g2319 ( 
.A(n_57),
.Y(n_2319)
);

INVx1_ASAP7_75t_L g2320 ( 
.A(n_2055),
.Y(n_2320)
);

CKINVDCx5p33_ASAP7_75t_R g2321 ( 
.A(n_527),
.Y(n_2321)
);

BUFx6f_ASAP7_75t_L g2322 ( 
.A(n_1859),
.Y(n_2322)
);

CKINVDCx20_ASAP7_75t_R g2323 ( 
.A(n_2123),
.Y(n_2323)
);

INVx1_ASAP7_75t_L g2324 ( 
.A(n_137),
.Y(n_2324)
);

CKINVDCx5p33_ASAP7_75t_R g2325 ( 
.A(n_2170),
.Y(n_2325)
);

CKINVDCx5p33_ASAP7_75t_R g2326 ( 
.A(n_1542),
.Y(n_2326)
);

CKINVDCx16_ASAP7_75t_R g2327 ( 
.A(n_533),
.Y(n_2327)
);

INVx1_ASAP7_75t_L g2328 ( 
.A(n_1606),
.Y(n_2328)
);

BUFx3_ASAP7_75t_L g2329 ( 
.A(n_606),
.Y(n_2329)
);

CKINVDCx5p33_ASAP7_75t_R g2330 ( 
.A(n_1900),
.Y(n_2330)
);

INVx1_ASAP7_75t_L g2331 ( 
.A(n_1200),
.Y(n_2331)
);

CKINVDCx5p33_ASAP7_75t_R g2332 ( 
.A(n_2099),
.Y(n_2332)
);

INVx1_ASAP7_75t_L g2333 ( 
.A(n_884),
.Y(n_2333)
);

INVx1_ASAP7_75t_SL g2334 ( 
.A(n_2061),
.Y(n_2334)
);

INVx1_ASAP7_75t_L g2335 ( 
.A(n_1858),
.Y(n_2335)
);

INVx1_ASAP7_75t_L g2336 ( 
.A(n_153),
.Y(n_2336)
);

BUFx5_ASAP7_75t_L g2337 ( 
.A(n_802),
.Y(n_2337)
);

CKINVDCx5p33_ASAP7_75t_R g2338 ( 
.A(n_327),
.Y(n_2338)
);

CKINVDCx5p33_ASAP7_75t_R g2339 ( 
.A(n_546),
.Y(n_2339)
);

INVx1_ASAP7_75t_L g2340 ( 
.A(n_1454),
.Y(n_2340)
);

CKINVDCx5p33_ASAP7_75t_R g2341 ( 
.A(n_2071),
.Y(n_2341)
);

INVx1_ASAP7_75t_L g2342 ( 
.A(n_1000),
.Y(n_2342)
);

CKINVDCx5p33_ASAP7_75t_R g2343 ( 
.A(n_1173),
.Y(n_2343)
);

CKINVDCx5p33_ASAP7_75t_R g2344 ( 
.A(n_1383),
.Y(n_2344)
);

BUFx10_ASAP7_75t_L g2345 ( 
.A(n_225),
.Y(n_2345)
);

CKINVDCx5p33_ASAP7_75t_R g2346 ( 
.A(n_301),
.Y(n_2346)
);

CKINVDCx20_ASAP7_75t_R g2347 ( 
.A(n_1956),
.Y(n_2347)
);

CKINVDCx5p33_ASAP7_75t_R g2348 ( 
.A(n_265),
.Y(n_2348)
);

CKINVDCx5p33_ASAP7_75t_R g2349 ( 
.A(n_2057),
.Y(n_2349)
);

HB1xp67_ASAP7_75t_L g2350 ( 
.A(n_1480),
.Y(n_2350)
);

INVx1_ASAP7_75t_L g2351 ( 
.A(n_1788),
.Y(n_2351)
);

BUFx6f_ASAP7_75t_L g2352 ( 
.A(n_1007),
.Y(n_2352)
);

CKINVDCx20_ASAP7_75t_R g2353 ( 
.A(n_2240),
.Y(n_2353)
);

BUFx3_ASAP7_75t_L g2354 ( 
.A(n_2159),
.Y(n_2354)
);

BUFx6f_ASAP7_75t_L g2355 ( 
.A(n_1899),
.Y(n_2355)
);

CKINVDCx5p33_ASAP7_75t_R g2356 ( 
.A(n_52),
.Y(n_2356)
);

CKINVDCx5p33_ASAP7_75t_R g2357 ( 
.A(n_2126),
.Y(n_2357)
);

BUFx5_ASAP7_75t_L g2358 ( 
.A(n_970),
.Y(n_2358)
);

INVx1_ASAP7_75t_L g2359 ( 
.A(n_520),
.Y(n_2359)
);

INVx1_ASAP7_75t_L g2360 ( 
.A(n_554),
.Y(n_2360)
);

CKINVDCx5p33_ASAP7_75t_R g2361 ( 
.A(n_907),
.Y(n_2361)
);

INVx1_ASAP7_75t_L g2362 ( 
.A(n_541),
.Y(n_2362)
);

CKINVDCx5p33_ASAP7_75t_R g2363 ( 
.A(n_1483),
.Y(n_2363)
);

BUFx6f_ASAP7_75t_L g2364 ( 
.A(n_1528),
.Y(n_2364)
);

BUFx2_ASAP7_75t_L g2365 ( 
.A(n_1125),
.Y(n_2365)
);

INVx1_ASAP7_75t_L g2366 ( 
.A(n_2065),
.Y(n_2366)
);

CKINVDCx5p33_ASAP7_75t_R g2367 ( 
.A(n_1642),
.Y(n_2367)
);

CKINVDCx5p33_ASAP7_75t_R g2368 ( 
.A(n_893),
.Y(n_2368)
);

CKINVDCx5p33_ASAP7_75t_R g2369 ( 
.A(n_2044),
.Y(n_2369)
);

CKINVDCx20_ASAP7_75t_R g2370 ( 
.A(n_283),
.Y(n_2370)
);

INVx1_ASAP7_75t_L g2371 ( 
.A(n_1691),
.Y(n_2371)
);

INVx1_ASAP7_75t_L g2372 ( 
.A(n_1420),
.Y(n_2372)
);

CKINVDCx5p33_ASAP7_75t_R g2373 ( 
.A(n_1111),
.Y(n_2373)
);

CKINVDCx5p33_ASAP7_75t_R g2374 ( 
.A(n_1065),
.Y(n_2374)
);

CKINVDCx5p33_ASAP7_75t_R g2375 ( 
.A(n_1452),
.Y(n_2375)
);

CKINVDCx5p33_ASAP7_75t_R g2376 ( 
.A(n_275),
.Y(n_2376)
);

INVx2_ASAP7_75t_L g2377 ( 
.A(n_1545),
.Y(n_2377)
);

CKINVDCx5p33_ASAP7_75t_R g2378 ( 
.A(n_738),
.Y(n_2378)
);

CKINVDCx20_ASAP7_75t_R g2379 ( 
.A(n_294),
.Y(n_2379)
);

CKINVDCx5p33_ASAP7_75t_R g2380 ( 
.A(n_1805),
.Y(n_2380)
);

INVx2_ASAP7_75t_L g2381 ( 
.A(n_1219),
.Y(n_2381)
);

CKINVDCx5p33_ASAP7_75t_R g2382 ( 
.A(n_438),
.Y(n_2382)
);

INVx1_ASAP7_75t_L g2383 ( 
.A(n_805),
.Y(n_2383)
);

CKINVDCx5p33_ASAP7_75t_R g2384 ( 
.A(n_974),
.Y(n_2384)
);

INVx1_ASAP7_75t_L g2385 ( 
.A(n_1052),
.Y(n_2385)
);

CKINVDCx5p33_ASAP7_75t_R g2386 ( 
.A(n_268),
.Y(n_2386)
);

INVx2_ASAP7_75t_L g2387 ( 
.A(n_627),
.Y(n_2387)
);

CKINVDCx20_ASAP7_75t_R g2388 ( 
.A(n_1433),
.Y(n_2388)
);

INVx1_ASAP7_75t_L g2389 ( 
.A(n_69),
.Y(n_2389)
);

CKINVDCx5p33_ASAP7_75t_R g2390 ( 
.A(n_2072),
.Y(n_2390)
);

CKINVDCx20_ASAP7_75t_R g2391 ( 
.A(n_1785),
.Y(n_2391)
);

CKINVDCx5p33_ASAP7_75t_R g2392 ( 
.A(n_860),
.Y(n_2392)
);

CKINVDCx5p33_ASAP7_75t_R g2393 ( 
.A(n_1760),
.Y(n_2393)
);

CKINVDCx5p33_ASAP7_75t_R g2394 ( 
.A(n_915),
.Y(n_2394)
);

CKINVDCx5p33_ASAP7_75t_R g2395 ( 
.A(n_1595),
.Y(n_2395)
);

INVx1_ASAP7_75t_L g2396 ( 
.A(n_762),
.Y(n_2396)
);

BUFx3_ASAP7_75t_L g2397 ( 
.A(n_859),
.Y(n_2397)
);

INVx1_ASAP7_75t_L g2398 ( 
.A(n_2067),
.Y(n_2398)
);

INVx1_ASAP7_75t_L g2399 ( 
.A(n_134),
.Y(n_2399)
);

INVx1_ASAP7_75t_SL g2400 ( 
.A(n_1344),
.Y(n_2400)
);

CKINVDCx5p33_ASAP7_75t_R g2401 ( 
.A(n_1260),
.Y(n_2401)
);

INVx2_ASAP7_75t_L g2402 ( 
.A(n_1059),
.Y(n_2402)
);

CKINVDCx5p33_ASAP7_75t_R g2403 ( 
.A(n_1192),
.Y(n_2403)
);

CKINVDCx20_ASAP7_75t_R g2404 ( 
.A(n_2085),
.Y(n_2404)
);

CKINVDCx5p33_ASAP7_75t_R g2405 ( 
.A(n_1591),
.Y(n_2405)
);

INVx1_ASAP7_75t_L g2406 ( 
.A(n_2050),
.Y(n_2406)
);

INVx1_ASAP7_75t_SL g2407 ( 
.A(n_1103),
.Y(n_2407)
);

INVx1_ASAP7_75t_L g2408 ( 
.A(n_1942),
.Y(n_2408)
);

BUFx2_ASAP7_75t_L g2409 ( 
.A(n_1527),
.Y(n_2409)
);

INVx1_ASAP7_75t_L g2410 ( 
.A(n_1285),
.Y(n_2410)
);

BUFx3_ASAP7_75t_L g2411 ( 
.A(n_2136),
.Y(n_2411)
);

CKINVDCx5p33_ASAP7_75t_R g2412 ( 
.A(n_2193),
.Y(n_2412)
);

INVx1_ASAP7_75t_L g2413 ( 
.A(n_850),
.Y(n_2413)
);

INVx1_ASAP7_75t_L g2414 ( 
.A(n_541),
.Y(n_2414)
);

INVx1_ASAP7_75t_L g2415 ( 
.A(n_2222),
.Y(n_2415)
);

BUFx3_ASAP7_75t_L g2416 ( 
.A(n_746),
.Y(n_2416)
);

INVx1_ASAP7_75t_L g2417 ( 
.A(n_1167),
.Y(n_2417)
);

CKINVDCx5p33_ASAP7_75t_R g2418 ( 
.A(n_2079),
.Y(n_2418)
);

CKINVDCx16_ASAP7_75t_R g2419 ( 
.A(n_548),
.Y(n_2419)
);

CKINVDCx5p33_ASAP7_75t_R g2420 ( 
.A(n_413),
.Y(n_2420)
);

CKINVDCx5p33_ASAP7_75t_R g2421 ( 
.A(n_124),
.Y(n_2421)
);

CKINVDCx5p33_ASAP7_75t_R g2422 ( 
.A(n_1308),
.Y(n_2422)
);

INVx1_ASAP7_75t_L g2423 ( 
.A(n_697),
.Y(n_2423)
);

INVx1_ASAP7_75t_L g2424 ( 
.A(n_2082),
.Y(n_2424)
);

CKINVDCx5p33_ASAP7_75t_R g2425 ( 
.A(n_598),
.Y(n_2425)
);

INVx1_ASAP7_75t_L g2426 ( 
.A(n_1426),
.Y(n_2426)
);

BUFx10_ASAP7_75t_L g2427 ( 
.A(n_751),
.Y(n_2427)
);

CKINVDCx5p33_ASAP7_75t_R g2428 ( 
.A(n_14),
.Y(n_2428)
);

CKINVDCx5p33_ASAP7_75t_R g2429 ( 
.A(n_609),
.Y(n_2429)
);

CKINVDCx5p33_ASAP7_75t_R g2430 ( 
.A(n_937),
.Y(n_2430)
);

INVx1_ASAP7_75t_L g2431 ( 
.A(n_1904),
.Y(n_2431)
);

CKINVDCx5p33_ASAP7_75t_R g2432 ( 
.A(n_1123),
.Y(n_2432)
);

INVx1_ASAP7_75t_L g2433 ( 
.A(n_1527),
.Y(n_2433)
);

CKINVDCx20_ASAP7_75t_R g2434 ( 
.A(n_373),
.Y(n_2434)
);

CKINVDCx5p33_ASAP7_75t_R g2435 ( 
.A(n_256),
.Y(n_2435)
);

CKINVDCx5p33_ASAP7_75t_R g2436 ( 
.A(n_1301),
.Y(n_2436)
);

BUFx10_ASAP7_75t_L g2437 ( 
.A(n_1506),
.Y(n_2437)
);

CKINVDCx5p33_ASAP7_75t_R g2438 ( 
.A(n_350),
.Y(n_2438)
);

CKINVDCx5p33_ASAP7_75t_R g2439 ( 
.A(n_396),
.Y(n_2439)
);

CKINVDCx5p33_ASAP7_75t_R g2440 ( 
.A(n_487),
.Y(n_2440)
);

INVx1_ASAP7_75t_L g2441 ( 
.A(n_1298),
.Y(n_2441)
);

BUFx3_ASAP7_75t_L g2442 ( 
.A(n_301),
.Y(n_2442)
);

BUFx2_ASAP7_75t_L g2443 ( 
.A(n_1597),
.Y(n_2443)
);

CKINVDCx5p33_ASAP7_75t_R g2444 ( 
.A(n_1098),
.Y(n_2444)
);

CKINVDCx5p33_ASAP7_75t_R g2445 ( 
.A(n_2110),
.Y(n_2445)
);

CKINVDCx5p33_ASAP7_75t_R g2446 ( 
.A(n_1891),
.Y(n_2446)
);

CKINVDCx5p33_ASAP7_75t_R g2447 ( 
.A(n_1386),
.Y(n_2447)
);

INVx1_ASAP7_75t_SL g2448 ( 
.A(n_853),
.Y(n_2448)
);

BUFx2_ASAP7_75t_L g2449 ( 
.A(n_2076),
.Y(n_2449)
);

INVx1_ASAP7_75t_L g2450 ( 
.A(n_1893),
.Y(n_2450)
);

INVx1_ASAP7_75t_L g2451 ( 
.A(n_543),
.Y(n_2451)
);

CKINVDCx5p33_ASAP7_75t_R g2452 ( 
.A(n_2061),
.Y(n_2452)
);

INVx1_ASAP7_75t_L g2453 ( 
.A(n_907),
.Y(n_2453)
);

BUFx8_ASAP7_75t_SL g2454 ( 
.A(n_1751),
.Y(n_2454)
);

CKINVDCx5p33_ASAP7_75t_R g2455 ( 
.A(n_352),
.Y(n_2455)
);

BUFx10_ASAP7_75t_L g2456 ( 
.A(n_1629),
.Y(n_2456)
);

CKINVDCx5p33_ASAP7_75t_R g2457 ( 
.A(n_1053),
.Y(n_2457)
);

CKINVDCx5p33_ASAP7_75t_R g2458 ( 
.A(n_752),
.Y(n_2458)
);

INVx1_ASAP7_75t_L g2459 ( 
.A(n_1916),
.Y(n_2459)
);

CKINVDCx5p33_ASAP7_75t_R g2460 ( 
.A(n_1486),
.Y(n_2460)
);

INVx1_ASAP7_75t_L g2461 ( 
.A(n_2155),
.Y(n_2461)
);

CKINVDCx5p33_ASAP7_75t_R g2462 ( 
.A(n_272),
.Y(n_2462)
);

INVx2_ASAP7_75t_SL g2463 ( 
.A(n_2205),
.Y(n_2463)
);

CKINVDCx5p33_ASAP7_75t_R g2464 ( 
.A(n_2208),
.Y(n_2464)
);

BUFx6f_ASAP7_75t_L g2465 ( 
.A(n_1342),
.Y(n_2465)
);

INVx2_ASAP7_75t_SL g2466 ( 
.A(n_538),
.Y(n_2466)
);

CKINVDCx5p33_ASAP7_75t_R g2467 ( 
.A(n_1229),
.Y(n_2467)
);

INVx1_ASAP7_75t_L g2468 ( 
.A(n_1444),
.Y(n_2468)
);

CKINVDCx5p33_ASAP7_75t_R g2469 ( 
.A(n_2024),
.Y(n_2469)
);

CKINVDCx5p33_ASAP7_75t_R g2470 ( 
.A(n_369),
.Y(n_2470)
);

BUFx6f_ASAP7_75t_L g2471 ( 
.A(n_2180),
.Y(n_2471)
);

CKINVDCx5p33_ASAP7_75t_R g2472 ( 
.A(n_2175),
.Y(n_2472)
);

CKINVDCx5p33_ASAP7_75t_R g2473 ( 
.A(n_77),
.Y(n_2473)
);

INVx1_ASAP7_75t_L g2474 ( 
.A(n_271),
.Y(n_2474)
);

CKINVDCx5p33_ASAP7_75t_R g2475 ( 
.A(n_714),
.Y(n_2475)
);

CKINVDCx5p33_ASAP7_75t_R g2476 ( 
.A(n_953),
.Y(n_2476)
);

INVx1_ASAP7_75t_L g2477 ( 
.A(n_2026),
.Y(n_2477)
);

BUFx5_ASAP7_75t_L g2478 ( 
.A(n_462),
.Y(n_2478)
);

CKINVDCx5p33_ASAP7_75t_R g2479 ( 
.A(n_1339),
.Y(n_2479)
);

CKINVDCx5p33_ASAP7_75t_R g2480 ( 
.A(n_2255),
.Y(n_2480)
);

BUFx3_ASAP7_75t_L g2481 ( 
.A(n_1433),
.Y(n_2481)
);

INVx1_ASAP7_75t_L g2482 ( 
.A(n_192),
.Y(n_2482)
);

INVx1_ASAP7_75t_L g2483 ( 
.A(n_843),
.Y(n_2483)
);

INVx2_ASAP7_75t_SL g2484 ( 
.A(n_1012),
.Y(n_2484)
);

CKINVDCx5p33_ASAP7_75t_R g2485 ( 
.A(n_1317),
.Y(n_2485)
);

CKINVDCx5p33_ASAP7_75t_R g2486 ( 
.A(n_246),
.Y(n_2486)
);

CKINVDCx5p33_ASAP7_75t_R g2487 ( 
.A(n_1973),
.Y(n_2487)
);

INVx1_ASAP7_75t_SL g2488 ( 
.A(n_2212),
.Y(n_2488)
);

INVx1_ASAP7_75t_L g2489 ( 
.A(n_1991),
.Y(n_2489)
);

CKINVDCx5p33_ASAP7_75t_R g2490 ( 
.A(n_1082),
.Y(n_2490)
);

CKINVDCx5p33_ASAP7_75t_R g2491 ( 
.A(n_1633),
.Y(n_2491)
);

INVx1_ASAP7_75t_L g2492 ( 
.A(n_1244),
.Y(n_2492)
);

CKINVDCx5p33_ASAP7_75t_R g2493 ( 
.A(n_2094),
.Y(n_2493)
);

INVx1_ASAP7_75t_SL g2494 ( 
.A(n_302),
.Y(n_2494)
);

INVx2_ASAP7_75t_SL g2495 ( 
.A(n_2151),
.Y(n_2495)
);

INVx1_ASAP7_75t_L g2496 ( 
.A(n_2008),
.Y(n_2496)
);

INVx2_ASAP7_75t_L g2497 ( 
.A(n_630),
.Y(n_2497)
);

CKINVDCx20_ASAP7_75t_R g2498 ( 
.A(n_1038),
.Y(n_2498)
);

CKINVDCx5p33_ASAP7_75t_R g2499 ( 
.A(n_2041),
.Y(n_2499)
);

INVx1_ASAP7_75t_L g2500 ( 
.A(n_526),
.Y(n_2500)
);

CKINVDCx5p33_ASAP7_75t_R g2501 ( 
.A(n_2066),
.Y(n_2501)
);

CKINVDCx5p33_ASAP7_75t_R g2502 ( 
.A(n_218),
.Y(n_2502)
);

INVx1_ASAP7_75t_L g2503 ( 
.A(n_655),
.Y(n_2503)
);

CKINVDCx5p33_ASAP7_75t_R g2504 ( 
.A(n_1411),
.Y(n_2504)
);

CKINVDCx5p33_ASAP7_75t_R g2505 ( 
.A(n_1347),
.Y(n_2505)
);

INVx2_ASAP7_75t_L g2506 ( 
.A(n_68),
.Y(n_2506)
);

INVx1_ASAP7_75t_L g2507 ( 
.A(n_617),
.Y(n_2507)
);

INVx1_ASAP7_75t_L g2508 ( 
.A(n_340),
.Y(n_2508)
);

CKINVDCx5p33_ASAP7_75t_R g2509 ( 
.A(n_1629),
.Y(n_2509)
);

INVx2_ASAP7_75t_L g2510 ( 
.A(n_437),
.Y(n_2510)
);

INVx1_ASAP7_75t_L g2511 ( 
.A(n_2096),
.Y(n_2511)
);

INVx1_ASAP7_75t_L g2512 ( 
.A(n_1001),
.Y(n_2512)
);

INVx1_ASAP7_75t_L g2513 ( 
.A(n_1732),
.Y(n_2513)
);

CKINVDCx5p33_ASAP7_75t_R g2514 ( 
.A(n_173),
.Y(n_2514)
);

CKINVDCx5p33_ASAP7_75t_R g2515 ( 
.A(n_1679),
.Y(n_2515)
);

INVx1_ASAP7_75t_L g2516 ( 
.A(n_495),
.Y(n_2516)
);

CKINVDCx5p33_ASAP7_75t_R g2517 ( 
.A(n_1067),
.Y(n_2517)
);

INVx2_ASAP7_75t_L g2518 ( 
.A(n_890),
.Y(n_2518)
);

INVx1_ASAP7_75t_L g2519 ( 
.A(n_361),
.Y(n_2519)
);

INVx1_ASAP7_75t_SL g2520 ( 
.A(n_1772),
.Y(n_2520)
);

CKINVDCx20_ASAP7_75t_R g2521 ( 
.A(n_208),
.Y(n_2521)
);

CKINVDCx5p33_ASAP7_75t_R g2522 ( 
.A(n_2164),
.Y(n_2522)
);

INVx1_ASAP7_75t_L g2523 ( 
.A(n_1461),
.Y(n_2523)
);

CKINVDCx5p33_ASAP7_75t_R g2524 ( 
.A(n_1440),
.Y(n_2524)
);

CKINVDCx5p33_ASAP7_75t_R g2525 ( 
.A(n_315),
.Y(n_2525)
);

CKINVDCx5p33_ASAP7_75t_R g2526 ( 
.A(n_2182),
.Y(n_2526)
);

CKINVDCx5p33_ASAP7_75t_R g2527 ( 
.A(n_2243),
.Y(n_2527)
);

CKINVDCx5p33_ASAP7_75t_R g2528 ( 
.A(n_1825),
.Y(n_2528)
);

CKINVDCx20_ASAP7_75t_R g2529 ( 
.A(n_148),
.Y(n_2529)
);

CKINVDCx5p33_ASAP7_75t_R g2530 ( 
.A(n_629),
.Y(n_2530)
);

BUFx6f_ASAP7_75t_L g2531 ( 
.A(n_16),
.Y(n_2531)
);

INVx1_ASAP7_75t_L g2532 ( 
.A(n_1385),
.Y(n_2532)
);

CKINVDCx5p33_ASAP7_75t_R g2533 ( 
.A(n_1941),
.Y(n_2533)
);

CKINVDCx5p33_ASAP7_75t_R g2534 ( 
.A(n_2236),
.Y(n_2534)
);

CKINVDCx5p33_ASAP7_75t_R g2535 ( 
.A(n_1597),
.Y(n_2535)
);

CKINVDCx5p33_ASAP7_75t_R g2536 ( 
.A(n_1179),
.Y(n_2536)
);

CKINVDCx5p33_ASAP7_75t_R g2537 ( 
.A(n_2169),
.Y(n_2537)
);

CKINVDCx5p33_ASAP7_75t_R g2538 ( 
.A(n_1546),
.Y(n_2538)
);

INVx1_ASAP7_75t_L g2539 ( 
.A(n_2245),
.Y(n_2539)
);

BUFx3_ASAP7_75t_L g2540 ( 
.A(n_331),
.Y(n_2540)
);

CKINVDCx5p33_ASAP7_75t_R g2541 ( 
.A(n_415),
.Y(n_2541)
);

CKINVDCx5p33_ASAP7_75t_R g2542 ( 
.A(n_1239),
.Y(n_2542)
);

BUFx10_ASAP7_75t_L g2543 ( 
.A(n_1486),
.Y(n_2543)
);

BUFx3_ASAP7_75t_L g2544 ( 
.A(n_1518),
.Y(n_2544)
);

INVx2_ASAP7_75t_L g2545 ( 
.A(n_958),
.Y(n_2545)
);

BUFx6f_ASAP7_75t_L g2546 ( 
.A(n_1113),
.Y(n_2546)
);

INVx1_ASAP7_75t_L g2547 ( 
.A(n_2032),
.Y(n_2547)
);

CKINVDCx5p33_ASAP7_75t_R g2548 ( 
.A(n_2140),
.Y(n_2548)
);

CKINVDCx20_ASAP7_75t_R g2549 ( 
.A(n_1677),
.Y(n_2549)
);

CKINVDCx5p33_ASAP7_75t_R g2550 ( 
.A(n_1273),
.Y(n_2550)
);

CKINVDCx5p33_ASAP7_75t_R g2551 ( 
.A(n_1452),
.Y(n_2551)
);

INVx1_ASAP7_75t_L g2552 ( 
.A(n_84),
.Y(n_2552)
);

INVx1_ASAP7_75t_L g2553 ( 
.A(n_396),
.Y(n_2553)
);

CKINVDCx5p33_ASAP7_75t_R g2554 ( 
.A(n_2056),
.Y(n_2554)
);

INVx1_ASAP7_75t_L g2555 ( 
.A(n_2010),
.Y(n_2555)
);

CKINVDCx20_ASAP7_75t_R g2556 ( 
.A(n_2130),
.Y(n_2556)
);

INVx1_ASAP7_75t_L g2557 ( 
.A(n_295),
.Y(n_2557)
);

CKINVDCx5p33_ASAP7_75t_R g2558 ( 
.A(n_445),
.Y(n_2558)
);

INVx1_ASAP7_75t_L g2559 ( 
.A(n_179),
.Y(n_2559)
);

CKINVDCx5p33_ASAP7_75t_R g2560 ( 
.A(n_745),
.Y(n_2560)
);

CKINVDCx5p33_ASAP7_75t_R g2561 ( 
.A(n_1299),
.Y(n_2561)
);

CKINVDCx5p33_ASAP7_75t_R g2562 ( 
.A(n_2021),
.Y(n_2562)
);

BUFx8_ASAP7_75t_SL g2563 ( 
.A(n_614),
.Y(n_2563)
);

CKINVDCx5p33_ASAP7_75t_R g2564 ( 
.A(n_1967),
.Y(n_2564)
);

CKINVDCx5p33_ASAP7_75t_R g2565 ( 
.A(n_2244),
.Y(n_2565)
);

INVx1_ASAP7_75t_L g2566 ( 
.A(n_183),
.Y(n_2566)
);

INVx1_ASAP7_75t_L g2567 ( 
.A(n_235),
.Y(n_2567)
);

BUFx3_ASAP7_75t_L g2568 ( 
.A(n_1830),
.Y(n_2568)
);

CKINVDCx5p33_ASAP7_75t_R g2569 ( 
.A(n_604),
.Y(n_2569)
);

CKINVDCx5p33_ASAP7_75t_R g2570 ( 
.A(n_1514),
.Y(n_2570)
);

INVx1_ASAP7_75t_L g2571 ( 
.A(n_2262),
.Y(n_2571)
);

BUFx6f_ASAP7_75t_L g2572 ( 
.A(n_1106),
.Y(n_2572)
);

INVx1_ASAP7_75t_L g2573 ( 
.A(n_2199),
.Y(n_2573)
);

CKINVDCx5p33_ASAP7_75t_R g2574 ( 
.A(n_2183),
.Y(n_2574)
);

CKINVDCx5p33_ASAP7_75t_R g2575 ( 
.A(n_2150),
.Y(n_2575)
);

CKINVDCx5p33_ASAP7_75t_R g2576 ( 
.A(n_2211),
.Y(n_2576)
);

CKINVDCx5p33_ASAP7_75t_R g2577 ( 
.A(n_2152),
.Y(n_2577)
);

CKINVDCx5p33_ASAP7_75t_R g2578 ( 
.A(n_1366),
.Y(n_2578)
);

CKINVDCx5p33_ASAP7_75t_R g2579 ( 
.A(n_333),
.Y(n_2579)
);

BUFx2_ASAP7_75t_L g2580 ( 
.A(n_1832),
.Y(n_2580)
);

INVx1_ASAP7_75t_L g2581 ( 
.A(n_397),
.Y(n_2581)
);

CKINVDCx5p33_ASAP7_75t_R g2582 ( 
.A(n_626),
.Y(n_2582)
);

CKINVDCx5p33_ASAP7_75t_R g2583 ( 
.A(n_456),
.Y(n_2583)
);

INVx1_ASAP7_75t_L g2584 ( 
.A(n_1460),
.Y(n_2584)
);

CKINVDCx5p33_ASAP7_75t_R g2585 ( 
.A(n_1064),
.Y(n_2585)
);

INVx1_ASAP7_75t_L g2586 ( 
.A(n_2188),
.Y(n_2586)
);

INVx1_ASAP7_75t_L g2587 ( 
.A(n_1596),
.Y(n_2587)
);

INVx1_ASAP7_75t_L g2588 ( 
.A(n_1028),
.Y(n_2588)
);

INVx1_ASAP7_75t_L g2589 ( 
.A(n_903),
.Y(n_2589)
);

INVx1_ASAP7_75t_L g2590 ( 
.A(n_1438),
.Y(n_2590)
);

CKINVDCx5p33_ASAP7_75t_R g2591 ( 
.A(n_1300),
.Y(n_2591)
);

CKINVDCx5p33_ASAP7_75t_R g2592 ( 
.A(n_2092),
.Y(n_2592)
);

CKINVDCx5p33_ASAP7_75t_R g2593 ( 
.A(n_2058),
.Y(n_2593)
);

CKINVDCx5p33_ASAP7_75t_R g2594 ( 
.A(n_1682),
.Y(n_2594)
);

CKINVDCx5p33_ASAP7_75t_R g2595 ( 
.A(n_1983),
.Y(n_2595)
);

BUFx3_ASAP7_75t_L g2596 ( 
.A(n_759),
.Y(n_2596)
);

CKINVDCx5p33_ASAP7_75t_R g2597 ( 
.A(n_1199),
.Y(n_2597)
);

INVx1_ASAP7_75t_L g2598 ( 
.A(n_2029),
.Y(n_2598)
);

INVx1_ASAP7_75t_L g2599 ( 
.A(n_1451),
.Y(n_2599)
);

CKINVDCx5p33_ASAP7_75t_R g2600 ( 
.A(n_1539),
.Y(n_2600)
);

BUFx3_ASAP7_75t_L g2601 ( 
.A(n_738),
.Y(n_2601)
);

INVx1_ASAP7_75t_SL g2602 ( 
.A(n_1351),
.Y(n_2602)
);

INVxp67_ASAP7_75t_SL g2603 ( 
.A(n_682),
.Y(n_2603)
);

CKINVDCx16_ASAP7_75t_R g2604 ( 
.A(n_1658),
.Y(n_2604)
);

BUFx6f_ASAP7_75t_L g2605 ( 
.A(n_116),
.Y(n_2605)
);

CKINVDCx20_ASAP7_75t_R g2606 ( 
.A(n_2084),
.Y(n_2606)
);

CKINVDCx5p33_ASAP7_75t_R g2607 ( 
.A(n_531),
.Y(n_2607)
);

CKINVDCx5p33_ASAP7_75t_R g2608 ( 
.A(n_405),
.Y(n_2608)
);

INVx2_ASAP7_75t_SL g2609 ( 
.A(n_170),
.Y(n_2609)
);

CKINVDCx5p33_ASAP7_75t_R g2610 ( 
.A(n_399),
.Y(n_2610)
);

INVx1_ASAP7_75t_L g2611 ( 
.A(n_83),
.Y(n_2611)
);

CKINVDCx5p33_ASAP7_75t_R g2612 ( 
.A(n_155),
.Y(n_2612)
);

CKINVDCx5p33_ASAP7_75t_R g2613 ( 
.A(n_1177),
.Y(n_2613)
);

CKINVDCx5p33_ASAP7_75t_R g2614 ( 
.A(n_949),
.Y(n_2614)
);

INVx1_ASAP7_75t_L g2615 ( 
.A(n_302),
.Y(n_2615)
);

INVx1_ASAP7_75t_L g2616 ( 
.A(n_886),
.Y(n_2616)
);

CKINVDCx5p33_ASAP7_75t_R g2617 ( 
.A(n_2235),
.Y(n_2617)
);

CKINVDCx5p33_ASAP7_75t_R g2618 ( 
.A(n_1923),
.Y(n_2618)
);

CKINVDCx20_ASAP7_75t_R g2619 ( 
.A(n_644),
.Y(n_2619)
);

CKINVDCx5p33_ASAP7_75t_R g2620 ( 
.A(n_2231),
.Y(n_2620)
);

CKINVDCx16_ASAP7_75t_R g2621 ( 
.A(n_1788),
.Y(n_2621)
);

CKINVDCx5p33_ASAP7_75t_R g2622 ( 
.A(n_1919),
.Y(n_2622)
);

CKINVDCx5p33_ASAP7_75t_R g2623 ( 
.A(n_669),
.Y(n_2623)
);

CKINVDCx5p33_ASAP7_75t_R g2624 ( 
.A(n_1374),
.Y(n_2624)
);

INVx1_ASAP7_75t_L g2625 ( 
.A(n_1386),
.Y(n_2625)
);

CKINVDCx5p33_ASAP7_75t_R g2626 ( 
.A(n_1623),
.Y(n_2626)
);

CKINVDCx5p33_ASAP7_75t_R g2627 ( 
.A(n_264),
.Y(n_2627)
);

CKINVDCx5p33_ASAP7_75t_R g2628 ( 
.A(n_318),
.Y(n_2628)
);

CKINVDCx20_ASAP7_75t_R g2629 ( 
.A(n_1925),
.Y(n_2629)
);

INVx1_ASAP7_75t_L g2630 ( 
.A(n_426),
.Y(n_2630)
);

CKINVDCx5p33_ASAP7_75t_R g2631 ( 
.A(n_1549),
.Y(n_2631)
);

INVx1_ASAP7_75t_L g2632 ( 
.A(n_2234),
.Y(n_2632)
);

INVx1_ASAP7_75t_L g2633 ( 
.A(n_1577),
.Y(n_2633)
);

CKINVDCx5p33_ASAP7_75t_R g2634 ( 
.A(n_1110),
.Y(n_2634)
);

CKINVDCx5p33_ASAP7_75t_R g2635 ( 
.A(n_798),
.Y(n_2635)
);

CKINVDCx5p33_ASAP7_75t_R g2636 ( 
.A(n_260),
.Y(n_2636)
);

HB1xp67_ASAP7_75t_L g2637 ( 
.A(n_774),
.Y(n_2637)
);

CKINVDCx5p33_ASAP7_75t_R g2638 ( 
.A(n_2204),
.Y(n_2638)
);

CKINVDCx5p33_ASAP7_75t_R g2639 ( 
.A(n_347),
.Y(n_2639)
);

INVx1_ASAP7_75t_L g2640 ( 
.A(n_1854),
.Y(n_2640)
);

CKINVDCx5p33_ASAP7_75t_R g2641 ( 
.A(n_955),
.Y(n_2641)
);

INVx2_ASAP7_75t_L g2642 ( 
.A(n_1160),
.Y(n_2642)
);

INVx1_ASAP7_75t_L g2643 ( 
.A(n_2212),
.Y(n_2643)
);

CKINVDCx5p33_ASAP7_75t_R g2644 ( 
.A(n_1890),
.Y(n_2644)
);

BUFx6f_ASAP7_75t_L g2645 ( 
.A(n_710),
.Y(n_2645)
);

CKINVDCx5p33_ASAP7_75t_R g2646 ( 
.A(n_1606),
.Y(n_2646)
);

INVx2_ASAP7_75t_L g2647 ( 
.A(n_1018),
.Y(n_2647)
);

CKINVDCx5p33_ASAP7_75t_R g2648 ( 
.A(n_2034),
.Y(n_2648)
);

INVx1_ASAP7_75t_L g2649 ( 
.A(n_2239),
.Y(n_2649)
);

CKINVDCx5p33_ASAP7_75t_R g2650 ( 
.A(n_1355),
.Y(n_2650)
);

CKINVDCx5p33_ASAP7_75t_R g2651 ( 
.A(n_2082),
.Y(n_2651)
);

INVx1_ASAP7_75t_L g2652 ( 
.A(n_495),
.Y(n_2652)
);

INVx1_ASAP7_75t_L g2653 ( 
.A(n_1716),
.Y(n_2653)
);

CKINVDCx5p33_ASAP7_75t_R g2654 ( 
.A(n_1935),
.Y(n_2654)
);

BUFx2_ASAP7_75t_L g2655 ( 
.A(n_2192),
.Y(n_2655)
);

BUFx10_ASAP7_75t_L g2656 ( 
.A(n_186),
.Y(n_2656)
);

CKINVDCx5p33_ASAP7_75t_R g2657 ( 
.A(n_225),
.Y(n_2657)
);

CKINVDCx5p33_ASAP7_75t_R g2658 ( 
.A(n_1202),
.Y(n_2658)
);

CKINVDCx16_ASAP7_75t_R g2659 ( 
.A(n_32),
.Y(n_2659)
);

INVx1_ASAP7_75t_L g2660 ( 
.A(n_1179),
.Y(n_2660)
);

CKINVDCx5p33_ASAP7_75t_R g2661 ( 
.A(n_1940),
.Y(n_2661)
);

INVx1_ASAP7_75t_SL g2662 ( 
.A(n_2127),
.Y(n_2662)
);

INVx1_ASAP7_75t_L g2663 ( 
.A(n_289),
.Y(n_2663)
);

INVx1_ASAP7_75t_L g2664 ( 
.A(n_365),
.Y(n_2664)
);

CKINVDCx5p33_ASAP7_75t_R g2665 ( 
.A(n_1038),
.Y(n_2665)
);

CKINVDCx5p33_ASAP7_75t_R g2666 ( 
.A(n_1219),
.Y(n_2666)
);

INVx1_ASAP7_75t_L g2667 ( 
.A(n_383),
.Y(n_2667)
);

INVx1_ASAP7_75t_L g2668 ( 
.A(n_2068),
.Y(n_2668)
);

CKINVDCx5p33_ASAP7_75t_R g2669 ( 
.A(n_547),
.Y(n_2669)
);

CKINVDCx14_ASAP7_75t_R g2670 ( 
.A(n_2200),
.Y(n_2670)
);

INVx1_ASAP7_75t_L g2671 ( 
.A(n_1881),
.Y(n_2671)
);

BUFx10_ASAP7_75t_L g2672 ( 
.A(n_2225),
.Y(n_2672)
);

CKINVDCx5p33_ASAP7_75t_R g2673 ( 
.A(n_1153),
.Y(n_2673)
);

CKINVDCx5p33_ASAP7_75t_R g2674 ( 
.A(n_655),
.Y(n_2674)
);

CKINVDCx5p33_ASAP7_75t_R g2675 ( 
.A(n_796),
.Y(n_2675)
);

BUFx6f_ASAP7_75t_L g2676 ( 
.A(n_1779),
.Y(n_2676)
);

CKINVDCx5p33_ASAP7_75t_R g2677 ( 
.A(n_1226),
.Y(n_2677)
);

INVx1_ASAP7_75t_L g2678 ( 
.A(n_1398),
.Y(n_2678)
);

CKINVDCx5p33_ASAP7_75t_R g2679 ( 
.A(n_1083),
.Y(n_2679)
);

CKINVDCx20_ASAP7_75t_R g2680 ( 
.A(n_747),
.Y(n_2680)
);

INVx1_ASAP7_75t_L g2681 ( 
.A(n_2240),
.Y(n_2681)
);

INVx2_ASAP7_75t_L g2682 ( 
.A(n_1626),
.Y(n_2682)
);

INVxp67_ASAP7_75t_SL g2683 ( 
.A(n_2064),
.Y(n_2683)
);

CKINVDCx5p33_ASAP7_75t_R g2684 ( 
.A(n_454),
.Y(n_2684)
);

CKINVDCx5p33_ASAP7_75t_R g2685 ( 
.A(n_1656),
.Y(n_2685)
);

INVx2_ASAP7_75t_L g2686 ( 
.A(n_2066),
.Y(n_2686)
);

INVx1_ASAP7_75t_L g2687 ( 
.A(n_2111),
.Y(n_2687)
);

CKINVDCx5p33_ASAP7_75t_R g2688 ( 
.A(n_2145),
.Y(n_2688)
);

INVx2_ASAP7_75t_L g2689 ( 
.A(n_823),
.Y(n_2689)
);

INVx1_ASAP7_75t_L g2690 ( 
.A(n_131),
.Y(n_2690)
);

INVx1_ASAP7_75t_L g2691 ( 
.A(n_586),
.Y(n_2691)
);

INVx1_ASAP7_75t_L g2692 ( 
.A(n_620),
.Y(n_2692)
);

CKINVDCx5p33_ASAP7_75t_R g2693 ( 
.A(n_583),
.Y(n_2693)
);

INVx1_ASAP7_75t_L g2694 ( 
.A(n_874),
.Y(n_2694)
);

CKINVDCx16_ASAP7_75t_R g2695 ( 
.A(n_581),
.Y(n_2695)
);

CKINVDCx5p33_ASAP7_75t_R g2696 ( 
.A(n_334),
.Y(n_2696)
);

CKINVDCx5p33_ASAP7_75t_R g2697 ( 
.A(n_715),
.Y(n_2697)
);

INVx1_ASAP7_75t_L g2698 ( 
.A(n_2116),
.Y(n_2698)
);

INVx1_ASAP7_75t_L g2699 ( 
.A(n_263),
.Y(n_2699)
);

CKINVDCx5p33_ASAP7_75t_R g2700 ( 
.A(n_1619),
.Y(n_2700)
);

CKINVDCx5p33_ASAP7_75t_R g2701 ( 
.A(n_1088),
.Y(n_2701)
);

CKINVDCx5p33_ASAP7_75t_R g2702 ( 
.A(n_2011),
.Y(n_2702)
);

CKINVDCx20_ASAP7_75t_R g2703 ( 
.A(n_2259),
.Y(n_2703)
);

CKINVDCx5p33_ASAP7_75t_R g2704 ( 
.A(n_1406),
.Y(n_2704)
);

CKINVDCx5p33_ASAP7_75t_R g2705 ( 
.A(n_2103),
.Y(n_2705)
);

CKINVDCx5p33_ASAP7_75t_R g2706 ( 
.A(n_2129),
.Y(n_2706)
);

CKINVDCx5p33_ASAP7_75t_R g2707 ( 
.A(n_2218),
.Y(n_2707)
);

BUFx6f_ASAP7_75t_L g2708 ( 
.A(n_2189),
.Y(n_2708)
);

INVx1_ASAP7_75t_L g2709 ( 
.A(n_8),
.Y(n_2709)
);

CKINVDCx5p33_ASAP7_75t_R g2710 ( 
.A(n_1706),
.Y(n_2710)
);

CKINVDCx20_ASAP7_75t_R g2711 ( 
.A(n_1435),
.Y(n_2711)
);

INVx1_ASAP7_75t_L g2712 ( 
.A(n_1406),
.Y(n_2712)
);

CKINVDCx20_ASAP7_75t_R g2713 ( 
.A(n_2015),
.Y(n_2713)
);

INVx1_ASAP7_75t_L g2714 ( 
.A(n_1814),
.Y(n_2714)
);

CKINVDCx5p33_ASAP7_75t_R g2715 ( 
.A(n_2138),
.Y(n_2715)
);

CKINVDCx5p33_ASAP7_75t_R g2716 ( 
.A(n_1202),
.Y(n_2716)
);

INVx1_ASAP7_75t_L g2717 ( 
.A(n_1690),
.Y(n_2717)
);

CKINVDCx5p33_ASAP7_75t_R g2718 ( 
.A(n_496),
.Y(n_2718)
);

CKINVDCx20_ASAP7_75t_R g2719 ( 
.A(n_265),
.Y(n_2719)
);

INVx4_ASAP7_75t_R g2720 ( 
.A(n_2028),
.Y(n_2720)
);

BUFx6f_ASAP7_75t_L g2721 ( 
.A(n_1095),
.Y(n_2721)
);

CKINVDCx5p33_ASAP7_75t_R g2722 ( 
.A(n_998),
.Y(n_2722)
);

CKINVDCx5p33_ASAP7_75t_R g2723 ( 
.A(n_2122),
.Y(n_2723)
);

INVx1_ASAP7_75t_L g2724 ( 
.A(n_2258),
.Y(n_2724)
);

INVx1_ASAP7_75t_L g2725 ( 
.A(n_1542),
.Y(n_2725)
);

CKINVDCx5p33_ASAP7_75t_R g2726 ( 
.A(n_779),
.Y(n_2726)
);

CKINVDCx5p33_ASAP7_75t_R g2727 ( 
.A(n_931),
.Y(n_2727)
);

CKINVDCx5p33_ASAP7_75t_R g2728 ( 
.A(n_158),
.Y(n_2728)
);

CKINVDCx5p33_ASAP7_75t_R g2729 ( 
.A(n_366),
.Y(n_2729)
);

INVx1_ASAP7_75t_L g2730 ( 
.A(n_112),
.Y(n_2730)
);

CKINVDCx5p33_ASAP7_75t_R g2731 ( 
.A(n_573),
.Y(n_2731)
);

INVx2_ASAP7_75t_SL g2732 ( 
.A(n_208),
.Y(n_2732)
);

CKINVDCx5p33_ASAP7_75t_R g2733 ( 
.A(n_1010),
.Y(n_2733)
);

INVx1_ASAP7_75t_L g2734 ( 
.A(n_1678),
.Y(n_2734)
);

CKINVDCx5p33_ASAP7_75t_R g2735 ( 
.A(n_1296),
.Y(n_2735)
);

CKINVDCx5p33_ASAP7_75t_R g2736 ( 
.A(n_203),
.Y(n_2736)
);

CKINVDCx5p33_ASAP7_75t_R g2737 ( 
.A(n_2030),
.Y(n_2737)
);

CKINVDCx5p33_ASAP7_75t_R g2738 ( 
.A(n_2039),
.Y(n_2738)
);

CKINVDCx20_ASAP7_75t_R g2739 ( 
.A(n_774),
.Y(n_2739)
);

CKINVDCx5p33_ASAP7_75t_R g2740 ( 
.A(n_1935),
.Y(n_2740)
);

CKINVDCx5p33_ASAP7_75t_R g2741 ( 
.A(n_2058),
.Y(n_2741)
);

CKINVDCx5p33_ASAP7_75t_R g2742 ( 
.A(n_1185),
.Y(n_2742)
);

CKINVDCx5p33_ASAP7_75t_R g2743 ( 
.A(n_749),
.Y(n_2743)
);

CKINVDCx5p33_ASAP7_75t_R g2744 ( 
.A(n_2077),
.Y(n_2744)
);

INVx1_ASAP7_75t_SL g2745 ( 
.A(n_1604),
.Y(n_2745)
);

CKINVDCx5p33_ASAP7_75t_R g2746 ( 
.A(n_1551),
.Y(n_2746)
);

BUFx10_ASAP7_75t_L g2747 ( 
.A(n_1186),
.Y(n_2747)
);

CKINVDCx5p33_ASAP7_75t_R g2748 ( 
.A(n_1387),
.Y(n_2748)
);

CKINVDCx5p33_ASAP7_75t_R g2749 ( 
.A(n_2036),
.Y(n_2749)
);

BUFx2_ASAP7_75t_L g2750 ( 
.A(n_573),
.Y(n_2750)
);

BUFx8_ASAP7_75t_SL g2751 ( 
.A(n_240),
.Y(n_2751)
);

CKINVDCx5p33_ASAP7_75t_R g2752 ( 
.A(n_1837),
.Y(n_2752)
);

CKINVDCx5p33_ASAP7_75t_R g2753 ( 
.A(n_1576),
.Y(n_2753)
);

BUFx3_ASAP7_75t_L g2754 ( 
.A(n_1425),
.Y(n_2754)
);

CKINVDCx5p33_ASAP7_75t_R g2755 ( 
.A(n_2197),
.Y(n_2755)
);

CKINVDCx5p33_ASAP7_75t_R g2756 ( 
.A(n_437),
.Y(n_2756)
);

INVx1_ASAP7_75t_L g2757 ( 
.A(n_159),
.Y(n_2757)
);

BUFx2_ASAP7_75t_L g2758 ( 
.A(n_1968),
.Y(n_2758)
);

INVx1_ASAP7_75t_L g2759 ( 
.A(n_1989),
.Y(n_2759)
);

CKINVDCx5p33_ASAP7_75t_R g2760 ( 
.A(n_2081),
.Y(n_2760)
);

BUFx2_ASAP7_75t_SL g2761 ( 
.A(n_212),
.Y(n_2761)
);

CKINVDCx5p33_ASAP7_75t_R g2762 ( 
.A(n_177),
.Y(n_2762)
);

BUFx3_ASAP7_75t_L g2763 ( 
.A(n_1838),
.Y(n_2763)
);

BUFx3_ASAP7_75t_L g2764 ( 
.A(n_152),
.Y(n_2764)
);

CKINVDCx5p33_ASAP7_75t_R g2765 ( 
.A(n_1423),
.Y(n_2765)
);

INVx1_ASAP7_75t_L g2766 ( 
.A(n_947),
.Y(n_2766)
);

CKINVDCx5p33_ASAP7_75t_R g2767 ( 
.A(n_2089),
.Y(n_2767)
);

CKINVDCx5p33_ASAP7_75t_R g2768 ( 
.A(n_17),
.Y(n_2768)
);

CKINVDCx5p33_ASAP7_75t_R g2769 ( 
.A(n_1508),
.Y(n_2769)
);

INVx1_ASAP7_75t_L g2770 ( 
.A(n_12),
.Y(n_2770)
);

BUFx5_ASAP7_75t_L g2771 ( 
.A(n_2198),
.Y(n_2771)
);

BUFx6f_ASAP7_75t_L g2772 ( 
.A(n_2011),
.Y(n_2772)
);

CKINVDCx5p33_ASAP7_75t_R g2773 ( 
.A(n_991),
.Y(n_2773)
);

CKINVDCx5p33_ASAP7_75t_R g2774 ( 
.A(n_406),
.Y(n_2774)
);

CKINVDCx5p33_ASAP7_75t_R g2775 ( 
.A(n_2166),
.Y(n_2775)
);

CKINVDCx5p33_ASAP7_75t_R g2776 ( 
.A(n_513),
.Y(n_2776)
);

CKINVDCx5p33_ASAP7_75t_R g2777 ( 
.A(n_2038),
.Y(n_2777)
);

INVx1_ASAP7_75t_L g2778 ( 
.A(n_1057),
.Y(n_2778)
);

CKINVDCx20_ASAP7_75t_R g2779 ( 
.A(n_2010),
.Y(n_2779)
);

CKINVDCx5p33_ASAP7_75t_R g2780 ( 
.A(n_2077),
.Y(n_2780)
);

INVx1_ASAP7_75t_L g2781 ( 
.A(n_2031),
.Y(n_2781)
);

CKINVDCx5p33_ASAP7_75t_R g2782 ( 
.A(n_916),
.Y(n_2782)
);

CKINVDCx5p33_ASAP7_75t_R g2783 ( 
.A(n_836),
.Y(n_2783)
);

CKINVDCx16_ASAP7_75t_R g2784 ( 
.A(n_1786),
.Y(n_2784)
);

INVx1_ASAP7_75t_L g2785 ( 
.A(n_2141),
.Y(n_2785)
);

CKINVDCx5p33_ASAP7_75t_R g2786 ( 
.A(n_947),
.Y(n_2786)
);

CKINVDCx5p33_ASAP7_75t_R g2787 ( 
.A(n_834),
.Y(n_2787)
);

CKINVDCx5p33_ASAP7_75t_R g2788 ( 
.A(n_340),
.Y(n_2788)
);

INVx1_ASAP7_75t_L g2789 ( 
.A(n_2181),
.Y(n_2789)
);

INVx1_ASAP7_75t_L g2790 ( 
.A(n_1232),
.Y(n_2790)
);

BUFx10_ASAP7_75t_L g2791 ( 
.A(n_84),
.Y(n_2791)
);

CKINVDCx5p33_ASAP7_75t_R g2792 ( 
.A(n_760),
.Y(n_2792)
);

CKINVDCx5p33_ASAP7_75t_R g2793 ( 
.A(n_2036),
.Y(n_2793)
);

BUFx3_ASAP7_75t_L g2794 ( 
.A(n_618),
.Y(n_2794)
);

CKINVDCx5p33_ASAP7_75t_R g2795 ( 
.A(n_1762),
.Y(n_2795)
);

CKINVDCx5p33_ASAP7_75t_R g2796 ( 
.A(n_514),
.Y(n_2796)
);

CKINVDCx5p33_ASAP7_75t_R g2797 ( 
.A(n_500),
.Y(n_2797)
);

CKINVDCx5p33_ASAP7_75t_R g2798 ( 
.A(n_237),
.Y(n_2798)
);

INVx1_ASAP7_75t_L g2799 ( 
.A(n_1538),
.Y(n_2799)
);

CKINVDCx5p33_ASAP7_75t_R g2800 ( 
.A(n_667),
.Y(n_2800)
);

CKINVDCx5p33_ASAP7_75t_R g2801 ( 
.A(n_1497),
.Y(n_2801)
);

CKINVDCx5p33_ASAP7_75t_R g2802 ( 
.A(n_196),
.Y(n_2802)
);

CKINVDCx5p33_ASAP7_75t_R g2803 ( 
.A(n_2209),
.Y(n_2803)
);

BUFx2_ASAP7_75t_L g2804 ( 
.A(n_1322),
.Y(n_2804)
);

CKINVDCx5p33_ASAP7_75t_R g2805 ( 
.A(n_2162),
.Y(n_2805)
);

CKINVDCx5p33_ASAP7_75t_R g2806 ( 
.A(n_308),
.Y(n_2806)
);

CKINVDCx5p33_ASAP7_75t_R g2807 ( 
.A(n_821),
.Y(n_2807)
);

CKINVDCx5p33_ASAP7_75t_R g2808 ( 
.A(n_775),
.Y(n_2808)
);

CKINVDCx5p33_ASAP7_75t_R g2809 ( 
.A(n_115),
.Y(n_2809)
);

CKINVDCx5p33_ASAP7_75t_R g2810 ( 
.A(n_76),
.Y(n_2810)
);

CKINVDCx5p33_ASAP7_75t_R g2811 ( 
.A(n_1096),
.Y(n_2811)
);

CKINVDCx5p33_ASAP7_75t_R g2812 ( 
.A(n_929),
.Y(n_2812)
);

CKINVDCx5p33_ASAP7_75t_R g2813 ( 
.A(n_379),
.Y(n_2813)
);

BUFx6f_ASAP7_75t_L g2814 ( 
.A(n_2075),
.Y(n_2814)
);

INVx1_ASAP7_75t_L g2815 ( 
.A(n_18),
.Y(n_2815)
);

CKINVDCx5p33_ASAP7_75t_R g2816 ( 
.A(n_1195),
.Y(n_2816)
);

INVx1_ASAP7_75t_L g2817 ( 
.A(n_1046),
.Y(n_2817)
);

CKINVDCx5p33_ASAP7_75t_R g2818 ( 
.A(n_117),
.Y(n_2818)
);

INVx1_ASAP7_75t_L g2819 ( 
.A(n_1403),
.Y(n_2819)
);

CKINVDCx16_ASAP7_75t_R g2820 ( 
.A(n_1901),
.Y(n_2820)
);

INVx2_ASAP7_75t_SL g2821 ( 
.A(n_1742),
.Y(n_2821)
);

CKINVDCx5p33_ASAP7_75t_R g2822 ( 
.A(n_1811),
.Y(n_2822)
);

INVx1_ASAP7_75t_L g2823 ( 
.A(n_1448),
.Y(n_2823)
);

INVx1_ASAP7_75t_L g2824 ( 
.A(n_1857),
.Y(n_2824)
);

CKINVDCx5p33_ASAP7_75t_R g2825 ( 
.A(n_851),
.Y(n_2825)
);

INVx1_ASAP7_75t_L g2826 ( 
.A(n_1153),
.Y(n_2826)
);

CKINVDCx5p33_ASAP7_75t_R g2827 ( 
.A(n_2123),
.Y(n_2827)
);

INVx1_ASAP7_75t_L g2828 ( 
.A(n_365),
.Y(n_2828)
);

BUFx3_ASAP7_75t_L g2829 ( 
.A(n_603),
.Y(n_2829)
);

CKINVDCx5p33_ASAP7_75t_R g2830 ( 
.A(n_2228),
.Y(n_2830)
);

CKINVDCx5p33_ASAP7_75t_R g2831 ( 
.A(n_2110),
.Y(n_2831)
);

INVx1_ASAP7_75t_L g2832 ( 
.A(n_293),
.Y(n_2832)
);

CKINVDCx5p33_ASAP7_75t_R g2833 ( 
.A(n_1291),
.Y(n_2833)
);

CKINVDCx5p33_ASAP7_75t_R g2834 ( 
.A(n_2178),
.Y(n_2834)
);

CKINVDCx5p33_ASAP7_75t_R g2835 ( 
.A(n_363),
.Y(n_2835)
);

CKINVDCx5p33_ASAP7_75t_R g2836 ( 
.A(n_1536),
.Y(n_2836)
);

INVx1_ASAP7_75t_SL g2837 ( 
.A(n_977),
.Y(n_2837)
);

CKINVDCx5p33_ASAP7_75t_R g2838 ( 
.A(n_758),
.Y(n_2838)
);

CKINVDCx5p33_ASAP7_75t_R g2839 ( 
.A(n_1560),
.Y(n_2839)
);

INVx2_ASAP7_75t_SL g2840 ( 
.A(n_2098),
.Y(n_2840)
);

INVx1_ASAP7_75t_L g2841 ( 
.A(n_1430),
.Y(n_2841)
);

CKINVDCx20_ASAP7_75t_R g2842 ( 
.A(n_2206),
.Y(n_2842)
);

BUFx2_ASAP7_75t_L g2843 ( 
.A(n_2133),
.Y(n_2843)
);

INVx2_ASAP7_75t_L g2844 ( 
.A(n_216),
.Y(n_2844)
);

CKINVDCx20_ASAP7_75t_R g2845 ( 
.A(n_426),
.Y(n_2845)
);

INVx1_ASAP7_75t_L g2846 ( 
.A(n_1684),
.Y(n_2846)
);

INVx1_ASAP7_75t_L g2847 ( 
.A(n_162),
.Y(n_2847)
);

INVx1_ASAP7_75t_L g2848 ( 
.A(n_679),
.Y(n_2848)
);

INVx1_ASAP7_75t_L g2849 ( 
.A(n_2187),
.Y(n_2849)
);

INVx1_ASAP7_75t_L g2850 ( 
.A(n_499),
.Y(n_2850)
);

INVxp33_ASAP7_75t_R g2851 ( 
.A(n_176),
.Y(n_2851)
);

INVx1_ASAP7_75t_L g2852 ( 
.A(n_761),
.Y(n_2852)
);

CKINVDCx5p33_ASAP7_75t_R g2853 ( 
.A(n_487),
.Y(n_2853)
);

CKINVDCx5p33_ASAP7_75t_R g2854 ( 
.A(n_820),
.Y(n_2854)
);

BUFx10_ASAP7_75t_L g2855 ( 
.A(n_1594),
.Y(n_2855)
);

INVx1_ASAP7_75t_L g2856 ( 
.A(n_296),
.Y(n_2856)
);

CKINVDCx5p33_ASAP7_75t_R g2857 ( 
.A(n_1464),
.Y(n_2857)
);

CKINVDCx5p33_ASAP7_75t_R g2858 ( 
.A(n_660),
.Y(n_2858)
);

CKINVDCx5p33_ASAP7_75t_R g2859 ( 
.A(n_2224),
.Y(n_2859)
);

CKINVDCx5p33_ASAP7_75t_R g2860 ( 
.A(n_1769),
.Y(n_2860)
);

CKINVDCx5p33_ASAP7_75t_R g2861 ( 
.A(n_423),
.Y(n_2861)
);

INVx2_ASAP7_75t_L g2862 ( 
.A(n_2101),
.Y(n_2862)
);

INVx1_ASAP7_75t_L g2863 ( 
.A(n_51),
.Y(n_2863)
);

CKINVDCx5p33_ASAP7_75t_R g2864 ( 
.A(n_2071),
.Y(n_2864)
);

INVx2_ASAP7_75t_SL g2865 ( 
.A(n_556),
.Y(n_2865)
);

CKINVDCx5p33_ASAP7_75t_R g2866 ( 
.A(n_747),
.Y(n_2866)
);

CKINVDCx5p33_ASAP7_75t_R g2867 ( 
.A(n_737),
.Y(n_2867)
);

CKINVDCx5p33_ASAP7_75t_R g2868 ( 
.A(n_1894),
.Y(n_2868)
);

INVx1_ASAP7_75t_L g2869 ( 
.A(n_1848),
.Y(n_2869)
);

INVx1_ASAP7_75t_L g2870 ( 
.A(n_313),
.Y(n_2870)
);

INVx2_ASAP7_75t_L g2871 ( 
.A(n_2117),
.Y(n_2871)
);

CKINVDCx5p33_ASAP7_75t_R g2872 ( 
.A(n_137),
.Y(n_2872)
);

BUFx5_ASAP7_75t_L g2873 ( 
.A(n_2165),
.Y(n_2873)
);

INVx2_ASAP7_75t_L g2874 ( 
.A(n_2201),
.Y(n_2874)
);

INVx1_ASAP7_75t_L g2875 ( 
.A(n_998),
.Y(n_2875)
);

INVx1_ASAP7_75t_L g2876 ( 
.A(n_389),
.Y(n_2876)
);

CKINVDCx5p33_ASAP7_75t_R g2877 ( 
.A(n_815),
.Y(n_2877)
);

CKINVDCx5p33_ASAP7_75t_R g2878 ( 
.A(n_2232),
.Y(n_2878)
);

CKINVDCx6p67_ASAP7_75t_R g2879 ( 
.A(n_1373),
.Y(n_2879)
);

CKINVDCx5p33_ASAP7_75t_R g2880 ( 
.A(n_1786),
.Y(n_2880)
);

CKINVDCx5p33_ASAP7_75t_R g2881 ( 
.A(n_1268),
.Y(n_2881)
);

BUFx2_ASAP7_75t_L g2882 ( 
.A(n_118),
.Y(n_2882)
);

INVx2_ASAP7_75t_SL g2883 ( 
.A(n_98),
.Y(n_2883)
);

INVxp67_ASAP7_75t_L g2884 ( 
.A(n_1357),
.Y(n_2884)
);

INVx1_ASAP7_75t_L g2885 ( 
.A(n_2054),
.Y(n_2885)
);

CKINVDCx5p33_ASAP7_75t_R g2886 ( 
.A(n_1801),
.Y(n_2886)
);

CKINVDCx5p33_ASAP7_75t_R g2887 ( 
.A(n_2195),
.Y(n_2887)
);

INVx1_ASAP7_75t_L g2888 ( 
.A(n_2093),
.Y(n_2888)
);

INVx1_ASAP7_75t_L g2889 ( 
.A(n_1638),
.Y(n_2889)
);

CKINVDCx20_ASAP7_75t_R g2890 ( 
.A(n_1120),
.Y(n_2890)
);

INVx2_ASAP7_75t_SL g2891 ( 
.A(n_145),
.Y(n_2891)
);

INVx1_ASAP7_75t_L g2892 ( 
.A(n_2168),
.Y(n_2892)
);

CKINVDCx5p33_ASAP7_75t_R g2893 ( 
.A(n_627),
.Y(n_2893)
);

CKINVDCx5p33_ASAP7_75t_R g2894 ( 
.A(n_395),
.Y(n_2894)
);

CKINVDCx5p33_ASAP7_75t_R g2895 ( 
.A(n_1279),
.Y(n_2895)
);

BUFx10_ASAP7_75t_L g2896 ( 
.A(n_1276),
.Y(n_2896)
);

CKINVDCx20_ASAP7_75t_R g2897 ( 
.A(n_688),
.Y(n_2897)
);

INVx1_ASAP7_75t_L g2898 ( 
.A(n_885),
.Y(n_2898)
);

INVx1_ASAP7_75t_L g2899 ( 
.A(n_611),
.Y(n_2899)
);

BUFx5_ASAP7_75t_L g2900 ( 
.A(n_1724),
.Y(n_2900)
);

CKINVDCx5p33_ASAP7_75t_R g2901 ( 
.A(n_1617),
.Y(n_2901)
);

INVx2_ASAP7_75t_SL g2902 ( 
.A(n_2087),
.Y(n_2902)
);

CKINVDCx5p33_ASAP7_75t_R g2903 ( 
.A(n_1329),
.Y(n_2903)
);

INVx2_ASAP7_75t_L g2904 ( 
.A(n_2176),
.Y(n_2904)
);

CKINVDCx5p33_ASAP7_75t_R g2905 ( 
.A(n_2134),
.Y(n_2905)
);

CKINVDCx5p33_ASAP7_75t_R g2906 ( 
.A(n_1813),
.Y(n_2906)
);

CKINVDCx5p33_ASAP7_75t_R g2907 ( 
.A(n_18),
.Y(n_2907)
);

CKINVDCx5p33_ASAP7_75t_R g2908 ( 
.A(n_1492),
.Y(n_2908)
);

CKINVDCx5p33_ASAP7_75t_R g2909 ( 
.A(n_986),
.Y(n_2909)
);

CKINVDCx5p33_ASAP7_75t_R g2910 ( 
.A(n_1154),
.Y(n_2910)
);

CKINVDCx5p33_ASAP7_75t_R g2911 ( 
.A(n_822),
.Y(n_2911)
);

CKINVDCx20_ASAP7_75t_R g2912 ( 
.A(n_1176),
.Y(n_2912)
);

INVx1_ASAP7_75t_L g2913 ( 
.A(n_797),
.Y(n_2913)
);

INVx1_ASAP7_75t_L g2914 ( 
.A(n_475),
.Y(n_2914)
);

INVx2_ASAP7_75t_L g2915 ( 
.A(n_1810),
.Y(n_2915)
);

CKINVDCx5p33_ASAP7_75t_R g2916 ( 
.A(n_942),
.Y(n_2916)
);

INVx2_ASAP7_75t_SL g2917 ( 
.A(n_478),
.Y(n_2917)
);

CKINVDCx5p33_ASAP7_75t_R g2918 ( 
.A(n_1136),
.Y(n_2918)
);

INVx1_ASAP7_75t_SL g2919 ( 
.A(n_2023),
.Y(n_2919)
);

INVx1_ASAP7_75t_L g2920 ( 
.A(n_564),
.Y(n_2920)
);

CKINVDCx5p33_ASAP7_75t_R g2921 ( 
.A(n_2216),
.Y(n_2921)
);

INVx1_ASAP7_75t_L g2922 ( 
.A(n_1178),
.Y(n_2922)
);

CKINVDCx5p33_ASAP7_75t_R g2923 ( 
.A(n_1105),
.Y(n_2923)
);

CKINVDCx5p33_ASAP7_75t_R g2924 ( 
.A(n_2227),
.Y(n_2924)
);

CKINVDCx5p33_ASAP7_75t_R g2925 ( 
.A(n_1087),
.Y(n_2925)
);

BUFx6f_ASAP7_75t_L g2926 ( 
.A(n_1583),
.Y(n_2926)
);

INVx1_ASAP7_75t_L g2927 ( 
.A(n_1608),
.Y(n_2927)
);

CKINVDCx5p33_ASAP7_75t_R g2928 ( 
.A(n_1533),
.Y(n_2928)
);

INVx1_ASAP7_75t_SL g2929 ( 
.A(n_2024),
.Y(n_2929)
);

CKINVDCx5p33_ASAP7_75t_R g2930 ( 
.A(n_2177),
.Y(n_2930)
);

CKINVDCx5p33_ASAP7_75t_R g2931 ( 
.A(n_1133),
.Y(n_2931)
);

BUFx10_ASAP7_75t_L g2932 ( 
.A(n_1409),
.Y(n_2932)
);

CKINVDCx5p33_ASAP7_75t_R g2933 ( 
.A(n_2200),
.Y(n_2933)
);

BUFx2_ASAP7_75t_L g2934 ( 
.A(n_514),
.Y(n_2934)
);

INVx1_ASAP7_75t_L g2935 ( 
.A(n_1460),
.Y(n_2935)
);

CKINVDCx5p33_ASAP7_75t_R g2936 ( 
.A(n_1734),
.Y(n_2936)
);

INVx1_ASAP7_75t_L g2937 ( 
.A(n_1550),
.Y(n_2937)
);

CKINVDCx5p33_ASAP7_75t_R g2938 ( 
.A(n_2243),
.Y(n_2938)
);

INVx1_ASAP7_75t_L g2939 ( 
.A(n_803),
.Y(n_2939)
);

CKINVDCx5p33_ASAP7_75t_R g2940 ( 
.A(n_2046),
.Y(n_2940)
);

INVx1_ASAP7_75t_L g2941 ( 
.A(n_295),
.Y(n_2941)
);

CKINVDCx5p33_ASAP7_75t_R g2942 ( 
.A(n_367),
.Y(n_2942)
);

CKINVDCx5p33_ASAP7_75t_R g2943 ( 
.A(n_17),
.Y(n_2943)
);

CKINVDCx5p33_ASAP7_75t_R g2944 ( 
.A(n_554),
.Y(n_2944)
);

CKINVDCx5p33_ASAP7_75t_R g2945 ( 
.A(n_2129),
.Y(n_2945)
);

INVx1_ASAP7_75t_L g2946 ( 
.A(n_1293),
.Y(n_2946)
);

INVx1_ASAP7_75t_L g2947 ( 
.A(n_14),
.Y(n_2947)
);

CKINVDCx5p33_ASAP7_75t_R g2948 ( 
.A(n_1809),
.Y(n_2948)
);

CKINVDCx5p33_ASAP7_75t_R g2949 ( 
.A(n_1105),
.Y(n_2949)
);

INVx2_ASAP7_75t_SL g2950 ( 
.A(n_2203),
.Y(n_2950)
);

CKINVDCx5p33_ASAP7_75t_R g2951 ( 
.A(n_588),
.Y(n_2951)
);

CKINVDCx5p33_ASAP7_75t_R g2952 ( 
.A(n_432),
.Y(n_2952)
);

CKINVDCx5p33_ASAP7_75t_R g2953 ( 
.A(n_878),
.Y(n_2953)
);

CKINVDCx20_ASAP7_75t_R g2954 ( 
.A(n_225),
.Y(n_2954)
);

BUFx3_ASAP7_75t_L g2955 ( 
.A(n_2107),
.Y(n_2955)
);

CKINVDCx5p33_ASAP7_75t_R g2956 ( 
.A(n_1796),
.Y(n_2956)
);

CKINVDCx5p33_ASAP7_75t_R g2957 ( 
.A(n_618),
.Y(n_2957)
);

CKINVDCx5p33_ASAP7_75t_R g2958 ( 
.A(n_1924),
.Y(n_2958)
);

CKINVDCx5p33_ASAP7_75t_R g2959 ( 
.A(n_1904),
.Y(n_2959)
);

INVx1_ASAP7_75t_L g2960 ( 
.A(n_2163),
.Y(n_2960)
);

INVx2_ASAP7_75t_L g2961 ( 
.A(n_931),
.Y(n_2961)
);

INVx1_ASAP7_75t_L g2962 ( 
.A(n_2116),
.Y(n_2962)
);

BUFx10_ASAP7_75t_L g2963 ( 
.A(n_988),
.Y(n_2963)
);

CKINVDCx5p33_ASAP7_75t_R g2964 ( 
.A(n_1802),
.Y(n_2964)
);

CKINVDCx5p33_ASAP7_75t_R g2965 ( 
.A(n_477),
.Y(n_2965)
);

CKINVDCx5p33_ASAP7_75t_R g2966 ( 
.A(n_382),
.Y(n_2966)
);

CKINVDCx5p33_ASAP7_75t_R g2967 ( 
.A(n_1893),
.Y(n_2967)
);

INVx1_ASAP7_75t_L g2968 ( 
.A(n_1107),
.Y(n_2968)
);

CKINVDCx5p33_ASAP7_75t_R g2969 ( 
.A(n_1536),
.Y(n_2969)
);

BUFx5_ASAP7_75t_L g2970 ( 
.A(n_2194),
.Y(n_2970)
);

INVx1_ASAP7_75t_L g2971 ( 
.A(n_2093),
.Y(n_2971)
);

CKINVDCx5p33_ASAP7_75t_R g2972 ( 
.A(n_1371),
.Y(n_2972)
);

CKINVDCx5p33_ASAP7_75t_R g2973 ( 
.A(n_972),
.Y(n_2973)
);

CKINVDCx5p33_ASAP7_75t_R g2974 ( 
.A(n_1559),
.Y(n_2974)
);

BUFx5_ASAP7_75t_L g2975 ( 
.A(n_1638),
.Y(n_2975)
);

CKINVDCx5p33_ASAP7_75t_R g2976 ( 
.A(n_1488),
.Y(n_2976)
);

CKINVDCx5p33_ASAP7_75t_R g2977 ( 
.A(n_2241),
.Y(n_2977)
);

CKINVDCx5p33_ASAP7_75t_R g2978 ( 
.A(n_458),
.Y(n_2978)
);

BUFx3_ASAP7_75t_L g2979 ( 
.A(n_863),
.Y(n_2979)
);

INVx1_ASAP7_75t_L g2980 ( 
.A(n_988),
.Y(n_2980)
);

CKINVDCx5p33_ASAP7_75t_R g2981 ( 
.A(n_2080),
.Y(n_2981)
);

INVx2_ASAP7_75t_L g2982 ( 
.A(n_2091),
.Y(n_2982)
);

INVx1_ASAP7_75t_SL g2983 ( 
.A(n_2208),
.Y(n_2983)
);

CKINVDCx5p33_ASAP7_75t_R g2984 ( 
.A(n_1774),
.Y(n_2984)
);

CKINVDCx20_ASAP7_75t_R g2985 ( 
.A(n_1869),
.Y(n_2985)
);

INVx2_ASAP7_75t_SL g2986 ( 
.A(n_447),
.Y(n_2986)
);

CKINVDCx5p33_ASAP7_75t_R g2987 ( 
.A(n_2092),
.Y(n_2987)
);

BUFx6f_ASAP7_75t_L g2988 ( 
.A(n_988),
.Y(n_2988)
);

INVx1_ASAP7_75t_L g2989 ( 
.A(n_984),
.Y(n_2989)
);

INVx1_ASAP7_75t_L g2990 ( 
.A(n_2227),
.Y(n_2990)
);

CKINVDCx5p33_ASAP7_75t_R g2991 ( 
.A(n_2179),
.Y(n_2991)
);

INVx1_ASAP7_75t_L g2992 ( 
.A(n_903),
.Y(n_2992)
);

CKINVDCx20_ASAP7_75t_R g2993 ( 
.A(n_2019),
.Y(n_2993)
);

CKINVDCx5p33_ASAP7_75t_R g2994 ( 
.A(n_674),
.Y(n_2994)
);

CKINVDCx20_ASAP7_75t_R g2995 ( 
.A(n_2042),
.Y(n_2995)
);

INVx1_ASAP7_75t_L g2996 ( 
.A(n_2080),
.Y(n_2996)
);

INVx1_ASAP7_75t_SL g2997 ( 
.A(n_1084),
.Y(n_2997)
);

CKINVDCx5p33_ASAP7_75t_R g2998 ( 
.A(n_1247),
.Y(n_2998)
);

CKINVDCx5p33_ASAP7_75t_R g2999 ( 
.A(n_0),
.Y(n_2999)
);

BUFx10_ASAP7_75t_L g3000 ( 
.A(n_2114),
.Y(n_3000)
);

INVx2_ASAP7_75t_L g3001 ( 
.A(n_1497),
.Y(n_3001)
);

INVx1_ASAP7_75t_L g3002 ( 
.A(n_1225),
.Y(n_3002)
);

INVx1_ASAP7_75t_L g3003 ( 
.A(n_2124),
.Y(n_3003)
);

CKINVDCx5p33_ASAP7_75t_R g3004 ( 
.A(n_503),
.Y(n_3004)
);

CKINVDCx20_ASAP7_75t_R g3005 ( 
.A(n_707),
.Y(n_3005)
);

INVx1_ASAP7_75t_L g3006 ( 
.A(n_1345),
.Y(n_3006)
);

INVx2_ASAP7_75t_L g3007 ( 
.A(n_1391),
.Y(n_3007)
);

CKINVDCx5p33_ASAP7_75t_R g3008 ( 
.A(n_2230),
.Y(n_3008)
);

BUFx6f_ASAP7_75t_L g3009 ( 
.A(n_591),
.Y(n_3009)
);

INVx1_ASAP7_75t_L g3010 ( 
.A(n_547),
.Y(n_3010)
);

CKINVDCx5p33_ASAP7_75t_R g3011 ( 
.A(n_965),
.Y(n_3011)
);

CKINVDCx5p33_ASAP7_75t_R g3012 ( 
.A(n_1423),
.Y(n_3012)
);

BUFx6f_ASAP7_75t_L g3013 ( 
.A(n_1942),
.Y(n_3013)
);

CKINVDCx5p33_ASAP7_75t_R g3014 ( 
.A(n_952),
.Y(n_3014)
);

CKINVDCx5p33_ASAP7_75t_R g3015 ( 
.A(n_1309),
.Y(n_3015)
);

INVx1_ASAP7_75t_SL g3016 ( 
.A(n_2223),
.Y(n_3016)
);

CKINVDCx5p33_ASAP7_75t_R g3017 ( 
.A(n_1817),
.Y(n_3017)
);

CKINVDCx5p33_ASAP7_75t_R g3018 ( 
.A(n_1632),
.Y(n_3018)
);

CKINVDCx20_ASAP7_75t_R g3019 ( 
.A(n_389),
.Y(n_3019)
);

INVx1_ASAP7_75t_L g3020 ( 
.A(n_1515),
.Y(n_3020)
);

INVx1_ASAP7_75t_L g3021 ( 
.A(n_2078),
.Y(n_3021)
);

CKINVDCx5p33_ASAP7_75t_R g3022 ( 
.A(n_1642),
.Y(n_3022)
);

CKINVDCx5p33_ASAP7_75t_R g3023 ( 
.A(n_2050),
.Y(n_3023)
);

CKINVDCx5p33_ASAP7_75t_R g3024 ( 
.A(n_1435),
.Y(n_3024)
);

INVx1_ASAP7_75t_L g3025 ( 
.A(n_151),
.Y(n_3025)
);

CKINVDCx5p33_ASAP7_75t_R g3026 ( 
.A(n_1177),
.Y(n_3026)
);

CKINVDCx5p33_ASAP7_75t_R g3027 ( 
.A(n_2063),
.Y(n_3027)
);

CKINVDCx5p33_ASAP7_75t_R g3028 ( 
.A(n_326),
.Y(n_3028)
);

CKINVDCx5p33_ASAP7_75t_R g3029 ( 
.A(n_164),
.Y(n_3029)
);

BUFx3_ASAP7_75t_L g3030 ( 
.A(n_2256),
.Y(n_3030)
);

CKINVDCx5p33_ASAP7_75t_R g3031 ( 
.A(n_1835),
.Y(n_3031)
);

CKINVDCx20_ASAP7_75t_R g3032 ( 
.A(n_653),
.Y(n_3032)
);

CKINVDCx5p33_ASAP7_75t_R g3033 ( 
.A(n_625),
.Y(n_3033)
);

CKINVDCx5p33_ASAP7_75t_R g3034 ( 
.A(n_1075),
.Y(n_3034)
);

INVx1_ASAP7_75t_L g3035 ( 
.A(n_1163),
.Y(n_3035)
);

CKINVDCx5p33_ASAP7_75t_R g3036 ( 
.A(n_70),
.Y(n_3036)
);

CKINVDCx5p33_ASAP7_75t_R g3037 ( 
.A(n_1327),
.Y(n_3037)
);

INVx1_ASAP7_75t_L g3038 ( 
.A(n_1248),
.Y(n_3038)
);

INVx1_ASAP7_75t_L g3039 ( 
.A(n_1774),
.Y(n_3039)
);

CKINVDCx20_ASAP7_75t_R g3040 ( 
.A(n_1489),
.Y(n_3040)
);

CKINVDCx5p33_ASAP7_75t_R g3041 ( 
.A(n_2237),
.Y(n_3041)
);

INVx1_ASAP7_75t_L g3042 ( 
.A(n_1045),
.Y(n_3042)
);

BUFx2_ASAP7_75t_L g3043 ( 
.A(n_653),
.Y(n_3043)
);

CKINVDCx5p33_ASAP7_75t_R g3044 ( 
.A(n_1581),
.Y(n_3044)
);

INVx1_ASAP7_75t_L g3045 ( 
.A(n_1411),
.Y(n_3045)
);

CKINVDCx5p33_ASAP7_75t_R g3046 ( 
.A(n_2259),
.Y(n_3046)
);

INVx1_ASAP7_75t_L g3047 ( 
.A(n_2018),
.Y(n_3047)
);

INVx1_ASAP7_75t_L g3048 ( 
.A(n_2037),
.Y(n_3048)
);

CKINVDCx5p33_ASAP7_75t_R g3049 ( 
.A(n_1733),
.Y(n_3049)
);

INVx1_ASAP7_75t_SL g3050 ( 
.A(n_2261),
.Y(n_3050)
);

INVx1_ASAP7_75t_L g3051 ( 
.A(n_924),
.Y(n_3051)
);

INVx1_ASAP7_75t_L g3052 ( 
.A(n_2079),
.Y(n_3052)
);

CKINVDCx20_ASAP7_75t_R g3053 ( 
.A(n_140),
.Y(n_3053)
);

CKINVDCx5p33_ASAP7_75t_R g3054 ( 
.A(n_2177),
.Y(n_3054)
);

CKINVDCx5p33_ASAP7_75t_R g3055 ( 
.A(n_1013),
.Y(n_3055)
);

CKINVDCx5p33_ASAP7_75t_R g3056 ( 
.A(n_2041),
.Y(n_3056)
);

INVx1_ASAP7_75t_L g3057 ( 
.A(n_546),
.Y(n_3057)
);

CKINVDCx5p33_ASAP7_75t_R g3058 ( 
.A(n_1751),
.Y(n_3058)
);

INVx1_ASAP7_75t_L g3059 ( 
.A(n_2153),
.Y(n_3059)
);

CKINVDCx5p33_ASAP7_75t_R g3060 ( 
.A(n_83),
.Y(n_3060)
);

CKINVDCx5p33_ASAP7_75t_R g3061 ( 
.A(n_1512),
.Y(n_3061)
);

CKINVDCx5p33_ASAP7_75t_R g3062 ( 
.A(n_2035),
.Y(n_3062)
);

BUFx3_ASAP7_75t_L g3063 ( 
.A(n_1367),
.Y(n_3063)
);

INVx1_ASAP7_75t_L g3064 ( 
.A(n_2070),
.Y(n_3064)
);

CKINVDCx5p33_ASAP7_75t_R g3065 ( 
.A(n_97),
.Y(n_3065)
);

INVx1_ASAP7_75t_L g3066 ( 
.A(n_1278),
.Y(n_3066)
);

BUFx10_ASAP7_75t_L g3067 ( 
.A(n_2218),
.Y(n_3067)
);

CKINVDCx20_ASAP7_75t_R g3068 ( 
.A(n_1670),
.Y(n_3068)
);

INVx1_ASAP7_75t_L g3069 ( 
.A(n_809),
.Y(n_3069)
);

CKINVDCx5p33_ASAP7_75t_R g3070 ( 
.A(n_2048),
.Y(n_3070)
);

INVx1_ASAP7_75t_L g3071 ( 
.A(n_2156),
.Y(n_3071)
);

BUFx10_ASAP7_75t_L g3072 ( 
.A(n_1879),
.Y(n_3072)
);

INVx2_ASAP7_75t_L g3073 ( 
.A(n_1773),
.Y(n_3073)
);

CKINVDCx5p33_ASAP7_75t_R g3074 ( 
.A(n_340),
.Y(n_3074)
);

CKINVDCx20_ASAP7_75t_R g3075 ( 
.A(n_1091),
.Y(n_3075)
);

CKINVDCx5p33_ASAP7_75t_R g3076 ( 
.A(n_2236),
.Y(n_3076)
);

CKINVDCx5p33_ASAP7_75t_R g3077 ( 
.A(n_1154),
.Y(n_3077)
);

CKINVDCx5p33_ASAP7_75t_R g3078 ( 
.A(n_1112),
.Y(n_3078)
);

BUFx3_ASAP7_75t_L g3079 ( 
.A(n_1363),
.Y(n_3079)
);

INVx1_ASAP7_75t_L g3080 ( 
.A(n_2229),
.Y(n_3080)
);

CKINVDCx16_ASAP7_75t_R g3081 ( 
.A(n_1847),
.Y(n_3081)
);

BUFx6f_ASAP7_75t_L g3082 ( 
.A(n_2151),
.Y(n_3082)
);

CKINVDCx5p33_ASAP7_75t_R g3083 ( 
.A(n_1758),
.Y(n_3083)
);

CKINVDCx20_ASAP7_75t_R g3084 ( 
.A(n_608),
.Y(n_3084)
);

INVx1_ASAP7_75t_L g3085 ( 
.A(n_1204),
.Y(n_3085)
);

CKINVDCx5p33_ASAP7_75t_R g3086 ( 
.A(n_418),
.Y(n_3086)
);

INVx1_ASAP7_75t_L g3087 ( 
.A(n_2221),
.Y(n_3087)
);

CKINVDCx5p33_ASAP7_75t_R g3088 ( 
.A(n_1528),
.Y(n_3088)
);

CKINVDCx5p33_ASAP7_75t_R g3089 ( 
.A(n_622),
.Y(n_3089)
);

CKINVDCx5p33_ASAP7_75t_R g3090 ( 
.A(n_387),
.Y(n_3090)
);

CKINVDCx5p33_ASAP7_75t_R g3091 ( 
.A(n_1899),
.Y(n_3091)
);

INVx1_ASAP7_75t_L g3092 ( 
.A(n_2017),
.Y(n_3092)
);

BUFx5_ASAP7_75t_L g3093 ( 
.A(n_1534),
.Y(n_3093)
);

CKINVDCx5p33_ASAP7_75t_R g3094 ( 
.A(n_2139),
.Y(n_3094)
);

CKINVDCx16_ASAP7_75t_R g3095 ( 
.A(n_1966),
.Y(n_3095)
);

INVx1_ASAP7_75t_SL g3096 ( 
.A(n_1743),
.Y(n_3096)
);

CKINVDCx5p33_ASAP7_75t_R g3097 ( 
.A(n_257),
.Y(n_3097)
);

INVx2_ASAP7_75t_L g3098 ( 
.A(n_842),
.Y(n_3098)
);

CKINVDCx20_ASAP7_75t_R g3099 ( 
.A(n_2135),
.Y(n_3099)
);

CKINVDCx5p33_ASAP7_75t_R g3100 ( 
.A(n_2167),
.Y(n_3100)
);

INVx1_ASAP7_75t_L g3101 ( 
.A(n_1986),
.Y(n_3101)
);

CKINVDCx5p33_ASAP7_75t_R g3102 ( 
.A(n_874),
.Y(n_3102)
);

CKINVDCx5p33_ASAP7_75t_R g3103 ( 
.A(n_1975),
.Y(n_3103)
);

INVx1_ASAP7_75t_L g3104 ( 
.A(n_330),
.Y(n_3104)
);

CKINVDCx5p33_ASAP7_75t_R g3105 ( 
.A(n_837),
.Y(n_3105)
);

CKINVDCx20_ASAP7_75t_R g3106 ( 
.A(n_786),
.Y(n_3106)
);

CKINVDCx5p33_ASAP7_75t_R g3107 ( 
.A(n_1651),
.Y(n_3107)
);

BUFx10_ASAP7_75t_L g3108 ( 
.A(n_2203),
.Y(n_3108)
);

BUFx6f_ASAP7_75t_L g3109 ( 
.A(n_38),
.Y(n_3109)
);

INVx1_ASAP7_75t_L g3110 ( 
.A(n_1816),
.Y(n_3110)
);

CKINVDCx5p33_ASAP7_75t_R g3111 ( 
.A(n_198),
.Y(n_3111)
);

BUFx5_ASAP7_75t_L g3112 ( 
.A(n_800),
.Y(n_3112)
);

BUFx10_ASAP7_75t_L g3113 ( 
.A(n_2146),
.Y(n_3113)
);

INVx1_ASAP7_75t_SL g3114 ( 
.A(n_2052),
.Y(n_3114)
);

CKINVDCx5p33_ASAP7_75t_R g3115 ( 
.A(n_1608),
.Y(n_3115)
);

CKINVDCx5p33_ASAP7_75t_R g3116 ( 
.A(n_2021),
.Y(n_3116)
);

INVx1_ASAP7_75t_L g3117 ( 
.A(n_35),
.Y(n_3117)
);

CKINVDCx5p33_ASAP7_75t_R g3118 ( 
.A(n_1821),
.Y(n_3118)
);

CKINVDCx5p33_ASAP7_75t_R g3119 ( 
.A(n_605),
.Y(n_3119)
);

CKINVDCx20_ASAP7_75t_R g3120 ( 
.A(n_700),
.Y(n_3120)
);

CKINVDCx5p33_ASAP7_75t_R g3121 ( 
.A(n_2207),
.Y(n_3121)
);

INVx2_ASAP7_75t_L g3122 ( 
.A(n_1419),
.Y(n_3122)
);

CKINVDCx5p33_ASAP7_75t_R g3123 ( 
.A(n_803),
.Y(n_3123)
);

INVx1_ASAP7_75t_L g3124 ( 
.A(n_1729),
.Y(n_3124)
);

CKINVDCx5p33_ASAP7_75t_R g3125 ( 
.A(n_2113),
.Y(n_3125)
);

INVx1_ASAP7_75t_SL g3126 ( 
.A(n_1659),
.Y(n_3126)
);

INVx1_ASAP7_75t_L g3127 ( 
.A(n_461),
.Y(n_3127)
);

CKINVDCx5p33_ASAP7_75t_R g3128 ( 
.A(n_726),
.Y(n_3128)
);

CKINVDCx5p33_ASAP7_75t_R g3129 ( 
.A(n_414),
.Y(n_3129)
);

INVx1_ASAP7_75t_L g3130 ( 
.A(n_1152),
.Y(n_3130)
);

CKINVDCx5p33_ASAP7_75t_R g3131 ( 
.A(n_2144),
.Y(n_3131)
);

CKINVDCx14_ASAP7_75t_R g3132 ( 
.A(n_2183),
.Y(n_3132)
);

INVx1_ASAP7_75t_L g3133 ( 
.A(n_2060),
.Y(n_3133)
);

CKINVDCx5p33_ASAP7_75t_R g3134 ( 
.A(n_1331),
.Y(n_3134)
);

CKINVDCx20_ASAP7_75t_R g3135 ( 
.A(n_1504),
.Y(n_3135)
);

CKINVDCx5p33_ASAP7_75t_R g3136 ( 
.A(n_1948),
.Y(n_3136)
);

INVx1_ASAP7_75t_L g3137 ( 
.A(n_503),
.Y(n_3137)
);

CKINVDCx5p33_ASAP7_75t_R g3138 ( 
.A(n_966),
.Y(n_3138)
);

CKINVDCx5p33_ASAP7_75t_R g3139 ( 
.A(n_1936),
.Y(n_3139)
);

CKINVDCx5p33_ASAP7_75t_R g3140 ( 
.A(n_1260),
.Y(n_3140)
);

INVx1_ASAP7_75t_L g3141 ( 
.A(n_1592),
.Y(n_3141)
);

INVx1_ASAP7_75t_L g3142 ( 
.A(n_1304),
.Y(n_3142)
);

INVx1_ASAP7_75t_SL g3143 ( 
.A(n_1259),
.Y(n_3143)
);

CKINVDCx5p33_ASAP7_75t_R g3144 ( 
.A(n_591),
.Y(n_3144)
);

INVx1_ASAP7_75t_L g3145 ( 
.A(n_2176),
.Y(n_3145)
);

INVx2_ASAP7_75t_L g3146 ( 
.A(n_1382),
.Y(n_3146)
);

BUFx2_ASAP7_75t_L g3147 ( 
.A(n_165),
.Y(n_3147)
);

CKINVDCx5p33_ASAP7_75t_R g3148 ( 
.A(n_2217),
.Y(n_3148)
);

CKINVDCx5p33_ASAP7_75t_R g3149 ( 
.A(n_578),
.Y(n_3149)
);

INVx1_ASAP7_75t_L g3150 ( 
.A(n_370),
.Y(n_3150)
);

CKINVDCx16_ASAP7_75t_R g3151 ( 
.A(n_2154),
.Y(n_3151)
);

BUFx10_ASAP7_75t_L g3152 ( 
.A(n_379),
.Y(n_3152)
);

CKINVDCx5p33_ASAP7_75t_R g3153 ( 
.A(n_1357),
.Y(n_3153)
);

CKINVDCx5p33_ASAP7_75t_R g3154 ( 
.A(n_2088),
.Y(n_3154)
);

CKINVDCx20_ASAP7_75t_R g3155 ( 
.A(n_246),
.Y(n_3155)
);

BUFx3_ASAP7_75t_L g3156 ( 
.A(n_1213),
.Y(n_3156)
);

CKINVDCx5p33_ASAP7_75t_R g3157 ( 
.A(n_754),
.Y(n_3157)
);

CKINVDCx5p33_ASAP7_75t_R g3158 ( 
.A(n_906),
.Y(n_3158)
);

CKINVDCx5p33_ASAP7_75t_R g3159 ( 
.A(n_983),
.Y(n_3159)
);

CKINVDCx5p33_ASAP7_75t_R g3160 ( 
.A(n_363),
.Y(n_3160)
);

INVx1_ASAP7_75t_SL g3161 ( 
.A(n_2202),
.Y(n_3161)
);

CKINVDCx5p33_ASAP7_75t_R g3162 ( 
.A(n_1115),
.Y(n_3162)
);

CKINVDCx5p33_ASAP7_75t_R g3163 ( 
.A(n_330),
.Y(n_3163)
);

INVx1_ASAP7_75t_L g3164 ( 
.A(n_275),
.Y(n_3164)
);

CKINVDCx20_ASAP7_75t_R g3165 ( 
.A(n_1308),
.Y(n_3165)
);

CKINVDCx20_ASAP7_75t_R g3166 ( 
.A(n_1894),
.Y(n_3166)
);

INVx2_ASAP7_75t_L g3167 ( 
.A(n_2120),
.Y(n_3167)
);

INVx1_ASAP7_75t_L g3168 ( 
.A(n_573),
.Y(n_3168)
);

CKINVDCx5p33_ASAP7_75t_R g3169 ( 
.A(n_1779),
.Y(n_3169)
);

BUFx2_ASAP7_75t_L g3170 ( 
.A(n_121),
.Y(n_3170)
);

INVx2_ASAP7_75t_L g3171 ( 
.A(n_550),
.Y(n_3171)
);

INVx2_ASAP7_75t_L g3172 ( 
.A(n_1024),
.Y(n_3172)
);

CKINVDCx5p33_ASAP7_75t_R g3173 ( 
.A(n_815),
.Y(n_3173)
);

CKINVDCx5p33_ASAP7_75t_R g3174 ( 
.A(n_1833),
.Y(n_3174)
);

BUFx3_ASAP7_75t_L g3175 ( 
.A(n_652),
.Y(n_3175)
);

CKINVDCx5p33_ASAP7_75t_R g3176 ( 
.A(n_1269),
.Y(n_3176)
);

CKINVDCx5p33_ASAP7_75t_R g3177 ( 
.A(n_1962),
.Y(n_3177)
);

CKINVDCx5p33_ASAP7_75t_R g3178 ( 
.A(n_1378),
.Y(n_3178)
);

BUFx3_ASAP7_75t_L g3179 ( 
.A(n_1832),
.Y(n_3179)
);

CKINVDCx5p33_ASAP7_75t_R g3180 ( 
.A(n_1670),
.Y(n_3180)
);

CKINVDCx5p33_ASAP7_75t_R g3181 ( 
.A(n_117),
.Y(n_3181)
);

CKINVDCx5p33_ASAP7_75t_R g3182 ( 
.A(n_1954),
.Y(n_3182)
);

CKINVDCx5p33_ASAP7_75t_R g3183 ( 
.A(n_2115),
.Y(n_3183)
);

INVx1_ASAP7_75t_L g3184 ( 
.A(n_586),
.Y(n_3184)
);

CKINVDCx20_ASAP7_75t_R g3185 ( 
.A(n_594),
.Y(n_3185)
);

CKINVDCx5p33_ASAP7_75t_R g3186 ( 
.A(n_2029),
.Y(n_3186)
);

INVx1_ASAP7_75t_L g3187 ( 
.A(n_205),
.Y(n_3187)
);

CKINVDCx5p33_ASAP7_75t_R g3188 ( 
.A(n_211),
.Y(n_3188)
);

CKINVDCx5p33_ASAP7_75t_R g3189 ( 
.A(n_1875),
.Y(n_3189)
);

CKINVDCx5p33_ASAP7_75t_R g3190 ( 
.A(n_1649),
.Y(n_3190)
);

INVx2_ASAP7_75t_L g3191 ( 
.A(n_2118),
.Y(n_3191)
);

CKINVDCx5p33_ASAP7_75t_R g3192 ( 
.A(n_922),
.Y(n_3192)
);

HB1xp67_ASAP7_75t_L g3193 ( 
.A(n_58),
.Y(n_3193)
);

INVx1_ASAP7_75t_L g3194 ( 
.A(n_329),
.Y(n_3194)
);

CKINVDCx5p33_ASAP7_75t_R g3195 ( 
.A(n_732),
.Y(n_3195)
);

INVx4_ASAP7_75t_R g3196 ( 
.A(n_1447),
.Y(n_3196)
);

INVx1_ASAP7_75t_L g3197 ( 
.A(n_261),
.Y(n_3197)
);

INVx1_ASAP7_75t_L g3198 ( 
.A(n_1304),
.Y(n_3198)
);

BUFx10_ASAP7_75t_L g3199 ( 
.A(n_1492),
.Y(n_3199)
);

CKINVDCx5p33_ASAP7_75t_R g3200 ( 
.A(n_1092),
.Y(n_3200)
);

INVx1_ASAP7_75t_L g3201 ( 
.A(n_2062),
.Y(n_3201)
);

INVx2_ASAP7_75t_L g3202 ( 
.A(n_1937),
.Y(n_3202)
);

CKINVDCx5p33_ASAP7_75t_R g3203 ( 
.A(n_1107),
.Y(n_3203)
);

CKINVDCx5p33_ASAP7_75t_R g3204 ( 
.A(n_427),
.Y(n_3204)
);

BUFx10_ASAP7_75t_L g3205 ( 
.A(n_508),
.Y(n_3205)
);

CKINVDCx5p33_ASAP7_75t_R g3206 ( 
.A(n_585),
.Y(n_3206)
);

CKINVDCx5p33_ASAP7_75t_R g3207 ( 
.A(n_2025),
.Y(n_3207)
);

CKINVDCx5p33_ASAP7_75t_R g3208 ( 
.A(n_144),
.Y(n_3208)
);

BUFx3_ASAP7_75t_L g3209 ( 
.A(n_1203),
.Y(n_3209)
);

CKINVDCx5p33_ASAP7_75t_R g3210 ( 
.A(n_927),
.Y(n_3210)
);

CKINVDCx5p33_ASAP7_75t_R g3211 ( 
.A(n_1973),
.Y(n_3211)
);

CKINVDCx5p33_ASAP7_75t_R g3212 ( 
.A(n_1167),
.Y(n_3212)
);

CKINVDCx5p33_ASAP7_75t_R g3213 ( 
.A(n_1845),
.Y(n_3213)
);

CKINVDCx5p33_ASAP7_75t_R g3214 ( 
.A(n_1473),
.Y(n_3214)
);

INVx1_ASAP7_75t_L g3215 ( 
.A(n_490),
.Y(n_3215)
);

CKINVDCx5p33_ASAP7_75t_R g3216 ( 
.A(n_1750),
.Y(n_3216)
);

INVx1_ASAP7_75t_SL g3217 ( 
.A(n_2043),
.Y(n_3217)
);

CKINVDCx5p33_ASAP7_75t_R g3218 ( 
.A(n_1484),
.Y(n_3218)
);

CKINVDCx5p33_ASAP7_75t_R g3219 ( 
.A(n_1450),
.Y(n_3219)
);

CKINVDCx20_ASAP7_75t_R g3220 ( 
.A(n_1495),
.Y(n_3220)
);

CKINVDCx5p33_ASAP7_75t_R g3221 ( 
.A(n_1963),
.Y(n_3221)
);

INVx1_ASAP7_75t_L g3222 ( 
.A(n_1036),
.Y(n_3222)
);

CKINVDCx20_ASAP7_75t_R g3223 ( 
.A(n_1222),
.Y(n_3223)
);

CKINVDCx5p33_ASAP7_75t_R g3224 ( 
.A(n_1771),
.Y(n_3224)
);

CKINVDCx5p33_ASAP7_75t_R g3225 ( 
.A(n_754),
.Y(n_3225)
);

CKINVDCx5p33_ASAP7_75t_R g3226 ( 
.A(n_1666),
.Y(n_3226)
);

INVx1_ASAP7_75t_L g3227 ( 
.A(n_1604),
.Y(n_3227)
);

INVx1_ASAP7_75t_L g3228 ( 
.A(n_4),
.Y(n_3228)
);

INVx1_ASAP7_75t_L g3229 ( 
.A(n_984),
.Y(n_3229)
);

CKINVDCx5p33_ASAP7_75t_R g3230 ( 
.A(n_2016),
.Y(n_3230)
);

CKINVDCx5p33_ASAP7_75t_R g3231 ( 
.A(n_2252),
.Y(n_3231)
);

INVx1_ASAP7_75t_L g3232 ( 
.A(n_1282),
.Y(n_3232)
);

INVx2_ASAP7_75t_L g3233 ( 
.A(n_789),
.Y(n_3233)
);

BUFx3_ASAP7_75t_L g3234 ( 
.A(n_1797),
.Y(n_3234)
);

CKINVDCx20_ASAP7_75t_R g3235 ( 
.A(n_861),
.Y(n_3235)
);

CKINVDCx5p33_ASAP7_75t_R g3236 ( 
.A(n_1507),
.Y(n_3236)
);

CKINVDCx5p33_ASAP7_75t_R g3237 ( 
.A(n_321),
.Y(n_3237)
);

CKINVDCx5p33_ASAP7_75t_R g3238 ( 
.A(n_968),
.Y(n_3238)
);

INVx2_ASAP7_75t_L g3239 ( 
.A(n_2143),
.Y(n_3239)
);

CKINVDCx5p33_ASAP7_75t_R g3240 ( 
.A(n_2173),
.Y(n_3240)
);

INVx1_ASAP7_75t_L g3241 ( 
.A(n_1728),
.Y(n_3241)
);

CKINVDCx5p33_ASAP7_75t_R g3242 ( 
.A(n_2047),
.Y(n_3242)
);

CKINVDCx5p33_ASAP7_75t_R g3243 ( 
.A(n_2209),
.Y(n_3243)
);

BUFx3_ASAP7_75t_L g3244 ( 
.A(n_1998),
.Y(n_3244)
);

CKINVDCx5p33_ASAP7_75t_R g3245 ( 
.A(n_396),
.Y(n_3245)
);

CKINVDCx5p33_ASAP7_75t_R g3246 ( 
.A(n_2125),
.Y(n_3246)
);

INVx1_ASAP7_75t_L g3247 ( 
.A(n_1383),
.Y(n_3247)
);

CKINVDCx5p33_ASAP7_75t_R g3248 ( 
.A(n_1639),
.Y(n_3248)
);

CKINVDCx5p33_ASAP7_75t_R g3249 ( 
.A(n_2160),
.Y(n_3249)
);

CKINVDCx5p33_ASAP7_75t_R g3250 ( 
.A(n_2104),
.Y(n_3250)
);

CKINVDCx5p33_ASAP7_75t_R g3251 ( 
.A(n_1004),
.Y(n_3251)
);

CKINVDCx20_ASAP7_75t_R g3252 ( 
.A(n_1210),
.Y(n_3252)
);

CKINVDCx20_ASAP7_75t_R g3253 ( 
.A(n_2020),
.Y(n_3253)
);

BUFx3_ASAP7_75t_L g3254 ( 
.A(n_1552),
.Y(n_3254)
);

CKINVDCx5p33_ASAP7_75t_R g3255 ( 
.A(n_397),
.Y(n_3255)
);

CKINVDCx5p33_ASAP7_75t_R g3256 ( 
.A(n_138),
.Y(n_3256)
);

INVx1_ASAP7_75t_L g3257 ( 
.A(n_354),
.Y(n_3257)
);

INVx1_ASAP7_75t_SL g3258 ( 
.A(n_410),
.Y(n_3258)
);

CKINVDCx5p33_ASAP7_75t_R g3259 ( 
.A(n_1174),
.Y(n_3259)
);

INVx1_ASAP7_75t_L g3260 ( 
.A(n_1080),
.Y(n_3260)
);

CKINVDCx5p33_ASAP7_75t_R g3261 ( 
.A(n_679),
.Y(n_3261)
);

CKINVDCx5p33_ASAP7_75t_R g3262 ( 
.A(n_1908),
.Y(n_3262)
);

CKINVDCx20_ASAP7_75t_R g3263 ( 
.A(n_2247),
.Y(n_3263)
);

BUFx6f_ASAP7_75t_L g3264 ( 
.A(n_2006),
.Y(n_3264)
);

CKINVDCx5p33_ASAP7_75t_R g3265 ( 
.A(n_307),
.Y(n_3265)
);

CKINVDCx5p33_ASAP7_75t_R g3266 ( 
.A(n_1425),
.Y(n_3266)
);

BUFx5_ASAP7_75t_L g3267 ( 
.A(n_514),
.Y(n_3267)
);

CKINVDCx5p33_ASAP7_75t_R g3268 ( 
.A(n_2095),
.Y(n_3268)
);

CKINVDCx5p33_ASAP7_75t_R g3269 ( 
.A(n_1573),
.Y(n_3269)
);

INVx1_ASAP7_75t_SL g3270 ( 
.A(n_1647),
.Y(n_3270)
);

CKINVDCx16_ASAP7_75t_R g3271 ( 
.A(n_115),
.Y(n_3271)
);

CKINVDCx20_ASAP7_75t_R g3272 ( 
.A(n_1505),
.Y(n_3272)
);

CKINVDCx5p33_ASAP7_75t_R g3273 ( 
.A(n_2132),
.Y(n_3273)
);

CKINVDCx5p33_ASAP7_75t_R g3274 ( 
.A(n_730),
.Y(n_3274)
);

CKINVDCx5p33_ASAP7_75t_R g3275 ( 
.A(n_743),
.Y(n_3275)
);

CKINVDCx5p33_ASAP7_75t_R g3276 ( 
.A(n_787),
.Y(n_3276)
);

INVx1_ASAP7_75t_L g3277 ( 
.A(n_1725),
.Y(n_3277)
);

CKINVDCx5p33_ASAP7_75t_R g3278 ( 
.A(n_1354),
.Y(n_3278)
);

CKINVDCx5p33_ASAP7_75t_R g3279 ( 
.A(n_640),
.Y(n_3279)
);

CKINVDCx5p33_ASAP7_75t_R g3280 ( 
.A(n_43),
.Y(n_3280)
);

CKINVDCx5p33_ASAP7_75t_R g3281 ( 
.A(n_1327),
.Y(n_3281)
);

CKINVDCx5p33_ASAP7_75t_R g3282 ( 
.A(n_1468),
.Y(n_3282)
);

CKINVDCx5p33_ASAP7_75t_R g3283 ( 
.A(n_188),
.Y(n_3283)
);

CKINVDCx5p33_ASAP7_75t_R g3284 ( 
.A(n_111),
.Y(n_3284)
);

CKINVDCx5p33_ASAP7_75t_R g3285 ( 
.A(n_1284),
.Y(n_3285)
);

INVx1_ASAP7_75t_L g3286 ( 
.A(n_431),
.Y(n_3286)
);

CKINVDCx5p33_ASAP7_75t_R g3287 ( 
.A(n_1890),
.Y(n_3287)
);

BUFx2_ASAP7_75t_L g3288 ( 
.A(n_1247),
.Y(n_3288)
);

INVx1_ASAP7_75t_L g3289 ( 
.A(n_1977),
.Y(n_3289)
);

CKINVDCx5p33_ASAP7_75t_R g3290 ( 
.A(n_112),
.Y(n_3290)
);

CKINVDCx5p33_ASAP7_75t_R g3291 ( 
.A(n_290),
.Y(n_3291)
);

INVx2_ASAP7_75t_L g3292 ( 
.A(n_1809),
.Y(n_3292)
);

CKINVDCx20_ASAP7_75t_R g3293 ( 
.A(n_1295),
.Y(n_3293)
);

BUFx5_ASAP7_75t_L g3294 ( 
.A(n_2219),
.Y(n_3294)
);

CKINVDCx5p33_ASAP7_75t_R g3295 ( 
.A(n_1475),
.Y(n_3295)
);

CKINVDCx5p33_ASAP7_75t_R g3296 ( 
.A(n_1537),
.Y(n_3296)
);

BUFx10_ASAP7_75t_L g3297 ( 
.A(n_404),
.Y(n_3297)
);

CKINVDCx5p33_ASAP7_75t_R g3298 ( 
.A(n_597),
.Y(n_3298)
);

BUFx8_ASAP7_75t_SL g3299 ( 
.A(n_291),
.Y(n_3299)
);

CKINVDCx5p33_ASAP7_75t_R g3300 ( 
.A(n_1367),
.Y(n_3300)
);

BUFx6f_ASAP7_75t_L g3301 ( 
.A(n_1160),
.Y(n_3301)
);

INVx1_ASAP7_75t_L g3302 ( 
.A(n_1869),
.Y(n_3302)
);

CKINVDCx5p33_ASAP7_75t_R g3303 ( 
.A(n_2155),
.Y(n_3303)
);

CKINVDCx20_ASAP7_75t_R g3304 ( 
.A(n_982),
.Y(n_3304)
);

INVx1_ASAP7_75t_L g3305 ( 
.A(n_450),
.Y(n_3305)
);

CKINVDCx5p33_ASAP7_75t_R g3306 ( 
.A(n_238),
.Y(n_3306)
);

INVx1_ASAP7_75t_L g3307 ( 
.A(n_873),
.Y(n_3307)
);

CKINVDCx5p33_ASAP7_75t_R g3308 ( 
.A(n_2214),
.Y(n_3308)
);

CKINVDCx16_ASAP7_75t_R g3309 ( 
.A(n_763),
.Y(n_3309)
);

CKINVDCx5p33_ASAP7_75t_R g3310 ( 
.A(n_1098),
.Y(n_3310)
);

BUFx5_ASAP7_75t_L g3311 ( 
.A(n_1051),
.Y(n_3311)
);

CKINVDCx5p33_ASAP7_75t_R g3312 ( 
.A(n_899),
.Y(n_3312)
);

CKINVDCx5p33_ASAP7_75t_R g3313 ( 
.A(n_1033),
.Y(n_3313)
);

CKINVDCx5p33_ASAP7_75t_R g3314 ( 
.A(n_2102),
.Y(n_3314)
);

CKINVDCx5p33_ASAP7_75t_R g3315 ( 
.A(n_2012),
.Y(n_3315)
);

CKINVDCx5p33_ASAP7_75t_R g3316 ( 
.A(n_1576),
.Y(n_3316)
);

CKINVDCx5p33_ASAP7_75t_R g3317 ( 
.A(n_1910),
.Y(n_3317)
);

INVx1_ASAP7_75t_L g3318 ( 
.A(n_2210),
.Y(n_3318)
);

CKINVDCx5p33_ASAP7_75t_R g3319 ( 
.A(n_1029),
.Y(n_3319)
);

CKINVDCx5p33_ASAP7_75t_R g3320 ( 
.A(n_1392),
.Y(n_3320)
);

CKINVDCx20_ASAP7_75t_R g3321 ( 
.A(n_1816),
.Y(n_3321)
);

CKINVDCx5p33_ASAP7_75t_R g3322 ( 
.A(n_1324),
.Y(n_3322)
);

INVx1_ASAP7_75t_L g3323 ( 
.A(n_2059),
.Y(n_3323)
);

INVx1_ASAP7_75t_L g3324 ( 
.A(n_1897),
.Y(n_3324)
);

INVx2_ASAP7_75t_L g3325 ( 
.A(n_874),
.Y(n_3325)
);

CKINVDCx5p33_ASAP7_75t_R g3326 ( 
.A(n_2242),
.Y(n_3326)
);

INVx1_ASAP7_75t_L g3327 ( 
.A(n_13),
.Y(n_3327)
);

CKINVDCx5p33_ASAP7_75t_R g3328 ( 
.A(n_641),
.Y(n_3328)
);

CKINVDCx5p33_ASAP7_75t_R g3329 ( 
.A(n_2089),
.Y(n_3329)
);

INVx1_ASAP7_75t_L g3330 ( 
.A(n_599),
.Y(n_3330)
);

CKINVDCx5p33_ASAP7_75t_R g3331 ( 
.A(n_1426),
.Y(n_3331)
);

CKINVDCx5p33_ASAP7_75t_R g3332 ( 
.A(n_1953),
.Y(n_3332)
);

CKINVDCx5p33_ASAP7_75t_R g3333 ( 
.A(n_1302),
.Y(n_3333)
);

INVx1_ASAP7_75t_L g3334 ( 
.A(n_803),
.Y(n_3334)
);

CKINVDCx5p33_ASAP7_75t_R g3335 ( 
.A(n_1185),
.Y(n_3335)
);

CKINVDCx5p33_ASAP7_75t_R g3336 ( 
.A(n_1489),
.Y(n_3336)
);

CKINVDCx5p33_ASAP7_75t_R g3337 ( 
.A(n_1340),
.Y(n_3337)
);

CKINVDCx5p33_ASAP7_75t_R g3338 ( 
.A(n_1104),
.Y(n_3338)
);

CKINVDCx5p33_ASAP7_75t_R g3339 ( 
.A(n_1238),
.Y(n_3339)
);

CKINVDCx5p33_ASAP7_75t_R g3340 ( 
.A(n_711),
.Y(n_3340)
);

INVx1_ASAP7_75t_L g3341 ( 
.A(n_1106),
.Y(n_3341)
);

INVxp67_ASAP7_75t_L g3342 ( 
.A(n_1592),
.Y(n_3342)
);

CKINVDCx5p33_ASAP7_75t_R g3343 ( 
.A(n_34),
.Y(n_3343)
);

CKINVDCx5p33_ASAP7_75t_R g3344 ( 
.A(n_692),
.Y(n_3344)
);

INVx1_ASAP7_75t_L g3345 ( 
.A(n_1494),
.Y(n_3345)
);

CKINVDCx5p33_ASAP7_75t_R g3346 ( 
.A(n_982),
.Y(n_3346)
);

INVx1_ASAP7_75t_L g3347 ( 
.A(n_705),
.Y(n_3347)
);

INVx1_ASAP7_75t_L g3348 ( 
.A(n_1852),
.Y(n_3348)
);

CKINVDCx5p33_ASAP7_75t_R g3349 ( 
.A(n_531),
.Y(n_3349)
);

CKINVDCx5p33_ASAP7_75t_R g3350 ( 
.A(n_1448),
.Y(n_3350)
);

CKINVDCx5p33_ASAP7_75t_R g3351 ( 
.A(n_1126),
.Y(n_3351)
);

CKINVDCx5p33_ASAP7_75t_R g3352 ( 
.A(n_1972),
.Y(n_3352)
);

INVx1_ASAP7_75t_L g3353 ( 
.A(n_2040),
.Y(n_3353)
);

CKINVDCx5p33_ASAP7_75t_R g3354 ( 
.A(n_487),
.Y(n_3354)
);

BUFx3_ASAP7_75t_L g3355 ( 
.A(n_899),
.Y(n_3355)
);

CKINVDCx5p33_ASAP7_75t_R g3356 ( 
.A(n_804),
.Y(n_3356)
);

CKINVDCx5p33_ASAP7_75t_R g3357 ( 
.A(n_2191),
.Y(n_3357)
);

BUFx10_ASAP7_75t_L g3358 ( 
.A(n_324),
.Y(n_3358)
);

INVx1_ASAP7_75t_L g3359 ( 
.A(n_2112),
.Y(n_3359)
);

CKINVDCx5p33_ASAP7_75t_R g3360 ( 
.A(n_1050),
.Y(n_3360)
);

CKINVDCx5p33_ASAP7_75t_R g3361 ( 
.A(n_770),
.Y(n_3361)
);

CKINVDCx5p33_ASAP7_75t_R g3362 ( 
.A(n_2190),
.Y(n_3362)
);

CKINVDCx5p33_ASAP7_75t_R g3363 ( 
.A(n_1500),
.Y(n_3363)
);

CKINVDCx5p33_ASAP7_75t_R g3364 ( 
.A(n_498),
.Y(n_3364)
);

CKINVDCx5p33_ASAP7_75t_R g3365 ( 
.A(n_580),
.Y(n_3365)
);

INVx1_ASAP7_75t_L g3366 ( 
.A(n_621),
.Y(n_3366)
);

CKINVDCx5p33_ASAP7_75t_R g3367 ( 
.A(n_1813),
.Y(n_3367)
);

CKINVDCx5p33_ASAP7_75t_R g3368 ( 
.A(n_1058),
.Y(n_3368)
);

INVx1_ASAP7_75t_L g3369 ( 
.A(n_1591),
.Y(n_3369)
);

CKINVDCx5p33_ASAP7_75t_R g3370 ( 
.A(n_1017),
.Y(n_3370)
);

INVx1_ASAP7_75t_L g3371 ( 
.A(n_1353),
.Y(n_3371)
);

CKINVDCx5p33_ASAP7_75t_R g3372 ( 
.A(n_1136),
.Y(n_3372)
);

INVx1_ASAP7_75t_L g3373 ( 
.A(n_1081),
.Y(n_3373)
);

CKINVDCx5p33_ASAP7_75t_R g3374 ( 
.A(n_435),
.Y(n_3374)
);

INVx1_ASAP7_75t_SL g3375 ( 
.A(n_416),
.Y(n_3375)
);

CKINVDCx20_ASAP7_75t_R g3376 ( 
.A(n_1756),
.Y(n_3376)
);

CKINVDCx5p33_ASAP7_75t_R g3377 ( 
.A(n_2006),
.Y(n_3377)
);

CKINVDCx5p33_ASAP7_75t_R g3378 ( 
.A(n_1163),
.Y(n_3378)
);

INVx1_ASAP7_75t_SL g3379 ( 
.A(n_366),
.Y(n_3379)
);

CKINVDCx5p33_ASAP7_75t_R g3380 ( 
.A(n_1000),
.Y(n_3380)
);

CKINVDCx20_ASAP7_75t_R g3381 ( 
.A(n_662),
.Y(n_3381)
);

INVx1_ASAP7_75t_L g3382 ( 
.A(n_2097),
.Y(n_3382)
);

INVx1_ASAP7_75t_L g3383 ( 
.A(n_618),
.Y(n_3383)
);

INVx1_ASAP7_75t_L g3384 ( 
.A(n_2040),
.Y(n_3384)
);

INVx1_ASAP7_75t_L g3385 ( 
.A(n_2149),
.Y(n_3385)
);

BUFx10_ASAP7_75t_L g3386 ( 
.A(n_1296),
.Y(n_3386)
);

CKINVDCx5p33_ASAP7_75t_R g3387 ( 
.A(n_430),
.Y(n_3387)
);

INVx2_ASAP7_75t_SL g3388 ( 
.A(n_1922),
.Y(n_3388)
);

INVx1_ASAP7_75t_L g3389 ( 
.A(n_682),
.Y(n_3389)
);

INVx1_ASAP7_75t_L g3390 ( 
.A(n_1970),
.Y(n_3390)
);

CKINVDCx14_ASAP7_75t_R g3391 ( 
.A(n_737),
.Y(n_3391)
);

CKINVDCx5p33_ASAP7_75t_R g3392 ( 
.A(n_2086),
.Y(n_3392)
);

CKINVDCx5p33_ASAP7_75t_R g3393 ( 
.A(n_436),
.Y(n_3393)
);

CKINVDCx5p33_ASAP7_75t_R g3394 ( 
.A(n_78),
.Y(n_3394)
);

CKINVDCx5p33_ASAP7_75t_R g3395 ( 
.A(n_341),
.Y(n_3395)
);

CKINVDCx5p33_ASAP7_75t_R g3396 ( 
.A(n_1158),
.Y(n_3396)
);

CKINVDCx5p33_ASAP7_75t_R g3397 ( 
.A(n_2172),
.Y(n_3397)
);

CKINVDCx5p33_ASAP7_75t_R g3398 ( 
.A(n_589),
.Y(n_3398)
);

CKINVDCx5p33_ASAP7_75t_R g3399 ( 
.A(n_1537),
.Y(n_3399)
);

CKINVDCx20_ASAP7_75t_R g3400 ( 
.A(n_403),
.Y(n_3400)
);

INVx1_ASAP7_75t_L g3401 ( 
.A(n_1658),
.Y(n_3401)
);

CKINVDCx5p33_ASAP7_75t_R g3402 ( 
.A(n_787),
.Y(n_3402)
);

INVx2_ASAP7_75t_SL g3403 ( 
.A(n_785),
.Y(n_3403)
);

CKINVDCx5p33_ASAP7_75t_R g3404 ( 
.A(n_2230),
.Y(n_3404)
);

CKINVDCx5p33_ASAP7_75t_R g3405 ( 
.A(n_1235),
.Y(n_3405)
);

CKINVDCx20_ASAP7_75t_R g3406 ( 
.A(n_358),
.Y(n_3406)
);

BUFx2_ASAP7_75t_L g3407 ( 
.A(n_1622),
.Y(n_3407)
);

CKINVDCx5p33_ASAP7_75t_R g3408 ( 
.A(n_2033),
.Y(n_3408)
);

BUFx3_ASAP7_75t_L g3409 ( 
.A(n_2027),
.Y(n_3409)
);

CKINVDCx5p33_ASAP7_75t_R g3410 ( 
.A(n_1660),
.Y(n_3410)
);

INVx2_ASAP7_75t_L g3411 ( 
.A(n_996),
.Y(n_3411)
);

BUFx10_ASAP7_75t_L g3412 ( 
.A(n_2142),
.Y(n_3412)
);

CKINVDCx16_ASAP7_75t_R g3413 ( 
.A(n_1472),
.Y(n_3413)
);

CKINVDCx20_ASAP7_75t_R g3414 ( 
.A(n_785),
.Y(n_3414)
);

INVx1_ASAP7_75t_L g3415 ( 
.A(n_1749),
.Y(n_3415)
);

INVx1_ASAP7_75t_L g3416 ( 
.A(n_706),
.Y(n_3416)
);

BUFx3_ASAP7_75t_L g3417 ( 
.A(n_2101),
.Y(n_3417)
);

INVx1_ASAP7_75t_L g3418 ( 
.A(n_1886),
.Y(n_3418)
);

CKINVDCx16_ASAP7_75t_R g3419 ( 
.A(n_2054),
.Y(n_3419)
);

CKINVDCx5p33_ASAP7_75t_R g3420 ( 
.A(n_1501),
.Y(n_3420)
);

CKINVDCx5p33_ASAP7_75t_R g3421 ( 
.A(n_2238),
.Y(n_3421)
);

CKINVDCx5p33_ASAP7_75t_R g3422 ( 
.A(n_1353),
.Y(n_3422)
);

CKINVDCx14_ASAP7_75t_R g3423 ( 
.A(n_1072),
.Y(n_3423)
);

INVx1_ASAP7_75t_L g3424 ( 
.A(n_2022),
.Y(n_3424)
);

CKINVDCx20_ASAP7_75t_R g3425 ( 
.A(n_641),
.Y(n_3425)
);

CKINVDCx5p33_ASAP7_75t_R g3426 ( 
.A(n_1347),
.Y(n_3426)
);

CKINVDCx5p33_ASAP7_75t_R g3427 ( 
.A(n_434),
.Y(n_3427)
);

CKINVDCx5p33_ASAP7_75t_R g3428 ( 
.A(n_29),
.Y(n_3428)
);

INVx1_ASAP7_75t_L g3429 ( 
.A(n_2085),
.Y(n_3429)
);

INVx1_ASAP7_75t_L g3430 ( 
.A(n_1317),
.Y(n_3430)
);

CKINVDCx5p33_ASAP7_75t_R g3431 ( 
.A(n_376),
.Y(n_3431)
);

CKINVDCx5p33_ASAP7_75t_R g3432 ( 
.A(n_1380),
.Y(n_3432)
);

CKINVDCx5p33_ASAP7_75t_R g3433 ( 
.A(n_2051),
.Y(n_3433)
);

INVx1_ASAP7_75t_L g3434 ( 
.A(n_1312),
.Y(n_3434)
);

CKINVDCx5p33_ASAP7_75t_R g3435 ( 
.A(n_2185),
.Y(n_3435)
);

CKINVDCx5p33_ASAP7_75t_R g3436 ( 
.A(n_2220),
.Y(n_3436)
);

INVx1_ASAP7_75t_L g3437 ( 
.A(n_2119),
.Y(n_3437)
);

CKINVDCx5p33_ASAP7_75t_R g3438 ( 
.A(n_87),
.Y(n_3438)
);

CKINVDCx20_ASAP7_75t_R g3439 ( 
.A(n_2161),
.Y(n_3439)
);

INVx1_ASAP7_75t_L g3440 ( 
.A(n_1238),
.Y(n_3440)
);

INVx1_ASAP7_75t_L g3441 ( 
.A(n_651),
.Y(n_3441)
);

INVx1_ASAP7_75t_L g3442 ( 
.A(n_1466),
.Y(n_3442)
);

INVx2_ASAP7_75t_SL g3443 ( 
.A(n_1438),
.Y(n_3443)
);

INVx1_ASAP7_75t_L g3444 ( 
.A(n_310),
.Y(n_3444)
);

INVx1_ASAP7_75t_L g3445 ( 
.A(n_946),
.Y(n_3445)
);

INVx1_ASAP7_75t_L g3446 ( 
.A(n_791),
.Y(n_3446)
);

CKINVDCx5p33_ASAP7_75t_R g3447 ( 
.A(n_1718),
.Y(n_3447)
);

INVx1_ASAP7_75t_L g3448 ( 
.A(n_1598),
.Y(n_3448)
);

CKINVDCx20_ASAP7_75t_R g3449 ( 
.A(n_223),
.Y(n_3449)
);

INVx1_ASAP7_75t_L g3450 ( 
.A(n_2107),
.Y(n_3450)
);

CKINVDCx5p33_ASAP7_75t_R g3451 ( 
.A(n_1416),
.Y(n_3451)
);

CKINVDCx5p33_ASAP7_75t_R g3452 ( 
.A(n_617),
.Y(n_3452)
);

CKINVDCx5p33_ASAP7_75t_R g3453 ( 
.A(n_2152),
.Y(n_3453)
);

CKINVDCx5p33_ASAP7_75t_R g3454 ( 
.A(n_59),
.Y(n_3454)
);

CKINVDCx5p33_ASAP7_75t_R g3455 ( 
.A(n_563),
.Y(n_3455)
);

CKINVDCx5p33_ASAP7_75t_R g3456 ( 
.A(n_2248),
.Y(n_3456)
);

INVx1_ASAP7_75t_L g3457 ( 
.A(n_2108),
.Y(n_3457)
);

CKINVDCx5p33_ASAP7_75t_R g3458 ( 
.A(n_1872),
.Y(n_3458)
);

CKINVDCx5p33_ASAP7_75t_R g3459 ( 
.A(n_910),
.Y(n_3459)
);

INVx1_ASAP7_75t_L g3460 ( 
.A(n_522),
.Y(n_3460)
);

CKINVDCx5p33_ASAP7_75t_R g3461 ( 
.A(n_458),
.Y(n_3461)
);

CKINVDCx5p33_ASAP7_75t_R g3462 ( 
.A(n_308),
.Y(n_3462)
);

CKINVDCx5p33_ASAP7_75t_R g3463 ( 
.A(n_221),
.Y(n_3463)
);

INVx1_ASAP7_75t_L g3464 ( 
.A(n_2091),
.Y(n_3464)
);

CKINVDCx5p33_ASAP7_75t_R g3465 ( 
.A(n_2103),
.Y(n_3465)
);

CKINVDCx20_ASAP7_75t_R g3466 ( 
.A(n_2073),
.Y(n_3466)
);

CKINVDCx5p33_ASAP7_75t_R g3467 ( 
.A(n_568),
.Y(n_3467)
);

INVx1_ASAP7_75t_L g3468 ( 
.A(n_251),
.Y(n_3468)
);

INVx1_ASAP7_75t_L g3469 ( 
.A(n_91),
.Y(n_3469)
);

CKINVDCx5p33_ASAP7_75t_R g3470 ( 
.A(n_2012),
.Y(n_3470)
);

INVx2_ASAP7_75t_L g3471 ( 
.A(n_2014),
.Y(n_3471)
);

BUFx3_ASAP7_75t_L g3472 ( 
.A(n_1927),
.Y(n_3472)
);

CKINVDCx20_ASAP7_75t_R g3473 ( 
.A(n_242),
.Y(n_3473)
);

CKINVDCx16_ASAP7_75t_R g3474 ( 
.A(n_652),
.Y(n_3474)
);

INVx1_ASAP7_75t_L g3475 ( 
.A(n_1270),
.Y(n_3475)
);

CKINVDCx5p33_ASAP7_75t_R g3476 ( 
.A(n_1300),
.Y(n_3476)
);

INVx1_ASAP7_75t_L g3477 ( 
.A(n_653),
.Y(n_3477)
);

INVx2_ASAP7_75t_L g3478 ( 
.A(n_1011),
.Y(n_3478)
);

BUFx6f_ASAP7_75t_L g3479 ( 
.A(n_504),
.Y(n_3479)
);

INVx1_ASAP7_75t_L g3480 ( 
.A(n_500),
.Y(n_3480)
);

CKINVDCx5p33_ASAP7_75t_R g3481 ( 
.A(n_574),
.Y(n_3481)
);

INVx1_ASAP7_75t_L g3482 ( 
.A(n_637),
.Y(n_3482)
);

CKINVDCx5p33_ASAP7_75t_R g3483 ( 
.A(n_404),
.Y(n_3483)
);

INVx1_ASAP7_75t_L g3484 ( 
.A(n_532),
.Y(n_3484)
);

CKINVDCx5p33_ASAP7_75t_R g3485 ( 
.A(n_1662),
.Y(n_3485)
);

CKINVDCx20_ASAP7_75t_R g3486 ( 
.A(n_2215),
.Y(n_3486)
);

INVx1_ASAP7_75t_L g3487 ( 
.A(n_1934),
.Y(n_3487)
);

CKINVDCx5p33_ASAP7_75t_R g3488 ( 
.A(n_10),
.Y(n_3488)
);

CKINVDCx5p33_ASAP7_75t_R g3489 ( 
.A(n_1224),
.Y(n_3489)
);

CKINVDCx5p33_ASAP7_75t_R g3490 ( 
.A(n_1080),
.Y(n_3490)
);

CKINVDCx5p33_ASAP7_75t_R g3491 ( 
.A(n_1127),
.Y(n_3491)
);

CKINVDCx5p33_ASAP7_75t_R g3492 ( 
.A(n_61),
.Y(n_3492)
);

INVx1_ASAP7_75t_L g3493 ( 
.A(n_1602),
.Y(n_3493)
);

CKINVDCx20_ASAP7_75t_R g3494 ( 
.A(n_1424),
.Y(n_3494)
);

INVx1_ASAP7_75t_L g3495 ( 
.A(n_2233),
.Y(n_3495)
);

CKINVDCx5p33_ASAP7_75t_R g3496 ( 
.A(n_1339),
.Y(n_3496)
);

CKINVDCx5p33_ASAP7_75t_R g3497 ( 
.A(n_265),
.Y(n_3497)
);

INVx2_ASAP7_75t_L g3498 ( 
.A(n_2105),
.Y(n_3498)
);

INVx1_ASAP7_75t_SL g3499 ( 
.A(n_722),
.Y(n_3499)
);

INVx1_ASAP7_75t_SL g3500 ( 
.A(n_1701),
.Y(n_3500)
);

INVx1_ASAP7_75t_L g3501 ( 
.A(n_1412),
.Y(n_3501)
);

HB1xp67_ASAP7_75t_L g3502 ( 
.A(n_1484),
.Y(n_3502)
);

INVx1_ASAP7_75t_L g3503 ( 
.A(n_504),
.Y(n_3503)
);

CKINVDCx5p33_ASAP7_75t_R g3504 ( 
.A(n_1735),
.Y(n_3504)
);

CKINVDCx5p33_ASAP7_75t_R g3505 ( 
.A(n_1767),
.Y(n_3505)
);

CKINVDCx20_ASAP7_75t_R g3506 ( 
.A(n_700),
.Y(n_3506)
);

CKINVDCx5p33_ASAP7_75t_R g3507 ( 
.A(n_2069),
.Y(n_3507)
);

CKINVDCx20_ASAP7_75t_R g3508 ( 
.A(n_1131),
.Y(n_3508)
);

CKINVDCx5p33_ASAP7_75t_R g3509 ( 
.A(n_668),
.Y(n_3509)
);

CKINVDCx5p33_ASAP7_75t_R g3510 ( 
.A(n_1445),
.Y(n_3510)
);

INVx1_ASAP7_75t_L g3511 ( 
.A(n_2049),
.Y(n_3511)
);

CKINVDCx5p33_ASAP7_75t_R g3512 ( 
.A(n_2099),
.Y(n_3512)
);

CKINVDCx20_ASAP7_75t_R g3513 ( 
.A(n_2083),
.Y(n_3513)
);

CKINVDCx16_ASAP7_75t_R g3514 ( 
.A(n_844),
.Y(n_3514)
);

CKINVDCx5p33_ASAP7_75t_R g3515 ( 
.A(n_2007),
.Y(n_3515)
);

CKINVDCx5p33_ASAP7_75t_R g3516 ( 
.A(n_875),
.Y(n_3516)
);

INVx2_ASAP7_75t_L g3517 ( 
.A(n_529),
.Y(n_3517)
);

INVx1_ASAP7_75t_L g3518 ( 
.A(n_718),
.Y(n_3518)
);

CKINVDCx5p33_ASAP7_75t_R g3519 ( 
.A(n_2109),
.Y(n_3519)
);

CKINVDCx16_ASAP7_75t_R g3520 ( 
.A(n_2100),
.Y(n_3520)
);

INVx1_ASAP7_75t_SL g3521 ( 
.A(n_435),
.Y(n_3521)
);

INVx1_ASAP7_75t_L g3522 ( 
.A(n_1323),
.Y(n_3522)
);

CKINVDCx16_ASAP7_75t_R g3523 ( 
.A(n_29),
.Y(n_3523)
);

INVx1_ASAP7_75t_L g3524 ( 
.A(n_1281),
.Y(n_3524)
);

CKINVDCx5p33_ASAP7_75t_R g3525 ( 
.A(n_1295),
.Y(n_3525)
);

CKINVDCx5p33_ASAP7_75t_R g3526 ( 
.A(n_566),
.Y(n_3526)
);

INVx1_ASAP7_75t_L g3527 ( 
.A(n_108),
.Y(n_3527)
);

CKINVDCx5p33_ASAP7_75t_R g3528 ( 
.A(n_2117),
.Y(n_3528)
);

CKINVDCx20_ASAP7_75t_R g3529 ( 
.A(n_1062),
.Y(n_3529)
);

INVx1_ASAP7_75t_L g3530 ( 
.A(n_1811),
.Y(n_3530)
);

BUFx10_ASAP7_75t_L g3531 ( 
.A(n_2090),
.Y(n_3531)
);

INVx1_ASAP7_75t_L g3532 ( 
.A(n_647),
.Y(n_3532)
);

INVx1_ASAP7_75t_L g3533 ( 
.A(n_51),
.Y(n_3533)
);

CKINVDCx5p33_ASAP7_75t_R g3534 ( 
.A(n_1338),
.Y(n_3534)
);

CKINVDCx5p33_ASAP7_75t_R g3535 ( 
.A(n_2158),
.Y(n_3535)
);

INVx1_ASAP7_75t_L g3536 ( 
.A(n_1555),
.Y(n_3536)
);

CKINVDCx5p33_ASAP7_75t_R g3537 ( 
.A(n_294),
.Y(n_3537)
);

INVx1_ASAP7_75t_L g3538 ( 
.A(n_1284),
.Y(n_3538)
);

CKINVDCx5p33_ASAP7_75t_R g3539 ( 
.A(n_2128),
.Y(n_3539)
);

BUFx6f_ASAP7_75t_L g3540 ( 
.A(n_1868),
.Y(n_3540)
);

CKINVDCx5p33_ASAP7_75t_R g3541 ( 
.A(n_1007),
.Y(n_3541)
);

INVx2_ASAP7_75t_L g3542 ( 
.A(n_2019),
.Y(n_3542)
);

CKINVDCx5p33_ASAP7_75t_R g3543 ( 
.A(n_2046),
.Y(n_3543)
);

BUFx10_ASAP7_75t_L g3544 ( 
.A(n_1741),
.Y(n_3544)
);

INVx1_ASAP7_75t_L g3545 ( 
.A(n_14),
.Y(n_3545)
);

CKINVDCx5p33_ASAP7_75t_R g3546 ( 
.A(n_1851),
.Y(n_3546)
);

BUFx2_ASAP7_75t_L g3547 ( 
.A(n_1849),
.Y(n_3547)
);

BUFx10_ASAP7_75t_L g3548 ( 
.A(n_1879),
.Y(n_3548)
);

INVx2_ASAP7_75t_L g3549 ( 
.A(n_70),
.Y(n_3549)
);

CKINVDCx5p33_ASAP7_75t_R g3550 ( 
.A(n_982),
.Y(n_3550)
);

CKINVDCx5p33_ASAP7_75t_R g3551 ( 
.A(n_1651),
.Y(n_3551)
);

CKINVDCx5p33_ASAP7_75t_R g3552 ( 
.A(n_1535),
.Y(n_3552)
);

INVx1_ASAP7_75t_L g3553 ( 
.A(n_201),
.Y(n_3553)
);

CKINVDCx5p33_ASAP7_75t_R g3554 ( 
.A(n_2087),
.Y(n_3554)
);

CKINVDCx20_ASAP7_75t_R g3555 ( 
.A(n_1461),
.Y(n_3555)
);

CKINVDCx5p33_ASAP7_75t_R g3556 ( 
.A(n_458),
.Y(n_3556)
);

INVx1_ASAP7_75t_L g3557 ( 
.A(n_2141),
.Y(n_3557)
);

CKINVDCx5p33_ASAP7_75t_R g3558 ( 
.A(n_1432),
.Y(n_3558)
);

INVx1_ASAP7_75t_L g3559 ( 
.A(n_1263),
.Y(n_3559)
);

INVx1_ASAP7_75t_L g3560 ( 
.A(n_1061),
.Y(n_3560)
);

CKINVDCx5p33_ASAP7_75t_R g3561 ( 
.A(n_1502),
.Y(n_3561)
);

CKINVDCx20_ASAP7_75t_R g3562 ( 
.A(n_178),
.Y(n_3562)
);

INVx1_ASAP7_75t_L g3563 ( 
.A(n_508),
.Y(n_3563)
);

CKINVDCx5p33_ASAP7_75t_R g3564 ( 
.A(n_143),
.Y(n_3564)
);

CKINVDCx5p33_ASAP7_75t_R g3565 ( 
.A(n_1201),
.Y(n_3565)
);

INVx1_ASAP7_75t_L g3566 ( 
.A(n_1645),
.Y(n_3566)
);

CKINVDCx16_ASAP7_75t_R g3567 ( 
.A(n_2045),
.Y(n_3567)
);

INVx1_ASAP7_75t_L g3568 ( 
.A(n_2171),
.Y(n_3568)
);

BUFx6f_ASAP7_75t_L g3569 ( 
.A(n_2106),
.Y(n_3569)
);

INVx2_ASAP7_75t_L g3570 ( 
.A(n_208),
.Y(n_3570)
);

CKINVDCx16_ASAP7_75t_R g3571 ( 
.A(n_1697),
.Y(n_3571)
);

CKINVDCx5p33_ASAP7_75t_R g3572 ( 
.A(n_478),
.Y(n_3572)
);

CKINVDCx5p33_ASAP7_75t_R g3573 ( 
.A(n_341),
.Y(n_3573)
);

INVx2_ASAP7_75t_L g3574 ( 
.A(n_798),
.Y(n_3574)
);

BUFx3_ASAP7_75t_L g3575 ( 
.A(n_1804),
.Y(n_3575)
);

CKINVDCx5p33_ASAP7_75t_R g3576 ( 
.A(n_2179),
.Y(n_3576)
);

CKINVDCx5p33_ASAP7_75t_R g3577 ( 
.A(n_1833),
.Y(n_3577)
);

INVx1_ASAP7_75t_L g3578 ( 
.A(n_128),
.Y(n_3578)
);

CKINVDCx5p33_ASAP7_75t_R g3579 ( 
.A(n_1958),
.Y(n_3579)
);

INVx1_ASAP7_75t_L g3580 ( 
.A(n_55),
.Y(n_3580)
);

CKINVDCx5p33_ASAP7_75t_R g3581 ( 
.A(n_1754),
.Y(n_3581)
);

CKINVDCx5p33_ASAP7_75t_R g3582 ( 
.A(n_864),
.Y(n_3582)
);

CKINVDCx5p33_ASAP7_75t_R g3583 ( 
.A(n_670),
.Y(n_3583)
);

CKINVDCx5p33_ASAP7_75t_R g3584 ( 
.A(n_1273),
.Y(n_3584)
);

BUFx10_ASAP7_75t_L g3585 ( 
.A(n_904),
.Y(n_3585)
);

CKINVDCx5p33_ASAP7_75t_R g3586 ( 
.A(n_2074),
.Y(n_3586)
);

CKINVDCx16_ASAP7_75t_R g3587 ( 
.A(n_616),
.Y(n_3587)
);

INVx1_ASAP7_75t_L g3588 ( 
.A(n_1402),
.Y(n_3588)
);

INVx2_ASAP7_75t_L g3589 ( 
.A(n_833),
.Y(n_3589)
);

CKINVDCx5p33_ASAP7_75t_R g3590 ( 
.A(n_173),
.Y(n_3590)
);

HB1xp67_ASAP7_75t_L g3591 ( 
.A(n_1352),
.Y(n_3591)
);

CKINVDCx5p33_ASAP7_75t_R g3592 ( 
.A(n_2184),
.Y(n_3592)
);

CKINVDCx5p33_ASAP7_75t_R g3593 ( 
.A(n_2076),
.Y(n_3593)
);

CKINVDCx5p33_ASAP7_75t_R g3594 ( 
.A(n_994),
.Y(n_3594)
);

INVx2_ASAP7_75t_SL g3595 ( 
.A(n_703),
.Y(n_3595)
);

INVx1_ASAP7_75t_L g3596 ( 
.A(n_1085),
.Y(n_3596)
);

BUFx3_ASAP7_75t_L g3597 ( 
.A(n_122),
.Y(n_3597)
);

CKINVDCx5p33_ASAP7_75t_R g3598 ( 
.A(n_925),
.Y(n_3598)
);

INVx2_ASAP7_75t_SL g3599 ( 
.A(n_455),
.Y(n_3599)
);

BUFx3_ASAP7_75t_L g3600 ( 
.A(n_799),
.Y(n_3600)
);

CKINVDCx5p33_ASAP7_75t_R g3601 ( 
.A(n_2162),
.Y(n_3601)
);

CKINVDCx5p33_ASAP7_75t_R g3602 ( 
.A(n_252),
.Y(n_3602)
);

INVx2_ASAP7_75t_L g3603 ( 
.A(n_940),
.Y(n_3603)
);

CKINVDCx5p33_ASAP7_75t_R g3604 ( 
.A(n_2174),
.Y(n_3604)
);

INVx2_ASAP7_75t_SL g3605 ( 
.A(n_676),
.Y(n_3605)
);

CKINVDCx5p33_ASAP7_75t_R g3606 ( 
.A(n_1030),
.Y(n_3606)
);

CKINVDCx5p33_ASAP7_75t_R g3607 ( 
.A(n_276),
.Y(n_3607)
);

INVx1_ASAP7_75t_SL g3608 ( 
.A(n_1948),
.Y(n_3608)
);

CKINVDCx5p33_ASAP7_75t_R g3609 ( 
.A(n_2213),
.Y(n_3609)
);

INVx2_ASAP7_75t_L g3610 ( 
.A(n_146),
.Y(n_3610)
);

CKINVDCx5p33_ASAP7_75t_R g3611 ( 
.A(n_2170),
.Y(n_3611)
);

INVx1_ASAP7_75t_L g3612 ( 
.A(n_1842),
.Y(n_3612)
);

INVx2_ASAP7_75t_SL g3613 ( 
.A(n_2191),
.Y(n_3613)
);

INVx1_ASAP7_75t_L g3614 ( 
.A(n_2148),
.Y(n_3614)
);

CKINVDCx5p33_ASAP7_75t_R g3615 ( 
.A(n_1737),
.Y(n_3615)
);

INVx1_ASAP7_75t_L g3616 ( 
.A(n_2137),
.Y(n_3616)
);

CKINVDCx5p33_ASAP7_75t_R g3617 ( 
.A(n_2216),
.Y(n_3617)
);

INVxp67_ASAP7_75t_L g3618 ( 
.A(n_450),
.Y(n_3618)
);

CKINVDCx5p33_ASAP7_75t_R g3619 ( 
.A(n_2196),
.Y(n_3619)
);

INVx2_ASAP7_75t_L g3620 ( 
.A(n_538),
.Y(n_3620)
);

CKINVDCx5p33_ASAP7_75t_R g3621 ( 
.A(n_171),
.Y(n_3621)
);

CKINVDCx16_ASAP7_75t_R g3622 ( 
.A(n_4),
.Y(n_3622)
);

INVx1_ASAP7_75t_L g3623 ( 
.A(n_2053),
.Y(n_3623)
);

CKINVDCx5p33_ASAP7_75t_R g3624 ( 
.A(n_1530),
.Y(n_3624)
);

CKINVDCx5p33_ASAP7_75t_R g3625 ( 
.A(n_1456),
.Y(n_3625)
);

BUFx6f_ASAP7_75t_L g3626 ( 
.A(n_2186),
.Y(n_3626)
);

BUFx2_ASAP7_75t_L g3627 ( 
.A(n_1329),
.Y(n_3627)
);

CKINVDCx5p33_ASAP7_75t_R g3628 ( 
.A(n_1783),
.Y(n_3628)
);

INVx2_ASAP7_75t_L g3629 ( 
.A(n_2337),
.Y(n_3629)
);

INVx3_ASAP7_75t_L g3630 ( 
.A(n_2354),
.Y(n_3630)
);

INVx1_ASAP7_75t_L g3631 ( 
.A(n_2337),
.Y(n_3631)
);

INVxp67_ASAP7_75t_SL g3632 ( 
.A(n_2294),
.Y(n_3632)
);

INVx1_ASAP7_75t_SL g3633 ( 
.A(n_2563),
.Y(n_3633)
);

INVx1_ASAP7_75t_L g3634 ( 
.A(n_2337),
.Y(n_3634)
);

INVxp67_ASAP7_75t_SL g3635 ( 
.A(n_2637),
.Y(n_3635)
);

INVx1_ASAP7_75t_L g3636 ( 
.A(n_2337),
.Y(n_3636)
);

INVxp33_ASAP7_75t_L g3637 ( 
.A(n_3193),
.Y(n_3637)
);

INVx1_ASAP7_75t_L g3638 ( 
.A(n_2337),
.Y(n_3638)
);

BUFx3_ASAP7_75t_L g3639 ( 
.A(n_2311),
.Y(n_3639)
);

CKINVDCx20_ASAP7_75t_R g3640 ( 
.A(n_2670),
.Y(n_3640)
);

INVx1_ASAP7_75t_L g3641 ( 
.A(n_2358),
.Y(n_3641)
);

INVx2_ASAP7_75t_L g3642 ( 
.A(n_2358),
.Y(n_3642)
);

CKINVDCx16_ASAP7_75t_R g3643 ( 
.A(n_3622),
.Y(n_3643)
);

INVxp67_ASAP7_75t_SL g3644 ( 
.A(n_2308),
.Y(n_3644)
);

INVx1_ASAP7_75t_L g3645 ( 
.A(n_2358),
.Y(n_3645)
);

INVx1_ASAP7_75t_L g3646 ( 
.A(n_2358),
.Y(n_3646)
);

CKINVDCx5p33_ASAP7_75t_R g3647 ( 
.A(n_2751),
.Y(n_3647)
);

INVx1_ASAP7_75t_L g3648 ( 
.A(n_2358),
.Y(n_3648)
);

BUFx6f_ASAP7_75t_SL g3649 ( 
.A(n_2345),
.Y(n_3649)
);

INVxp67_ASAP7_75t_SL g3650 ( 
.A(n_2308),
.Y(n_3650)
);

INVxp67_ASAP7_75t_SL g3651 ( 
.A(n_2308),
.Y(n_3651)
);

BUFx2_ASAP7_75t_L g3652 ( 
.A(n_3299),
.Y(n_3652)
);

INVx1_ASAP7_75t_L g3653 ( 
.A(n_2478),
.Y(n_3653)
);

INVx1_ASAP7_75t_L g3654 ( 
.A(n_2478),
.Y(n_3654)
);

INVxp67_ASAP7_75t_SL g3655 ( 
.A(n_2352),
.Y(n_3655)
);

INVx1_ASAP7_75t_L g3656 ( 
.A(n_2478),
.Y(n_3656)
);

INVx1_ASAP7_75t_L g3657 ( 
.A(n_2478),
.Y(n_3657)
);

HB1xp67_ASAP7_75t_L g3658 ( 
.A(n_3391),
.Y(n_3658)
);

INVx1_ASAP7_75t_L g3659 ( 
.A(n_2478),
.Y(n_3659)
);

CKINVDCx5p33_ASAP7_75t_R g3660 ( 
.A(n_2454),
.Y(n_3660)
);

INVx1_ASAP7_75t_L g3661 ( 
.A(n_3112),
.Y(n_3661)
);

CKINVDCx16_ASAP7_75t_R g3662 ( 
.A(n_2327),
.Y(n_3662)
);

INVxp67_ASAP7_75t_L g3663 ( 
.A(n_2750),
.Y(n_3663)
);

CKINVDCx20_ASAP7_75t_R g3664 ( 
.A(n_3132),
.Y(n_3664)
);

INVxp33_ASAP7_75t_L g3665 ( 
.A(n_2882),
.Y(n_3665)
);

INVx1_ASAP7_75t_L g3666 ( 
.A(n_3112),
.Y(n_3666)
);

INVx2_ASAP7_75t_L g3667 ( 
.A(n_3112),
.Y(n_3667)
);

INVx1_ASAP7_75t_L g3668 ( 
.A(n_3112),
.Y(n_3668)
);

INVx2_ASAP7_75t_L g3669 ( 
.A(n_3112),
.Y(n_3669)
);

INVx2_ASAP7_75t_L g3670 ( 
.A(n_3267),
.Y(n_3670)
);

CKINVDCx5p33_ASAP7_75t_R g3671 ( 
.A(n_2419),
.Y(n_3671)
);

CKINVDCx5p33_ASAP7_75t_R g3672 ( 
.A(n_2659),
.Y(n_3672)
);

INVx1_ASAP7_75t_L g3673 ( 
.A(n_3267),
.Y(n_3673)
);

INVx1_ASAP7_75t_L g3674 ( 
.A(n_3267),
.Y(n_3674)
);

INVx1_ASAP7_75t_L g3675 ( 
.A(n_3267),
.Y(n_3675)
);

INVx2_ASAP7_75t_L g3676 ( 
.A(n_3267),
.Y(n_3676)
);

INVx1_ASAP7_75t_L g3677 ( 
.A(n_2771),
.Y(n_3677)
);

INVx1_ASAP7_75t_L g3678 ( 
.A(n_2771),
.Y(n_3678)
);

INVx1_ASAP7_75t_L g3679 ( 
.A(n_2771),
.Y(n_3679)
);

INVxp67_ASAP7_75t_SL g3680 ( 
.A(n_2352),
.Y(n_3680)
);

HB1xp67_ASAP7_75t_L g3681 ( 
.A(n_2695),
.Y(n_3681)
);

INVx1_ASAP7_75t_L g3682 ( 
.A(n_2771),
.Y(n_3682)
);

INVx1_ASAP7_75t_L g3683 ( 
.A(n_2771),
.Y(n_3683)
);

INVx1_ASAP7_75t_L g3684 ( 
.A(n_2873),
.Y(n_3684)
);

INVx1_ASAP7_75t_L g3685 ( 
.A(n_2873),
.Y(n_3685)
);

INVx2_ASAP7_75t_L g3686 ( 
.A(n_2873),
.Y(n_3686)
);

INVx1_ASAP7_75t_L g3687 ( 
.A(n_2873),
.Y(n_3687)
);

CKINVDCx5p33_ASAP7_75t_R g3688 ( 
.A(n_3271),
.Y(n_3688)
);

INVx1_ASAP7_75t_L g3689 ( 
.A(n_2873),
.Y(n_3689)
);

BUFx2_ASAP7_75t_L g3690 ( 
.A(n_2934),
.Y(n_3690)
);

BUFx2_ASAP7_75t_L g3691 ( 
.A(n_3043),
.Y(n_3691)
);

INVx1_ASAP7_75t_L g3692 ( 
.A(n_2900),
.Y(n_3692)
);

INVx1_ASAP7_75t_L g3693 ( 
.A(n_2900),
.Y(n_3693)
);

INVx1_ASAP7_75t_L g3694 ( 
.A(n_2900),
.Y(n_3694)
);

INVx1_ASAP7_75t_L g3695 ( 
.A(n_2900),
.Y(n_3695)
);

INVx1_ASAP7_75t_L g3696 ( 
.A(n_2900),
.Y(n_3696)
);

INVx1_ASAP7_75t_L g3697 ( 
.A(n_2970),
.Y(n_3697)
);

CKINVDCx14_ASAP7_75t_R g3698 ( 
.A(n_3423),
.Y(n_3698)
);

INVx1_ASAP7_75t_L g3699 ( 
.A(n_2970),
.Y(n_3699)
);

INVxp33_ASAP7_75t_SL g3700 ( 
.A(n_2350),
.Y(n_3700)
);

INVx2_ASAP7_75t_L g3701 ( 
.A(n_2970),
.Y(n_3701)
);

INVx1_ASAP7_75t_L g3702 ( 
.A(n_2970),
.Y(n_3702)
);

INVx1_ASAP7_75t_L g3703 ( 
.A(n_2970),
.Y(n_3703)
);

INVx1_ASAP7_75t_L g3704 ( 
.A(n_2975),
.Y(n_3704)
);

INVx1_ASAP7_75t_L g3705 ( 
.A(n_2975),
.Y(n_3705)
);

INVxp67_ASAP7_75t_SL g3706 ( 
.A(n_2352),
.Y(n_3706)
);

INVx1_ASAP7_75t_L g3707 ( 
.A(n_2975),
.Y(n_3707)
);

INVx1_ASAP7_75t_L g3708 ( 
.A(n_2975),
.Y(n_3708)
);

INVxp67_ASAP7_75t_SL g3709 ( 
.A(n_2531),
.Y(n_3709)
);

CKINVDCx5p33_ASAP7_75t_R g3710 ( 
.A(n_3309),
.Y(n_3710)
);

INVx1_ASAP7_75t_L g3711 ( 
.A(n_2975),
.Y(n_3711)
);

INVx1_ASAP7_75t_L g3712 ( 
.A(n_3093),
.Y(n_3712)
);

INVx1_ASAP7_75t_L g3713 ( 
.A(n_3093),
.Y(n_3713)
);

INVxp67_ASAP7_75t_L g3714 ( 
.A(n_3147),
.Y(n_3714)
);

CKINVDCx5p33_ASAP7_75t_R g3715 ( 
.A(n_3474),
.Y(n_3715)
);

HB1xp67_ASAP7_75t_L g3716 ( 
.A(n_3514),
.Y(n_3716)
);

INVx1_ASAP7_75t_L g3717 ( 
.A(n_3093),
.Y(n_3717)
);

BUFx6f_ASAP7_75t_L g3718 ( 
.A(n_2531),
.Y(n_3718)
);

INVxp67_ASAP7_75t_L g3719 ( 
.A(n_3170),
.Y(n_3719)
);

INVxp67_ASAP7_75t_SL g3720 ( 
.A(n_2531),
.Y(n_3720)
);

INVx1_ASAP7_75t_L g3721 ( 
.A(n_3093),
.Y(n_3721)
);

CKINVDCx5p33_ASAP7_75t_R g3722 ( 
.A(n_3523),
.Y(n_3722)
);

CKINVDCx5p33_ASAP7_75t_R g3723 ( 
.A(n_3587),
.Y(n_3723)
);

INVx1_ASAP7_75t_L g3724 ( 
.A(n_3093),
.Y(n_3724)
);

INVx2_ASAP7_75t_L g3725 ( 
.A(n_3294),
.Y(n_3725)
);

INVx1_ASAP7_75t_SL g3726 ( 
.A(n_2365),
.Y(n_3726)
);

INVx1_ASAP7_75t_L g3727 ( 
.A(n_3294),
.Y(n_3727)
);

INVxp67_ASAP7_75t_SL g3728 ( 
.A(n_2605),
.Y(n_3728)
);

INVxp67_ASAP7_75t_L g3729 ( 
.A(n_2409),
.Y(n_3729)
);

INVx1_ASAP7_75t_L g3730 ( 
.A(n_3294),
.Y(n_3730)
);

INVx1_ASAP7_75t_L g3731 ( 
.A(n_3294),
.Y(n_3731)
);

INVxp67_ASAP7_75t_SL g3732 ( 
.A(n_2605),
.Y(n_3732)
);

CKINVDCx16_ASAP7_75t_R g3733 ( 
.A(n_2604),
.Y(n_3733)
);

AND2x4_ASAP7_75t_L g3734 ( 
.A(n_2329),
.B(n_0),
.Y(n_3734)
);

INVxp67_ASAP7_75t_SL g3735 ( 
.A(n_2605),
.Y(n_3735)
);

INVx1_ASAP7_75t_L g3736 ( 
.A(n_3294),
.Y(n_3736)
);

INVxp67_ASAP7_75t_L g3737 ( 
.A(n_2443),
.Y(n_3737)
);

INVxp67_ASAP7_75t_SL g3738 ( 
.A(n_2645),
.Y(n_3738)
);

INVx1_ASAP7_75t_L g3739 ( 
.A(n_3311),
.Y(n_3739)
);

INVx1_ASAP7_75t_L g3740 ( 
.A(n_3311),
.Y(n_3740)
);

INVxp33_ASAP7_75t_SL g3741 ( 
.A(n_3502),
.Y(n_3741)
);

INVxp67_ASAP7_75t_L g3742 ( 
.A(n_2449),
.Y(n_3742)
);

INVxp33_ASAP7_75t_SL g3743 ( 
.A(n_3591),
.Y(n_3743)
);

INVx1_ASAP7_75t_L g3744 ( 
.A(n_3311),
.Y(n_3744)
);

INVx1_ASAP7_75t_L g3745 ( 
.A(n_3311),
.Y(n_3745)
);

INVx2_ASAP7_75t_L g3746 ( 
.A(n_3311),
.Y(n_3746)
);

INVx1_ASAP7_75t_L g3747 ( 
.A(n_2272),
.Y(n_3747)
);

INVx1_ASAP7_75t_L g3748 ( 
.A(n_2277),
.Y(n_3748)
);

INVx1_ASAP7_75t_L g3749 ( 
.A(n_2278),
.Y(n_3749)
);

INVx1_ASAP7_75t_L g3750 ( 
.A(n_2297),
.Y(n_3750)
);

CKINVDCx16_ASAP7_75t_R g3751 ( 
.A(n_2621),
.Y(n_3751)
);

INVxp67_ASAP7_75t_L g3752 ( 
.A(n_2580),
.Y(n_3752)
);

INVx1_ASAP7_75t_L g3753 ( 
.A(n_2314),
.Y(n_3753)
);

CKINVDCx16_ASAP7_75t_R g3754 ( 
.A(n_2784),
.Y(n_3754)
);

INVx1_ASAP7_75t_L g3755 ( 
.A(n_2324),
.Y(n_3755)
);

BUFx2_ASAP7_75t_L g3756 ( 
.A(n_2655),
.Y(n_3756)
);

INVx1_ASAP7_75t_L g3757 ( 
.A(n_2333),
.Y(n_3757)
);

CKINVDCx20_ASAP7_75t_R g3758 ( 
.A(n_2820),
.Y(n_3758)
);

INVx1_ASAP7_75t_L g3759 ( 
.A(n_2336),
.Y(n_3759)
);

INVxp33_ASAP7_75t_SL g3760 ( 
.A(n_2268),
.Y(n_3760)
);

INVxp33_ASAP7_75t_SL g3761 ( 
.A(n_2287),
.Y(n_3761)
);

CKINVDCx14_ASAP7_75t_R g3762 ( 
.A(n_2758),
.Y(n_3762)
);

INVx1_ASAP7_75t_L g3763 ( 
.A(n_2342),
.Y(n_3763)
);

INVx1_ASAP7_75t_L g3764 ( 
.A(n_2359),
.Y(n_3764)
);

INVx1_ASAP7_75t_L g3765 ( 
.A(n_2360),
.Y(n_3765)
);

INVx1_ASAP7_75t_L g3766 ( 
.A(n_2362),
.Y(n_3766)
);

CKINVDCx14_ASAP7_75t_R g3767 ( 
.A(n_2804),
.Y(n_3767)
);

INVxp33_ASAP7_75t_SL g3768 ( 
.A(n_2288),
.Y(n_3768)
);

CKINVDCx20_ASAP7_75t_R g3769 ( 
.A(n_3081),
.Y(n_3769)
);

INVx1_ASAP7_75t_L g3770 ( 
.A(n_2383),
.Y(n_3770)
);

INVx1_ASAP7_75t_L g3771 ( 
.A(n_2389),
.Y(n_3771)
);

INVx1_ASAP7_75t_L g3772 ( 
.A(n_2396),
.Y(n_3772)
);

INVx3_ASAP7_75t_L g3773 ( 
.A(n_2411),
.Y(n_3773)
);

INVx3_ASAP7_75t_L g3774 ( 
.A(n_2481),
.Y(n_3774)
);

INVx2_ASAP7_75t_SL g3775 ( 
.A(n_2345),
.Y(n_3775)
);

INVx1_ASAP7_75t_L g3776 ( 
.A(n_2399),
.Y(n_3776)
);

CKINVDCx20_ASAP7_75t_R g3777 ( 
.A(n_3095),
.Y(n_3777)
);

INVxp67_ASAP7_75t_SL g3778 ( 
.A(n_2645),
.Y(n_3778)
);

INVx1_ASAP7_75t_L g3779 ( 
.A(n_2413),
.Y(n_3779)
);

INVx1_ASAP7_75t_L g3780 ( 
.A(n_2414),
.Y(n_3780)
);

INVx1_ASAP7_75t_L g3781 ( 
.A(n_2423),
.Y(n_3781)
);

CKINVDCx5p33_ASAP7_75t_R g3782 ( 
.A(n_3151),
.Y(n_3782)
);

INVx1_ASAP7_75t_L g3783 ( 
.A(n_2451),
.Y(n_3783)
);

INVxp67_ASAP7_75t_L g3784 ( 
.A(n_2843),
.Y(n_3784)
);

INVx1_ASAP7_75t_L g3785 ( 
.A(n_2453),
.Y(n_3785)
);

BUFx6f_ASAP7_75t_L g3786 ( 
.A(n_2645),
.Y(n_3786)
);

INVx1_ASAP7_75t_L g3787 ( 
.A(n_2474),
.Y(n_3787)
);

CKINVDCx20_ASAP7_75t_R g3788 ( 
.A(n_3413),
.Y(n_3788)
);

CKINVDCx20_ASAP7_75t_R g3789 ( 
.A(n_3419),
.Y(n_3789)
);

INVx2_ASAP7_75t_L g3790 ( 
.A(n_2482),
.Y(n_3790)
);

CKINVDCx20_ASAP7_75t_R g3791 ( 
.A(n_3520),
.Y(n_3791)
);

INVx1_ASAP7_75t_L g3792 ( 
.A(n_2483),
.Y(n_3792)
);

INVxp33_ASAP7_75t_SL g3793 ( 
.A(n_2289),
.Y(n_3793)
);

INVx1_ASAP7_75t_L g3794 ( 
.A(n_2500),
.Y(n_3794)
);

CKINVDCx5p33_ASAP7_75t_R g3795 ( 
.A(n_3567),
.Y(n_3795)
);

INVx1_ASAP7_75t_L g3796 ( 
.A(n_2503),
.Y(n_3796)
);

INVx2_ASAP7_75t_L g3797 ( 
.A(n_2507),
.Y(n_3797)
);

CKINVDCx5p33_ASAP7_75t_R g3798 ( 
.A(n_3571),
.Y(n_3798)
);

INVx2_ASAP7_75t_L g3799 ( 
.A(n_2508),
.Y(n_3799)
);

INVx1_ASAP7_75t_L g3800 ( 
.A(n_2512),
.Y(n_3800)
);

CKINVDCx5p33_ASAP7_75t_R g3801 ( 
.A(n_2879),
.Y(n_3801)
);

INVx1_ASAP7_75t_L g3802 ( 
.A(n_2516),
.Y(n_3802)
);

INVx1_ASAP7_75t_L g3803 ( 
.A(n_2519),
.Y(n_3803)
);

CKINVDCx20_ASAP7_75t_R g3804 ( 
.A(n_2276),
.Y(n_3804)
);

INVxp67_ASAP7_75t_L g3805 ( 
.A(n_3288),
.Y(n_3805)
);

INVx1_ASAP7_75t_L g3806 ( 
.A(n_2552),
.Y(n_3806)
);

INVx2_ASAP7_75t_L g3807 ( 
.A(n_2553),
.Y(n_3807)
);

INVxp33_ASAP7_75t_SL g3808 ( 
.A(n_2290),
.Y(n_3808)
);

INVx1_ASAP7_75t_L g3809 ( 
.A(n_2557),
.Y(n_3809)
);

INVx1_ASAP7_75t_L g3810 ( 
.A(n_2559),
.Y(n_3810)
);

INVx1_ASAP7_75t_L g3811 ( 
.A(n_2566),
.Y(n_3811)
);

CKINVDCx14_ASAP7_75t_R g3812 ( 
.A(n_3407),
.Y(n_3812)
);

INVx1_ASAP7_75t_L g3813 ( 
.A(n_2567),
.Y(n_3813)
);

CKINVDCx5p33_ASAP7_75t_R g3814 ( 
.A(n_2293),
.Y(n_3814)
);

INVxp33_ASAP7_75t_SL g3815 ( 
.A(n_2298),
.Y(n_3815)
);

HB1xp67_ASAP7_75t_L g3816 ( 
.A(n_3621),
.Y(n_3816)
);

INVxp67_ASAP7_75t_SL g3817 ( 
.A(n_2988),
.Y(n_3817)
);

INVxp33_ASAP7_75t_L g3818 ( 
.A(n_3547),
.Y(n_3818)
);

INVx1_ASAP7_75t_L g3819 ( 
.A(n_2581),
.Y(n_3819)
);

INVx1_ASAP7_75t_L g3820 ( 
.A(n_2588),
.Y(n_3820)
);

INVx1_ASAP7_75t_L g3821 ( 
.A(n_2589),
.Y(n_3821)
);

INVx1_ASAP7_75t_L g3822 ( 
.A(n_2611),
.Y(n_3822)
);

INVx1_ASAP7_75t_L g3823 ( 
.A(n_2615),
.Y(n_3823)
);

INVx1_ASAP7_75t_L g3824 ( 
.A(n_2616),
.Y(n_3824)
);

INVx1_ASAP7_75t_L g3825 ( 
.A(n_2630),
.Y(n_3825)
);

INVx1_ASAP7_75t_L g3826 ( 
.A(n_2652),
.Y(n_3826)
);

BUFx6f_ASAP7_75t_L g3827 ( 
.A(n_2988),
.Y(n_3827)
);

INVx1_ASAP7_75t_L g3828 ( 
.A(n_2663),
.Y(n_3828)
);

INVx1_ASAP7_75t_L g3829 ( 
.A(n_2664),
.Y(n_3829)
);

INVx1_ASAP7_75t_L g3830 ( 
.A(n_2667),
.Y(n_3830)
);

CKINVDCx5p33_ASAP7_75t_R g3831 ( 
.A(n_2301),
.Y(n_3831)
);

INVx1_ASAP7_75t_SL g3832 ( 
.A(n_3627),
.Y(n_3832)
);

INVx1_ASAP7_75t_L g3833 ( 
.A(n_2690),
.Y(n_3833)
);

INVxp67_ASAP7_75t_SL g3834 ( 
.A(n_2988),
.Y(n_3834)
);

INVx1_ASAP7_75t_L g3835 ( 
.A(n_2691),
.Y(n_3835)
);

INVx1_ASAP7_75t_L g3836 ( 
.A(n_2692),
.Y(n_3836)
);

CKINVDCx5p33_ASAP7_75t_R g3837 ( 
.A(n_2305),
.Y(n_3837)
);

INVxp33_ASAP7_75t_SL g3838 ( 
.A(n_2307),
.Y(n_3838)
);

INVx1_ASAP7_75t_L g3839 ( 
.A(n_2694),
.Y(n_3839)
);

INVxp33_ASAP7_75t_SL g3840 ( 
.A(n_2315),
.Y(n_3840)
);

INVx1_ASAP7_75t_L g3841 ( 
.A(n_2699),
.Y(n_3841)
);

NOR2xp67_ASAP7_75t_L g3842 ( 
.A(n_2312),
.B(n_0),
.Y(n_3842)
);

INVx1_ASAP7_75t_L g3843 ( 
.A(n_2709),
.Y(n_3843)
);

CKINVDCx20_ASAP7_75t_R g3844 ( 
.A(n_2280),
.Y(n_3844)
);

CKINVDCx20_ASAP7_75t_R g3845 ( 
.A(n_2323),
.Y(n_3845)
);

CKINVDCx5p33_ASAP7_75t_R g3846 ( 
.A(n_2316),
.Y(n_3846)
);

INVx1_ASAP7_75t_L g3847 ( 
.A(n_2730),
.Y(n_3847)
);

BUFx3_ASAP7_75t_L g3848 ( 
.A(n_2397),
.Y(n_3848)
);

CKINVDCx5p33_ASAP7_75t_R g3849 ( 
.A(n_2319),
.Y(n_3849)
);

INVxp67_ASAP7_75t_SL g3850 ( 
.A(n_3009),
.Y(n_3850)
);

BUFx6f_ASAP7_75t_L g3851 ( 
.A(n_3009),
.Y(n_3851)
);

INVx1_ASAP7_75t_L g3852 ( 
.A(n_2757),
.Y(n_3852)
);

INVx1_ASAP7_75t_L g3853 ( 
.A(n_2766),
.Y(n_3853)
);

INVx1_ASAP7_75t_L g3854 ( 
.A(n_2770),
.Y(n_3854)
);

CKINVDCx5p33_ASAP7_75t_R g3855 ( 
.A(n_2321),
.Y(n_3855)
);

NOR2xp67_ASAP7_75t_L g3856 ( 
.A(n_2884),
.B(n_1),
.Y(n_3856)
);

INVx1_ASAP7_75t_SL g3857 ( 
.A(n_2370),
.Y(n_3857)
);

CKINVDCx5p33_ASAP7_75t_R g3858 ( 
.A(n_2338),
.Y(n_3858)
);

INVxp67_ASAP7_75t_L g3859 ( 
.A(n_3152),
.Y(n_3859)
);

BUFx2_ASAP7_75t_L g3860 ( 
.A(n_2416),
.Y(n_3860)
);

INVx2_ASAP7_75t_L g3861 ( 
.A(n_2815),
.Y(n_3861)
);

INVx1_ASAP7_75t_L g3862 ( 
.A(n_2817),
.Y(n_3862)
);

BUFx10_ASAP7_75t_L g3863 ( 
.A(n_2361),
.Y(n_3863)
);

INVx1_ASAP7_75t_L g3864 ( 
.A(n_2828),
.Y(n_3864)
);

CKINVDCx5p33_ASAP7_75t_R g3865 ( 
.A(n_2339),
.Y(n_3865)
);

INVx1_ASAP7_75t_SL g3866 ( 
.A(n_2434),
.Y(n_3866)
);

INVx1_ASAP7_75t_L g3867 ( 
.A(n_2832),
.Y(n_3867)
);

CKINVDCx5p33_ASAP7_75t_R g3868 ( 
.A(n_2346),
.Y(n_3868)
);

INVx1_ASAP7_75t_L g3869 ( 
.A(n_2847),
.Y(n_3869)
);

INVxp33_ASAP7_75t_L g3870 ( 
.A(n_2848),
.Y(n_3870)
);

CKINVDCx20_ASAP7_75t_R g3871 ( 
.A(n_2347),
.Y(n_3871)
);

BUFx2_ASAP7_75t_L g3872 ( 
.A(n_2442),
.Y(n_3872)
);

CKINVDCx5p33_ASAP7_75t_R g3873 ( 
.A(n_2348),
.Y(n_3873)
);

INVx1_ASAP7_75t_L g3874 ( 
.A(n_2850),
.Y(n_3874)
);

CKINVDCx16_ASAP7_75t_R g3875 ( 
.A(n_2427),
.Y(n_3875)
);

CKINVDCx16_ASAP7_75t_R g3876 ( 
.A(n_2427),
.Y(n_3876)
);

CKINVDCx16_ASAP7_75t_R g3877 ( 
.A(n_2656),
.Y(n_3877)
);

INVx1_ASAP7_75t_L g3878 ( 
.A(n_2852),
.Y(n_3878)
);

INVx1_ASAP7_75t_L g3879 ( 
.A(n_2856),
.Y(n_3879)
);

BUFx2_ASAP7_75t_L g3880 ( 
.A(n_2540),
.Y(n_3880)
);

BUFx6f_ASAP7_75t_L g3881 ( 
.A(n_3009),
.Y(n_3881)
);

CKINVDCx5p33_ASAP7_75t_R g3882 ( 
.A(n_2356),
.Y(n_3882)
);

INVx1_ASAP7_75t_L g3883 ( 
.A(n_2863),
.Y(n_3883)
);

CKINVDCx5p33_ASAP7_75t_R g3884 ( 
.A(n_2368),
.Y(n_3884)
);

CKINVDCx14_ASAP7_75t_R g3885 ( 
.A(n_2656),
.Y(n_3885)
);

CKINVDCx14_ASAP7_75t_R g3886 ( 
.A(n_2791),
.Y(n_3886)
);

INVxp67_ASAP7_75t_SL g3887 ( 
.A(n_3109),
.Y(n_3887)
);

INVx1_ASAP7_75t_L g3888 ( 
.A(n_2870),
.Y(n_3888)
);

CKINVDCx14_ASAP7_75t_R g3889 ( 
.A(n_2791),
.Y(n_3889)
);

INVx1_ASAP7_75t_L g3890 ( 
.A(n_2875),
.Y(n_3890)
);

INVx1_ASAP7_75t_L g3891 ( 
.A(n_2876),
.Y(n_3891)
);

INVx1_ASAP7_75t_L g3892 ( 
.A(n_2898),
.Y(n_3892)
);

INVx2_ASAP7_75t_L g3893 ( 
.A(n_2899),
.Y(n_3893)
);

CKINVDCx20_ASAP7_75t_R g3894 ( 
.A(n_2353),
.Y(n_3894)
);

INVx1_ASAP7_75t_L g3895 ( 
.A(n_2913),
.Y(n_3895)
);

INVx1_ASAP7_75t_L g3896 ( 
.A(n_2914),
.Y(n_3896)
);

INVxp67_ASAP7_75t_SL g3897 ( 
.A(n_3109),
.Y(n_3897)
);

CKINVDCx20_ASAP7_75t_R g3898 ( 
.A(n_2388),
.Y(n_3898)
);

INVx2_ASAP7_75t_L g3899 ( 
.A(n_2920),
.Y(n_3899)
);

INVx2_ASAP7_75t_L g3900 ( 
.A(n_2939),
.Y(n_3900)
);

BUFx3_ASAP7_75t_L g3901 ( 
.A(n_2596),
.Y(n_3901)
);

INVx1_ASAP7_75t_L g3902 ( 
.A(n_2941),
.Y(n_3902)
);

INVxp67_ASAP7_75t_L g3903 ( 
.A(n_2963),
.Y(n_3903)
);

INVx1_ASAP7_75t_L g3904 ( 
.A(n_2947),
.Y(n_3904)
);

BUFx3_ASAP7_75t_L g3905 ( 
.A(n_2601),
.Y(n_3905)
);

INVx1_ASAP7_75t_L g3906 ( 
.A(n_2980),
.Y(n_3906)
);

INVx2_ASAP7_75t_L g3907 ( 
.A(n_2989),
.Y(n_3907)
);

INVx1_ASAP7_75t_L g3908 ( 
.A(n_2992),
.Y(n_3908)
);

INVx1_ASAP7_75t_L g3909 ( 
.A(n_3010),
.Y(n_3909)
);

CKINVDCx20_ASAP7_75t_R g3910 ( 
.A(n_2391),
.Y(n_3910)
);

INVx1_ASAP7_75t_L g3911 ( 
.A(n_3025),
.Y(n_3911)
);

CKINVDCx5p33_ASAP7_75t_R g3912 ( 
.A(n_2376),
.Y(n_3912)
);

INVx1_ASAP7_75t_L g3913 ( 
.A(n_3042),
.Y(n_3913)
);

CKINVDCx5p33_ASAP7_75t_R g3914 ( 
.A(n_2378),
.Y(n_3914)
);

INVx1_ASAP7_75t_L g3915 ( 
.A(n_3051),
.Y(n_3915)
);

INVx1_ASAP7_75t_L g3916 ( 
.A(n_3057),
.Y(n_3916)
);

INVx1_ASAP7_75t_L g3917 ( 
.A(n_3069),
.Y(n_3917)
);

INVx1_ASAP7_75t_L g3918 ( 
.A(n_3104),
.Y(n_3918)
);

CKINVDCx5p33_ASAP7_75t_R g3919 ( 
.A(n_2382),
.Y(n_3919)
);

INVx1_ASAP7_75t_L g3920 ( 
.A(n_3117),
.Y(n_3920)
);

INVx1_ASAP7_75t_L g3921 ( 
.A(n_3127),
.Y(n_3921)
);

CKINVDCx5p33_ASAP7_75t_R g3922 ( 
.A(n_2384),
.Y(n_3922)
);

INVx1_ASAP7_75t_L g3923 ( 
.A(n_3137),
.Y(n_3923)
);

INVx1_ASAP7_75t_L g3924 ( 
.A(n_3150),
.Y(n_3924)
);

CKINVDCx5p33_ASAP7_75t_R g3925 ( 
.A(n_2386),
.Y(n_3925)
);

INVx1_ASAP7_75t_L g3926 ( 
.A(n_3164),
.Y(n_3926)
);

INVxp67_ASAP7_75t_L g3927 ( 
.A(n_3358),
.Y(n_3927)
);

CKINVDCx5p33_ASAP7_75t_R g3928 ( 
.A(n_2392),
.Y(n_3928)
);

INVx1_ASAP7_75t_L g3929 ( 
.A(n_3168),
.Y(n_3929)
);

INVx1_ASAP7_75t_L g3930 ( 
.A(n_3184),
.Y(n_3930)
);

INVx1_ASAP7_75t_L g3931 ( 
.A(n_3187),
.Y(n_3931)
);

CKINVDCx5p33_ASAP7_75t_R g3932 ( 
.A(n_2394),
.Y(n_3932)
);

INVxp67_ASAP7_75t_L g3933 ( 
.A(n_2963),
.Y(n_3933)
);

INVx1_ASAP7_75t_L g3934 ( 
.A(n_3194),
.Y(n_3934)
);

INVx1_ASAP7_75t_L g3935 ( 
.A(n_3197),
.Y(n_3935)
);

INVx2_ASAP7_75t_L g3936 ( 
.A(n_3215),
.Y(n_3936)
);

CKINVDCx5p33_ASAP7_75t_R g3937 ( 
.A(n_2420),
.Y(n_3937)
);

CKINVDCx20_ASAP7_75t_R g3938 ( 
.A(n_2404),
.Y(n_3938)
);

INVx1_ASAP7_75t_L g3939 ( 
.A(n_3222),
.Y(n_3939)
);

INVx1_ASAP7_75t_L g3940 ( 
.A(n_3228),
.Y(n_3940)
);

INVx2_ASAP7_75t_L g3941 ( 
.A(n_3229),
.Y(n_3941)
);

INVxp67_ASAP7_75t_SL g3942 ( 
.A(n_3109),
.Y(n_3942)
);

INVx2_ASAP7_75t_L g3943 ( 
.A(n_3257),
.Y(n_3943)
);

INVx1_ASAP7_75t_L g3944 ( 
.A(n_3286),
.Y(n_3944)
);

INVx2_ASAP7_75t_L g3945 ( 
.A(n_3305),
.Y(n_3945)
);

INVxp33_ASAP7_75t_SL g3946 ( 
.A(n_2421),
.Y(n_3946)
);

INVx1_ASAP7_75t_L g3947 ( 
.A(n_3307),
.Y(n_3947)
);

CKINVDCx5p33_ASAP7_75t_R g3948 ( 
.A(n_2425),
.Y(n_3948)
);

CKINVDCx16_ASAP7_75t_R g3949 ( 
.A(n_3152),
.Y(n_3949)
);

INVx1_ASAP7_75t_L g3950 ( 
.A(n_3327),
.Y(n_3950)
);

CKINVDCx20_ASAP7_75t_R g3951 ( 
.A(n_2549),
.Y(n_3951)
);

INVx4_ASAP7_75t_R g3952 ( 
.A(n_2544),
.Y(n_3952)
);

INVx2_ASAP7_75t_L g3953 ( 
.A(n_3330),
.Y(n_3953)
);

INVx2_ASAP7_75t_L g3954 ( 
.A(n_3334),
.Y(n_3954)
);

INVx1_ASAP7_75t_L g3955 ( 
.A(n_3347),
.Y(n_3955)
);

INVx1_ASAP7_75t_L g3956 ( 
.A(n_3366),
.Y(n_3956)
);

INVx1_ASAP7_75t_L g3957 ( 
.A(n_3383),
.Y(n_3957)
);

INVx1_ASAP7_75t_L g3958 ( 
.A(n_3389),
.Y(n_3958)
);

INVx1_ASAP7_75t_L g3959 ( 
.A(n_3416),
.Y(n_3959)
);

INVx1_ASAP7_75t_L g3960 ( 
.A(n_3441),
.Y(n_3960)
);

INVx1_ASAP7_75t_L g3961 ( 
.A(n_3444),
.Y(n_3961)
);

CKINVDCx5p33_ASAP7_75t_R g3962 ( 
.A(n_2428),
.Y(n_3962)
);

INVx1_ASAP7_75t_L g3963 ( 
.A(n_3445),
.Y(n_3963)
);

INVx1_ASAP7_75t_L g3964 ( 
.A(n_3446),
.Y(n_3964)
);

INVxp67_ASAP7_75t_L g3965 ( 
.A(n_3205),
.Y(n_3965)
);

INVx1_ASAP7_75t_L g3966 ( 
.A(n_3460),
.Y(n_3966)
);

INVx1_ASAP7_75t_L g3967 ( 
.A(n_3468),
.Y(n_3967)
);

INVx1_ASAP7_75t_L g3968 ( 
.A(n_3469),
.Y(n_3968)
);

CKINVDCx20_ASAP7_75t_R g3969 ( 
.A(n_2556),
.Y(n_3969)
);

HB1xp67_ASAP7_75t_L g3970 ( 
.A(n_2429),
.Y(n_3970)
);

CKINVDCx5p33_ASAP7_75t_R g3971 ( 
.A(n_2430),
.Y(n_3971)
);

INVxp33_ASAP7_75t_SL g3972 ( 
.A(n_2435),
.Y(n_3972)
);

INVxp33_ASAP7_75t_L g3973 ( 
.A(n_3477),
.Y(n_3973)
);

INVx1_ASAP7_75t_L g3974 ( 
.A(n_3480),
.Y(n_3974)
);

INVx1_ASAP7_75t_L g3975 ( 
.A(n_3482),
.Y(n_3975)
);

INVx1_ASAP7_75t_L g3976 ( 
.A(n_3484),
.Y(n_3976)
);

INVx1_ASAP7_75t_L g3977 ( 
.A(n_3503),
.Y(n_3977)
);

INVx1_ASAP7_75t_L g3978 ( 
.A(n_3518),
.Y(n_3978)
);

CKINVDCx20_ASAP7_75t_R g3979 ( 
.A(n_2606),
.Y(n_3979)
);

INVx1_ASAP7_75t_L g3980 ( 
.A(n_3527),
.Y(n_3980)
);

INVxp67_ASAP7_75t_SL g3981 ( 
.A(n_3479),
.Y(n_3981)
);

INVx1_ASAP7_75t_L g3982 ( 
.A(n_3532),
.Y(n_3982)
);

INVx1_ASAP7_75t_L g3983 ( 
.A(n_3533),
.Y(n_3983)
);

INVx1_ASAP7_75t_L g3984 ( 
.A(n_3545),
.Y(n_3984)
);

INVx1_ASAP7_75t_L g3985 ( 
.A(n_3553),
.Y(n_3985)
);

BUFx6f_ASAP7_75t_L g3986 ( 
.A(n_3479),
.Y(n_3986)
);

CKINVDCx20_ASAP7_75t_R g3987 ( 
.A(n_2629),
.Y(n_3987)
);

INVx1_ASAP7_75t_L g3988 ( 
.A(n_3563),
.Y(n_3988)
);

CKINVDCx5p33_ASAP7_75t_R g3989 ( 
.A(n_2438),
.Y(n_3989)
);

INVx1_ASAP7_75t_L g3990 ( 
.A(n_3578),
.Y(n_3990)
);

BUFx3_ASAP7_75t_L g3991 ( 
.A(n_2764),
.Y(n_3991)
);

INVx3_ASAP7_75t_L g3992 ( 
.A(n_2568),
.Y(n_3992)
);

INVx1_ASAP7_75t_L g3993 ( 
.A(n_3580),
.Y(n_3993)
);

INVx1_ASAP7_75t_L g3994 ( 
.A(n_2794),
.Y(n_3994)
);

INVx1_ASAP7_75t_L g3995 ( 
.A(n_2829),
.Y(n_3995)
);

INVx1_ASAP7_75t_L g3996 ( 
.A(n_2979),
.Y(n_3996)
);

CKINVDCx20_ASAP7_75t_R g3997 ( 
.A(n_2703),
.Y(n_3997)
);

CKINVDCx20_ASAP7_75t_R g3998 ( 
.A(n_2711),
.Y(n_3998)
);

INVx2_ASAP7_75t_L g3999 ( 
.A(n_2387),
.Y(n_3999)
);

INVx1_ASAP7_75t_L g4000 ( 
.A(n_3175),
.Y(n_4000)
);

INVx1_ASAP7_75t_L g4001 ( 
.A(n_3355),
.Y(n_4001)
);

INVx1_ASAP7_75t_L g4002 ( 
.A(n_3597),
.Y(n_4002)
);

HB1xp67_ASAP7_75t_L g4003 ( 
.A(n_2439),
.Y(n_4003)
);

BUFx3_ASAP7_75t_L g4004 ( 
.A(n_3600),
.Y(n_4004)
);

INVx1_ASAP7_75t_L g4005 ( 
.A(n_3479),
.Y(n_4005)
);

CKINVDCx14_ASAP7_75t_R g4006 ( 
.A(n_3205),
.Y(n_4006)
);

CKINVDCx20_ASAP7_75t_R g4007 ( 
.A(n_2713),
.Y(n_4007)
);

INVx1_ASAP7_75t_L g4008 ( 
.A(n_2497),
.Y(n_4008)
);

INVxp67_ASAP7_75t_SL g4009 ( 
.A(n_2322),
.Y(n_4009)
);

INVx2_ASAP7_75t_L g4010 ( 
.A(n_2506),
.Y(n_4010)
);

BUFx6f_ASAP7_75t_L g4011 ( 
.A(n_2322),
.Y(n_4011)
);

CKINVDCx5p33_ASAP7_75t_R g4012 ( 
.A(n_2440),
.Y(n_4012)
);

INVx1_ASAP7_75t_L g4013 ( 
.A(n_2510),
.Y(n_4013)
);

INVx1_ASAP7_75t_L g4014 ( 
.A(n_2518),
.Y(n_4014)
);

INVx2_ASAP7_75t_L g4015 ( 
.A(n_2545),
.Y(n_4015)
);

INVx1_ASAP7_75t_L g4016 ( 
.A(n_2647),
.Y(n_4016)
);

INVx1_ASAP7_75t_L g4017 ( 
.A(n_2689),
.Y(n_4017)
);

INVx1_ASAP7_75t_L g4018 ( 
.A(n_2844),
.Y(n_4018)
);

HB1xp67_ASAP7_75t_L g4019 ( 
.A(n_2455),
.Y(n_4019)
);

INVx1_ASAP7_75t_L g4020 ( 
.A(n_2961),
.Y(n_4020)
);

INVx1_ASAP7_75t_L g4021 ( 
.A(n_3098),
.Y(n_4021)
);

INVxp67_ASAP7_75t_SL g4022 ( 
.A(n_2322),
.Y(n_4022)
);

AND2x2_ASAP7_75t_L g4023 ( 
.A(n_2754),
.B(n_1),
.Y(n_4023)
);

NAND2xp5_ASAP7_75t_L g4024 ( 
.A(n_2466),
.B(n_1),
.Y(n_4024)
);

INVx1_ASAP7_75t_L g4025 ( 
.A(n_3171),
.Y(n_4025)
);

INVx1_ASAP7_75t_L g4026 ( 
.A(n_3172),
.Y(n_4026)
);

CKINVDCx16_ASAP7_75t_R g4027 ( 
.A(n_3297),
.Y(n_4027)
);

INVx2_ASAP7_75t_L g4028 ( 
.A(n_3233),
.Y(n_4028)
);

INVx1_ASAP7_75t_L g4029 ( 
.A(n_3325),
.Y(n_4029)
);

INVxp33_ASAP7_75t_L g4030 ( 
.A(n_3411),
.Y(n_4030)
);

INVxp67_ASAP7_75t_L g4031 ( 
.A(n_3297),
.Y(n_4031)
);

INVx1_ASAP7_75t_L g4032 ( 
.A(n_3478),
.Y(n_4032)
);

CKINVDCx5p33_ASAP7_75t_R g4033 ( 
.A(n_2458),
.Y(n_4033)
);

CKINVDCx20_ASAP7_75t_R g4034 ( 
.A(n_2779),
.Y(n_4034)
);

INVx1_ASAP7_75t_L g4035 ( 
.A(n_3517),
.Y(n_4035)
);

CKINVDCx16_ASAP7_75t_R g4036 ( 
.A(n_3358),
.Y(n_4036)
);

INVx1_ASAP7_75t_L g4037 ( 
.A(n_3549),
.Y(n_4037)
);

INVx1_ASAP7_75t_L g4038 ( 
.A(n_3570),
.Y(n_4038)
);

INVx1_ASAP7_75t_L g4039 ( 
.A(n_3574),
.Y(n_4039)
);

INVx1_ASAP7_75t_L g4040 ( 
.A(n_3589),
.Y(n_4040)
);

INVx1_ASAP7_75t_L g4041 ( 
.A(n_3603),
.Y(n_4041)
);

INVxp33_ASAP7_75t_L g4042 ( 
.A(n_3610),
.Y(n_4042)
);

INVx1_ASAP7_75t_L g4043 ( 
.A(n_3620),
.Y(n_4043)
);

INVx1_ASAP7_75t_L g4044 ( 
.A(n_2355),
.Y(n_4044)
);

INVx2_ASAP7_75t_L g4045 ( 
.A(n_3626),
.Y(n_4045)
);

BUFx8_ASAP7_75t_SL g4046 ( 
.A(n_3652),
.Y(n_4046)
);

BUFx8_ASAP7_75t_SL g4047 ( 
.A(n_3660),
.Y(n_4047)
);

INVx2_ASAP7_75t_L g4048 ( 
.A(n_4045),
.Y(n_4048)
);

NAND2xp5_ASAP7_75t_L g4049 ( 
.A(n_3644),
.B(n_2355),
.Y(n_4049)
);

BUFx8_ASAP7_75t_SL g4050 ( 
.A(n_3647),
.Y(n_4050)
);

INVx1_ASAP7_75t_L g4051 ( 
.A(n_4009),
.Y(n_4051)
);

INVx2_ASAP7_75t_SL g4052 ( 
.A(n_3863),
.Y(n_4052)
);

AND2x2_ASAP7_75t_L g4053 ( 
.A(n_3698),
.B(n_2763),
.Y(n_4053)
);

NOR2xp33_ASAP7_75t_L g4054 ( 
.A(n_3760),
.B(n_3761),
.Y(n_4054)
);

BUFx8_ASAP7_75t_SL g4055 ( 
.A(n_3804),
.Y(n_4055)
);

INVx4_ASAP7_75t_L g4056 ( 
.A(n_3814),
.Y(n_4056)
);

INVx1_ASAP7_75t_L g4057 ( 
.A(n_4022),
.Y(n_4057)
);

BUFx2_ASAP7_75t_L g4058 ( 
.A(n_3758),
.Y(n_4058)
);

BUFx8_ASAP7_75t_SL g4059 ( 
.A(n_3844),
.Y(n_4059)
);

NAND2xp5_ASAP7_75t_L g4060 ( 
.A(n_3650),
.B(n_2355),
.Y(n_4060)
);

AND2x4_ASAP7_75t_L g4061 ( 
.A(n_3658),
.B(n_2955),
.Y(n_4061)
);

OAI21x1_ASAP7_75t_L g4062 ( 
.A1(n_3629),
.A2(n_2317),
.B(n_2281),
.Y(n_4062)
);

INVx1_ASAP7_75t_L g4063 ( 
.A(n_3651),
.Y(n_4063)
);

BUFx6f_ASAP7_75t_L g4064 ( 
.A(n_3986),
.Y(n_4064)
);

INVx1_ASAP7_75t_L g4065 ( 
.A(n_3655),
.Y(n_4065)
);

BUFx6f_ASAP7_75t_L g4066 ( 
.A(n_3986),
.Y(n_4066)
);

INVx5_ASAP7_75t_L g4067 ( 
.A(n_3775),
.Y(n_4067)
);

BUFx6f_ASAP7_75t_L g4068 ( 
.A(n_3986),
.Y(n_4068)
);

INVx5_ASAP7_75t_L g4069 ( 
.A(n_3875),
.Y(n_4069)
);

BUFx6f_ASAP7_75t_L g4070 ( 
.A(n_3718),
.Y(n_4070)
);

HB1xp67_ASAP7_75t_L g4071 ( 
.A(n_3782),
.Y(n_4071)
);

BUFx6f_ASAP7_75t_L g4072 ( 
.A(n_3718),
.Y(n_4072)
);

BUFx8_ASAP7_75t_SL g4073 ( 
.A(n_3845),
.Y(n_4073)
);

BUFx8_ASAP7_75t_L g4074 ( 
.A(n_3649),
.Y(n_4074)
);

BUFx6f_ASAP7_75t_L g4075 ( 
.A(n_3786),
.Y(n_4075)
);

HB1xp67_ASAP7_75t_L g4076 ( 
.A(n_3795),
.Y(n_4076)
);

BUFx3_ASAP7_75t_L g4077 ( 
.A(n_3639),
.Y(n_4077)
);

BUFx2_ASAP7_75t_L g4078 ( 
.A(n_3769),
.Y(n_4078)
);

BUFx6f_ASAP7_75t_L g4079 ( 
.A(n_3786),
.Y(n_4079)
);

CKINVDCx5p33_ASAP7_75t_R g4080 ( 
.A(n_3831),
.Y(n_4080)
);

BUFx8_ASAP7_75t_SL g4081 ( 
.A(n_3871),
.Y(n_4081)
);

BUFx6f_ASAP7_75t_L g4082 ( 
.A(n_3827),
.Y(n_4082)
);

INVx2_ASAP7_75t_L g4083 ( 
.A(n_3827),
.Y(n_4083)
);

INVx5_ASAP7_75t_L g4084 ( 
.A(n_3876),
.Y(n_4084)
);

AND2x4_ASAP7_75t_L g4085 ( 
.A(n_3632),
.B(n_3030),
.Y(n_4085)
);

AND2x4_ASAP7_75t_L g4086 ( 
.A(n_3635),
.B(n_3063),
.Y(n_4086)
);

INVx1_ASAP7_75t_L g4087 ( 
.A(n_3680),
.Y(n_4087)
);

INVx1_ASAP7_75t_L g4088 ( 
.A(n_3706),
.Y(n_4088)
);

BUFx6f_ASAP7_75t_L g4089 ( 
.A(n_3851),
.Y(n_4089)
);

BUFx3_ASAP7_75t_L g4090 ( 
.A(n_3848),
.Y(n_4090)
);

NAND2xp5_ASAP7_75t_L g4091 ( 
.A(n_3709),
.B(n_2364),
.Y(n_4091)
);

INVx1_ASAP7_75t_L g4092 ( 
.A(n_3720),
.Y(n_4092)
);

AOI22xp5_ASAP7_75t_SL g4093 ( 
.A1(n_3777),
.A2(n_2282),
.B1(n_2498),
.B2(n_2379),
.Y(n_4093)
);

CKINVDCx20_ASAP7_75t_R g4094 ( 
.A(n_3894),
.Y(n_4094)
);

AND2x2_ASAP7_75t_L g4095 ( 
.A(n_3860),
.B(n_3079),
.Y(n_4095)
);

AND2x4_ASAP7_75t_L g4096 ( 
.A(n_3663),
.B(n_3156),
.Y(n_4096)
);

NAND2xp5_ASAP7_75t_L g4097 ( 
.A(n_3728),
.B(n_2364),
.Y(n_4097)
);

INVx1_ASAP7_75t_L g4098 ( 
.A(n_3732),
.Y(n_4098)
);

AOI22xp5_ASAP7_75t_SL g4099 ( 
.A1(n_3788),
.A2(n_2529),
.B1(n_2619),
.B2(n_2521),
.Y(n_4099)
);

INVx1_ASAP7_75t_L g4100 ( 
.A(n_3735),
.Y(n_4100)
);

BUFx6f_ASAP7_75t_L g4101 ( 
.A(n_3851),
.Y(n_4101)
);

BUFx3_ASAP7_75t_L g4102 ( 
.A(n_3901),
.Y(n_4102)
);

INVx1_ASAP7_75t_L g4103 ( 
.A(n_3738),
.Y(n_4103)
);

CKINVDCx5p33_ASAP7_75t_R g4104 ( 
.A(n_3837),
.Y(n_4104)
);

INVx1_ASAP7_75t_L g4105 ( 
.A(n_3778),
.Y(n_4105)
);

CKINVDCx5p33_ASAP7_75t_R g4106 ( 
.A(n_3846),
.Y(n_4106)
);

NOR2x1_ASAP7_75t_L g4107 ( 
.A(n_3631),
.B(n_3179),
.Y(n_4107)
);

AOI22x1_ASAP7_75t_SL g4108 ( 
.A1(n_3789),
.A2(n_2719),
.B1(n_2739),
.B2(n_2680),
.Y(n_4108)
);

INVx1_ASAP7_75t_L g4109 ( 
.A(n_3817),
.Y(n_4109)
);

AND2x4_ASAP7_75t_L g4110 ( 
.A(n_3714),
.B(n_3719),
.Y(n_4110)
);

INVx1_ASAP7_75t_L g4111 ( 
.A(n_3834),
.Y(n_4111)
);

CKINVDCx5p33_ASAP7_75t_R g4112 ( 
.A(n_3849),
.Y(n_4112)
);

INVx5_ASAP7_75t_L g4113 ( 
.A(n_3877),
.Y(n_4113)
);

BUFx8_ASAP7_75t_SL g4114 ( 
.A(n_3898),
.Y(n_4114)
);

AOI22xp5_ASAP7_75t_L g4115 ( 
.A1(n_3700),
.A2(n_2470),
.B1(n_2473),
.B2(n_2462),
.Y(n_4115)
);

OAI22xp5_ASAP7_75t_SL g4116 ( 
.A1(n_3791),
.A2(n_2845),
.B1(n_2954),
.B2(n_2897),
.Y(n_4116)
);

INVx2_ASAP7_75t_L g4117 ( 
.A(n_3881),
.Y(n_4117)
);

INVx3_ASAP7_75t_L g4118 ( 
.A(n_3881),
.Y(n_4118)
);

INVx1_ASAP7_75t_L g4119 ( 
.A(n_3850),
.Y(n_4119)
);

INVx2_ASAP7_75t_L g4120 ( 
.A(n_4011),
.Y(n_4120)
);

AND2x4_ASAP7_75t_L g4121 ( 
.A(n_3729),
.B(n_3209),
.Y(n_4121)
);

BUFx6f_ASAP7_75t_L g4122 ( 
.A(n_4011),
.Y(n_4122)
);

AND2x4_ASAP7_75t_L g4123 ( 
.A(n_3737),
.B(n_3234),
.Y(n_4123)
);

BUFx2_ASAP7_75t_L g4124 ( 
.A(n_3640),
.Y(n_4124)
);

INVx3_ASAP7_75t_L g4125 ( 
.A(n_3905),
.Y(n_4125)
);

BUFx6f_ASAP7_75t_L g4126 ( 
.A(n_3991),
.Y(n_4126)
);

AND2x2_ASAP7_75t_L g4127 ( 
.A(n_3872),
.B(n_3880),
.Y(n_4127)
);

INVx1_ASAP7_75t_L g4128 ( 
.A(n_3887),
.Y(n_4128)
);

INVx2_ASAP7_75t_L g4129 ( 
.A(n_3642),
.Y(n_4129)
);

BUFx3_ASAP7_75t_L g4130 ( 
.A(n_4004),
.Y(n_4130)
);

AOI22x1_ASAP7_75t_SL g4131 ( 
.A1(n_3910),
.A2(n_3019),
.B1(n_3032),
.B2(n_3005),
.Y(n_4131)
);

AND2x2_ASAP7_75t_L g4132 ( 
.A(n_3816),
.B(n_3244),
.Y(n_4132)
);

BUFx2_ASAP7_75t_L g4133 ( 
.A(n_3664),
.Y(n_4133)
);

CKINVDCx5p33_ASAP7_75t_R g4134 ( 
.A(n_3855),
.Y(n_4134)
);

CKINVDCx5p33_ASAP7_75t_R g4135 ( 
.A(n_3858),
.Y(n_4135)
);

INVx1_ASAP7_75t_L g4136 ( 
.A(n_3897),
.Y(n_4136)
);

INVx2_ASAP7_75t_SL g4137 ( 
.A(n_3865),
.Y(n_4137)
);

INVx1_ASAP7_75t_L g4138 ( 
.A(n_3942),
.Y(n_4138)
);

BUFx6f_ASAP7_75t_L g4139 ( 
.A(n_3790),
.Y(n_4139)
);

BUFx8_ASAP7_75t_L g4140 ( 
.A(n_3690),
.Y(n_4140)
);

OAI22x1_ASAP7_75t_R g4141 ( 
.A1(n_3938),
.A2(n_3084),
.B1(n_3106),
.B2(n_3053),
.Y(n_4141)
);

BUFx2_ASAP7_75t_L g4142 ( 
.A(n_3798),
.Y(n_4142)
);

BUFx8_ASAP7_75t_SL g4143 ( 
.A(n_3951),
.Y(n_4143)
);

BUFx2_ASAP7_75t_L g4144 ( 
.A(n_3671),
.Y(n_4144)
);

INVx2_ASAP7_75t_L g4145 ( 
.A(n_3667),
.Y(n_4145)
);

INVx2_ASAP7_75t_L g4146 ( 
.A(n_3669),
.Y(n_4146)
);

INVx1_ASAP7_75t_L g4147 ( 
.A(n_3981),
.Y(n_4147)
);

BUFx3_ASAP7_75t_L g4148 ( 
.A(n_3630),
.Y(n_4148)
);

INVx2_ASAP7_75t_SL g4149 ( 
.A(n_3868),
.Y(n_4149)
);

BUFx6f_ASAP7_75t_L g4150 ( 
.A(n_3797),
.Y(n_4150)
);

INVx2_ASAP7_75t_L g4151 ( 
.A(n_3670),
.Y(n_4151)
);

INVx2_ASAP7_75t_L g4152 ( 
.A(n_3676),
.Y(n_4152)
);

BUFx6f_ASAP7_75t_L g4153 ( 
.A(n_3799),
.Y(n_4153)
);

INVx1_ASAP7_75t_L g4154 ( 
.A(n_3634),
.Y(n_4154)
);

INVx2_ASAP7_75t_L g4155 ( 
.A(n_4005),
.Y(n_4155)
);

INVx5_ASAP7_75t_L g4156 ( 
.A(n_3949),
.Y(n_4156)
);

OA21x2_ASAP7_75t_L g4157 ( 
.A1(n_3636),
.A2(n_3641),
.B(n_3638),
.Y(n_4157)
);

CKINVDCx6p67_ASAP7_75t_R g4158 ( 
.A(n_3643),
.Y(n_4158)
);

INVx3_ASAP7_75t_L g4159 ( 
.A(n_3773),
.Y(n_4159)
);

BUFx6f_ASAP7_75t_L g4160 ( 
.A(n_3807),
.Y(n_4160)
);

AND2x4_ASAP7_75t_L g4161 ( 
.A(n_3742),
.B(n_3254),
.Y(n_4161)
);

AND2x2_ASAP7_75t_L g4162 ( 
.A(n_3970),
.B(n_3409),
.Y(n_4162)
);

INVx2_ASAP7_75t_L g4163 ( 
.A(n_3645),
.Y(n_4163)
);

HB1xp67_ASAP7_75t_L g4164 ( 
.A(n_3672),
.Y(n_4164)
);

OA21x2_ASAP7_75t_L g4165 ( 
.A1(n_3646),
.A2(n_2603),
.B(n_2381),
.Y(n_4165)
);

INVx1_ASAP7_75t_L g4166 ( 
.A(n_3648),
.Y(n_4166)
);

BUFx3_ASAP7_75t_L g4167 ( 
.A(n_3774),
.Y(n_4167)
);

INVx2_ASAP7_75t_L g4168 ( 
.A(n_3653),
.Y(n_4168)
);

OAI21x1_ASAP7_75t_L g4169 ( 
.A1(n_3654),
.A2(n_2402),
.B(n_2377),
.Y(n_4169)
);

INVx2_ASAP7_75t_L g4170 ( 
.A(n_3656),
.Y(n_4170)
);

INVx1_ASAP7_75t_L g4171 ( 
.A(n_3657),
.Y(n_4171)
);

BUFx3_ASAP7_75t_L g4172 ( 
.A(n_3992),
.Y(n_4172)
);

XNOR2xp5_ASAP7_75t_L g4173 ( 
.A(n_3969),
.B(n_3120),
.Y(n_4173)
);

AND2x2_ASAP7_75t_L g4174 ( 
.A(n_4003),
.B(n_3417),
.Y(n_4174)
);

BUFx8_ASAP7_75t_L g4175 ( 
.A(n_3691),
.Y(n_4175)
);

AOI22xp5_ASAP7_75t_L g4176 ( 
.A1(n_3741),
.A2(n_2476),
.B1(n_2486),
.B2(n_2475),
.Y(n_4176)
);

HB1xp67_ASAP7_75t_L g4177 ( 
.A(n_3688),
.Y(n_4177)
);

INVx2_ASAP7_75t_L g4178 ( 
.A(n_3659),
.Y(n_4178)
);

INVx2_ASAP7_75t_SL g4179 ( 
.A(n_3873),
.Y(n_4179)
);

AND2x4_ASAP7_75t_L g4180 ( 
.A(n_3752),
.B(n_3472),
.Y(n_4180)
);

INVx1_ASAP7_75t_L g4181 ( 
.A(n_3661),
.Y(n_4181)
);

INVxp67_ASAP7_75t_L g4182 ( 
.A(n_3681),
.Y(n_4182)
);

BUFx2_ASAP7_75t_L g4183 ( 
.A(n_3710),
.Y(n_4183)
);

BUFx6f_ASAP7_75t_L g4184 ( 
.A(n_3861),
.Y(n_4184)
);

INVx2_ASAP7_75t_L g4185 ( 
.A(n_3666),
.Y(n_4185)
);

INVx1_ASAP7_75t_L g4186 ( 
.A(n_3668),
.Y(n_4186)
);

INVxp33_ASAP7_75t_SL g4187 ( 
.A(n_3801),
.Y(n_4187)
);

AND2x2_ASAP7_75t_L g4188 ( 
.A(n_4019),
.B(n_3575),
.Y(n_4188)
);

BUFx12f_ASAP7_75t_L g4189 ( 
.A(n_3715),
.Y(n_4189)
);

INVx3_ASAP7_75t_L g4190 ( 
.A(n_3999),
.Y(n_4190)
);

HB1xp67_ASAP7_75t_L g4191 ( 
.A(n_3722),
.Y(n_4191)
);

INVx1_ASAP7_75t_L g4192 ( 
.A(n_3673),
.Y(n_4192)
);

CKINVDCx5p33_ASAP7_75t_R g4193 ( 
.A(n_3882),
.Y(n_4193)
);

INVx2_ASAP7_75t_L g4194 ( 
.A(n_3674),
.Y(n_4194)
);

INVx3_ASAP7_75t_L g4195 ( 
.A(n_4010),
.Y(n_4195)
);

HB1xp67_ASAP7_75t_L g4196 ( 
.A(n_3723),
.Y(n_4196)
);

INVx5_ASAP7_75t_L g4197 ( 
.A(n_4027),
.Y(n_4197)
);

INVx1_ASAP7_75t_L g4198 ( 
.A(n_3675),
.Y(n_4198)
);

INVx1_ASAP7_75t_L g4199 ( 
.A(n_4044),
.Y(n_4199)
);

BUFx6f_ASAP7_75t_L g4200 ( 
.A(n_3893),
.Y(n_4200)
);

HB1xp67_ASAP7_75t_L g4201 ( 
.A(n_3884),
.Y(n_4201)
);

OAI21x1_ASAP7_75t_L g4202 ( 
.A1(n_3686),
.A2(n_2682),
.B(n_2642),
.Y(n_4202)
);

INVx2_ASAP7_75t_L g4203 ( 
.A(n_3701),
.Y(n_4203)
);

INVxp67_ASAP7_75t_L g4204 ( 
.A(n_3716),
.Y(n_4204)
);

CKINVDCx5p33_ASAP7_75t_R g4205 ( 
.A(n_3912),
.Y(n_4205)
);

OAI22x1_ASAP7_75t_R g4206 ( 
.A1(n_3979),
.A2(n_3185),
.B1(n_3235),
.B2(n_3155),
.Y(n_4206)
);

INVx5_ASAP7_75t_L g4207 ( 
.A(n_4036),
.Y(n_4207)
);

BUFx3_ASAP7_75t_L g4208 ( 
.A(n_3994),
.Y(n_4208)
);

NAND2xp5_ASAP7_75t_L g4209 ( 
.A(n_3914),
.B(n_2364),
.Y(n_4209)
);

INVx1_ASAP7_75t_L g4210 ( 
.A(n_3677),
.Y(n_4210)
);

INVx5_ASAP7_75t_L g4211 ( 
.A(n_3662),
.Y(n_4211)
);

INVx5_ASAP7_75t_L g4212 ( 
.A(n_3756),
.Y(n_4212)
);

BUFx6f_ASAP7_75t_L g4213 ( 
.A(n_3899),
.Y(n_4213)
);

BUFx3_ASAP7_75t_L g4214 ( 
.A(n_3995),
.Y(n_4214)
);

CKINVDCx6p67_ASAP7_75t_R g4215 ( 
.A(n_3733),
.Y(n_4215)
);

BUFx6f_ASAP7_75t_L g4216 ( 
.A(n_3900),
.Y(n_4216)
);

OAI22xp5_ASAP7_75t_L g4217 ( 
.A1(n_3743),
.A2(n_2502),
.B1(n_2525),
.B2(n_2514),
.Y(n_4217)
);

AND2x4_ASAP7_75t_L g4218 ( 
.A(n_3784),
.B(n_2484),
.Y(n_4218)
);

BUFx6f_ASAP7_75t_L g4219 ( 
.A(n_3907),
.Y(n_4219)
);

NOR2xp33_ASAP7_75t_L g4220 ( 
.A(n_3768),
.B(n_3793),
.Y(n_4220)
);

INVx1_ASAP7_75t_L g4221 ( 
.A(n_3678),
.Y(n_4221)
);

AND2x4_ASAP7_75t_L g4222 ( 
.A(n_3805),
.B(n_2609),
.Y(n_4222)
);

INVx5_ASAP7_75t_L g4223 ( 
.A(n_3751),
.Y(n_4223)
);

INVx2_ASAP7_75t_L g4224 ( 
.A(n_3725),
.Y(n_4224)
);

BUFx8_ASAP7_75t_L g4225 ( 
.A(n_3996),
.Y(n_4225)
);

INVx2_ASAP7_75t_L g4226 ( 
.A(n_3746),
.Y(n_4226)
);

AND2x4_ASAP7_75t_L g4227 ( 
.A(n_4023),
.B(n_2732),
.Y(n_4227)
);

INVx5_ASAP7_75t_L g4228 ( 
.A(n_3754),
.Y(n_4228)
);

INVx3_ASAP7_75t_L g4229 ( 
.A(n_4015),
.Y(n_4229)
);

INVx5_ASAP7_75t_L g4230 ( 
.A(n_3734),
.Y(n_4230)
);

INVx1_ASAP7_75t_L g4231 ( 
.A(n_3679),
.Y(n_4231)
);

BUFx3_ASAP7_75t_L g4232 ( 
.A(n_4000),
.Y(n_4232)
);

BUFx3_ASAP7_75t_L g4233 ( 
.A(n_4001),
.Y(n_4233)
);

BUFx12f_ASAP7_75t_L g4234 ( 
.A(n_3919),
.Y(n_4234)
);

HB1xp67_ASAP7_75t_L g4235 ( 
.A(n_3922),
.Y(n_4235)
);

AND2x2_ASAP7_75t_L g4236 ( 
.A(n_3762),
.B(n_3585),
.Y(n_4236)
);

INVx2_ASAP7_75t_L g4237 ( 
.A(n_3936),
.Y(n_4237)
);

NAND2xp5_ASAP7_75t_L g4238 ( 
.A(n_3925),
.B(n_2465),
.Y(n_4238)
);

AOI22xp5_ASAP7_75t_L g4239 ( 
.A1(n_3726),
.A2(n_2541),
.B1(n_2558),
.B2(n_2530),
.Y(n_4239)
);

BUFx12f_ASAP7_75t_L g4240 ( 
.A(n_3928),
.Y(n_4240)
);

INVx2_ASAP7_75t_L g4241 ( 
.A(n_3941),
.Y(n_4241)
);

AOI22xp5_ASAP7_75t_SL g4242 ( 
.A1(n_3818),
.A2(n_3381),
.B1(n_3400),
.B2(n_3304),
.Y(n_4242)
);

BUFx3_ASAP7_75t_L g4243 ( 
.A(n_4002),
.Y(n_4243)
);

INVx3_ASAP7_75t_L g4244 ( 
.A(n_4028),
.Y(n_4244)
);

INVx1_ASAP7_75t_L g4245 ( 
.A(n_3682),
.Y(n_4245)
);

AOI22x1_ASAP7_75t_SL g4246 ( 
.A1(n_3987),
.A2(n_3414),
.B1(n_3425),
.B2(n_3406),
.Y(n_4246)
);

AND2x4_ASAP7_75t_L g4247 ( 
.A(n_3859),
.B(n_2865),
.Y(n_4247)
);

INVx1_ASAP7_75t_L g4248 ( 
.A(n_3683),
.Y(n_4248)
);

INVx1_ASAP7_75t_L g4249 ( 
.A(n_3684),
.Y(n_4249)
);

BUFx3_ASAP7_75t_L g4250 ( 
.A(n_3685),
.Y(n_4250)
);

INVx2_ASAP7_75t_L g4251 ( 
.A(n_3943),
.Y(n_4251)
);

AND2x2_ASAP7_75t_L g4252 ( 
.A(n_3767),
.B(n_3812),
.Y(n_4252)
);

INVx2_ASAP7_75t_L g4253 ( 
.A(n_3945),
.Y(n_4253)
);

INVx1_ASAP7_75t_L g4254 ( 
.A(n_3687),
.Y(n_4254)
);

NAND2xp5_ASAP7_75t_L g4255 ( 
.A(n_3932),
.B(n_2465),
.Y(n_4255)
);

AND2x2_ASAP7_75t_L g4256 ( 
.A(n_3937),
.B(n_3585),
.Y(n_4256)
);

INVx1_ASAP7_75t_L g4257 ( 
.A(n_3689),
.Y(n_4257)
);

NOR2x1_ASAP7_75t_L g4258 ( 
.A(n_3692),
.B(n_2686),
.Y(n_4258)
);

OAI21x1_ASAP7_75t_L g4259 ( 
.A1(n_3693),
.A2(n_2871),
.B(n_2862),
.Y(n_4259)
);

INVx1_ASAP7_75t_L g4260 ( 
.A(n_3694),
.Y(n_4260)
);

INVx2_ASAP7_75t_SL g4261 ( 
.A(n_3948),
.Y(n_4261)
);

INVx1_ASAP7_75t_L g4262 ( 
.A(n_3695),
.Y(n_4262)
);

INVx2_ASAP7_75t_L g4263 ( 
.A(n_3953),
.Y(n_4263)
);

BUFx6f_ASAP7_75t_L g4264 ( 
.A(n_3954),
.Y(n_4264)
);

INVx1_ASAP7_75t_L g4265 ( 
.A(n_3696),
.Y(n_4265)
);

INVx2_ASAP7_75t_L g4266 ( 
.A(n_3697),
.Y(n_4266)
);

NAND2xp5_ASAP7_75t_L g4267 ( 
.A(n_3962),
.B(n_2465),
.Y(n_4267)
);

AOI22xp5_ASAP7_75t_L g4268 ( 
.A1(n_3832),
.A2(n_2569),
.B1(n_2579),
.B2(n_2560),
.Y(n_4268)
);

HB1xp67_ASAP7_75t_L g4269 ( 
.A(n_3971),
.Y(n_4269)
);

INVx2_ASAP7_75t_L g4270 ( 
.A(n_3699),
.Y(n_4270)
);

BUFx6f_ASAP7_75t_L g4271 ( 
.A(n_3747),
.Y(n_4271)
);

BUFx6f_ASAP7_75t_L g4272 ( 
.A(n_3748),
.Y(n_4272)
);

INVx1_ASAP7_75t_L g4273 ( 
.A(n_3702),
.Y(n_4273)
);

HB1xp67_ASAP7_75t_L g4274 ( 
.A(n_3989),
.Y(n_4274)
);

NAND2xp5_ASAP7_75t_L g4275 ( 
.A(n_4012),
.B(n_4033),
.Y(n_4275)
);

INVxp67_ASAP7_75t_L g4276 ( 
.A(n_3857),
.Y(n_4276)
);

INVx1_ASAP7_75t_L g4277 ( 
.A(n_3703),
.Y(n_4277)
);

INVx2_ASAP7_75t_L g4278 ( 
.A(n_3704),
.Y(n_4278)
);

INVx1_ASAP7_75t_L g4279 ( 
.A(n_3705),
.Y(n_4279)
);

INVx2_ASAP7_75t_L g4280 ( 
.A(n_3707),
.Y(n_4280)
);

CKINVDCx20_ASAP7_75t_R g4281 ( 
.A(n_3997),
.Y(n_4281)
);

INVx2_ASAP7_75t_L g4282 ( 
.A(n_3708),
.Y(n_4282)
);

AND2x4_ASAP7_75t_L g4283 ( 
.A(n_3903),
.B(n_3927),
.Y(n_4283)
);

INVx2_ASAP7_75t_L g4284 ( 
.A(n_3711),
.Y(n_4284)
);

INVxp67_ASAP7_75t_L g4285 ( 
.A(n_3866),
.Y(n_4285)
);

HB1xp67_ASAP7_75t_L g4286 ( 
.A(n_3885),
.Y(n_4286)
);

INVx1_ASAP7_75t_L g4287 ( 
.A(n_3712),
.Y(n_4287)
);

BUFx8_ASAP7_75t_SL g4288 ( 
.A(n_3998),
.Y(n_4288)
);

BUFx6f_ASAP7_75t_L g4289 ( 
.A(n_3749),
.Y(n_4289)
);

INVx1_ASAP7_75t_L g4290 ( 
.A(n_3713),
.Y(n_4290)
);

OR2x2_ASAP7_75t_L g4291 ( 
.A(n_3933),
.B(n_2295),
.Y(n_4291)
);

BUFx6f_ASAP7_75t_L g4292 ( 
.A(n_3750),
.Y(n_4292)
);

BUFx8_ASAP7_75t_SL g4293 ( 
.A(n_4007),
.Y(n_4293)
);

OAI22xp5_ASAP7_75t_L g4294 ( 
.A1(n_3665),
.A2(n_2582),
.B1(n_2607),
.B2(n_2583),
.Y(n_4294)
);

AND2x4_ASAP7_75t_L g4295 ( 
.A(n_3965),
.B(n_2883),
.Y(n_4295)
);

INVx1_ASAP7_75t_L g4296 ( 
.A(n_3717),
.Y(n_4296)
);

BUFx6f_ASAP7_75t_L g4297 ( 
.A(n_3753),
.Y(n_4297)
);

INVx5_ASAP7_75t_L g4298 ( 
.A(n_3886),
.Y(n_4298)
);

BUFx6f_ASAP7_75t_L g4299 ( 
.A(n_3755),
.Y(n_4299)
);

OAI22xp5_ASAP7_75t_L g4300 ( 
.A1(n_3637),
.A2(n_2608),
.B1(n_2612),
.B2(n_2610),
.Y(n_4300)
);

BUFx12f_ASAP7_75t_L g4301 ( 
.A(n_3889),
.Y(n_4301)
);

INVx5_ASAP7_75t_L g4302 ( 
.A(n_4006),
.Y(n_4302)
);

CKINVDCx11_ASAP7_75t_R g4303 ( 
.A(n_4034),
.Y(n_4303)
);

INVx3_ASAP7_75t_L g4304 ( 
.A(n_3757),
.Y(n_4304)
);

BUFx6f_ASAP7_75t_L g4305 ( 
.A(n_3759),
.Y(n_4305)
);

BUFx6f_ASAP7_75t_L g4306 ( 
.A(n_3763),
.Y(n_4306)
);

AND2x2_ASAP7_75t_L g4307 ( 
.A(n_4030),
.B(n_2683),
.Y(n_4307)
);

INVx2_ASAP7_75t_L g4308 ( 
.A(n_3721),
.Y(n_4308)
);

INVx2_ASAP7_75t_L g4309 ( 
.A(n_3724),
.Y(n_4309)
);

NAND2xp5_ASAP7_75t_L g4310 ( 
.A(n_3727),
.B(n_2471),
.Y(n_4310)
);

NAND2xp5_ASAP7_75t_L g4311 ( 
.A(n_3730),
.B(n_2471),
.Y(n_4311)
);

INVx1_ASAP7_75t_L g4312 ( 
.A(n_3731),
.Y(n_4312)
);

BUFx6f_ASAP7_75t_L g4313 ( 
.A(n_3764),
.Y(n_4313)
);

OAI21x1_ASAP7_75t_L g4314 ( 
.A1(n_3736),
.A2(n_2904),
.B(n_2874),
.Y(n_4314)
);

CKINVDCx20_ASAP7_75t_R g4315 ( 
.A(n_3633),
.Y(n_4315)
);

BUFx3_ASAP7_75t_L g4316 ( 
.A(n_3739),
.Y(n_4316)
);

BUFx6f_ASAP7_75t_L g4317 ( 
.A(n_3765),
.Y(n_4317)
);

OAI21x1_ASAP7_75t_L g4318 ( 
.A1(n_3740),
.A2(n_3745),
.B(n_3744),
.Y(n_4318)
);

BUFx6f_ASAP7_75t_L g4319 ( 
.A(n_3766),
.Y(n_4319)
);

INVx2_ASAP7_75t_L g4320 ( 
.A(n_3770),
.Y(n_4320)
);

INVx3_ASAP7_75t_L g4321 ( 
.A(n_3771),
.Y(n_4321)
);

INVx1_ASAP7_75t_L g4322 ( 
.A(n_3772),
.Y(n_4322)
);

BUFx6f_ASAP7_75t_L g4323 ( 
.A(n_3776),
.Y(n_4323)
);

INVx1_ASAP7_75t_L g4324 ( 
.A(n_3779),
.Y(n_4324)
);

INVx2_ASAP7_75t_L g4325 ( 
.A(n_3780),
.Y(n_4325)
);

INVx2_ASAP7_75t_L g4326 ( 
.A(n_3781),
.Y(n_4326)
);

OAI21x1_ASAP7_75t_L g4327 ( 
.A1(n_4024),
.A2(n_2982),
.B(n_2915),
.Y(n_4327)
);

OAI22xp5_ASAP7_75t_SL g4328 ( 
.A1(n_3808),
.A2(n_3473),
.B1(n_3506),
.B2(n_3449),
.Y(n_4328)
);

OA21x2_ASAP7_75t_L g4329 ( 
.A1(n_3783),
.A2(n_3007),
.B(n_3001),
.Y(n_4329)
);

CKINVDCx5p33_ASAP7_75t_R g4330 ( 
.A(n_3815),
.Y(n_4330)
);

BUFx6f_ASAP7_75t_L g4331 ( 
.A(n_3785),
.Y(n_4331)
);

NAND2xp5_ASAP7_75t_L g4332 ( 
.A(n_3838),
.B(n_2471),
.Y(n_4332)
);

BUFx12f_ASAP7_75t_L g4333 ( 
.A(n_3952),
.Y(n_4333)
);

BUFx6f_ASAP7_75t_L g4334 ( 
.A(n_3787),
.Y(n_4334)
);

INVx1_ASAP7_75t_L g4335 ( 
.A(n_3792),
.Y(n_4335)
);

INVx2_ASAP7_75t_L g4336 ( 
.A(n_3794),
.Y(n_4336)
);

INVx1_ASAP7_75t_L g4337 ( 
.A(n_3796),
.Y(n_4337)
);

OAI22x1_ASAP7_75t_R g4338 ( 
.A1(n_3800),
.A2(n_3562),
.B1(n_2890),
.B2(n_2912),
.Y(n_4338)
);

INVxp67_ASAP7_75t_L g4339 ( 
.A(n_4031),
.Y(n_4339)
);

AOI22x1_ASAP7_75t_SL g4340 ( 
.A1(n_3802),
.A2(n_2985),
.B1(n_2993),
.B2(n_2842),
.Y(n_4340)
);

OA21x2_ASAP7_75t_L g4341 ( 
.A1(n_3803),
.A2(n_3122),
.B(n_3073),
.Y(n_4341)
);

INVx1_ASAP7_75t_L g4342 ( 
.A(n_3806),
.Y(n_4342)
);

AND2x4_ASAP7_75t_L g4343 ( 
.A(n_3842),
.B(n_2891),
.Y(n_4343)
);

OAI22xp5_ASAP7_75t_L g4344 ( 
.A1(n_3840),
.A2(n_2614),
.B1(n_2627),
.B2(n_2623),
.Y(n_4344)
);

AND2x4_ASAP7_75t_L g4345 ( 
.A(n_3856),
.B(n_2917),
.Y(n_4345)
);

AOI22x1_ASAP7_75t_SL g4346 ( 
.A1(n_3809),
.A2(n_3040),
.B1(n_3068),
.B2(n_2995),
.Y(n_4346)
);

INVxp67_ASAP7_75t_L g4347 ( 
.A(n_3810),
.Y(n_4347)
);

BUFx3_ASAP7_75t_L g4348 ( 
.A(n_3811),
.Y(n_4348)
);

BUFx6f_ASAP7_75t_L g4349 ( 
.A(n_3813),
.Y(n_4349)
);

NAND2xp5_ASAP7_75t_L g4350 ( 
.A(n_3946),
.B(n_2546),
.Y(n_4350)
);

BUFx6f_ASAP7_75t_L g4351 ( 
.A(n_3819),
.Y(n_4351)
);

INVx3_ASAP7_75t_L g4352 ( 
.A(n_3820),
.Y(n_4352)
);

INVx3_ASAP7_75t_L g4353 ( 
.A(n_3821),
.Y(n_4353)
);

AND2x2_ASAP7_75t_L g4354 ( 
.A(n_4042),
.B(n_3870),
.Y(n_4354)
);

BUFx6f_ASAP7_75t_L g4355 ( 
.A(n_3822),
.Y(n_4355)
);

BUFx12f_ASAP7_75t_L g4356 ( 
.A(n_3972),
.Y(n_4356)
);

INVx5_ASAP7_75t_L g4357 ( 
.A(n_3973),
.Y(n_4357)
);

INVx3_ASAP7_75t_L g4358 ( 
.A(n_3823),
.Y(n_4358)
);

NOR2xp33_ASAP7_75t_L g4359 ( 
.A(n_3824),
.B(n_2986),
.Y(n_4359)
);

BUFx2_ASAP7_75t_L g4360 ( 
.A(n_3825),
.Y(n_4360)
);

INVx6_ASAP7_75t_L g4361 ( 
.A(n_3826),
.Y(n_4361)
);

BUFx6f_ASAP7_75t_L g4362 ( 
.A(n_3828),
.Y(n_4362)
);

INVx1_ASAP7_75t_L g4363 ( 
.A(n_3829),
.Y(n_4363)
);

CKINVDCx5p33_ASAP7_75t_R g4364 ( 
.A(n_3830),
.Y(n_4364)
);

INVx3_ASAP7_75t_L g4365 ( 
.A(n_3833),
.Y(n_4365)
);

INVx2_ASAP7_75t_L g4366 ( 
.A(n_3835),
.Y(n_4366)
);

INVx2_ASAP7_75t_L g4367 ( 
.A(n_3836),
.Y(n_4367)
);

INVx3_ASAP7_75t_L g4368 ( 
.A(n_3839),
.Y(n_4368)
);

INVxp67_ASAP7_75t_L g4369 ( 
.A(n_3841),
.Y(n_4369)
);

CKINVDCx16_ASAP7_75t_R g4370 ( 
.A(n_3843),
.Y(n_4370)
);

HB1xp67_ASAP7_75t_L g4371 ( 
.A(n_3847),
.Y(n_4371)
);

AND2x2_ASAP7_75t_SL g4372 ( 
.A(n_3852),
.B(n_2546),
.Y(n_4372)
);

HB1xp67_ASAP7_75t_L g4373 ( 
.A(n_3853),
.Y(n_4373)
);

NAND2xp5_ASAP7_75t_L g4374 ( 
.A(n_3854),
.B(n_2546),
.Y(n_4374)
);

INVx1_ASAP7_75t_L g4375 ( 
.A(n_3862),
.Y(n_4375)
);

BUFx12f_ASAP7_75t_L g4376 ( 
.A(n_3864),
.Y(n_4376)
);

HB1xp67_ASAP7_75t_L g4377 ( 
.A(n_3867),
.Y(n_4377)
);

OA21x2_ASAP7_75t_L g4378 ( 
.A1(n_3869),
.A2(n_3167),
.B(n_3146),
.Y(n_4378)
);

INVx1_ASAP7_75t_L g4379 ( 
.A(n_3874),
.Y(n_4379)
);

INVx1_ASAP7_75t_L g4380 ( 
.A(n_3878),
.Y(n_4380)
);

HB1xp67_ASAP7_75t_L g4381 ( 
.A(n_3879),
.Y(n_4381)
);

OA21x2_ASAP7_75t_L g4382 ( 
.A1(n_3883),
.A2(n_3202),
.B(n_3191),
.Y(n_4382)
);

INVx5_ASAP7_75t_L g4383 ( 
.A(n_3888),
.Y(n_4383)
);

INVx1_ASAP7_75t_L g4384 ( 
.A(n_3890),
.Y(n_4384)
);

INVx2_ASAP7_75t_SL g4385 ( 
.A(n_3891),
.Y(n_4385)
);

BUFx2_ASAP7_75t_L g4386 ( 
.A(n_3892),
.Y(n_4386)
);

BUFx2_ASAP7_75t_L g4387 ( 
.A(n_3895),
.Y(n_4387)
);

OAI22xp5_ASAP7_75t_R g4388 ( 
.A1(n_3896),
.A2(n_2851),
.B1(n_2635),
.B2(n_2636),
.Y(n_4388)
);

INVx2_ASAP7_75t_L g4389 ( 
.A(n_3902),
.Y(n_4389)
);

BUFx12f_ASAP7_75t_L g4390 ( 
.A(n_3904),
.Y(n_4390)
);

CKINVDCx5p33_ASAP7_75t_R g4391 ( 
.A(n_3906),
.Y(n_4391)
);

AND2x6_ASAP7_75t_L g4392 ( 
.A(n_3908),
.B(n_2306),
.Y(n_4392)
);

NOR2xp33_ASAP7_75t_L g4393 ( 
.A(n_3909),
.B(n_3911),
.Y(n_4393)
);

INVx1_ASAP7_75t_L g4394 ( 
.A(n_3913),
.Y(n_4394)
);

NAND2xp5_ASAP7_75t_L g4395 ( 
.A(n_3915),
.B(n_2572),
.Y(n_4395)
);

OA21x2_ASAP7_75t_L g4396 ( 
.A1(n_3916),
.A2(n_3918),
.B(n_3917),
.Y(n_4396)
);

INVxp67_ASAP7_75t_L g4397 ( 
.A(n_3920),
.Y(n_4397)
);

INVx5_ASAP7_75t_L g4398 ( 
.A(n_3921),
.Y(n_4398)
);

INVx1_ASAP7_75t_L g4399 ( 
.A(n_3923),
.Y(n_4399)
);

OA21x2_ASAP7_75t_L g4400 ( 
.A1(n_3924),
.A2(n_3292),
.B(n_3239),
.Y(n_4400)
);

INVx5_ASAP7_75t_L g4401 ( 
.A(n_3926),
.Y(n_4401)
);

NAND2xp5_ASAP7_75t_L g4402 ( 
.A(n_3929),
.B(n_2572),
.Y(n_4402)
);

NOR2xp33_ASAP7_75t_L g4403 ( 
.A(n_3930),
.B(n_3931),
.Y(n_4403)
);

INVx1_ASAP7_75t_L g4404 ( 
.A(n_3934),
.Y(n_4404)
);

INVx1_ASAP7_75t_L g4405 ( 
.A(n_3935),
.Y(n_4405)
);

INVx5_ASAP7_75t_L g4406 ( 
.A(n_3939),
.Y(n_4406)
);

CKINVDCx5p33_ASAP7_75t_R g4407 ( 
.A(n_3940),
.Y(n_4407)
);

BUFx8_ASAP7_75t_SL g4408 ( 
.A(n_3944),
.Y(n_4408)
);

INVx2_ASAP7_75t_L g4409 ( 
.A(n_3947),
.Y(n_4409)
);

INVx3_ASAP7_75t_L g4410 ( 
.A(n_3950),
.Y(n_4410)
);

INVx5_ASAP7_75t_L g4411 ( 
.A(n_3955),
.Y(n_4411)
);

CKINVDCx5p33_ASAP7_75t_R g4412 ( 
.A(n_3956),
.Y(n_4412)
);

BUFx6f_ASAP7_75t_L g4413 ( 
.A(n_3957),
.Y(n_4413)
);

BUFx2_ASAP7_75t_L g4414 ( 
.A(n_3958),
.Y(n_4414)
);

BUFx12f_ASAP7_75t_L g4415 ( 
.A(n_3959),
.Y(n_4415)
);

BUFx6f_ASAP7_75t_L g4416 ( 
.A(n_3960),
.Y(n_4416)
);

BUFx12f_ASAP7_75t_L g4417 ( 
.A(n_3961),
.Y(n_4417)
);

NAND2xp5_ASAP7_75t_L g4418 ( 
.A(n_3963),
.B(n_2572),
.Y(n_4418)
);

HB1xp67_ASAP7_75t_L g4419 ( 
.A(n_3964),
.Y(n_4419)
);

INVx1_ASAP7_75t_L g4420 ( 
.A(n_3966),
.Y(n_4420)
);

INVx1_ASAP7_75t_L g4421 ( 
.A(n_3967),
.Y(n_4421)
);

BUFx3_ASAP7_75t_L g4422 ( 
.A(n_3968),
.Y(n_4422)
);

INVx2_ASAP7_75t_L g4423 ( 
.A(n_3974),
.Y(n_4423)
);

BUFx6f_ASAP7_75t_L g4424 ( 
.A(n_3975),
.Y(n_4424)
);

INVx2_ASAP7_75t_L g4425 ( 
.A(n_3976),
.Y(n_4425)
);

OAI21x1_ASAP7_75t_L g4426 ( 
.A1(n_3977),
.A2(n_3498),
.B(n_3471),
.Y(n_4426)
);

BUFx2_ASAP7_75t_L g4427 ( 
.A(n_3978),
.Y(n_4427)
);

BUFx12f_ASAP7_75t_L g4428 ( 
.A(n_3980),
.Y(n_4428)
);

INVx3_ASAP7_75t_L g4429 ( 
.A(n_3982),
.Y(n_4429)
);

HB1xp67_ASAP7_75t_L g4430 ( 
.A(n_3983),
.Y(n_4430)
);

INVx5_ASAP7_75t_L g4431 ( 
.A(n_3984),
.Y(n_4431)
);

INVx2_ASAP7_75t_L g4432 ( 
.A(n_3985),
.Y(n_4432)
);

INVx2_ASAP7_75t_L g4433 ( 
.A(n_3988),
.Y(n_4433)
);

OAI22x1_ASAP7_75t_SL g4434 ( 
.A1(n_3990),
.A2(n_3099),
.B1(n_3135),
.B2(n_3075),
.Y(n_4434)
);

BUFx6f_ASAP7_75t_L g4435 ( 
.A(n_3993),
.Y(n_4435)
);

BUFx2_ASAP7_75t_L g4436 ( 
.A(n_4008),
.Y(n_4436)
);

AND2x2_ASAP7_75t_L g4437 ( 
.A(n_4013),
.B(n_2463),
.Y(n_4437)
);

BUFx6f_ASAP7_75t_L g4438 ( 
.A(n_4014),
.Y(n_4438)
);

NOR2x1_ASAP7_75t_L g4439 ( 
.A(n_4016),
.B(n_3542),
.Y(n_4439)
);

INVx2_ASAP7_75t_L g4440 ( 
.A(n_4017),
.Y(n_4440)
);

INVx2_ASAP7_75t_L g4441 ( 
.A(n_4018),
.Y(n_4441)
);

INVx1_ASAP7_75t_L g4442 ( 
.A(n_4020),
.Y(n_4442)
);

BUFx6f_ASAP7_75t_L g4443 ( 
.A(n_4021),
.Y(n_4443)
);

BUFx6f_ASAP7_75t_L g4444 ( 
.A(n_4025),
.Y(n_4444)
);

NOR2xp33_ASAP7_75t_L g4445 ( 
.A(n_4026),
.B(n_3403),
.Y(n_4445)
);

INVx5_ASAP7_75t_L g4446 ( 
.A(n_4029),
.Y(n_4446)
);

BUFx6f_ASAP7_75t_L g4447 ( 
.A(n_4032),
.Y(n_4447)
);

BUFx6f_ASAP7_75t_L g4448 ( 
.A(n_4035),
.Y(n_4448)
);

INVx5_ASAP7_75t_L g4449 ( 
.A(n_4037),
.Y(n_4449)
);

INVx2_ASAP7_75t_L g4450 ( 
.A(n_4038),
.Y(n_4450)
);

INVx2_ASAP7_75t_L g4451 ( 
.A(n_4039),
.Y(n_4451)
);

CKINVDCx5p33_ASAP7_75t_R g4452 ( 
.A(n_4040),
.Y(n_4452)
);

NAND2xp5_ASAP7_75t_L g4453 ( 
.A(n_4041),
.B(n_4043),
.Y(n_4453)
);

BUFx2_ASAP7_75t_L g4454 ( 
.A(n_3758),
.Y(n_4454)
);

NAND2xp5_ASAP7_75t_L g4455 ( 
.A(n_3644),
.B(n_2676),
.Y(n_4455)
);

BUFx6f_ASAP7_75t_L g4456 ( 
.A(n_3986),
.Y(n_4456)
);

BUFx8_ASAP7_75t_SL g4457 ( 
.A(n_3652),
.Y(n_4457)
);

BUFx2_ASAP7_75t_L g4458 ( 
.A(n_3758),
.Y(n_4458)
);

BUFx6f_ASAP7_75t_L g4459 ( 
.A(n_3986),
.Y(n_4459)
);

OAI22x1_ASAP7_75t_R g4460 ( 
.A1(n_3804),
.A2(n_3166),
.B1(n_3220),
.B2(n_3165),
.Y(n_4460)
);

BUFx3_ASAP7_75t_L g4461 ( 
.A(n_3639),
.Y(n_4461)
);

AND2x4_ASAP7_75t_L g4462 ( 
.A(n_3658),
.B(n_3595),
.Y(n_4462)
);

AND2x2_ASAP7_75t_L g4463 ( 
.A(n_3698),
.B(n_2495),
.Y(n_4463)
);

BUFx6f_ASAP7_75t_L g4464 ( 
.A(n_3986),
.Y(n_4464)
);

BUFx6f_ASAP7_75t_L g4465 ( 
.A(n_3986),
.Y(n_4465)
);

HB1xp67_ASAP7_75t_L g4466 ( 
.A(n_3782),
.Y(n_4466)
);

AND2x2_ASAP7_75t_L g4467 ( 
.A(n_3698),
.B(n_2821),
.Y(n_4467)
);

HB1xp67_ASAP7_75t_L g4468 ( 
.A(n_3782),
.Y(n_4468)
);

INVx5_ASAP7_75t_L g4469 ( 
.A(n_3863),
.Y(n_4469)
);

INVx2_ASAP7_75t_L g4470 ( 
.A(n_4045),
.Y(n_4470)
);

INVxp67_ASAP7_75t_L g4471 ( 
.A(n_3681),
.Y(n_4471)
);

INVx1_ASAP7_75t_L g4472 ( 
.A(n_4009),
.Y(n_4472)
);

AOI22x1_ASAP7_75t_SL g4473 ( 
.A1(n_3758),
.A2(n_3252),
.B1(n_3253),
.B2(n_3223),
.Y(n_4473)
);

BUFx2_ASAP7_75t_L g4474 ( 
.A(n_3758),
.Y(n_4474)
);

NOR2xp33_ASAP7_75t_L g4475 ( 
.A(n_3760),
.B(n_3599),
.Y(n_4475)
);

BUFx2_ASAP7_75t_L g4476 ( 
.A(n_3758),
.Y(n_4476)
);

AND2x4_ASAP7_75t_L g4477 ( 
.A(n_3658),
.B(n_3605),
.Y(n_4477)
);

BUFx6f_ASAP7_75t_L g4478 ( 
.A(n_3986),
.Y(n_4478)
);

HB1xp67_ASAP7_75t_L g4479 ( 
.A(n_3782),
.Y(n_4479)
);

INVx2_ASAP7_75t_L g4480 ( 
.A(n_4045),
.Y(n_4480)
);

INVx5_ASAP7_75t_L g4481 ( 
.A(n_3863),
.Y(n_4481)
);

INVx2_ASAP7_75t_L g4482 ( 
.A(n_4045),
.Y(n_4482)
);

INVx1_ASAP7_75t_L g4483 ( 
.A(n_4009),
.Y(n_4483)
);

INVx1_ASAP7_75t_L g4484 ( 
.A(n_4009),
.Y(n_4484)
);

BUFx6f_ASAP7_75t_L g4485 ( 
.A(n_3986),
.Y(n_4485)
);

INVx5_ASAP7_75t_L g4486 ( 
.A(n_3863),
.Y(n_4486)
);

AND2x4_ASAP7_75t_L g4487 ( 
.A(n_3658),
.B(n_2840),
.Y(n_4487)
);

NAND2xp5_ASAP7_75t_L g4488 ( 
.A(n_3644),
.B(n_2676),
.Y(n_4488)
);

INVx3_ASAP7_75t_L g4489 ( 
.A(n_3718),
.Y(n_4489)
);

INVx3_ASAP7_75t_L g4490 ( 
.A(n_3718),
.Y(n_4490)
);

AOI22x1_ASAP7_75t_SL g4491 ( 
.A1(n_3758),
.A2(n_3272),
.B1(n_3293),
.B2(n_3263),
.Y(n_4491)
);

NAND2xp5_ASAP7_75t_SL g4492 ( 
.A(n_3733),
.B(n_2676),
.Y(n_4492)
);

AND2x4_ASAP7_75t_L g4493 ( 
.A(n_3658),
.B(n_2902),
.Y(n_4493)
);

CKINVDCx20_ASAP7_75t_R g4494 ( 
.A(n_3804),
.Y(n_4494)
);

INVx5_ASAP7_75t_L g4495 ( 
.A(n_3863),
.Y(n_4495)
);

NOR2xp33_ASAP7_75t_L g4496 ( 
.A(n_3760),
.B(n_2628),
.Y(n_4496)
);

CKINVDCx5p33_ASAP7_75t_R g4497 ( 
.A(n_3660),
.Y(n_4497)
);

CKINVDCx5p33_ASAP7_75t_R g4498 ( 
.A(n_3660),
.Y(n_4498)
);

CKINVDCx5p33_ASAP7_75t_R g4499 ( 
.A(n_3660),
.Y(n_4499)
);

AND2x4_ASAP7_75t_L g4500 ( 
.A(n_3658),
.B(n_2950),
.Y(n_4500)
);

INVx6_ASAP7_75t_L g4501 ( 
.A(n_3863),
.Y(n_4501)
);

INVx2_ASAP7_75t_L g4502 ( 
.A(n_4045),
.Y(n_4502)
);

INVx2_ASAP7_75t_L g4503 ( 
.A(n_4045),
.Y(n_4503)
);

AOI22x1_ASAP7_75t_SL g4504 ( 
.A1(n_3758),
.A2(n_3376),
.B1(n_3439),
.B2(n_3321),
.Y(n_4504)
);

BUFx3_ASAP7_75t_L g4505 ( 
.A(n_3639),
.Y(n_4505)
);

AOI22x1_ASAP7_75t_SL g4506 ( 
.A1(n_3758),
.A2(n_3486),
.B1(n_3494),
.B2(n_3466),
.Y(n_4506)
);

BUFx6f_ASAP7_75t_L g4507 ( 
.A(n_3986),
.Y(n_4507)
);

BUFx12f_ASAP7_75t_L g4508 ( 
.A(n_3660),
.Y(n_4508)
);

BUFx3_ASAP7_75t_L g4509 ( 
.A(n_3639),
.Y(n_4509)
);

INVx1_ASAP7_75t_L g4510 ( 
.A(n_4009),
.Y(n_4510)
);

INVx1_ASAP7_75t_L g4511 ( 
.A(n_4009),
.Y(n_4511)
);

BUFx8_ASAP7_75t_SL g4512 ( 
.A(n_3652),
.Y(n_4512)
);

BUFx8_ASAP7_75t_SL g4513 ( 
.A(n_3652),
.Y(n_4513)
);

BUFx8_ASAP7_75t_SL g4514 ( 
.A(n_3652),
.Y(n_4514)
);

HB1xp67_ASAP7_75t_L g4515 ( 
.A(n_3782),
.Y(n_4515)
);

BUFx3_ASAP7_75t_L g4516 ( 
.A(n_3639),
.Y(n_4516)
);

BUFx3_ASAP7_75t_L g4517 ( 
.A(n_3639),
.Y(n_4517)
);

INVx3_ASAP7_75t_L g4518 ( 
.A(n_3718),
.Y(n_4518)
);

BUFx6f_ASAP7_75t_L g4519 ( 
.A(n_3986),
.Y(n_4519)
);

INVx1_ASAP7_75t_L g4520 ( 
.A(n_4009),
.Y(n_4520)
);

INVx2_ASAP7_75t_L g4521 ( 
.A(n_4045),
.Y(n_4521)
);

BUFx2_ASAP7_75t_L g4522 ( 
.A(n_3758),
.Y(n_4522)
);

AND2x6_ASAP7_75t_L g4523 ( 
.A(n_4023),
.B(n_2448),
.Y(n_4523)
);

BUFx6f_ASAP7_75t_L g4524 ( 
.A(n_3986),
.Y(n_4524)
);

AOI22xp5_ASAP7_75t_L g4525 ( 
.A1(n_3700),
.A2(n_2641),
.B1(n_2657),
.B2(n_2639),
.Y(n_4525)
);

NAND2xp5_ASAP7_75t_L g4526 ( 
.A(n_3644),
.B(n_2708),
.Y(n_4526)
);

INVx2_ASAP7_75t_L g4527 ( 
.A(n_4045),
.Y(n_4527)
);

AND2x6_ASAP7_75t_L g4528 ( 
.A(n_4023),
.B(n_2494),
.Y(n_4528)
);

BUFx3_ASAP7_75t_L g4529 ( 
.A(n_3639),
.Y(n_4529)
);

CKINVDCx20_ASAP7_75t_R g4530 ( 
.A(n_3804),
.Y(n_4530)
);

BUFx12f_ASAP7_75t_L g4531 ( 
.A(n_3660),
.Y(n_4531)
);

INVx2_ASAP7_75t_L g4532 ( 
.A(n_4045),
.Y(n_4532)
);

BUFx3_ASAP7_75t_L g4533 ( 
.A(n_3639),
.Y(n_4533)
);

BUFx8_ASAP7_75t_SL g4534 ( 
.A(n_3652),
.Y(n_4534)
);

HB1xp67_ASAP7_75t_L g4535 ( 
.A(n_3782),
.Y(n_4535)
);

BUFx6f_ASAP7_75t_L g4536 ( 
.A(n_3986),
.Y(n_4536)
);

BUFx6f_ASAP7_75t_L g4537 ( 
.A(n_3986),
.Y(n_4537)
);

CKINVDCx5p33_ASAP7_75t_R g4538 ( 
.A(n_3660),
.Y(n_4538)
);

CKINVDCx5p33_ASAP7_75t_R g4539 ( 
.A(n_3660),
.Y(n_4539)
);

OAI21x1_ASAP7_75t_L g4540 ( 
.A1(n_3629),
.A2(n_2267),
.B(n_2266),
.Y(n_4540)
);

INVx1_ASAP7_75t_L g4541 ( 
.A(n_4009),
.Y(n_4541)
);

AND2x2_ASAP7_75t_L g4542 ( 
.A(n_3698),
.B(n_3388),
.Y(n_4542)
);

INVx2_ASAP7_75t_L g4543 ( 
.A(n_4048),
.Y(n_4543)
);

INVx2_ASAP7_75t_L g4544 ( 
.A(n_4470),
.Y(n_4544)
);

AND2x2_ASAP7_75t_L g4545 ( 
.A(n_4354),
.B(n_2437),
.Y(n_4545)
);

BUFx6f_ASAP7_75t_L g4546 ( 
.A(n_4064),
.Y(n_4546)
);

INVx1_ASAP7_75t_L g4547 ( 
.A(n_4348),
.Y(n_4547)
);

NAND2xp33_ASAP7_75t_L g4548 ( 
.A(n_4523),
.B(n_2708),
.Y(n_4548)
);

INVx1_ASAP7_75t_L g4549 ( 
.A(n_4422),
.Y(n_4549)
);

CKINVDCx5p33_ASAP7_75t_R g4550 ( 
.A(n_4055),
.Y(n_4550)
);

NAND2xp5_ASAP7_75t_L g4551 ( 
.A(n_4372),
.B(n_2708),
.Y(n_4551)
);

AND2x2_ASAP7_75t_L g4552 ( 
.A(n_4127),
.B(n_2437),
.Y(n_4552)
);

NOR2xp33_ASAP7_75t_L g4553 ( 
.A(n_4275),
.B(n_2665),
.Y(n_4553)
);

INVx1_ASAP7_75t_L g4554 ( 
.A(n_4322),
.Y(n_4554)
);

INVx1_ASAP7_75t_L g4555 ( 
.A(n_4324),
.Y(n_4555)
);

INVx1_ASAP7_75t_L g4556 ( 
.A(n_4335),
.Y(n_4556)
);

INVx2_ASAP7_75t_L g4557 ( 
.A(n_4480),
.Y(n_4557)
);

CKINVDCx5p33_ASAP7_75t_R g4558 ( 
.A(n_4059),
.Y(n_4558)
);

INVx1_ASAP7_75t_L g4559 ( 
.A(n_4337),
.Y(n_4559)
);

AND2x4_ASAP7_75t_L g4560 ( 
.A(n_4230),
.B(n_3443),
.Y(n_4560)
);

INVx1_ASAP7_75t_L g4561 ( 
.A(n_4342),
.Y(n_4561)
);

INVx1_ASAP7_75t_L g4562 ( 
.A(n_4363),
.Y(n_4562)
);

AND2x2_ASAP7_75t_L g4563 ( 
.A(n_4357),
.B(n_4252),
.Y(n_4563)
);

INVx2_ASAP7_75t_L g4564 ( 
.A(n_4482),
.Y(n_4564)
);

HB1xp67_ASAP7_75t_L g4565 ( 
.A(n_4276),
.Y(n_4565)
);

BUFx2_ASAP7_75t_L g4566 ( 
.A(n_4285),
.Y(n_4566)
);

INVx3_ASAP7_75t_L g4567 ( 
.A(n_4126),
.Y(n_4567)
);

INVx2_ASAP7_75t_L g4568 ( 
.A(n_4502),
.Y(n_4568)
);

INVx1_ASAP7_75t_L g4569 ( 
.A(n_4375),
.Y(n_4569)
);

INVx1_ASAP7_75t_L g4570 ( 
.A(n_4379),
.Y(n_4570)
);

NAND2xp5_ASAP7_75t_L g4571 ( 
.A(n_4209),
.B(n_4238),
.Y(n_4571)
);

INVx2_ASAP7_75t_L g4572 ( 
.A(n_4503),
.Y(n_4572)
);

INVx3_ASAP7_75t_L g4573 ( 
.A(n_4122),
.Y(n_4573)
);

INVx2_ASAP7_75t_L g4574 ( 
.A(n_4521),
.Y(n_4574)
);

HB1xp67_ASAP7_75t_L g4575 ( 
.A(n_4125),
.Y(n_4575)
);

NOR2x1_ASAP7_75t_L g4576 ( 
.A(n_4056),
.B(n_2275),
.Y(n_4576)
);

NAND2xp5_ASAP7_75t_SL g4577 ( 
.A(n_4469),
.B(n_2721),
.Y(n_4577)
);

NAND2xp5_ASAP7_75t_L g4578 ( 
.A(n_4255),
.B(n_4267),
.Y(n_4578)
);

NAND2xp5_ASAP7_75t_SL g4579 ( 
.A(n_4481),
.B(n_4486),
.Y(n_4579)
);

INVx2_ASAP7_75t_L g4580 ( 
.A(n_4527),
.Y(n_4580)
);

NAND2xp5_ASAP7_75t_L g4581 ( 
.A(n_4250),
.B(n_2721),
.Y(n_4581)
);

BUFx6f_ASAP7_75t_L g4582 ( 
.A(n_4066),
.Y(n_4582)
);

BUFx6f_ASAP7_75t_L g4583 ( 
.A(n_4068),
.Y(n_4583)
);

AND2x2_ASAP7_75t_L g4584 ( 
.A(n_4236),
.B(n_2456),
.Y(n_4584)
);

NAND2xp5_ASAP7_75t_L g4585 ( 
.A(n_4316),
.B(n_2721),
.Y(n_4585)
);

INVx4_ASAP7_75t_L g4586 ( 
.A(n_4333),
.Y(n_4586)
);

INVx1_ASAP7_75t_L g4587 ( 
.A(n_4380),
.Y(n_4587)
);

CKINVDCx5p33_ASAP7_75t_R g4588 ( 
.A(n_4073),
.Y(n_4588)
);

INVxp67_ASAP7_75t_L g4589 ( 
.A(n_4291),
.Y(n_4589)
);

INVx1_ASAP7_75t_L g4590 ( 
.A(n_4384),
.Y(n_4590)
);

NAND2xp5_ASAP7_75t_SL g4591 ( 
.A(n_4495),
.B(n_2772),
.Y(n_4591)
);

INVx1_ASAP7_75t_L g4592 ( 
.A(n_4394),
.Y(n_4592)
);

INVx1_ASAP7_75t_L g4593 ( 
.A(n_4399),
.Y(n_4593)
);

INVx2_ASAP7_75t_L g4594 ( 
.A(n_4532),
.Y(n_4594)
);

NAND2xp5_ASAP7_75t_L g4595 ( 
.A(n_4154),
.B(n_2772),
.Y(n_4595)
);

HB1xp67_ASAP7_75t_L g4596 ( 
.A(n_4148),
.Y(n_4596)
);

INVx1_ASAP7_75t_L g4597 ( 
.A(n_4404),
.Y(n_4597)
);

AND2x4_ASAP7_75t_L g4598 ( 
.A(n_4077),
.B(n_3613),
.Y(n_4598)
);

INVx1_ASAP7_75t_L g4599 ( 
.A(n_4405),
.Y(n_4599)
);

INVx2_ASAP7_75t_L g4600 ( 
.A(n_4129),
.Y(n_4600)
);

INVx4_ASAP7_75t_L g4601 ( 
.A(n_4211),
.Y(n_4601)
);

HB1xp67_ASAP7_75t_L g4602 ( 
.A(n_4167),
.Y(n_4602)
);

INVx2_ASAP7_75t_L g4603 ( 
.A(n_4145),
.Y(n_4603)
);

INVx1_ASAP7_75t_L g4604 ( 
.A(n_4420),
.Y(n_4604)
);

BUFx3_ASAP7_75t_L g4605 ( 
.A(n_4090),
.Y(n_4605)
);

INVx1_ASAP7_75t_L g4606 ( 
.A(n_4421),
.Y(n_4606)
);

OA21x2_ASAP7_75t_L g4607 ( 
.A1(n_4318),
.A2(n_3618),
.B(n_2273),
.Y(n_4607)
);

NAND2xp5_ASAP7_75t_L g4608 ( 
.A(n_4166),
.B(n_2772),
.Y(n_4608)
);

BUFx2_ASAP7_75t_L g4609 ( 
.A(n_4140),
.Y(n_4609)
);

BUFx8_ASAP7_75t_L g4610 ( 
.A(n_4301),
.Y(n_4610)
);

INVx1_ASAP7_75t_L g4611 ( 
.A(n_4271),
.Y(n_4611)
);

INVx1_ASAP7_75t_L g4612 ( 
.A(n_4272),
.Y(n_4612)
);

INVx2_ASAP7_75t_L g4613 ( 
.A(n_4146),
.Y(n_4613)
);

INVx1_ASAP7_75t_L g4614 ( 
.A(n_4289),
.Y(n_4614)
);

INVx3_ASAP7_75t_L g4615 ( 
.A(n_4070),
.Y(n_4615)
);

INVx2_ASAP7_75t_L g4616 ( 
.A(n_4151),
.Y(n_4616)
);

BUFx6f_ASAP7_75t_L g4617 ( 
.A(n_4456),
.Y(n_4617)
);

NAND2x1_ASAP7_75t_L g4618 ( 
.A(n_4157),
.B(n_2720),
.Y(n_4618)
);

INVx1_ASAP7_75t_L g4619 ( 
.A(n_4292),
.Y(n_4619)
);

BUFx3_ASAP7_75t_L g4620 ( 
.A(n_4102),
.Y(n_4620)
);

INVx2_ASAP7_75t_SL g4621 ( 
.A(n_4053),
.Y(n_4621)
);

BUFx8_ASAP7_75t_L g4622 ( 
.A(n_4058),
.Y(n_4622)
);

BUFx6f_ASAP7_75t_L g4623 ( 
.A(n_4459),
.Y(n_4623)
);

NOR2xp33_ASAP7_75t_L g4624 ( 
.A(n_4496),
.B(n_2669),
.Y(n_4624)
);

OAI22xp5_ASAP7_75t_SL g4625 ( 
.A1(n_4328),
.A2(n_3513),
.B1(n_3529),
.B2(n_3508),
.Y(n_4625)
);

AND2x2_ASAP7_75t_L g4626 ( 
.A(n_4307),
.B(n_2456),
.Y(n_4626)
);

NAND2x1p5_ASAP7_75t_L g4627 ( 
.A(n_4298),
.B(n_2814),
.Y(n_4627)
);

BUFx2_ASAP7_75t_L g4628 ( 
.A(n_4175),
.Y(n_4628)
);

INVx1_ASAP7_75t_L g4629 ( 
.A(n_4297),
.Y(n_4629)
);

AND2x2_ASAP7_75t_L g4630 ( 
.A(n_4370),
.B(n_2543),
.Y(n_4630)
);

BUFx2_ASAP7_75t_L g4631 ( 
.A(n_4130),
.Y(n_4631)
);

INVx1_ASAP7_75t_L g4632 ( 
.A(n_4299),
.Y(n_4632)
);

INVx5_ASAP7_75t_L g4633 ( 
.A(n_4408),
.Y(n_4633)
);

AND2x4_ASAP7_75t_L g4634 ( 
.A(n_4461),
.B(n_3342),
.Y(n_4634)
);

INVx1_ASAP7_75t_L g4635 ( 
.A(n_4305),
.Y(n_4635)
);

INVx1_ASAP7_75t_L g4636 ( 
.A(n_4306),
.Y(n_4636)
);

INVx1_ASAP7_75t_L g4637 ( 
.A(n_4313),
.Y(n_4637)
);

BUFx6f_ASAP7_75t_L g4638 ( 
.A(n_4464),
.Y(n_4638)
);

INVx3_ASAP7_75t_L g4639 ( 
.A(n_4072),
.Y(n_4639)
);

INVx1_ASAP7_75t_L g4640 ( 
.A(n_4317),
.Y(n_4640)
);

INVx3_ASAP7_75t_L g4641 ( 
.A(n_4075),
.Y(n_4641)
);

INVx1_ASAP7_75t_L g4642 ( 
.A(n_4319),
.Y(n_4642)
);

INVx1_ASAP7_75t_L g4643 ( 
.A(n_4323),
.Y(n_4643)
);

INVx3_ASAP7_75t_L g4644 ( 
.A(n_4079),
.Y(n_4644)
);

INVx1_ASAP7_75t_L g4645 ( 
.A(n_4331),
.Y(n_4645)
);

INVx1_ASAP7_75t_L g4646 ( 
.A(n_4334),
.Y(n_4646)
);

INVx1_ASAP7_75t_L g4647 ( 
.A(n_4349),
.Y(n_4647)
);

AND2x6_ASAP7_75t_L g4648 ( 
.A(n_4463),
.B(n_2837),
.Y(n_4648)
);

INVx2_ASAP7_75t_L g4649 ( 
.A(n_4152),
.Y(n_4649)
);

CKINVDCx5p33_ASAP7_75t_R g4650 ( 
.A(n_4081),
.Y(n_4650)
);

INVx1_ASAP7_75t_L g4651 ( 
.A(n_4351),
.Y(n_4651)
);

HB1xp67_ASAP7_75t_L g4652 ( 
.A(n_4172),
.Y(n_4652)
);

AND2x2_ASAP7_75t_L g4653 ( 
.A(n_4095),
.B(n_4302),
.Y(n_4653)
);

CKINVDCx5p33_ASAP7_75t_R g4654 ( 
.A(n_4114),
.Y(n_4654)
);

AND2x2_ASAP7_75t_L g4655 ( 
.A(n_4132),
.B(n_2543),
.Y(n_4655)
);

BUFx6f_ASAP7_75t_L g4656 ( 
.A(n_4465),
.Y(n_4656)
);

INVx1_ASAP7_75t_L g4657 ( 
.A(n_4355),
.Y(n_4657)
);

INVx2_ASAP7_75t_L g4658 ( 
.A(n_4203),
.Y(n_4658)
);

NOR2xp33_ASAP7_75t_L g4659 ( 
.A(n_4332),
.B(n_2674),
.Y(n_4659)
);

NOR2xp33_ASAP7_75t_L g4660 ( 
.A(n_4350),
.B(n_2675),
.Y(n_4660)
);

BUFx3_ASAP7_75t_L g4661 ( 
.A(n_4505),
.Y(n_4661)
);

INVx1_ASAP7_75t_L g4662 ( 
.A(n_4362),
.Y(n_4662)
);

INVx1_ASAP7_75t_L g4663 ( 
.A(n_4413),
.Y(n_4663)
);

BUFx8_ASAP7_75t_L g4664 ( 
.A(n_4078),
.Y(n_4664)
);

BUFx6f_ASAP7_75t_L g4665 ( 
.A(n_4478),
.Y(n_4665)
);

INVx2_ASAP7_75t_L g4666 ( 
.A(n_4224),
.Y(n_4666)
);

NAND2xp5_ASAP7_75t_L g4667 ( 
.A(n_4171),
.B(n_2814),
.Y(n_4667)
);

BUFx6f_ASAP7_75t_L g4668 ( 
.A(n_4485),
.Y(n_4668)
);

INVx4_ASAP7_75t_L g4669 ( 
.A(n_4223),
.Y(n_4669)
);

INVx1_ASAP7_75t_L g4670 ( 
.A(n_4416),
.Y(n_4670)
);

INVx1_ASAP7_75t_L g4671 ( 
.A(n_4424),
.Y(n_4671)
);

BUFx6f_ASAP7_75t_L g4672 ( 
.A(n_4507),
.Y(n_4672)
);

AND2x2_ASAP7_75t_L g4673 ( 
.A(n_4162),
.B(n_2672),
.Y(n_4673)
);

AND2x2_ASAP7_75t_SL g4674 ( 
.A(n_4144),
.B(n_2814),
.Y(n_4674)
);

INVx2_ASAP7_75t_L g4675 ( 
.A(n_4226),
.Y(n_4675)
);

INVx1_ASAP7_75t_L g4676 ( 
.A(n_4435),
.Y(n_4676)
);

INVx2_ASAP7_75t_L g4677 ( 
.A(n_4237),
.Y(n_4677)
);

INVx1_ASAP7_75t_L g4678 ( 
.A(n_4181),
.Y(n_4678)
);

INVx2_ASAP7_75t_L g4679 ( 
.A(n_4241),
.Y(n_4679)
);

INVx1_ASAP7_75t_L g4680 ( 
.A(n_4186),
.Y(n_4680)
);

INVx2_ASAP7_75t_L g4681 ( 
.A(n_4251),
.Y(n_4681)
);

NAND2xp5_ASAP7_75t_L g4682 ( 
.A(n_4192),
.B(n_2926),
.Y(n_4682)
);

BUFx6f_ASAP7_75t_L g4683 ( 
.A(n_4519),
.Y(n_4683)
);

INVx5_ASAP7_75t_L g4684 ( 
.A(n_4376),
.Y(n_4684)
);

NAND2xp33_ASAP7_75t_L g4685 ( 
.A(n_4523),
.B(n_2926),
.Y(n_4685)
);

INVx2_ASAP7_75t_L g4686 ( 
.A(n_4253),
.Y(n_4686)
);

INVx2_ASAP7_75t_L g4687 ( 
.A(n_4263),
.Y(n_4687)
);

AND2x2_ASAP7_75t_L g4688 ( 
.A(n_4174),
.B(n_2672),
.Y(n_4688)
);

NAND2xp5_ASAP7_75t_L g4689 ( 
.A(n_4198),
.B(n_2926),
.Y(n_4689)
);

INVx2_ASAP7_75t_L g4690 ( 
.A(n_4139),
.Y(n_4690)
);

INVx2_ASAP7_75t_L g4691 ( 
.A(n_4150),
.Y(n_4691)
);

AND2x4_ASAP7_75t_L g4692 ( 
.A(n_4509),
.B(n_2279),
.Y(n_4692)
);

INVx2_ASAP7_75t_L g4693 ( 
.A(n_4153),
.Y(n_4693)
);

INVxp67_ASAP7_75t_L g4694 ( 
.A(n_4283),
.Y(n_4694)
);

INVx1_ASAP7_75t_L g4695 ( 
.A(n_4210),
.Y(n_4695)
);

INVx1_ASAP7_75t_L g4696 ( 
.A(n_4221),
.Y(n_4696)
);

INVx1_ASAP7_75t_L g4697 ( 
.A(n_4231),
.Y(n_4697)
);

INVx1_ASAP7_75t_L g4698 ( 
.A(n_4245),
.Y(n_4698)
);

INVx1_ASAP7_75t_L g4699 ( 
.A(n_4248),
.Y(n_4699)
);

INVx6_ASAP7_75t_L g4700 ( 
.A(n_4074),
.Y(n_4700)
);

INVx1_ASAP7_75t_SL g4701 ( 
.A(n_4094),
.Y(n_4701)
);

INVx3_ASAP7_75t_L g4702 ( 
.A(n_4082),
.Y(n_4702)
);

INVx4_ASAP7_75t_L g4703 ( 
.A(n_4228),
.Y(n_4703)
);

INVx2_ASAP7_75t_L g4704 ( 
.A(n_4160),
.Y(n_4704)
);

BUFx2_ASAP7_75t_L g4705 ( 
.A(n_4516),
.Y(n_4705)
);

INVx1_ASAP7_75t_L g4706 ( 
.A(n_4249),
.Y(n_4706)
);

INVx1_ASAP7_75t_L g4707 ( 
.A(n_4254),
.Y(n_4707)
);

INVx1_ASAP7_75t_L g4708 ( 
.A(n_4257),
.Y(n_4708)
);

INVx2_ASAP7_75t_L g4709 ( 
.A(n_4184),
.Y(n_4709)
);

HB1xp67_ASAP7_75t_L g4710 ( 
.A(n_4159),
.Y(n_4710)
);

OAI22xp5_ASAP7_75t_L g4711 ( 
.A1(n_4115),
.A2(n_4525),
.B1(n_4176),
.B2(n_4475),
.Y(n_4711)
);

INVx1_ASAP7_75t_L g4712 ( 
.A(n_4260),
.Y(n_4712)
);

BUFx6f_ASAP7_75t_L g4713 ( 
.A(n_4524),
.Y(n_4713)
);

BUFx6f_ASAP7_75t_L g4714 ( 
.A(n_4536),
.Y(n_4714)
);

BUFx6f_ASAP7_75t_L g4715 ( 
.A(n_4537),
.Y(n_4715)
);

INVx1_ASAP7_75t_L g4716 ( 
.A(n_4262),
.Y(n_4716)
);

BUFx6f_ASAP7_75t_L g4717 ( 
.A(n_4089),
.Y(n_4717)
);

INVx1_ASAP7_75t_L g4718 ( 
.A(n_4265),
.Y(n_4718)
);

AND2x4_ASAP7_75t_L g4719 ( 
.A(n_4517),
.B(n_2296),
.Y(n_4719)
);

NAND2xp5_ASAP7_75t_SL g4720 ( 
.A(n_4137),
.B(n_3013),
.Y(n_4720)
);

INVx1_ASAP7_75t_L g4721 ( 
.A(n_4273),
.Y(n_4721)
);

CKINVDCx8_ASAP7_75t_R g4722 ( 
.A(n_4069),
.Y(n_4722)
);

BUFx6f_ASAP7_75t_L g4723 ( 
.A(n_4101),
.Y(n_4723)
);

AND2x4_ASAP7_75t_L g4724 ( 
.A(n_4529),
.B(n_2320),
.Y(n_4724)
);

INVx1_ASAP7_75t_L g4725 ( 
.A(n_4277),
.Y(n_4725)
);

INVx2_ASAP7_75t_L g4726 ( 
.A(n_4200),
.Y(n_4726)
);

NAND2xp33_ASAP7_75t_L g4727 ( 
.A(n_4528),
.B(n_3013),
.Y(n_4727)
);

INVx1_ASAP7_75t_L g4728 ( 
.A(n_4279),
.Y(n_4728)
);

OAI22xp5_ASAP7_75t_SL g4729 ( 
.A1(n_4116),
.A2(n_3555),
.B1(n_3375),
.B2(n_3379),
.Y(n_4729)
);

BUFx6f_ASAP7_75t_L g4730 ( 
.A(n_4533),
.Y(n_4730)
);

AND2x6_ASAP7_75t_L g4731 ( 
.A(n_4467),
.B(n_3258),
.Y(n_4731)
);

INVx1_ASAP7_75t_L g4732 ( 
.A(n_4287),
.Y(n_4732)
);

HB1xp67_ASAP7_75t_L g4733 ( 
.A(n_4542),
.Y(n_4733)
);

CKINVDCx8_ASAP7_75t_R g4734 ( 
.A(n_4084),
.Y(n_4734)
);

INVx3_ASAP7_75t_L g4735 ( 
.A(n_4213),
.Y(n_4735)
);

INVx2_ASAP7_75t_L g4736 ( 
.A(n_4216),
.Y(n_4736)
);

INVxp67_ASAP7_75t_L g4737 ( 
.A(n_4256),
.Y(n_4737)
);

AND2x2_ASAP7_75t_L g4738 ( 
.A(n_4188),
.B(n_2747),
.Y(n_4738)
);

INVx1_ASAP7_75t_L g4739 ( 
.A(n_4290),
.Y(n_4739)
);

INVx1_ASAP7_75t_L g4740 ( 
.A(n_4296),
.Y(n_4740)
);

OA21x2_ASAP7_75t_L g4741 ( 
.A1(n_4327),
.A2(n_2331),
.B(n_2328),
.Y(n_4741)
);

INVx1_ASAP7_75t_L g4742 ( 
.A(n_4312),
.Y(n_4742)
);

HB1xp67_ASAP7_75t_L g4743 ( 
.A(n_4182),
.Y(n_4743)
);

OR2x2_ASAP7_75t_L g4744 ( 
.A(n_4344),
.B(n_2761),
.Y(n_4744)
);

BUFx6f_ASAP7_75t_L g4745 ( 
.A(n_4426),
.Y(n_4745)
);

INVx1_ASAP7_75t_L g4746 ( 
.A(n_4163),
.Y(n_4746)
);

AND2x4_ASAP7_75t_L g4747 ( 
.A(n_4061),
.B(n_2335),
.Y(n_4747)
);

INVx1_ASAP7_75t_L g4748 ( 
.A(n_4168),
.Y(n_4748)
);

INVx3_ASAP7_75t_L g4749 ( 
.A(n_4219),
.Y(n_4749)
);

BUFx2_ASAP7_75t_L g4750 ( 
.A(n_4528),
.Y(n_4750)
);

INVx2_ASAP7_75t_L g4751 ( 
.A(n_4264),
.Y(n_4751)
);

OA21x2_ASAP7_75t_L g4752 ( 
.A1(n_4062),
.A2(n_2351),
.B(n_2340),
.Y(n_4752)
);

INVx1_ASAP7_75t_L g4753 ( 
.A(n_4170),
.Y(n_4753)
);

AND2x2_ASAP7_75t_L g4754 ( 
.A(n_4067),
.B(n_2747),
.Y(n_4754)
);

INVx1_ASAP7_75t_L g4755 ( 
.A(n_4178),
.Y(n_4755)
);

BUFx6f_ASAP7_75t_L g4756 ( 
.A(n_4540),
.Y(n_4756)
);

INVx2_ASAP7_75t_L g4757 ( 
.A(n_4155),
.Y(n_4757)
);

BUFx6f_ASAP7_75t_L g4758 ( 
.A(n_4259),
.Y(n_4758)
);

INVx3_ASAP7_75t_L g4759 ( 
.A(n_4118),
.Y(n_4759)
);

BUFx6f_ASAP7_75t_L g4760 ( 
.A(n_4314),
.Y(n_4760)
);

INVx2_ASAP7_75t_L g4761 ( 
.A(n_4440),
.Y(n_4761)
);

INVx1_ASAP7_75t_L g4762 ( 
.A(n_4185),
.Y(n_4762)
);

HB1xp67_ASAP7_75t_L g4763 ( 
.A(n_4204),
.Y(n_4763)
);

INVx4_ASAP7_75t_L g4764 ( 
.A(n_4452),
.Y(n_4764)
);

INVx2_ASAP7_75t_L g4765 ( 
.A(n_4441),
.Y(n_4765)
);

INVx1_ASAP7_75t_L g4766 ( 
.A(n_4194),
.Y(n_4766)
);

INVx4_ASAP7_75t_L g4767 ( 
.A(n_4080),
.Y(n_4767)
);

INVx2_ASAP7_75t_L g4768 ( 
.A(n_4450),
.Y(n_4768)
);

BUFx2_ASAP7_75t_L g4769 ( 
.A(n_4315),
.Y(n_4769)
);

NOR2xp33_ASAP7_75t_L g4770 ( 
.A(n_4492),
.B(n_2684),
.Y(n_4770)
);

AND2x2_ASAP7_75t_SL g4771 ( 
.A(n_4183),
.B(n_3013),
.Y(n_4771)
);

INVx1_ASAP7_75t_L g4772 ( 
.A(n_4266),
.Y(n_4772)
);

INVx1_ASAP7_75t_L g4773 ( 
.A(n_4270),
.Y(n_4773)
);

BUFx3_ASAP7_75t_L g4774 ( 
.A(n_4436),
.Y(n_4774)
);

INVxp33_ASAP7_75t_L g4775 ( 
.A(n_4173),
.Y(n_4775)
);

INVx3_ASAP7_75t_L g4776 ( 
.A(n_4489),
.Y(n_4776)
);

INVx1_ASAP7_75t_L g4777 ( 
.A(n_4278),
.Y(n_4777)
);

BUFx2_ASAP7_75t_L g4778 ( 
.A(n_4454),
.Y(n_4778)
);

BUFx6f_ASAP7_75t_L g4779 ( 
.A(n_4169),
.Y(n_4779)
);

INVx1_ASAP7_75t_L g4780 ( 
.A(n_4280),
.Y(n_4780)
);

NAND2xp5_ASAP7_75t_L g4781 ( 
.A(n_4051),
.B(n_3082),
.Y(n_4781)
);

INVx2_ASAP7_75t_L g4782 ( 
.A(n_4451),
.Y(n_4782)
);

AND2x2_ASAP7_75t_L g4783 ( 
.A(n_4110),
.B(n_2855),
.Y(n_4783)
);

BUFx6f_ASAP7_75t_L g4784 ( 
.A(n_4202),
.Y(n_4784)
);

INVx2_ASAP7_75t_L g4785 ( 
.A(n_4083),
.Y(n_4785)
);

INVx1_ASAP7_75t_L g4786 ( 
.A(n_4282),
.Y(n_4786)
);

INVx1_ASAP7_75t_L g4787 ( 
.A(n_4284),
.Y(n_4787)
);

INVx1_ASAP7_75t_L g4788 ( 
.A(n_4308),
.Y(n_4788)
);

INVx1_ASAP7_75t_L g4789 ( 
.A(n_4309),
.Y(n_4789)
);

CKINVDCx5p33_ASAP7_75t_R g4790 ( 
.A(n_4143),
.Y(n_4790)
);

NAND2xp5_ASAP7_75t_SL g4791 ( 
.A(n_4149),
.B(n_3082),
.Y(n_4791)
);

BUFx6f_ASAP7_75t_L g4792 ( 
.A(n_4208),
.Y(n_4792)
);

INVx2_ASAP7_75t_L g4793 ( 
.A(n_4117),
.Y(n_4793)
);

BUFx2_ASAP7_75t_L g4794 ( 
.A(n_4458),
.Y(n_4794)
);

BUFx8_ASAP7_75t_L g4795 ( 
.A(n_4474),
.Y(n_4795)
);

INVx2_ASAP7_75t_L g4796 ( 
.A(n_4120),
.Y(n_4796)
);

INVx1_ASAP7_75t_L g4797 ( 
.A(n_4214),
.Y(n_4797)
);

INVx1_ASAP7_75t_L g4798 ( 
.A(n_4232),
.Y(n_4798)
);

INVx1_ASAP7_75t_L g4799 ( 
.A(n_4233),
.Y(n_4799)
);

INVx1_ASAP7_75t_L g4800 ( 
.A(n_4243),
.Y(n_4800)
);

INVx1_ASAP7_75t_L g4801 ( 
.A(n_4361),
.Y(n_4801)
);

INVx2_ASAP7_75t_L g4802 ( 
.A(n_4438),
.Y(n_4802)
);

AND2x2_ASAP7_75t_L g4803 ( 
.A(n_4054),
.B(n_2855),
.Y(n_4803)
);

INVx1_ASAP7_75t_L g4804 ( 
.A(n_4371),
.Y(n_4804)
);

AND2x2_ASAP7_75t_L g4805 ( 
.A(n_4220),
.B(n_2896),
.Y(n_4805)
);

AND2x6_ASAP7_75t_L g4806 ( 
.A(n_4343),
.B(n_3499),
.Y(n_4806)
);

INVx3_ASAP7_75t_L g4807 ( 
.A(n_4490),
.Y(n_4807)
);

INVx1_ASAP7_75t_L g4808 ( 
.A(n_4373),
.Y(n_4808)
);

NAND2xp5_ASAP7_75t_SL g4809 ( 
.A(n_4179),
.B(n_3082),
.Y(n_4809)
);

INVx3_ASAP7_75t_L g4810 ( 
.A(n_4518),
.Y(n_4810)
);

INVx1_ASAP7_75t_L g4811 ( 
.A(n_4377),
.Y(n_4811)
);

INVx1_ASAP7_75t_L g4812 ( 
.A(n_4381),
.Y(n_4812)
);

NAND2xp5_ASAP7_75t_L g4813 ( 
.A(n_4057),
.B(n_3264),
.Y(n_4813)
);

BUFx6f_ASAP7_75t_L g4814 ( 
.A(n_4443),
.Y(n_4814)
);

AND2x6_ASAP7_75t_L g4815 ( 
.A(n_4345),
.B(n_3521),
.Y(n_4815)
);

INVx1_ASAP7_75t_L g4816 ( 
.A(n_4419),
.Y(n_4816)
);

INVx1_ASAP7_75t_L g4817 ( 
.A(n_4430),
.Y(n_4817)
);

INVx1_ASAP7_75t_L g4818 ( 
.A(n_4063),
.Y(n_4818)
);

AND2x4_ASAP7_75t_L g4819 ( 
.A(n_4227),
.B(n_2366),
.Y(n_4819)
);

INVx4_ASAP7_75t_L g4820 ( 
.A(n_4104),
.Y(n_4820)
);

INVx1_ASAP7_75t_L g4821 ( 
.A(n_4065),
.Y(n_4821)
);

INVx2_ASAP7_75t_L g4822 ( 
.A(n_4444),
.Y(n_4822)
);

AND2x2_ASAP7_75t_L g4823 ( 
.A(n_4247),
.B(n_2896),
.Y(n_4823)
);

NOR2xp33_ASAP7_75t_L g4824 ( 
.A(n_4261),
.B(n_4472),
.Y(n_4824)
);

INVx1_ASAP7_75t_L g4825 ( 
.A(n_4087),
.Y(n_4825)
);

INVx1_ASAP7_75t_L g4826 ( 
.A(n_4088),
.Y(n_4826)
);

INVx1_ASAP7_75t_L g4827 ( 
.A(n_4092),
.Y(n_4827)
);

INVx2_ASAP7_75t_L g4828 ( 
.A(n_4447),
.Y(n_4828)
);

BUFx6f_ASAP7_75t_L g4829 ( 
.A(n_4448),
.Y(n_4829)
);

INVx1_ASAP7_75t_L g4830 ( 
.A(n_4098),
.Y(n_4830)
);

INVx4_ASAP7_75t_L g4831 ( 
.A(n_4106),
.Y(n_4831)
);

INVxp33_ASAP7_75t_SL g4832 ( 
.A(n_4286),
.Y(n_4832)
);

BUFx6f_ASAP7_75t_L g4833 ( 
.A(n_4165),
.Y(n_4833)
);

AND2x6_ASAP7_75t_L g4834 ( 
.A(n_4462),
.B(n_2300),
.Y(n_4834)
);

INVx3_ASAP7_75t_L g4835 ( 
.A(n_4190),
.Y(n_4835)
);

INVx1_ASAP7_75t_L g4836 ( 
.A(n_4100),
.Y(n_4836)
);

INVxp67_ASAP7_75t_L g4837 ( 
.A(n_4392),
.Y(n_4837)
);

INVx1_ASAP7_75t_L g4838 ( 
.A(n_4103),
.Y(n_4838)
);

BUFx6f_ASAP7_75t_L g4839 ( 
.A(n_4390),
.Y(n_4839)
);

INVx2_ASAP7_75t_L g4840 ( 
.A(n_4199),
.Y(n_4840)
);

AND2x2_ASAP7_75t_L g4841 ( 
.A(n_4295),
.B(n_2932),
.Y(n_4841)
);

INVx2_ASAP7_75t_L g4842 ( 
.A(n_4320),
.Y(n_4842)
);

INVx1_ASAP7_75t_L g4843 ( 
.A(n_4105),
.Y(n_4843)
);

OAI22xp5_ASAP7_75t_SL g4844 ( 
.A1(n_4281),
.A2(n_2696),
.B1(n_2697),
.B2(n_2693),
.Y(n_4844)
);

INVx1_ASAP7_75t_L g4845 ( 
.A(n_4109),
.Y(n_4845)
);

INVx3_ASAP7_75t_L g4846 ( 
.A(n_4195),
.Y(n_4846)
);

INVx1_ASAP7_75t_L g4847 ( 
.A(n_4111),
.Y(n_4847)
);

INVx2_ASAP7_75t_L g4848 ( 
.A(n_4325),
.Y(n_4848)
);

INVx2_ASAP7_75t_L g4849 ( 
.A(n_4326),
.Y(n_4849)
);

INVx1_ASAP7_75t_L g4850 ( 
.A(n_4119),
.Y(n_4850)
);

INVx2_ASAP7_75t_L g4851 ( 
.A(n_4336),
.Y(n_4851)
);

INVx1_ASAP7_75t_L g4852 ( 
.A(n_4128),
.Y(n_4852)
);

INVx1_ASAP7_75t_L g4853 ( 
.A(n_4136),
.Y(n_4853)
);

AND2x2_ASAP7_75t_L g4854 ( 
.A(n_4138),
.B(n_2932),
.Y(n_4854)
);

INVx1_ASAP7_75t_L g4855 ( 
.A(n_4147),
.Y(n_4855)
);

NOR2xp33_ASAP7_75t_SL g4856 ( 
.A(n_4187),
.B(n_2334),
.Y(n_4856)
);

BUFx8_ASAP7_75t_L g4857 ( 
.A(n_4476),
.Y(n_4857)
);

BUFx6f_ASAP7_75t_L g4858 ( 
.A(n_4415),
.Y(n_4858)
);

NOR2xp33_ASAP7_75t_L g4859 ( 
.A(n_4483),
.B(n_2718),
.Y(n_4859)
);

INVx1_ASAP7_75t_L g4860 ( 
.A(n_4385),
.Y(n_4860)
);

INVx2_ASAP7_75t_L g4861 ( 
.A(n_4366),
.Y(n_4861)
);

INVx2_ASAP7_75t_L g4862 ( 
.A(n_4367),
.Y(n_4862)
);

INVx1_ASAP7_75t_L g4863 ( 
.A(n_4389),
.Y(n_4863)
);

AND2x4_ASAP7_75t_L g4864 ( 
.A(n_4085),
.B(n_2371),
.Y(n_4864)
);

AND3x2_ASAP7_75t_L g4865 ( 
.A(n_4142),
.B(n_2385),
.C(n_2372),
.Y(n_4865)
);

INVx1_ASAP7_75t_L g4866 ( 
.A(n_4409),
.Y(n_4866)
);

NAND2xp5_ASAP7_75t_L g4867 ( 
.A(n_4484),
.B(n_3264),
.Y(n_4867)
);

INVx2_ASAP7_75t_L g4868 ( 
.A(n_4423),
.Y(n_4868)
);

AND2x4_ASAP7_75t_L g4869 ( 
.A(n_4086),
.B(n_2398),
.Y(n_4869)
);

NAND2xp5_ASAP7_75t_L g4870 ( 
.A(n_4510),
.B(n_3264),
.Y(n_4870)
);

INVx4_ASAP7_75t_L g4871 ( 
.A(n_4112),
.Y(n_4871)
);

INVx2_ASAP7_75t_L g4872 ( 
.A(n_4425),
.Y(n_4872)
);

INVx1_ASAP7_75t_L g4873 ( 
.A(n_4432),
.Y(n_4873)
);

INVx2_ASAP7_75t_L g4874 ( 
.A(n_4433),
.Y(n_4874)
);

NAND2xp5_ASAP7_75t_SL g4875 ( 
.A(n_4364),
.B(n_3301),
.Y(n_4875)
);

INVx1_ASAP7_75t_L g4876 ( 
.A(n_4511),
.Y(n_4876)
);

INVx1_ASAP7_75t_L g4877 ( 
.A(n_4520),
.Y(n_4877)
);

INVx2_ASAP7_75t_L g4878 ( 
.A(n_4442),
.Y(n_4878)
);

BUFx6f_ASAP7_75t_L g4879 ( 
.A(n_4417),
.Y(n_4879)
);

AND2x2_ASAP7_75t_L g4880 ( 
.A(n_4391),
.B(n_3000),
.Y(n_4880)
);

OA21x2_ASAP7_75t_L g4881 ( 
.A1(n_4310),
.A2(n_2408),
.B(n_2406),
.Y(n_4881)
);

INVx2_ASAP7_75t_L g4882 ( 
.A(n_4229),
.Y(n_4882)
);

INVx1_ASAP7_75t_L g4883 ( 
.A(n_4541),
.Y(n_4883)
);

INVx2_ASAP7_75t_L g4884 ( 
.A(n_4244),
.Y(n_4884)
);

AND2x4_ASAP7_75t_L g4885 ( 
.A(n_4096),
.B(n_2410),
.Y(n_4885)
);

INVx1_ASAP7_75t_L g4886 ( 
.A(n_4049),
.Y(n_4886)
);

AND2x4_ASAP7_75t_L g4887 ( 
.A(n_4121),
.B(n_2415),
.Y(n_4887)
);

INVx2_ASAP7_75t_L g4888 ( 
.A(n_4396),
.Y(n_4888)
);

AOI22xp5_ASAP7_75t_L g4889 ( 
.A1(n_4407),
.A2(n_2407),
.B1(n_2488),
.B2(n_2400),
.Y(n_4889)
);

AND2x2_ASAP7_75t_L g4890 ( 
.A(n_4412),
.B(n_3000),
.Y(n_4890)
);

INVx1_ASAP7_75t_L g4891 ( 
.A(n_4060),
.Y(n_4891)
);

BUFx2_ASAP7_75t_L g4892 ( 
.A(n_4522),
.Y(n_4892)
);

INVx4_ASAP7_75t_L g4893 ( 
.A(n_4134),
.Y(n_4893)
);

BUFx6f_ASAP7_75t_L g4894 ( 
.A(n_4428),
.Y(n_4894)
);

AOI22xp5_ASAP7_75t_L g4895 ( 
.A1(n_4471),
.A2(n_2602),
.B1(n_2662),
.B2(n_2520),
.Y(n_4895)
);

AND3x2_ASAP7_75t_L g4896 ( 
.A(n_4164),
.B(n_2424),
.C(n_2417),
.Y(n_4896)
);

AND2x6_ASAP7_75t_L g4897 ( 
.A(n_4477),
.B(n_2745),
.Y(n_4897)
);

NOR2xp33_ASAP7_75t_L g4898 ( 
.A(n_4339),
.B(n_2722),
.Y(n_4898)
);

INVx1_ASAP7_75t_L g4899 ( 
.A(n_4091),
.Y(n_4899)
);

INVx1_ASAP7_75t_L g4900 ( 
.A(n_4097),
.Y(n_4900)
);

INVx1_ASAP7_75t_L g4901 ( 
.A(n_4455),
.Y(n_4901)
);

INVx1_ASAP7_75t_L g4902 ( 
.A(n_4488),
.Y(n_4902)
);

INVx1_ASAP7_75t_L g4903 ( 
.A(n_4526),
.Y(n_4903)
);

AND2x2_ASAP7_75t_L g4904 ( 
.A(n_4487),
.B(n_3067),
.Y(n_4904)
);

INVx1_ASAP7_75t_L g4905 ( 
.A(n_4304),
.Y(n_4905)
);

NAND2xp5_ASAP7_75t_SL g4906 ( 
.A(n_4052),
.B(n_3301),
.Y(n_4906)
);

INVx2_ASAP7_75t_L g4907 ( 
.A(n_4321),
.Y(n_4907)
);

INVx2_ASAP7_75t_L g4908 ( 
.A(n_4352),
.Y(n_4908)
);

INVx3_ASAP7_75t_L g4909 ( 
.A(n_4353),
.Y(n_4909)
);

AND2x2_ASAP7_75t_L g4910 ( 
.A(n_4493),
.B(n_3067),
.Y(n_4910)
);

INVx1_ASAP7_75t_L g4911 ( 
.A(n_4358),
.Y(n_4911)
);

INVx2_ASAP7_75t_L g4912 ( 
.A(n_4365),
.Y(n_4912)
);

INVx2_ASAP7_75t_SL g4913 ( 
.A(n_4212),
.Y(n_4913)
);

INVx3_ASAP7_75t_L g4914 ( 
.A(n_4368),
.Y(n_4914)
);

CKINVDCx5p33_ASAP7_75t_R g4915 ( 
.A(n_4288),
.Y(n_4915)
);

INVx2_ASAP7_75t_L g4916 ( 
.A(n_4410),
.Y(n_4916)
);

NAND2xp33_ASAP7_75t_L g4917 ( 
.A(n_4107),
.B(n_3301),
.Y(n_4917)
);

INVx3_ASAP7_75t_L g4918 ( 
.A(n_4429),
.Y(n_4918)
);

INVx2_ASAP7_75t_L g4919 ( 
.A(n_4329),
.Y(n_4919)
);

BUFx8_ASAP7_75t_L g4920 ( 
.A(n_4189),
.Y(n_4920)
);

BUFx6f_ASAP7_75t_L g4921 ( 
.A(n_4341),
.Y(n_4921)
);

INVx1_ASAP7_75t_L g4922 ( 
.A(n_4311),
.Y(n_4922)
);

BUFx8_ASAP7_75t_L g4923 ( 
.A(n_4508),
.Y(n_4923)
);

XOR2xp5_ASAP7_75t_L g4924 ( 
.A(n_4494),
.B(n_2264),
.Y(n_4924)
);

INVx2_ASAP7_75t_L g4925 ( 
.A(n_4378),
.Y(n_4925)
);

CKINVDCx5p33_ASAP7_75t_R g4926 ( 
.A(n_4293),
.Y(n_4926)
);

INVx2_ASAP7_75t_L g4927 ( 
.A(n_4382),
.Y(n_4927)
);

INVx1_ASAP7_75t_L g4928 ( 
.A(n_4360),
.Y(n_4928)
);

INVx1_ASAP7_75t_L g4929 ( 
.A(n_4386),
.Y(n_4929)
);

INVx1_ASAP7_75t_L g4930 ( 
.A(n_4387),
.Y(n_4930)
);

INVx2_ASAP7_75t_L g4931 ( 
.A(n_4400),
.Y(n_4931)
);

INVx2_ASAP7_75t_L g4932 ( 
.A(n_4453),
.Y(n_4932)
);

INVx2_ASAP7_75t_L g4933 ( 
.A(n_4258),
.Y(n_4933)
);

INVx1_ASAP7_75t_L g4934 ( 
.A(n_4414),
.Y(n_4934)
);

AND2x4_ASAP7_75t_L g4935 ( 
.A(n_4123),
.B(n_2426),
.Y(n_4935)
);

INVx3_ASAP7_75t_L g4936 ( 
.A(n_4446),
.Y(n_4936)
);

INVx1_ASAP7_75t_L g4937 ( 
.A(n_4427),
.Y(n_4937)
);

AND2x6_ASAP7_75t_L g4938 ( 
.A(n_4500),
.B(n_4437),
.Y(n_4938)
);

INVx1_ASAP7_75t_L g4939 ( 
.A(n_4347),
.Y(n_4939)
);

NAND2xp5_ASAP7_75t_L g4940 ( 
.A(n_4369),
.B(n_3540),
.Y(n_4940)
);

NAND2xp5_ASAP7_75t_L g4941 ( 
.A(n_4397),
.B(n_4161),
.Y(n_4941)
);

INVx1_ASAP7_75t_L g4942 ( 
.A(n_4374),
.Y(n_4942)
);

NOR2xp33_ASAP7_75t_L g4943 ( 
.A(n_4135),
.B(n_2726),
.Y(n_4943)
);

INVx2_ASAP7_75t_L g4944 ( 
.A(n_4439),
.Y(n_4944)
);

INVx2_ASAP7_75t_L g4945 ( 
.A(n_4395),
.Y(n_4945)
);

INVx2_ASAP7_75t_L g4946 ( 
.A(n_4402),
.Y(n_4946)
);

INVx1_ASAP7_75t_L g4947 ( 
.A(n_4418),
.Y(n_4947)
);

INVx2_ASAP7_75t_L g4948 ( 
.A(n_4449),
.Y(n_4948)
);

INVx1_ASAP7_75t_L g4949 ( 
.A(n_4393),
.Y(n_4949)
);

BUFx6f_ASAP7_75t_L g4950 ( 
.A(n_4180),
.Y(n_4950)
);

HB1xp67_ASAP7_75t_L g4951 ( 
.A(n_4218),
.Y(n_4951)
);

INVx1_ASAP7_75t_L g4952 ( 
.A(n_4403),
.Y(n_4952)
);

INVx1_ASAP7_75t_SL g4953 ( 
.A(n_4530),
.Y(n_4953)
);

INVx1_ASAP7_75t_L g4954 ( 
.A(n_4383),
.Y(n_4954)
);

BUFx6f_ASAP7_75t_L g4955 ( 
.A(n_4222),
.Y(n_4955)
);

INVx1_ASAP7_75t_L g4956 ( 
.A(n_4398),
.Y(n_4956)
);

NAND2xp5_ASAP7_75t_L g4957 ( 
.A(n_4359),
.B(n_4445),
.Y(n_4957)
);

AND2x2_ASAP7_75t_L g4958 ( 
.A(n_4201),
.B(n_3072),
.Y(n_4958)
);

NAND2xp5_ASAP7_75t_L g4959 ( 
.A(n_4193),
.B(n_3540),
.Y(n_4959)
);

NAND2xp5_ASAP7_75t_L g4960 ( 
.A(n_4205),
.B(n_3540),
.Y(n_4960)
);

INVx2_ASAP7_75t_L g4961 ( 
.A(n_4401),
.Y(n_4961)
);

NAND2xp5_ASAP7_75t_L g4962 ( 
.A(n_4392),
.B(n_3569),
.Y(n_4962)
);

BUFx6f_ASAP7_75t_L g4963 ( 
.A(n_4406),
.Y(n_4963)
);

AND2x2_ASAP7_75t_L g4964 ( 
.A(n_4235),
.B(n_4269),
.Y(n_4964)
);

INVx2_ASAP7_75t_L g4965 ( 
.A(n_4411),
.Y(n_4965)
);

INVx1_ASAP7_75t_L g4966 ( 
.A(n_4431),
.Y(n_4966)
);

BUFx2_ASAP7_75t_L g4967 ( 
.A(n_4124),
.Y(n_4967)
);

INVx1_ASAP7_75t_L g4968 ( 
.A(n_4274),
.Y(n_4968)
);

BUFx6f_ASAP7_75t_L g4969 ( 
.A(n_4113),
.Y(n_4969)
);

OA21x2_ASAP7_75t_L g4970 ( 
.A1(n_4239),
.A2(n_2433),
.B(n_2431),
.Y(n_4970)
);

CKINVDCx5p33_ASAP7_75t_R g4971 ( 
.A(n_4303),
.Y(n_4971)
);

INVx1_ASAP7_75t_L g4972 ( 
.A(n_4177),
.Y(n_4972)
);

AND2x2_ASAP7_75t_L g4973 ( 
.A(n_4268),
.B(n_3072),
.Y(n_4973)
);

INVx1_ASAP7_75t_L g4974 ( 
.A(n_4191),
.Y(n_4974)
);

BUFx6f_ASAP7_75t_L g4975 ( 
.A(n_4156),
.Y(n_4975)
);

INVx2_ASAP7_75t_L g4976 ( 
.A(n_4071),
.Y(n_4976)
);

BUFx6f_ASAP7_75t_L g4977 ( 
.A(n_4197),
.Y(n_4977)
);

CKINVDCx5p33_ASAP7_75t_R g4978 ( 
.A(n_4047),
.Y(n_4978)
);

AND2x4_ASAP7_75t_L g4979 ( 
.A(n_4196),
.B(n_2441),
.Y(n_4979)
);

BUFx2_ASAP7_75t_L g4980 ( 
.A(n_4133),
.Y(n_4980)
);

INVx1_ASAP7_75t_L g4981 ( 
.A(n_4076),
.Y(n_4981)
);

INVx2_ASAP7_75t_L g4982 ( 
.A(n_4466),
.Y(n_4982)
);

BUFx2_ASAP7_75t_L g4983 ( 
.A(n_4330),
.Y(n_4983)
);

INVx1_ASAP7_75t_L g4984 ( 
.A(n_4468),
.Y(n_4984)
);

INVx1_ASAP7_75t_L g4985 ( 
.A(n_4479),
.Y(n_4985)
);

INVx1_ASAP7_75t_L g4986 ( 
.A(n_4515),
.Y(n_4986)
);

INVx1_ASAP7_75t_L g4987 ( 
.A(n_4535),
.Y(n_4987)
);

INVx2_ASAP7_75t_L g4988 ( 
.A(n_4217),
.Y(n_4988)
);

INVx1_ASAP7_75t_L g4989 ( 
.A(n_4294),
.Y(n_4989)
);

INVx2_ASAP7_75t_L g4990 ( 
.A(n_4225),
.Y(n_4990)
);

INVx1_ASAP7_75t_L g4991 ( 
.A(n_4300),
.Y(n_4991)
);

INVx1_ASAP7_75t_L g4992 ( 
.A(n_4501),
.Y(n_4992)
);

INVx1_ASAP7_75t_L g4993 ( 
.A(n_4234),
.Y(n_4993)
);

INVx2_ASAP7_75t_L g4994 ( 
.A(n_4240),
.Y(n_4994)
);

INVx1_ASAP7_75t_L g4995 ( 
.A(n_4356),
.Y(n_4995)
);

HB1xp67_ASAP7_75t_L g4996 ( 
.A(n_4207),
.Y(n_4996)
);

INVx2_ASAP7_75t_L g4997 ( 
.A(n_4497),
.Y(n_4997)
);

INVx2_ASAP7_75t_L g4998 ( 
.A(n_4498),
.Y(n_4998)
);

BUFx12f_ASAP7_75t_L g4999 ( 
.A(n_4499),
.Y(n_4999)
);

INVx2_ASAP7_75t_L g5000 ( 
.A(n_4538),
.Y(n_5000)
);

AND3x2_ASAP7_75t_L g5001 ( 
.A(n_4388),
.B(n_2459),
.C(n_2450),
.Y(n_5001)
);

INVx2_ASAP7_75t_L g5002 ( 
.A(n_4539),
.Y(n_5002)
);

INVx2_ASAP7_75t_L g5003 ( 
.A(n_4340),
.Y(n_5003)
);

INVx2_ASAP7_75t_L g5004 ( 
.A(n_4346),
.Y(n_5004)
);

AND2x2_ASAP7_75t_L g5005 ( 
.A(n_4158),
.B(n_3108),
.Y(n_5005)
);

BUFx3_ASAP7_75t_L g5006 ( 
.A(n_4531),
.Y(n_5006)
);

OAI21x1_ASAP7_75t_L g5007 ( 
.A1(n_4215),
.A2(n_2468),
.B(n_2461),
.Y(n_5007)
);

BUFx6f_ASAP7_75t_L g5008 ( 
.A(n_4046),
.Y(n_5008)
);

INVx2_ASAP7_75t_L g5009 ( 
.A(n_4434),
.Y(n_5009)
);

AND2x4_ASAP7_75t_L g5010 ( 
.A(n_4242),
.B(n_2477),
.Y(n_5010)
);

INVx2_ASAP7_75t_L g5011 ( 
.A(n_4473),
.Y(n_5011)
);

INVx1_ASAP7_75t_L g5012 ( 
.A(n_4338),
.Y(n_5012)
);

INVx1_ASAP7_75t_L g5013 ( 
.A(n_4093),
.Y(n_5013)
);

AND2x2_ASAP7_75t_L g5014 ( 
.A(n_4099),
.B(n_3108),
.Y(n_5014)
);

NAND2xp5_ASAP7_75t_L g5015 ( 
.A(n_4050),
.B(n_3569),
.Y(n_5015)
);

INVx1_ASAP7_75t_L g5016 ( 
.A(n_4460),
.Y(n_5016)
);

BUFx3_ASAP7_75t_L g5017 ( 
.A(n_4457),
.Y(n_5017)
);

NAND2xp5_ASAP7_75t_L g5018 ( 
.A(n_4491),
.B(n_3569),
.Y(n_5018)
);

OAI21x1_ASAP7_75t_L g5019 ( 
.A1(n_4504),
.A2(n_2492),
.B(n_2489),
.Y(n_5019)
);

INVx3_ASAP7_75t_L g5020 ( 
.A(n_4512),
.Y(n_5020)
);

INVx2_ASAP7_75t_L g5021 ( 
.A(n_4506),
.Y(n_5021)
);

INVx1_ASAP7_75t_L g5022 ( 
.A(n_4108),
.Y(n_5022)
);

INVx1_ASAP7_75t_L g5023 ( 
.A(n_4141),
.Y(n_5023)
);

INVx1_ASAP7_75t_L g5024 ( 
.A(n_4206),
.Y(n_5024)
);

BUFx6f_ASAP7_75t_L g5025 ( 
.A(n_4513),
.Y(n_5025)
);

AND2x4_ASAP7_75t_L g5026 ( 
.A(n_4131),
.B(n_2496),
.Y(n_5026)
);

INVx1_ASAP7_75t_L g5027 ( 
.A(n_4246),
.Y(n_5027)
);

INVx2_ASAP7_75t_L g5028 ( 
.A(n_4514),
.Y(n_5028)
);

OR2x6_ASAP7_75t_L g5029 ( 
.A(n_4534),
.B(n_3626),
.Y(n_5029)
);

INVx1_ASAP7_75t_L g5030 ( 
.A(n_4348),
.Y(n_5030)
);

INVx1_ASAP7_75t_L g5031 ( 
.A(n_4348),
.Y(n_5031)
);

NAND2xp5_ASAP7_75t_L g5032 ( 
.A(n_4372),
.B(n_3626),
.Y(n_5032)
);

HB1xp67_ASAP7_75t_L g5033 ( 
.A(n_4354),
.Y(n_5033)
);

INVx1_ASAP7_75t_L g5034 ( 
.A(n_4348),
.Y(n_5034)
);

INVx1_ASAP7_75t_L g5035 ( 
.A(n_4348),
.Y(n_5035)
);

INVx2_ASAP7_75t_L g5036 ( 
.A(n_4048),
.Y(n_5036)
);

INVx2_ASAP7_75t_L g5037 ( 
.A(n_4048),
.Y(n_5037)
);

OAI21x1_ASAP7_75t_L g5038 ( 
.A1(n_4318),
.A2(n_2513),
.B(n_2511),
.Y(n_5038)
);

INVx1_ASAP7_75t_L g5039 ( 
.A(n_4348),
.Y(n_5039)
);

BUFx6f_ASAP7_75t_L g5040 ( 
.A(n_4064),
.Y(n_5040)
);

NOR2xp33_ASAP7_75t_L g5041 ( 
.A(n_4275),
.B(n_2727),
.Y(n_5041)
);

INVx1_ASAP7_75t_L g5042 ( 
.A(n_4348),
.Y(n_5042)
);

INVx1_ASAP7_75t_L g5043 ( 
.A(n_4348),
.Y(n_5043)
);

NAND2xp33_ASAP7_75t_L g5044 ( 
.A(n_4523),
.B(n_2728),
.Y(n_5044)
);

INVx1_ASAP7_75t_L g5045 ( 
.A(n_4348),
.Y(n_5045)
);

INVx2_ASAP7_75t_L g5046 ( 
.A(n_4048),
.Y(n_5046)
);

INVx2_ASAP7_75t_L g5047 ( 
.A(n_4048),
.Y(n_5047)
);

AND2x6_ASAP7_75t_L g5048 ( 
.A(n_4252),
.B(n_2919),
.Y(n_5048)
);

AND2x2_ASAP7_75t_L g5049 ( 
.A(n_4354),
.B(n_3113),
.Y(n_5049)
);

BUFx6f_ASAP7_75t_L g5050 ( 
.A(n_4064),
.Y(n_5050)
);

AND2x4_ASAP7_75t_L g5051 ( 
.A(n_4354),
.B(n_2523),
.Y(n_5051)
);

AND2x4_ASAP7_75t_L g5052 ( 
.A(n_4354),
.B(n_2532),
.Y(n_5052)
);

INVx3_ASAP7_75t_L g5053 ( 
.A(n_4126),
.Y(n_5053)
);

INVx1_ASAP7_75t_L g5054 ( 
.A(n_4348),
.Y(n_5054)
);

NOR2xp33_ASAP7_75t_L g5055 ( 
.A(n_4275),
.B(n_2729),
.Y(n_5055)
);

INVx2_ASAP7_75t_L g5056 ( 
.A(n_4048),
.Y(n_5056)
);

INVx1_ASAP7_75t_L g5057 ( 
.A(n_4348),
.Y(n_5057)
);

NAND2xp5_ASAP7_75t_SL g5058 ( 
.A(n_4354),
.B(n_2731),
.Y(n_5058)
);

AND3x2_ASAP7_75t_L g5059 ( 
.A(n_4286),
.B(n_2547),
.C(n_2539),
.Y(n_5059)
);

INVx1_ASAP7_75t_L g5060 ( 
.A(n_4348),
.Y(n_5060)
);

INVx2_ASAP7_75t_L g5061 ( 
.A(n_4048),
.Y(n_5061)
);

INVx2_ASAP7_75t_L g5062 ( 
.A(n_4048),
.Y(n_5062)
);

INVx1_ASAP7_75t_L g5063 ( 
.A(n_4348),
.Y(n_5063)
);

INVx1_ASAP7_75t_L g5064 ( 
.A(n_4348),
.Y(n_5064)
);

OR2x6_ASAP7_75t_L g5065 ( 
.A(n_4333),
.B(n_2555),
.Y(n_5065)
);

INVx1_ASAP7_75t_L g5066 ( 
.A(n_4348),
.Y(n_5066)
);

BUFx6f_ASAP7_75t_L g5067 ( 
.A(n_4064),
.Y(n_5067)
);

INVx2_ASAP7_75t_L g5068 ( 
.A(n_4048),
.Y(n_5068)
);

INVx1_ASAP7_75t_L g5069 ( 
.A(n_4348),
.Y(n_5069)
);

BUFx3_ASAP7_75t_L g5070 ( 
.A(n_4333),
.Y(n_5070)
);

INVx1_ASAP7_75t_L g5071 ( 
.A(n_4348),
.Y(n_5071)
);

INVxp67_ASAP7_75t_L g5072 ( 
.A(n_4354),
.Y(n_5072)
);

INVx3_ASAP7_75t_L g5073 ( 
.A(n_4126),
.Y(n_5073)
);

BUFx6f_ASAP7_75t_L g5074 ( 
.A(n_4064),
.Y(n_5074)
);

INVx2_ASAP7_75t_L g5075 ( 
.A(n_4048),
.Y(n_5075)
);

INVx1_ASAP7_75t_L g5076 ( 
.A(n_4348),
.Y(n_5076)
);

INVx1_ASAP7_75t_L g5077 ( 
.A(n_4348),
.Y(n_5077)
);

CKINVDCx20_ASAP7_75t_R g5078 ( 
.A(n_4094),
.Y(n_5078)
);

AND2x2_ASAP7_75t_L g5079 ( 
.A(n_4354),
.B(n_3113),
.Y(n_5079)
);

INVx1_ASAP7_75t_L g5080 ( 
.A(n_4348),
.Y(n_5080)
);

INVx1_ASAP7_75t_L g5081 ( 
.A(n_4348),
.Y(n_5081)
);

OAI21x1_ASAP7_75t_L g5082 ( 
.A1(n_4318),
.A2(n_2573),
.B(n_2571),
.Y(n_5082)
);

HB1xp67_ASAP7_75t_L g5083 ( 
.A(n_4354),
.Y(n_5083)
);

INVx3_ASAP7_75t_L g5084 ( 
.A(n_4126),
.Y(n_5084)
);

INVx1_ASAP7_75t_L g5085 ( 
.A(n_4348),
.Y(n_5085)
);

INVx1_ASAP7_75t_L g5086 ( 
.A(n_4348),
.Y(n_5086)
);

INVx1_ASAP7_75t_L g5087 ( 
.A(n_4348),
.Y(n_5087)
);

INVx1_ASAP7_75t_L g5088 ( 
.A(n_4348),
.Y(n_5088)
);

INVx1_ASAP7_75t_L g5089 ( 
.A(n_4348),
.Y(n_5089)
);

INVxp67_ASAP7_75t_L g5090 ( 
.A(n_4354),
.Y(n_5090)
);

AND2x4_ASAP7_75t_L g5091 ( 
.A(n_4354),
.B(n_2584),
.Y(n_5091)
);

INVx1_ASAP7_75t_L g5092 ( 
.A(n_4348),
.Y(n_5092)
);

INVx1_ASAP7_75t_L g5093 ( 
.A(n_4348),
.Y(n_5093)
);

NAND2xp5_ASAP7_75t_L g5094 ( 
.A(n_4372),
.B(n_2586),
.Y(n_5094)
);

INVx1_ASAP7_75t_L g5095 ( 
.A(n_4348),
.Y(n_5095)
);

INVx1_ASAP7_75t_L g5096 ( 
.A(n_4348),
.Y(n_5096)
);

CKINVDCx8_ASAP7_75t_R g5097 ( 
.A(n_4069),
.Y(n_5097)
);

INVx1_ASAP7_75t_L g5098 ( 
.A(n_4348),
.Y(n_5098)
);

NAND2xp5_ASAP7_75t_L g5099 ( 
.A(n_4372),
.B(n_2587),
.Y(n_5099)
);

NAND2xp5_ASAP7_75t_SL g5100 ( 
.A(n_4354),
.B(n_2733),
.Y(n_5100)
);

BUFx6f_ASAP7_75t_L g5101 ( 
.A(n_4064),
.Y(n_5101)
);

BUFx6f_ASAP7_75t_L g5102 ( 
.A(n_4064),
.Y(n_5102)
);

NAND2xp5_ASAP7_75t_L g5103 ( 
.A(n_4372),
.B(n_2590),
.Y(n_5103)
);

NOR2xp33_ASAP7_75t_L g5104 ( 
.A(n_4275),
.B(n_2736),
.Y(n_5104)
);

BUFx6f_ASAP7_75t_L g5105 ( 
.A(n_4064),
.Y(n_5105)
);

INVx1_ASAP7_75t_L g5106 ( 
.A(n_4348),
.Y(n_5106)
);

INVx1_ASAP7_75t_L g5107 ( 
.A(n_4348),
.Y(n_5107)
);

INVx2_ASAP7_75t_L g5108 ( 
.A(n_4048),
.Y(n_5108)
);

CKINVDCx5p33_ASAP7_75t_R g5109 ( 
.A(n_4055),
.Y(n_5109)
);

NAND2xp5_ASAP7_75t_L g5110 ( 
.A(n_4372),
.B(n_2598),
.Y(n_5110)
);

INVx1_ASAP7_75t_L g5111 ( 
.A(n_4348),
.Y(n_5111)
);

INVx3_ASAP7_75t_L g5112 ( 
.A(n_4717),
.Y(n_5112)
);

INVx2_ASAP7_75t_L g5113 ( 
.A(n_4600),
.Y(n_5113)
);

INVx2_ASAP7_75t_L g5114 ( 
.A(n_4603),
.Y(n_5114)
);

INVx3_ASAP7_75t_L g5115 ( 
.A(n_4717),
.Y(n_5115)
);

INVx1_ASAP7_75t_L g5116 ( 
.A(n_4554),
.Y(n_5116)
);

BUFx10_ASAP7_75t_L g5117 ( 
.A(n_5008),
.Y(n_5117)
);

NAND2xp5_ASAP7_75t_SL g5118 ( 
.A(n_4624),
.B(n_2265),
.Y(n_5118)
);

INVx1_ASAP7_75t_L g5119 ( 
.A(n_4555),
.Y(n_5119)
);

INVx3_ASAP7_75t_L g5120 ( 
.A(n_4723),
.Y(n_5120)
);

INVx1_ASAP7_75t_L g5121 ( 
.A(n_4556),
.Y(n_5121)
);

INVx1_ASAP7_75t_L g5122 ( 
.A(n_4559),
.Y(n_5122)
);

INVx1_ASAP7_75t_L g5123 ( 
.A(n_4561),
.Y(n_5123)
);

NAND2xp5_ASAP7_75t_L g5124 ( 
.A(n_4571),
.B(n_2269),
.Y(n_5124)
);

BUFx3_ASAP7_75t_L g5125 ( 
.A(n_4605),
.Y(n_5125)
);

INVx1_ASAP7_75t_L g5126 ( 
.A(n_4562),
.Y(n_5126)
);

INVx1_ASAP7_75t_L g5127 ( 
.A(n_4569),
.Y(n_5127)
);

INVx3_ASAP7_75t_L g5128 ( 
.A(n_4723),
.Y(n_5128)
);

INVx1_ASAP7_75t_L g5129 ( 
.A(n_4570),
.Y(n_5129)
);

NAND2xp5_ASAP7_75t_SL g5130 ( 
.A(n_4674),
.B(n_2270),
.Y(n_5130)
);

INVx3_ASAP7_75t_L g5131 ( 
.A(n_4546),
.Y(n_5131)
);

INVx2_ASAP7_75t_L g5132 ( 
.A(n_4613),
.Y(n_5132)
);

OR2x2_ASAP7_75t_L g5133 ( 
.A(n_4589),
.B(n_2929),
.Y(n_5133)
);

INVx2_ASAP7_75t_L g5134 ( 
.A(n_4616),
.Y(n_5134)
);

OR2x6_ASAP7_75t_L g5135 ( 
.A(n_4839),
.B(n_2599),
.Y(n_5135)
);

INVx1_ASAP7_75t_L g5136 ( 
.A(n_4587),
.Y(n_5136)
);

CKINVDCx5p33_ASAP7_75t_R g5137 ( 
.A(n_4550),
.Y(n_5137)
);

BUFx10_ASAP7_75t_L g5138 ( 
.A(n_5008),
.Y(n_5138)
);

NAND2xp5_ASAP7_75t_SL g5139 ( 
.A(n_4771),
.B(n_2271),
.Y(n_5139)
);

INVx1_ASAP7_75t_L g5140 ( 
.A(n_4590),
.Y(n_5140)
);

INVxp33_ASAP7_75t_SL g5141 ( 
.A(n_4558),
.Y(n_5141)
);

INVx5_ASAP7_75t_L g5142 ( 
.A(n_4969),
.Y(n_5142)
);

INVx1_ASAP7_75t_L g5143 ( 
.A(n_4592),
.Y(n_5143)
);

INVx2_ASAP7_75t_L g5144 ( 
.A(n_4649),
.Y(n_5144)
);

BUFx2_ASAP7_75t_L g5145 ( 
.A(n_4566),
.Y(n_5145)
);

NAND2xp5_ASAP7_75t_L g5146 ( 
.A(n_4578),
.B(n_2274),
.Y(n_5146)
);

INVx3_ASAP7_75t_L g5147 ( 
.A(n_4546),
.Y(n_5147)
);

INVx2_ASAP7_75t_L g5148 ( 
.A(n_4658),
.Y(n_5148)
);

INVx2_ASAP7_75t_L g5149 ( 
.A(n_4666),
.Y(n_5149)
);

INVx1_ASAP7_75t_L g5150 ( 
.A(n_4593),
.Y(n_5150)
);

AOI22xp5_ASAP7_75t_L g5151 ( 
.A1(n_4989),
.A2(n_2997),
.B1(n_3016),
.B2(n_2983),
.Y(n_5151)
);

OAI22xp5_ASAP7_75t_L g5152 ( 
.A1(n_4991),
.A2(n_3096),
.B1(n_3114),
.B2(n_3050),
.Y(n_5152)
);

INVx2_ASAP7_75t_L g5153 ( 
.A(n_4675),
.Y(n_5153)
);

OR2x2_ASAP7_75t_L g5154 ( 
.A(n_5033),
.B(n_3126),
.Y(n_5154)
);

INVx3_ASAP7_75t_L g5155 ( 
.A(n_4582),
.Y(n_5155)
);

INVx3_ASAP7_75t_L g5156 ( 
.A(n_4582),
.Y(n_5156)
);

AOI22xp33_ASAP7_75t_L g5157 ( 
.A1(n_4888),
.A2(n_2632),
.B1(n_2633),
.B2(n_2625),
.Y(n_5157)
);

INVx2_ASAP7_75t_L g5158 ( 
.A(n_4677),
.Y(n_5158)
);

INVx1_ASAP7_75t_L g5159 ( 
.A(n_4597),
.Y(n_5159)
);

INVx1_ASAP7_75t_L g5160 ( 
.A(n_4599),
.Y(n_5160)
);

INVx1_ASAP7_75t_L g5161 ( 
.A(n_4604),
.Y(n_5161)
);

NAND3xp33_ASAP7_75t_L g5162 ( 
.A(n_4659),
.B(n_2756),
.C(n_2743),
.Y(n_5162)
);

AOI22xp33_ASAP7_75t_L g5163 ( 
.A1(n_4833),
.A2(n_4925),
.B1(n_4927),
.B2(n_4919),
.Y(n_5163)
);

INVx2_ASAP7_75t_L g5164 ( 
.A(n_4679),
.Y(n_5164)
);

INVx1_ASAP7_75t_L g5165 ( 
.A(n_4606),
.Y(n_5165)
);

NAND2xp5_ASAP7_75t_SL g5166 ( 
.A(n_4955),
.B(n_2283),
.Y(n_5166)
);

NAND2xp5_ASAP7_75t_SL g5167 ( 
.A(n_4955),
.B(n_2284),
.Y(n_5167)
);

INVx2_ASAP7_75t_SL g5168 ( 
.A(n_4565),
.Y(n_5168)
);

NAND2xp33_ASAP7_75t_L g5169 ( 
.A(n_4833),
.B(n_2762),
.Y(n_5169)
);

INVx4_ASAP7_75t_L g5170 ( 
.A(n_4814),
.Y(n_5170)
);

INVx2_ASAP7_75t_SL g5171 ( 
.A(n_4774),
.Y(n_5171)
);

INVx1_ASAP7_75t_L g5172 ( 
.A(n_4681),
.Y(n_5172)
);

AOI22xp33_ASAP7_75t_L g5173 ( 
.A1(n_4931),
.A2(n_2643),
.B1(n_2649),
.B2(n_2640),
.Y(n_5173)
);

AND2x6_ASAP7_75t_L g5174 ( 
.A(n_4745),
.B(n_2653),
.Y(n_5174)
);

INVx3_ASAP7_75t_L g5175 ( 
.A(n_4583),
.Y(n_5175)
);

NAND2xp33_ASAP7_75t_SL g5176 ( 
.A(n_4750),
.B(n_2768),
.Y(n_5176)
);

INVx2_ASAP7_75t_L g5177 ( 
.A(n_4686),
.Y(n_5177)
);

INVx3_ASAP7_75t_L g5178 ( 
.A(n_4583),
.Y(n_5178)
);

INVx2_ASAP7_75t_L g5179 ( 
.A(n_4687),
.Y(n_5179)
);

INVx2_ASAP7_75t_L g5180 ( 
.A(n_4543),
.Y(n_5180)
);

AOI21x1_ASAP7_75t_L g5181 ( 
.A1(n_4618),
.A2(n_2668),
.B(n_2660),
.Y(n_5181)
);

BUFx2_ASAP7_75t_L g5182 ( 
.A(n_4648),
.Y(n_5182)
);

INVx2_ASAP7_75t_SL g5183 ( 
.A(n_4545),
.Y(n_5183)
);

INVx2_ASAP7_75t_L g5184 ( 
.A(n_4544),
.Y(n_5184)
);

INVx1_ASAP7_75t_L g5185 ( 
.A(n_4882),
.Y(n_5185)
);

INVx2_ASAP7_75t_L g5186 ( 
.A(n_4557),
.Y(n_5186)
);

INVx2_ASAP7_75t_L g5187 ( 
.A(n_4564),
.Y(n_5187)
);

INVx2_ASAP7_75t_L g5188 ( 
.A(n_4568),
.Y(n_5188)
);

INVx1_ASAP7_75t_L g5189 ( 
.A(n_4884),
.Y(n_5189)
);

INVx1_ASAP7_75t_L g5190 ( 
.A(n_4572),
.Y(n_5190)
);

AOI22xp5_ASAP7_75t_L g5191 ( 
.A1(n_4711),
.A2(n_3161),
.B1(n_3217),
.B2(n_3143),
.Y(n_5191)
);

NAND2xp5_ASAP7_75t_L g5192 ( 
.A(n_4553),
.B(n_2285),
.Y(n_5192)
);

NOR2xp33_ASAP7_75t_L g5193 ( 
.A(n_5041),
.B(n_5055),
.Y(n_5193)
);

NOR2xp33_ASAP7_75t_L g5194 ( 
.A(n_5104),
.B(n_3270),
.Y(n_5194)
);

BUFx6f_ASAP7_75t_L g5195 ( 
.A(n_4617),
.Y(n_5195)
);

CKINVDCx5p33_ASAP7_75t_R g5196 ( 
.A(n_4588),
.Y(n_5196)
);

INVx2_ASAP7_75t_L g5197 ( 
.A(n_4574),
.Y(n_5197)
);

NAND2xp5_ASAP7_75t_L g5198 ( 
.A(n_4886),
.B(n_2286),
.Y(n_5198)
);

AOI22xp33_ASAP7_75t_L g5199 ( 
.A1(n_4921),
.A2(n_2678),
.B1(n_2681),
.B2(n_2671),
.Y(n_5199)
);

INVx2_ASAP7_75t_L g5200 ( 
.A(n_4580),
.Y(n_5200)
);

INVx3_ASAP7_75t_L g5201 ( 
.A(n_4617),
.Y(n_5201)
);

INVx1_ASAP7_75t_L g5202 ( 
.A(n_4594),
.Y(n_5202)
);

INVx2_ASAP7_75t_L g5203 ( 
.A(n_5036),
.Y(n_5203)
);

AOI22xp33_ASAP7_75t_SL g5204 ( 
.A1(n_4856),
.A2(n_3386),
.B1(n_3412),
.B2(n_3199),
.Y(n_5204)
);

INVx2_ASAP7_75t_L g5205 ( 
.A(n_5037),
.Y(n_5205)
);

INVx1_ASAP7_75t_L g5206 ( 
.A(n_5046),
.Y(n_5206)
);

INVx2_ASAP7_75t_L g5207 ( 
.A(n_5047),
.Y(n_5207)
);

BUFx3_ASAP7_75t_L g5208 ( 
.A(n_4620),
.Y(n_5208)
);

AND2x4_ASAP7_75t_L g5209 ( 
.A(n_4661),
.B(n_2687),
.Y(n_5209)
);

INVx2_ASAP7_75t_L g5210 ( 
.A(n_5056),
.Y(n_5210)
);

OAI22xp33_ASAP7_75t_L g5211 ( 
.A1(n_4988),
.A2(n_3608),
.B1(n_3500),
.B2(n_2774),
.Y(n_5211)
);

AOI22xp33_ASAP7_75t_L g5212 ( 
.A1(n_4921),
.A2(n_2712),
.B1(n_2714),
.B2(n_2698),
.Y(n_5212)
);

INVx2_ASAP7_75t_L g5213 ( 
.A(n_5061),
.Y(n_5213)
);

INVx2_ASAP7_75t_L g5214 ( 
.A(n_5062),
.Y(n_5214)
);

AO21x2_ASAP7_75t_L g5215 ( 
.A1(n_5038),
.A2(n_2724),
.B(n_2717),
.Y(n_5215)
);

NOR2xp33_ASAP7_75t_L g5216 ( 
.A(n_5072),
.B(n_2773),
.Y(n_5216)
);

AND2x2_ASAP7_75t_L g5217 ( 
.A(n_4626),
.B(n_3199),
.Y(n_5217)
);

INVx1_ASAP7_75t_L g5218 ( 
.A(n_5068),
.Y(n_5218)
);

NAND2xp5_ASAP7_75t_SL g5219 ( 
.A(n_4803),
.B(n_4805),
.Y(n_5219)
);

INVx1_ASAP7_75t_L g5220 ( 
.A(n_5075),
.Y(n_5220)
);

BUFx6f_ASAP7_75t_L g5221 ( 
.A(n_4623),
.Y(n_5221)
);

AND2x2_ASAP7_75t_SL g5222 ( 
.A(n_4548),
.B(n_2725),
.Y(n_5222)
);

NOR2xp33_ASAP7_75t_L g5223 ( 
.A(n_5090),
.B(n_2776),
.Y(n_5223)
);

NOR2xp33_ASAP7_75t_L g5224 ( 
.A(n_4943),
.B(n_2782),
.Y(n_5224)
);

NAND2xp5_ASAP7_75t_L g5225 ( 
.A(n_4891),
.B(n_2291),
.Y(n_5225)
);

INVx1_ASAP7_75t_L g5226 ( 
.A(n_5108),
.Y(n_5226)
);

AND2x6_ASAP7_75t_L g5227 ( 
.A(n_4745),
.B(n_2734),
.Y(n_5227)
);

NAND2xp5_ASAP7_75t_L g5228 ( 
.A(n_4899),
.B(n_2292),
.Y(n_5228)
);

BUFx6f_ASAP7_75t_L g5229 ( 
.A(n_4623),
.Y(n_5229)
);

NAND2xp5_ASAP7_75t_SL g5230 ( 
.A(n_4824),
.B(n_2299),
.Y(n_5230)
);

NAND2xp5_ASAP7_75t_SL g5231 ( 
.A(n_4737),
.B(n_2302),
.Y(n_5231)
);

INVx3_ASAP7_75t_L g5232 ( 
.A(n_4638),
.Y(n_5232)
);

INVx1_ASAP7_75t_L g5233 ( 
.A(n_4842),
.Y(n_5233)
);

INVxp33_ASAP7_75t_L g5234 ( 
.A(n_4898),
.Y(n_5234)
);

INVx2_ASAP7_75t_L g5235 ( 
.A(n_4848),
.Y(n_5235)
);

INVx2_ASAP7_75t_L g5236 ( 
.A(n_4849),
.Y(n_5236)
);

INVx2_ASAP7_75t_L g5237 ( 
.A(n_4851),
.Y(n_5237)
);

INVx2_ASAP7_75t_L g5238 ( 
.A(n_4861),
.Y(n_5238)
);

INVx2_ASAP7_75t_L g5239 ( 
.A(n_4862),
.Y(n_5239)
);

INVx2_ASAP7_75t_L g5240 ( 
.A(n_4868),
.Y(n_5240)
);

BUFx2_ASAP7_75t_L g5241 ( 
.A(n_4648),
.Y(n_5241)
);

BUFx6f_ASAP7_75t_L g5242 ( 
.A(n_4638),
.Y(n_5242)
);

OAI22xp33_ASAP7_75t_SL g5243 ( 
.A1(n_4744),
.A2(n_2786),
.B1(n_2787),
.B2(n_2783),
.Y(n_5243)
);

AOI22xp33_ASAP7_75t_L g5244 ( 
.A1(n_4607),
.A2(n_2778),
.B1(n_2781),
.B2(n_2759),
.Y(n_5244)
);

NOR2xp33_ASAP7_75t_L g5245 ( 
.A(n_4949),
.B(n_2788),
.Y(n_5245)
);

INVx2_ASAP7_75t_L g5246 ( 
.A(n_4872),
.Y(n_5246)
);

NAND2xp5_ASAP7_75t_L g5247 ( 
.A(n_4900),
.B(n_4901),
.Y(n_5247)
);

INVx4_ASAP7_75t_L g5248 ( 
.A(n_4814),
.Y(n_5248)
);

INVx1_ASAP7_75t_L g5249 ( 
.A(n_4874),
.Y(n_5249)
);

NAND2xp5_ASAP7_75t_L g5250 ( 
.A(n_4902),
.B(n_2303),
.Y(n_5250)
);

INVx1_ASAP7_75t_L g5251 ( 
.A(n_4835),
.Y(n_5251)
);

INVx2_ASAP7_75t_L g5252 ( 
.A(n_4761),
.Y(n_5252)
);

INVx2_ASAP7_75t_L g5253 ( 
.A(n_4765),
.Y(n_5253)
);

NAND2xp5_ASAP7_75t_SL g5254 ( 
.A(n_4764),
.B(n_2304),
.Y(n_5254)
);

NAND2xp5_ASAP7_75t_SL g5255 ( 
.A(n_4957),
.B(n_2309),
.Y(n_5255)
);

INVx2_ASAP7_75t_SL g5256 ( 
.A(n_5049),
.Y(n_5256)
);

INVx3_ASAP7_75t_L g5257 ( 
.A(n_4656),
.Y(n_5257)
);

INVx1_ASAP7_75t_L g5258 ( 
.A(n_4846),
.Y(n_5258)
);

OAI22xp33_ASAP7_75t_L g5259 ( 
.A1(n_4551),
.A2(n_5032),
.B1(n_5099),
.B2(n_5094),
.Y(n_5259)
);

INVx2_ASAP7_75t_L g5260 ( 
.A(n_4768),
.Y(n_5260)
);

NAND2xp5_ASAP7_75t_SL g5261 ( 
.A(n_4621),
.B(n_2310),
.Y(n_5261)
);

INVxp33_ASAP7_75t_L g5262 ( 
.A(n_4924),
.Y(n_5262)
);

INVx2_ASAP7_75t_L g5263 ( 
.A(n_4782),
.Y(n_5263)
);

AOI22xp5_ASAP7_75t_L g5264 ( 
.A1(n_4660),
.A2(n_2318),
.B1(n_2325),
.B2(n_2313),
.Y(n_5264)
);

INVx2_ASAP7_75t_L g5265 ( 
.A(n_4757),
.Y(n_5265)
);

INVx3_ASAP7_75t_L g5266 ( 
.A(n_4656),
.Y(n_5266)
);

NAND2xp5_ASAP7_75t_SL g5267 ( 
.A(n_4584),
.B(n_2326),
.Y(n_5267)
);

BUFx6f_ASAP7_75t_L g5268 ( 
.A(n_4665),
.Y(n_5268)
);

NAND2xp33_ASAP7_75t_L g5269 ( 
.A(n_4938),
.B(n_2792),
.Y(n_5269)
);

NAND2xp5_ASAP7_75t_SL g5270 ( 
.A(n_4655),
.B(n_2330),
.Y(n_5270)
);

INVx1_ASAP7_75t_L g5271 ( 
.A(n_4678),
.Y(n_5271)
);

NAND2xp5_ASAP7_75t_SL g5272 ( 
.A(n_4673),
.B(n_2332),
.Y(n_5272)
);

INVx2_ASAP7_75t_L g5273 ( 
.A(n_4746),
.Y(n_5273)
);

CKINVDCx6p67_ASAP7_75t_R g5274 ( 
.A(n_4633),
.Y(n_5274)
);

INVx2_ASAP7_75t_L g5275 ( 
.A(n_4748),
.Y(n_5275)
);

OR2x6_ASAP7_75t_L g5276 ( 
.A(n_4839),
.B(n_2785),
.Y(n_5276)
);

INVx2_ASAP7_75t_L g5277 ( 
.A(n_4753),
.Y(n_5277)
);

INVx2_ASAP7_75t_L g5278 ( 
.A(n_4755),
.Y(n_5278)
);

INVx3_ASAP7_75t_L g5279 ( 
.A(n_4665),
.Y(n_5279)
);

NAND2xp33_ASAP7_75t_SL g5280 ( 
.A(n_4973),
.B(n_2796),
.Y(n_5280)
);

INVx1_ASAP7_75t_L g5281 ( 
.A(n_4680),
.Y(n_5281)
);

INVx2_ASAP7_75t_L g5282 ( 
.A(n_4762),
.Y(n_5282)
);

INVx1_ASAP7_75t_L g5283 ( 
.A(n_4695),
.Y(n_5283)
);

INVx2_ASAP7_75t_L g5284 ( 
.A(n_4766),
.Y(n_5284)
);

INVx1_ASAP7_75t_L g5285 ( 
.A(n_4696),
.Y(n_5285)
);

INVx1_ASAP7_75t_L g5286 ( 
.A(n_4697),
.Y(n_5286)
);

INVx2_ASAP7_75t_L g5287 ( 
.A(n_4772),
.Y(n_5287)
);

AOI22xp5_ASAP7_75t_L g5288 ( 
.A1(n_4903),
.A2(n_2343),
.B1(n_2344),
.B2(n_2341),
.Y(n_5288)
);

AOI21x1_ASAP7_75t_L g5289 ( 
.A1(n_4781),
.A2(n_4867),
.B(n_4813),
.Y(n_5289)
);

INVx2_ASAP7_75t_L g5290 ( 
.A(n_4773),
.Y(n_5290)
);

NAND2xp5_ASAP7_75t_SL g5291 ( 
.A(n_4688),
.B(n_2349),
.Y(n_5291)
);

NOR2x1p5_ASAP7_75t_L g5292 ( 
.A(n_5070),
.B(n_2797),
.Y(n_5292)
);

INVx8_ASAP7_75t_L g5293 ( 
.A(n_4999),
.Y(n_5293)
);

INVx3_ASAP7_75t_L g5294 ( 
.A(n_4668),
.Y(n_5294)
);

INVxp33_ASAP7_75t_L g5295 ( 
.A(n_5079),
.Y(n_5295)
);

AND2x2_ASAP7_75t_L g5296 ( 
.A(n_4738),
.B(n_3386),
.Y(n_5296)
);

INVx2_ASAP7_75t_L g5297 ( 
.A(n_4777),
.Y(n_5297)
);

INVx4_ASAP7_75t_L g5298 ( 
.A(n_4829),
.Y(n_5298)
);

INVx2_ASAP7_75t_L g5299 ( 
.A(n_4780),
.Y(n_5299)
);

NAND3xp33_ASAP7_75t_L g5300 ( 
.A(n_4770),
.B(n_2800),
.C(n_2798),
.Y(n_5300)
);

INVx1_ASAP7_75t_L g5301 ( 
.A(n_4698),
.Y(n_5301)
);

AND2x4_ASAP7_75t_L g5302 ( 
.A(n_4567),
.B(n_2789),
.Y(n_5302)
);

BUFx3_ASAP7_75t_L g5303 ( 
.A(n_4730),
.Y(n_5303)
);

INVx2_ASAP7_75t_L g5304 ( 
.A(n_4786),
.Y(n_5304)
);

CKINVDCx5p33_ASAP7_75t_R g5305 ( 
.A(n_4650),
.Y(n_5305)
);

OAI22xp5_ASAP7_75t_L g5306 ( 
.A1(n_4952),
.A2(n_2363),
.B1(n_2367),
.B2(n_2357),
.Y(n_5306)
);

INVx1_ASAP7_75t_SL g5307 ( 
.A(n_4769),
.Y(n_5307)
);

BUFx10_ASAP7_75t_L g5308 ( 
.A(n_5025),
.Y(n_5308)
);

INVx2_ASAP7_75t_SL g5309 ( 
.A(n_4598),
.Y(n_5309)
);

INVx2_ASAP7_75t_L g5310 ( 
.A(n_4787),
.Y(n_5310)
);

INVx1_ASAP7_75t_L g5311 ( 
.A(n_4699),
.Y(n_5311)
);

INVx2_ASAP7_75t_L g5312 ( 
.A(n_4788),
.Y(n_5312)
);

INVx2_ASAP7_75t_SL g5313 ( 
.A(n_4634),
.Y(n_5313)
);

INVx2_ASAP7_75t_L g5314 ( 
.A(n_4789),
.Y(n_5314)
);

NAND2xp5_ASAP7_75t_SL g5315 ( 
.A(n_4950),
.B(n_2369),
.Y(n_5315)
);

INVx2_ASAP7_75t_L g5316 ( 
.A(n_4840),
.Y(n_5316)
);

INVx1_ASAP7_75t_L g5317 ( 
.A(n_4706),
.Y(n_5317)
);

INVx2_ASAP7_75t_L g5318 ( 
.A(n_4878),
.Y(n_5318)
);

INVx2_ASAP7_75t_L g5319 ( 
.A(n_4863),
.Y(n_5319)
);

INVx1_ASAP7_75t_L g5320 ( 
.A(n_4707),
.Y(n_5320)
);

INVx1_ASAP7_75t_L g5321 ( 
.A(n_4708),
.Y(n_5321)
);

NAND2xp5_ASAP7_75t_L g5322 ( 
.A(n_4922),
.B(n_4932),
.Y(n_5322)
);

NAND2xp5_ASAP7_75t_SL g5323 ( 
.A(n_4950),
.B(n_4959),
.Y(n_5323)
);

INVx4_ASAP7_75t_L g5324 ( 
.A(n_4829),
.Y(n_5324)
);

NOR2xp33_ASAP7_75t_L g5325 ( 
.A(n_4960),
.B(n_2802),
.Y(n_5325)
);

INVx2_ASAP7_75t_L g5326 ( 
.A(n_4866),
.Y(n_5326)
);

INVx2_ASAP7_75t_L g5327 ( 
.A(n_4873),
.Y(n_5327)
);

NAND2xp5_ASAP7_75t_L g5328 ( 
.A(n_4942),
.B(n_2373),
.Y(n_5328)
);

CKINVDCx5p33_ASAP7_75t_R g5329 ( 
.A(n_4654),
.Y(n_5329)
);

INVx1_ASAP7_75t_L g5330 ( 
.A(n_4712),
.Y(n_5330)
);

INVx1_ASAP7_75t_L g5331 ( 
.A(n_4716),
.Y(n_5331)
);

INVx2_ASAP7_75t_L g5332 ( 
.A(n_4718),
.Y(n_5332)
);

INVx4_ASAP7_75t_L g5333 ( 
.A(n_4730),
.Y(n_5333)
);

AOI22xp33_ASAP7_75t_SL g5334 ( 
.A1(n_4729),
.A2(n_3531),
.B1(n_3544),
.B2(n_3412),
.Y(n_5334)
);

INVx1_ASAP7_75t_L g5335 ( 
.A(n_4721),
.Y(n_5335)
);

INVx1_ASAP7_75t_L g5336 ( 
.A(n_4725),
.Y(n_5336)
);

INVx4_ASAP7_75t_L g5337 ( 
.A(n_4969),
.Y(n_5337)
);

AO21x2_ASAP7_75t_L g5338 ( 
.A1(n_5082),
.A2(n_2799),
.B(n_2790),
.Y(n_5338)
);

NAND2xp33_ASAP7_75t_R g5339 ( 
.A(n_4778),
.B(n_2806),
.Y(n_5339)
);

NAND2xp5_ASAP7_75t_L g5340 ( 
.A(n_4947),
.B(n_2374),
.Y(n_5340)
);

BUFx10_ASAP7_75t_L g5341 ( 
.A(n_5025),
.Y(n_5341)
);

INVx2_ASAP7_75t_L g5342 ( 
.A(n_4728),
.Y(n_5342)
);

INVx3_ASAP7_75t_L g5343 ( 
.A(n_4668),
.Y(n_5343)
);

NAND2xp5_ASAP7_75t_SL g5344 ( 
.A(n_4733),
.B(n_2375),
.Y(n_5344)
);

BUFx6f_ASAP7_75t_L g5345 ( 
.A(n_4672),
.Y(n_5345)
);

INVx4_ASAP7_75t_L g5346 ( 
.A(n_4975),
.Y(n_5346)
);

NAND2xp5_ASAP7_75t_L g5347 ( 
.A(n_4732),
.B(n_2380),
.Y(n_5347)
);

CKINVDCx5p33_ASAP7_75t_R g5348 ( 
.A(n_4790),
.Y(n_5348)
);

INVx3_ASAP7_75t_L g5349 ( 
.A(n_4672),
.Y(n_5349)
);

INVx1_ASAP7_75t_L g5350 ( 
.A(n_4739),
.Y(n_5350)
);

NAND2xp5_ASAP7_75t_L g5351 ( 
.A(n_4740),
.B(n_2390),
.Y(n_5351)
);

INVx2_ASAP7_75t_SL g5352 ( 
.A(n_5083),
.Y(n_5352)
);

INVx2_ASAP7_75t_L g5353 ( 
.A(n_4742),
.Y(n_5353)
);

INVx1_ASAP7_75t_L g5354 ( 
.A(n_4818),
.Y(n_5354)
);

BUFx10_ASAP7_75t_L g5355 ( 
.A(n_4978),
.Y(n_5355)
);

INVx1_ASAP7_75t_L g5356 ( 
.A(n_4821),
.Y(n_5356)
);

INVx1_ASAP7_75t_L g5357 ( 
.A(n_4825),
.Y(n_5357)
);

AND2x4_ASAP7_75t_L g5358 ( 
.A(n_5053),
.B(n_2819),
.Y(n_5358)
);

NAND2xp5_ASAP7_75t_L g5359 ( 
.A(n_4945),
.B(n_2393),
.Y(n_5359)
);

INVx1_ASAP7_75t_L g5360 ( 
.A(n_4826),
.Y(n_5360)
);

INVx1_ASAP7_75t_L g5361 ( 
.A(n_4827),
.Y(n_5361)
);

NAND2xp33_ASAP7_75t_L g5362 ( 
.A(n_4938),
.B(n_4576),
.Y(n_5362)
);

AND2x4_ASAP7_75t_L g5363 ( 
.A(n_5073),
.B(n_5084),
.Y(n_5363)
);

INVx3_ASAP7_75t_L g5364 ( 
.A(n_4683),
.Y(n_5364)
);

INVx4_ASAP7_75t_L g5365 ( 
.A(n_4975),
.Y(n_5365)
);

INVx2_ASAP7_75t_L g5366 ( 
.A(n_4785),
.Y(n_5366)
);

BUFx3_ASAP7_75t_L g5367 ( 
.A(n_5078),
.Y(n_5367)
);

BUFx3_ASAP7_75t_L g5368 ( 
.A(n_4792),
.Y(n_5368)
);

AND2x2_ASAP7_75t_L g5369 ( 
.A(n_4552),
.B(n_3531),
.Y(n_5369)
);

NOR2xp33_ASAP7_75t_L g5370 ( 
.A(n_4743),
.B(n_2807),
.Y(n_5370)
);

NAND2xp5_ASAP7_75t_L g5371 ( 
.A(n_4946),
.B(n_2395),
.Y(n_5371)
);

NAND3xp33_ASAP7_75t_L g5372 ( 
.A(n_5103),
.B(n_2809),
.C(n_2808),
.Y(n_5372)
);

AOI22xp33_ASAP7_75t_L g5373 ( 
.A1(n_5110),
.A2(n_2824),
.B1(n_2826),
.B2(n_2823),
.Y(n_5373)
);

INVxp67_ASAP7_75t_SL g5374 ( 
.A(n_4830),
.Y(n_5374)
);

AOI22xp5_ASAP7_75t_L g5375 ( 
.A1(n_4933),
.A2(n_2403),
.B1(n_2405),
.B2(n_2401),
.Y(n_5375)
);

INVx2_ASAP7_75t_L g5376 ( 
.A(n_4793),
.Y(n_5376)
);

INVx4_ASAP7_75t_L g5377 ( 
.A(n_4977),
.Y(n_5377)
);

AOI22xp5_ASAP7_75t_L g5378 ( 
.A1(n_4837),
.A2(n_2418),
.B1(n_2422),
.B2(n_2412),
.Y(n_5378)
);

NAND2xp5_ASAP7_75t_SL g5379 ( 
.A(n_4909),
.B(n_2432),
.Y(n_5379)
);

AND2x2_ASAP7_75t_L g5380 ( 
.A(n_4964),
.B(n_3544),
.Y(n_5380)
);

INVx2_ASAP7_75t_L g5381 ( 
.A(n_4796),
.Y(n_5381)
);

AND2x2_ASAP7_75t_L g5382 ( 
.A(n_4854),
.B(n_3548),
.Y(n_5382)
);

INVxp67_ASAP7_75t_SL g5383 ( 
.A(n_4836),
.Y(n_5383)
);

NAND2xp5_ASAP7_75t_SL g5384 ( 
.A(n_4914),
.B(n_2436),
.Y(n_5384)
);

NAND2xp5_ASAP7_75t_L g5385 ( 
.A(n_4838),
.B(n_2444),
.Y(n_5385)
);

NAND2xp5_ASAP7_75t_L g5386 ( 
.A(n_4843),
.B(n_2445),
.Y(n_5386)
);

INVx2_ASAP7_75t_L g5387 ( 
.A(n_4752),
.Y(n_5387)
);

INVx2_ASAP7_75t_L g5388 ( 
.A(n_4845),
.Y(n_5388)
);

NAND2xp5_ASAP7_75t_SL g5389 ( 
.A(n_4918),
.B(n_2446),
.Y(n_5389)
);

NAND2xp5_ASAP7_75t_L g5390 ( 
.A(n_4847),
.B(n_2447),
.Y(n_5390)
);

AOI22xp5_ASAP7_75t_L g5391 ( 
.A1(n_4850),
.A2(n_2457),
.B1(n_2460),
.B2(n_2452),
.Y(n_5391)
);

BUFx3_ASAP7_75t_L g5392 ( 
.A(n_4792),
.Y(n_5392)
);

INVx3_ASAP7_75t_L g5393 ( 
.A(n_4683),
.Y(n_5393)
);

INVx2_ASAP7_75t_L g5394 ( 
.A(n_4852),
.Y(n_5394)
);

INVx2_ASAP7_75t_SL g5395 ( 
.A(n_4560),
.Y(n_5395)
);

INVx1_ASAP7_75t_L g5396 ( 
.A(n_4853),
.Y(n_5396)
);

NAND2xp5_ASAP7_75t_SL g5397 ( 
.A(n_4939),
.B(n_2464),
.Y(n_5397)
);

INVx2_ASAP7_75t_L g5398 ( 
.A(n_4855),
.Y(n_5398)
);

AOI22xp33_ASAP7_75t_L g5399 ( 
.A1(n_4876),
.A2(n_2846),
.B1(n_2849),
.B2(n_2841),
.Y(n_5399)
);

NOR2xp33_ASAP7_75t_L g5400 ( 
.A(n_4763),
.B(n_4941),
.Y(n_5400)
);

INVx1_ASAP7_75t_L g5401 ( 
.A(n_4877),
.Y(n_5401)
);

INVx2_ASAP7_75t_L g5402 ( 
.A(n_4883),
.Y(n_5402)
);

CKINVDCx5p33_ASAP7_75t_R g5403 ( 
.A(n_4915),
.Y(n_5403)
);

INVx1_ASAP7_75t_L g5404 ( 
.A(n_4907),
.Y(n_5404)
);

INVx2_ASAP7_75t_L g5405 ( 
.A(n_4908),
.Y(n_5405)
);

INVx2_ASAP7_75t_L g5406 ( 
.A(n_4912),
.Y(n_5406)
);

NAND2xp5_ASAP7_75t_SL g5407 ( 
.A(n_4880),
.B(n_2467),
.Y(n_5407)
);

INVx2_ASAP7_75t_L g5408 ( 
.A(n_4916),
.Y(n_5408)
);

INVx1_ASAP7_75t_L g5409 ( 
.A(n_4905),
.Y(n_5409)
);

INVx3_ASAP7_75t_L g5410 ( 
.A(n_4713),
.Y(n_5410)
);

AND2x2_ASAP7_75t_L g5411 ( 
.A(n_4630),
.B(n_3548),
.Y(n_5411)
);

INVx1_ASAP7_75t_L g5412 ( 
.A(n_4911),
.Y(n_5412)
);

INVx1_ASAP7_75t_L g5413 ( 
.A(n_4881),
.Y(n_5413)
);

NAND2xp5_ASAP7_75t_SL g5414 ( 
.A(n_4890),
.B(n_4958),
.Y(n_5414)
);

NAND2xp5_ASAP7_75t_SL g5415 ( 
.A(n_4860),
.B(n_2469),
.Y(n_5415)
);

INVx1_ASAP7_75t_L g5416 ( 
.A(n_4547),
.Y(n_5416)
);

INVx1_ASAP7_75t_L g5417 ( 
.A(n_4549),
.Y(n_5417)
);

NOR2xp33_ASAP7_75t_L g5418 ( 
.A(n_4928),
.B(n_2810),
.Y(n_5418)
);

INVx2_ASAP7_75t_SL g5419 ( 
.A(n_5051),
.Y(n_5419)
);

INVx1_ASAP7_75t_L g5420 ( 
.A(n_5030),
.Y(n_5420)
);

AOI22xp33_ASAP7_75t_SL g5421 ( 
.A1(n_4625),
.A2(n_2813),
.B1(n_2818),
.B2(n_2812),
.Y(n_5421)
);

NAND2xp5_ASAP7_75t_SL g5422 ( 
.A(n_5031),
.B(n_2472),
.Y(n_5422)
);

BUFx2_ASAP7_75t_L g5423 ( 
.A(n_4731),
.Y(n_5423)
);

INVx2_ASAP7_75t_L g5424 ( 
.A(n_4784),
.Y(n_5424)
);

OR2x2_ASAP7_75t_L g5425 ( 
.A(n_5058),
.B(n_5100),
.Y(n_5425)
);

CKINVDCx5p33_ASAP7_75t_R g5426 ( 
.A(n_4926),
.Y(n_5426)
);

INVx2_ASAP7_75t_L g5427 ( 
.A(n_4784),
.Y(n_5427)
);

OR2x6_ASAP7_75t_L g5428 ( 
.A(n_4858),
.B(n_2869),
.Y(n_5428)
);

INVx1_ASAP7_75t_L g5429 ( 
.A(n_5034),
.Y(n_5429)
);

INVx1_ASAP7_75t_L g5430 ( 
.A(n_5035),
.Y(n_5430)
);

BUFx10_ASAP7_75t_L g5431 ( 
.A(n_4700),
.Y(n_5431)
);

NAND2xp5_ASAP7_75t_SL g5432 ( 
.A(n_5039),
.B(n_2479),
.Y(n_5432)
);

INVx4_ASAP7_75t_L g5433 ( 
.A(n_4977),
.Y(n_5433)
);

INVx1_ASAP7_75t_L g5434 ( 
.A(n_5042),
.Y(n_5434)
);

BUFx6f_ASAP7_75t_L g5435 ( 
.A(n_4713),
.Y(n_5435)
);

INVx2_ASAP7_75t_L g5436 ( 
.A(n_4758),
.Y(n_5436)
);

OAI22xp33_ASAP7_75t_L g5437 ( 
.A1(n_4889),
.A2(n_2835),
.B1(n_2838),
.B2(n_2825),
.Y(n_5437)
);

NAND2xp5_ASAP7_75t_SL g5438 ( 
.A(n_5043),
.B(n_2480),
.Y(n_5438)
);

INVx1_ASAP7_75t_L g5439 ( 
.A(n_5045),
.Y(n_5439)
);

INVx1_ASAP7_75t_L g5440 ( 
.A(n_5054),
.Y(n_5440)
);

INVx2_ASAP7_75t_L g5441 ( 
.A(n_4758),
.Y(n_5441)
);

INVx1_ASAP7_75t_L g5442 ( 
.A(n_5057),
.Y(n_5442)
);

NOR2xp33_ASAP7_75t_L g5443 ( 
.A(n_4929),
.B(n_2853),
.Y(n_5443)
);

INVx1_ASAP7_75t_L g5444 ( 
.A(n_5060),
.Y(n_5444)
);

INVx2_ASAP7_75t_L g5445 ( 
.A(n_4760),
.Y(n_5445)
);

INVx3_ASAP7_75t_L g5446 ( 
.A(n_4714),
.Y(n_5446)
);

INVx1_ASAP7_75t_L g5447 ( 
.A(n_5063),
.Y(n_5447)
);

INVx1_ASAP7_75t_L g5448 ( 
.A(n_5064),
.Y(n_5448)
);

NAND2xp5_ASAP7_75t_L g5449 ( 
.A(n_4859),
.B(n_2485),
.Y(n_5449)
);

INVx3_ASAP7_75t_L g5450 ( 
.A(n_4714),
.Y(n_5450)
);

AND3x1_ASAP7_75t_L g5451 ( 
.A(n_5014),
.B(n_2888),
.C(n_2885),
.Y(n_5451)
);

INVx2_ASAP7_75t_L g5452 ( 
.A(n_4760),
.Y(n_5452)
);

NAND2xp33_ASAP7_75t_R g5453 ( 
.A(n_4794),
.B(n_2854),
.Y(n_5453)
);

INVx2_ASAP7_75t_L g5454 ( 
.A(n_4779),
.Y(n_5454)
);

AOI22xp33_ASAP7_75t_L g5455 ( 
.A1(n_5052),
.A2(n_2892),
.B1(n_2922),
.B2(n_2889),
.Y(n_5455)
);

NAND2xp5_ASAP7_75t_L g5456 ( 
.A(n_4944),
.B(n_4581),
.Y(n_5456)
);

AND2x6_ASAP7_75t_L g5457 ( 
.A(n_4779),
.B(n_2927),
.Y(n_5457)
);

INVx5_ASAP7_75t_L g5458 ( 
.A(n_4858),
.Y(n_5458)
);

INVx2_ASAP7_75t_SL g5459 ( 
.A(n_5091),
.Y(n_5459)
);

AO21x2_ASAP7_75t_L g5460 ( 
.A1(n_4585),
.A2(n_2937),
.B(n_2935),
.Y(n_5460)
);

INVxp67_ASAP7_75t_SL g5461 ( 
.A(n_4575),
.Y(n_5461)
);

INVx2_ASAP7_75t_SL g5462 ( 
.A(n_4692),
.Y(n_5462)
);

OAI22x1_ASAP7_75t_L g5463 ( 
.A1(n_5013),
.A2(n_2861),
.B1(n_2866),
.B2(n_2858),
.Y(n_5463)
);

NAND2xp5_ASAP7_75t_SL g5464 ( 
.A(n_5066),
.B(n_5069),
.Y(n_5464)
);

NOR2xp33_ASAP7_75t_L g5465 ( 
.A(n_4930),
.B(n_2867),
.Y(n_5465)
);

OAI21xp33_ASAP7_75t_SL g5466 ( 
.A1(n_4962),
.A2(n_2960),
.B(n_2946),
.Y(n_5466)
);

INVx2_ASAP7_75t_L g5467 ( 
.A(n_4756),
.Y(n_5467)
);

NAND2xp5_ASAP7_75t_SL g5468 ( 
.A(n_5071),
.B(n_5076),
.Y(n_5468)
);

INVx2_ASAP7_75t_L g5469 ( 
.A(n_4756),
.Y(n_5469)
);

INVx4_ASAP7_75t_L g5470 ( 
.A(n_4879),
.Y(n_5470)
);

NAND2xp33_ASAP7_75t_SL g5471 ( 
.A(n_5018),
.B(n_2872),
.Y(n_5471)
);

NOR2xp33_ASAP7_75t_L g5472 ( 
.A(n_4934),
.B(n_2877),
.Y(n_5472)
);

NOR2xp33_ASAP7_75t_L g5473 ( 
.A(n_4937),
.B(n_2893),
.Y(n_5473)
);

INVx2_ASAP7_75t_SL g5474 ( 
.A(n_4719),
.Y(n_5474)
);

INVx2_ASAP7_75t_L g5475 ( 
.A(n_5077),
.Y(n_5475)
);

NAND2xp5_ASAP7_75t_L g5476 ( 
.A(n_4870),
.B(n_4940),
.Y(n_5476)
);

CKINVDCx5p33_ASAP7_75t_R g5477 ( 
.A(n_5109),
.Y(n_5477)
);

INVx1_ASAP7_75t_L g5478 ( 
.A(n_5080),
.Y(n_5478)
);

AND3x2_ASAP7_75t_L g5479 ( 
.A(n_4609),
.B(n_2968),
.C(n_2962),
.Y(n_5479)
);

AND2x2_ASAP7_75t_L g5480 ( 
.A(n_4754),
.B(n_2894),
.Y(n_5480)
);

INVx1_ASAP7_75t_SL g5481 ( 
.A(n_4892),
.Y(n_5481)
);

INVx3_ASAP7_75t_L g5482 ( 
.A(n_4715),
.Y(n_5482)
);

INVx4_ASAP7_75t_L g5483 ( 
.A(n_4879),
.Y(n_5483)
);

INVx3_ASAP7_75t_L g5484 ( 
.A(n_4715),
.Y(n_5484)
);

INVx2_ASAP7_75t_SL g5485 ( 
.A(n_4724),
.Y(n_5485)
);

INVx2_ASAP7_75t_L g5486 ( 
.A(n_5081),
.Y(n_5486)
);

BUFx3_ASAP7_75t_L g5487 ( 
.A(n_4631),
.Y(n_5487)
);

NAND2xp5_ASAP7_75t_SL g5488 ( 
.A(n_5085),
.B(n_2487),
.Y(n_5488)
);

INVx4_ASAP7_75t_L g5489 ( 
.A(n_4894),
.Y(n_5489)
);

INVx1_ASAP7_75t_L g5490 ( 
.A(n_5086),
.Y(n_5490)
);

BUFx3_ASAP7_75t_L g5491 ( 
.A(n_4705),
.Y(n_5491)
);

NAND2xp5_ASAP7_75t_L g5492 ( 
.A(n_4864),
.B(n_2490),
.Y(n_5492)
);

INVx2_ASAP7_75t_L g5493 ( 
.A(n_5087),
.Y(n_5493)
);

NAND2xp5_ASAP7_75t_SL g5494 ( 
.A(n_5088),
.B(n_2491),
.Y(n_5494)
);

AND2x4_ASAP7_75t_L g5495 ( 
.A(n_4735),
.B(n_2971),
.Y(n_5495)
);

INVx1_ASAP7_75t_L g5496 ( 
.A(n_5089),
.Y(n_5496)
);

BUFx6f_ASAP7_75t_L g5497 ( 
.A(n_5040),
.Y(n_5497)
);

INVx2_ASAP7_75t_L g5498 ( 
.A(n_5092),
.Y(n_5498)
);

NOR2xp33_ASAP7_75t_L g5499 ( 
.A(n_4804),
.B(n_2907),
.Y(n_5499)
);

NOR2xp33_ASAP7_75t_L g5500 ( 
.A(n_4808),
.B(n_2909),
.Y(n_5500)
);

OAI22xp33_ASAP7_75t_L g5501 ( 
.A1(n_4895),
.A2(n_2916),
.B1(n_2942),
.B2(n_2911),
.Y(n_5501)
);

INVx2_ASAP7_75t_L g5502 ( 
.A(n_5093),
.Y(n_5502)
);

INVx8_ASAP7_75t_L g5503 ( 
.A(n_4731),
.Y(n_5503)
);

AND2x6_ASAP7_75t_L g5504 ( 
.A(n_5027),
.B(n_2990),
.Y(n_5504)
);

NAND3xp33_ASAP7_75t_L g5505 ( 
.A(n_5044),
.B(n_2944),
.C(n_2943),
.Y(n_5505)
);

AND2x2_ASAP7_75t_SL g5506 ( 
.A(n_4685),
.B(n_2996),
.Y(n_5506)
);

CKINVDCx20_ASAP7_75t_R g5507 ( 
.A(n_4971),
.Y(n_5507)
);

INVx1_ASAP7_75t_SL g5508 ( 
.A(n_4967),
.Y(n_5508)
);

NOR2xp33_ASAP7_75t_L g5509 ( 
.A(n_4811),
.B(n_2951),
.Y(n_5509)
);

INVx3_ASAP7_75t_L g5510 ( 
.A(n_5040),
.Y(n_5510)
);

BUFx10_ASAP7_75t_L g5511 ( 
.A(n_4894),
.Y(n_5511)
);

INVx1_ASAP7_75t_L g5512 ( 
.A(n_5095),
.Y(n_5512)
);

INVx2_ASAP7_75t_L g5513 ( 
.A(n_5096),
.Y(n_5513)
);

CKINVDCx5p33_ASAP7_75t_R g5514 ( 
.A(n_4767),
.Y(n_5514)
);

AOI22xp33_ASAP7_75t_L g5515 ( 
.A1(n_4970),
.A2(n_3003),
.B1(n_3006),
.B2(n_3002),
.Y(n_5515)
);

INVx1_ASAP7_75t_L g5516 ( 
.A(n_5098),
.Y(n_5516)
);

CKINVDCx5p33_ASAP7_75t_R g5517 ( 
.A(n_4820),
.Y(n_5517)
);

INVx2_ASAP7_75t_L g5518 ( 
.A(n_5106),
.Y(n_5518)
);

AOI22xp33_ASAP7_75t_L g5519 ( 
.A1(n_4741),
.A2(n_3021),
.B1(n_3035),
.B2(n_3020),
.Y(n_5519)
);

INVx2_ASAP7_75t_L g5520 ( 
.A(n_5107),
.Y(n_5520)
);

INVx2_ASAP7_75t_L g5521 ( 
.A(n_5111),
.Y(n_5521)
);

OR2x2_ASAP7_75t_L g5522 ( 
.A(n_4951),
.B(n_4812),
.Y(n_5522)
);

NAND2xp33_ASAP7_75t_SL g5523 ( 
.A(n_5012),
.B(n_4968),
.Y(n_5523)
);

AOI22xp33_ASAP7_75t_L g5524 ( 
.A1(n_4819),
.A2(n_3039),
.B1(n_3045),
.B2(n_3038),
.Y(n_5524)
);

INVx2_ASAP7_75t_L g5525 ( 
.A(n_4802),
.Y(n_5525)
);

NOR2x1p5_ASAP7_75t_L g5526 ( 
.A(n_4586),
.B(n_2952),
.Y(n_5526)
);

BUFx6f_ASAP7_75t_SL g5527 ( 
.A(n_5017),
.Y(n_5527)
);

NOR2xp33_ASAP7_75t_L g5528 ( 
.A(n_4816),
.B(n_2953),
.Y(n_5528)
);

XNOR2xp5_ASAP7_75t_L g5529 ( 
.A(n_4701),
.B(n_2493),
.Y(n_5529)
);

CKINVDCx5p33_ASAP7_75t_R g5530 ( 
.A(n_4831),
.Y(n_5530)
);

INVx2_ASAP7_75t_L g5531 ( 
.A(n_4822),
.Y(n_5531)
);

INVx1_ASAP7_75t_L g5532 ( 
.A(n_4710),
.Y(n_5532)
);

INVx2_ASAP7_75t_L g5533 ( 
.A(n_4828),
.Y(n_5533)
);

BUFx3_ASAP7_75t_L g5534 ( 
.A(n_4801),
.Y(n_5534)
);

INVx1_ASAP7_75t_L g5535 ( 
.A(n_4759),
.Y(n_5535)
);

INVx1_ASAP7_75t_L g5536 ( 
.A(n_4776),
.Y(n_5536)
);

BUFx4f_ASAP7_75t_L g5537 ( 
.A(n_5048),
.Y(n_5537)
);

INVx2_ASAP7_75t_L g5538 ( 
.A(n_4690),
.Y(n_5538)
);

INVx3_ASAP7_75t_L g5539 ( 
.A(n_5050),
.Y(n_5539)
);

INVx1_ASAP7_75t_L g5540 ( 
.A(n_4807),
.Y(n_5540)
);

INVx3_ASAP7_75t_L g5541 ( 
.A(n_5050),
.Y(n_5541)
);

INVx2_ASAP7_75t_L g5542 ( 
.A(n_4691),
.Y(n_5542)
);

OAI22xp33_ASAP7_75t_L g5543 ( 
.A1(n_4817),
.A2(n_2965),
.B1(n_2966),
.B2(n_2957),
.Y(n_5543)
);

AOI22xp5_ASAP7_75t_L g5544 ( 
.A1(n_4979),
.A2(n_2501),
.B1(n_2504),
.B2(n_2499),
.Y(n_5544)
);

INVx1_ASAP7_75t_L g5545 ( 
.A(n_4810),
.Y(n_5545)
);

AOI22xp33_ASAP7_75t_L g5546 ( 
.A1(n_4869),
.A2(n_5010),
.B1(n_4887),
.B2(n_4935),
.Y(n_5546)
);

BUFx3_ASAP7_75t_L g5547 ( 
.A(n_4749),
.Y(n_5547)
);

INVx1_ASAP7_75t_L g5548 ( 
.A(n_4797),
.Y(n_5548)
);

INVx2_ASAP7_75t_L g5549 ( 
.A(n_4693),
.Y(n_5549)
);

AOI22xp5_ASAP7_75t_L g5550 ( 
.A1(n_4727),
.A2(n_2509),
.B1(n_2515),
.B2(n_2505),
.Y(n_5550)
);

NAND3xp33_ASAP7_75t_L g5551 ( 
.A(n_4875),
.B(n_2978),
.C(n_2973),
.Y(n_5551)
);

INVx1_ASAP7_75t_L g5552 ( 
.A(n_4798),
.Y(n_5552)
);

INVx1_ASAP7_75t_L g5553 ( 
.A(n_4799),
.Y(n_5553)
);

AOI22xp33_ASAP7_75t_L g5554 ( 
.A1(n_4885),
.A2(n_3048),
.B1(n_3052),
.B2(n_3047),
.Y(n_5554)
);

INVx2_ASAP7_75t_L g5555 ( 
.A(n_4704),
.Y(n_5555)
);

NAND2xp5_ASAP7_75t_L g5556 ( 
.A(n_4595),
.B(n_2517),
.Y(n_5556)
);

INVx1_ASAP7_75t_L g5557 ( 
.A(n_4800),
.Y(n_5557)
);

BUFx3_ASAP7_75t_L g5558 ( 
.A(n_5067),
.Y(n_5558)
);

NOR2xp33_ASAP7_75t_L g5559 ( 
.A(n_4694),
.B(n_2994),
.Y(n_5559)
);

INVx1_ASAP7_75t_L g5560 ( 
.A(n_4611),
.Y(n_5560)
);

NOR2xp33_ASAP7_75t_R g5561 ( 
.A(n_4722),
.B(n_2999),
.Y(n_5561)
);

NOR2xp33_ASAP7_75t_L g5562 ( 
.A(n_4976),
.B(n_3004),
.Y(n_5562)
);

INVx1_ASAP7_75t_L g5563 ( 
.A(n_4612),
.Y(n_5563)
);

INVx2_ASAP7_75t_L g5564 ( 
.A(n_4709),
.Y(n_5564)
);

INVx2_ASAP7_75t_L g5565 ( 
.A(n_4726),
.Y(n_5565)
);

NAND2xp5_ASAP7_75t_L g5566 ( 
.A(n_4608),
.B(n_2522),
.Y(n_5566)
);

NAND2xp5_ASAP7_75t_SL g5567 ( 
.A(n_4653),
.B(n_2524),
.Y(n_5567)
);

INVx2_ASAP7_75t_L g5568 ( 
.A(n_4736),
.Y(n_5568)
);

BUFx3_ASAP7_75t_L g5569 ( 
.A(n_5067),
.Y(n_5569)
);

INVx1_ASAP7_75t_L g5570 ( 
.A(n_4614),
.Y(n_5570)
);

INVx2_ASAP7_75t_SL g5571 ( 
.A(n_4783),
.Y(n_5571)
);

NOR2xp33_ASAP7_75t_L g5572 ( 
.A(n_4982),
.B(n_3011),
.Y(n_5572)
);

INVx1_ASAP7_75t_L g5573 ( 
.A(n_4619),
.Y(n_5573)
);

BUFx4f_ASAP7_75t_L g5574 ( 
.A(n_5048),
.Y(n_5574)
);

INVx3_ASAP7_75t_L g5575 ( 
.A(n_5074),
.Y(n_5575)
);

INVx1_ASAP7_75t_L g5576 ( 
.A(n_4629),
.Y(n_5576)
);

INVx2_ASAP7_75t_L g5577 ( 
.A(n_4751),
.Y(n_5577)
);

NAND2xp5_ASAP7_75t_L g5578 ( 
.A(n_4667),
.B(n_2526),
.Y(n_5578)
);

INVx2_ASAP7_75t_L g5579 ( 
.A(n_4682),
.Y(n_5579)
);

INVx2_ASAP7_75t_L g5580 ( 
.A(n_4689),
.Y(n_5580)
);

INVx3_ASAP7_75t_L g5581 ( 
.A(n_5074),
.Y(n_5581)
);

INVx1_ASAP7_75t_L g5582 ( 
.A(n_4632),
.Y(n_5582)
);

INVx2_ASAP7_75t_L g5583 ( 
.A(n_4635),
.Y(n_5583)
);

NAND2xp5_ASAP7_75t_L g5584 ( 
.A(n_4904),
.B(n_2527),
.Y(n_5584)
);

NOR2xp33_ASAP7_75t_L g5585 ( 
.A(n_4972),
.B(n_3014),
.Y(n_5585)
);

NAND2xp33_ASAP7_75t_R g5586 ( 
.A(n_4980),
.B(n_3028),
.Y(n_5586)
);

INVx3_ASAP7_75t_L g5587 ( 
.A(n_5101),
.Y(n_5587)
);

NAND2xp5_ASAP7_75t_L g5588 ( 
.A(n_4910),
.B(n_2528),
.Y(n_5588)
);

INVx1_ASAP7_75t_L g5589 ( 
.A(n_4636),
.Y(n_5589)
);

INVx1_ASAP7_75t_L g5590 ( 
.A(n_4637),
.Y(n_5590)
);

CKINVDCx11_ASAP7_75t_R g5591 ( 
.A(n_4734),
.Y(n_5591)
);

INVx1_ASAP7_75t_L g5592 ( 
.A(n_4640),
.Y(n_5592)
);

INVxp67_ASAP7_75t_SL g5593 ( 
.A(n_4596),
.Y(n_5593)
);

NAND2xp5_ASAP7_75t_SL g5594 ( 
.A(n_4871),
.B(n_2533),
.Y(n_5594)
);

INVx1_ASAP7_75t_L g5595 ( 
.A(n_4642),
.Y(n_5595)
);

NAND2xp33_ASAP7_75t_L g5596 ( 
.A(n_4834),
.B(n_3029),
.Y(n_5596)
);

INVx1_ASAP7_75t_L g5597 ( 
.A(n_4643),
.Y(n_5597)
);

INVx3_ASAP7_75t_L g5598 ( 
.A(n_5101),
.Y(n_5598)
);

NAND3xp33_ASAP7_75t_L g5599 ( 
.A(n_4974),
.B(n_3036),
.C(n_3033),
.Y(n_5599)
);

INVx2_ASAP7_75t_L g5600 ( 
.A(n_4645),
.Y(n_5600)
);

INVx4_ASAP7_75t_L g5601 ( 
.A(n_5102),
.Y(n_5601)
);

INVx2_ASAP7_75t_L g5602 ( 
.A(n_4646),
.Y(n_5602)
);

NAND2xp5_ASAP7_75t_SL g5603 ( 
.A(n_4893),
.B(n_2534),
.Y(n_5603)
);

CKINVDCx5p33_ASAP7_75t_R g5604 ( 
.A(n_4983),
.Y(n_5604)
);

INVx2_ASAP7_75t_L g5605 ( 
.A(n_4647),
.Y(n_5605)
);

INVx2_ASAP7_75t_L g5606 ( 
.A(n_4651),
.Y(n_5606)
);

INVx2_ASAP7_75t_L g5607 ( 
.A(n_4657),
.Y(n_5607)
);

INVx2_ASAP7_75t_L g5608 ( 
.A(n_4662),
.Y(n_5608)
);

INVx2_ASAP7_75t_L g5609 ( 
.A(n_4663),
.Y(n_5609)
);

INVx2_ASAP7_75t_SL g5610 ( 
.A(n_4563),
.Y(n_5610)
);

INVx2_ASAP7_75t_L g5611 ( 
.A(n_4670),
.Y(n_5611)
);

INVx2_ASAP7_75t_SL g5612 ( 
.A(n_4823),
.Y(n_5612)
);

NAND2xp5_ASAP7_75t_SL g5613 ( 
.A(n_4684),
.B(n_4981),
.Y(n_5613)
);

BUFx10_ASAP7_75t_L g5614 ( 
.A(n_4995),
.Y(n_5614)
);

INVx2_ASAP7_75t_L g5615 ( 
.A(n_4671),
.Y(n_5615)
);

AO22x2_ASAP7_75t_L g5616 ( 
.A1(n_5023),
.A2(n_3064),
.B1(n_3066),
.B2(n_3059),
.Y(n_5616)
);

NAND2xp5_ASAP7_75t_L g5617 ( 
.A(n_4841),
.B(n_2535),
.Y(n_5617)
);

INVx2_ASAP7_75t_L g5618 ( 
.A(n_4676),
.Y(n_5618)
);

NAND2xp5_ASAP7_75t_L g5619 ( 
.A(n_4747),
.B(n_2536),
.Y(n_5619)
);

INVx3_ASAP7_75t_L g5620 ( 
.A(n_5102),
.Y(n_5620)
);

NOR2xp33_ASAP7_75t_L g5621 ( 
.A(n_4984),
.B(n_3055),
.Y(n_5621)
);

INVx2_ASAP7_75t_L g5622 ( 
.A(n_5105),
.Y(n_5622)
);

INVx1_ASAP7_75t_L g5623 ( 
.A(n_4602),
.Y(n_5623)
);

INVx5_ASAP7_75t_L g5624 ( 
.A(n_4963),
.Y(n_5624)
);

INVxp67_ASAP7_75t_L g5625 ( 
.A(n_4806),
.Y(n_5625)
);

INVx1_ASAP7_75t_L g5626 ( 
.A(n_4652),
.Y(n_5626)
);

INVx1_ASAP7_75t_L g5627 ( 
.A(n_5105),
.Y(n_5627)
);

NOR2xp67_ASAP7_75t_L g5628 ( 
.A(n_4684),
.B(n_2537),
.Y(n_5628)
);

INVx1_ASAP7_75t_L g5629 ( 
.A(n_4917),
.Y(n_5629)
);

INVx8_ASAP7_75t_L g5630 ( 
.A(n_5065),
.Y(n_5630)
);

INVx1_ASAP7_75t_L g5631 ( 
.A(n_4573),
.Y(n_5631)
);

INVx2_ASAP7_75t_L g5632 ( 
.A(n_4615),
.Y(n_5632)
);

INVx2_ASAP7_75t_L g5633 ( 
.A(n_4639),
.Y(n_5633)
);

NAND2xp5_ASAP7_75t_SL g5634 ( 
.A(n_4985),
.B(n_2538),
.Y(n_5634)
);

INVx2_ASAP7_75t_SL g5635 ( 
.A(n_4986),
.Y(n_5635)
);

NAND2xp5_ASAP7_75t_SL g5636 ( 
.A(n_4987),
.B(n_2542),
.Y(n_5636)
);

INVx1_ASAP7_75t_L g5637 ( 
.A(n_4641),
.Y(n_5637)
);

INVx1_ASAP7_75t_L g5638 ( 
.A(n_4644),
.Y(n_5638)
);

INVx1_ASAP7_75t_L g5639 ( 
.A(n_4702),
.Y(n_5639)
);

NOR3xp33_ASAP7_75t_L g5640 ( 
.A(n_4844),
.B(n_2550),
.C(n_2548),
.Y(n_5640)
);

INVx3_ASAP7_75t_L g5641 ( 
.A(n_4948),
.Y(n_5641)
);

INVx2_ASAP7_75t_SL g5642 ( 
.A(n_4865),
.Y(n_5642)
);

INVx2_ASAP7_75t_L g5643 ( 
.A(n_5007),
.Y(n_5643)
);

BUFx6f_ASAP7_75t_L g5644 ( 
.A(n_4963),
.Y(n_5644)
);

INVx2_ASAP7_75t_L g5645 ( 
.A(n_4896),
.Y(n_5645)
);

INVxp67_ASAP7_75t_SL g5646 ( 
.A(n_4720),
.Y(n_5646)
);

INVx1_ASAP7_75t_L g5647 ( 
.A(n_4791),
.Y(n_5647)
);

INVx3_ASAP7_75t_L g5648 ( 
.A(n_4961),
.Y(n_5648)
);

NAND2xp5_ASAP7_75t_SL g5649 ( 
.A(n_4997),
.B(n_2551),
.Y(n_5649)
);

INVx4_ASAP7_75t_L g5650 ( 
.A(n_4601),
.Y(n_5650)
);

INVx2_ASAP7_75t_L g5651 ( 
.A(n_4965),
.Y(n_5651)
);

OR2x2_ASAP7_75t_L g5652 ( 
.A(n_4953),
.B(n_3060),
.Y(n_5652)
);

INVx2_ASAP7_75t_SL g5653 ( 
.A(n_5059),
.Y(n_5653)
);

NAND2xp5_ASAP7_75t_L g5654 ( 
.A(n_4809),
.B(n_2554),
.Y(n_5654)
);

INVx2_ASAP7_75t_L g5655 ( 
.A(n_4954),
.Y(n_5655)
);

INVx2_ASAP7_75t_L g5656 ( 
.A(n_4956),
.Y(n_5656)
);

INVx2_ASAP7_75t_L g5657 ( 
.A(n_4966),
.Y(n_5657)
);

BUFx6f_ASAP7_75t_L g5658 ( 
.A(n_5097),
.Y(n_5658)
);

INVx2_ASAP7_75t_L g5659 ( 
.A(n_5388),
.Y(n_5659)
);

INVx1_ASAP7_75t_L g5660 ( 
.A(n_5116),
.Y(n_5660)
);

AND2x2_ASAP7_75t_L g5661 ( 
.A(n_5194),
.B(n_4998),
.Y(n_5661)
);

INVx1_ASAP7_75t_L g5662 ( 
.A(n_5119),
.Y(n_5662)
);

INVx1_ASAP7_75t_L g5663 ( 
.A(n_5121),
.Y(n_5663)
);

AND2x6_ASAP7_75t_L g5664 ( 
.A(n_5217),
.B(n_5000),
.Y(n_5664)
);

OAI22xp5_ASAP7_75t_L g5665 ( 
.A1(n_5193),
.A2(n_5002),
.B1(n_5016),
.B2(n_4832),
.Y(n_5665)
);

INVx1_ASAP7_75t_L g5666 ( 
.A(n_5122),
.Y(n_5666)
);

INVx1_ASAP7_75t_L g5667 ( 
.A(n_5123),
.Y(n_5667)
);

INVxp67_ASAP7_75t_SL g5668 ( 
.A(n_5163),
.Y(n_5668)
);

NAND2xp5_ASAP7_75t_L g5669 ( 
.A(n_5247),
.B(n_5322),
.Y(n_5669)
);

BUFx6f_ASAP7_75t_L g5670 ( 
.A(n_5644),
.Y(n_5670)
);

AND3x4_ASAP7_75t_L g5671 ( 
.A(n_5640),
.B(n_5026),
.C(n_5009),
.Y(n_5671)
);

INVx1_ASAP7_75t_L g5672 ( 
.A(n_5126),
.Y(n_5672)
);

CKINVDCx5p33_ASAP7_75t_R g5673 ( 
.A(n_5137),
.Y(n_5673)
);

INVx1_ASAP7_75t_L g5674 ( 
.A(n_5127),
.Y(n_5674)
);

INVx5_ASAP7_75t_L g5675 ( 
.A(n_5658),
.Y(n_5675)
);

INVx1_ASAP7_75t_L g5676 ( 
.A(n_5129),
.Y(n_5676)
);

INVx2_ASAP7_75t_L g5677 ( 
.A(n_5394),
.Y(n_5677)
);

INVx2_ASAP7_75t_SL g5678 ( 
.A(n_5145),
.Y(n_5678)
);

INVx1_ASAP7_75t_L g5679 ( 
.A(n_5136),
.Y(n_5679)
);

INVx2_ASAP7_75t_L g5680 ( 
.A(n_5398),
.Y(n_5680)
);

INVx1_ASAP7_75t_L g5681 ( 
.A(n_5140),
.Y(n_5681)
);

INVxp67_ASAP7_75t_SL g5682 ( 
.A(n_5436),
.Y(n_5682)
);

NOR2xp33_ASAP7_75t_L g5683 ( 
.A(n_5234),
.B(n_4775),
.Y(n_5683)
);

NAND2xp5_ASAP7_75t_L g5684 ( 
.A(n_5224),
.B(n_4834),
.Y(n_5684)
);

BUFx3_ASAP7_75t_L g5685 ( 
.A(n_5644),
.Y(n_5685)
);

INVx1_ASAP7_75t_L g5686 ( 
.A(n_5143),
.Y(n_5686)
);

INVx1_ASAP7_75t_L g5687 ( 
.A(n_5150),
.Y(n_5687)
);

BUFx6f_ASAP7_75t_L g5688 ( 
.A(n_5195),
.Y(n_5688)
);

NAND2x1p5_ASAP7_75t_L g5689 ( 
.A(n_5333),
.B(n_4669),
.Y(n_5689)
);

NOR2xp33_ASAP7_75t_L g5690 ( 
.A(n_5295),
.B(n_5024),
.Y(n_5690)
);

NAND2xp5_ASAP7_75t_L g5691 ( 
.A(n_5124),
.B(n_4897),
.Y(n_5691)
);

INVx3_ASAP7_75t_L g5692 ( 
.A(n_5195),
.Y(n_5692)
);

INVx2_ASAP7_75t_L g5693 ( 
.A(n_5402),
.Y(n_5693)
);

INVx4_ASAP7_75t_L g5694 ( 
.A(n_5458),
.Y(n_5694)
);

AND2x2_ASAP7_75t_L g5695 ( 
.A(n_5380),
.B(n_5005),
.Y(n_5695)
);

NAND2xp5_ASAP7_75t_L g5696 ( 
.A(n_5146),
.B(n_4897),
.Y(n_5696)
);

NOR2xp33_ASAP7_75t_L g5697 ( 
.A(n_5219),
.B(n_5400),
.Y(n_5697)
);

INVx1_ASAP7_75t_SL g5698 ( 
.A(n_5481),
.Y(n_5698)
);

INVx1_ASAP7_75t_SL g5699 ( 
.A(n_5508),
.Y(n_5699)
);

BUFx3_ASAP7_75t_L g5700 ( 
.A(n_5303),
.Y(n_5700)
);

INVx3_ASAP7_75t_L g5701 ( 
.A(n_5221),
.Y(n_5701)
);

INVx1_ASAP7_75t_L g5702 ( 
.A(n_5159),
.Y(n_5702)
);

INVx2_ASAP7_75t_L g5703 ( 
.A(n_5113),
.Y(n_5703)
);

INVx1_ASAP7_75t_L g5704 ( 
.A(n_5160),
.Y(n_5704)
);

INVx1_ASAP7_75t_SL g5705 ( 
.A(n_5307),
.Y(n_5705)
);

INVxp67_ASAP7_75t_L g5706 ( 
.A(n_5296),
.Y(n_5706)
);

INVx1_ASAP7_75t_L g5707 ( 
.A(n_5161),
.Y(n_5707)
);

NAND2xp5_ASAP7_75t_SL g5708 ( 
.A(n_5183),
.B(n_5015),
.Y(n_5708)
);

BUFx6f_ASAP7_75t_L g5709 ( 
.A(n_5221),
.Y(n_5709)
);

INVx2_ASAP7_75t_L g5710 ( 
.A(n_5114),
.Y(n_5710)
);

NAND2xp5_ASAP7_75t_L g5711 ( 
.A(n_5192),
.B(n_4806),
.Y(n_5711)
);

INVx2_ASAP7_75t_L g5712 ( 
.A(n_5132),
.Y(n_5712)
);

BUFx6f_ASAP7_75t_L g5713 ( 
.A(n_5229),
.Y(n_5713)
);

INVx1_ASAP7_75t_L g5714 ( 
.A(n_5165),
.Y(n_5714)
);

BUFx6f_ASAP7_75t_L g5715 ( 
.A(n_5229),
.Y(n_5715)
);

INVx3_ASAP7_75t_L g5716 ( 
.A(n_5242),
.Y(n_5716)
);

AND2x4_ASAP7_75t_L g5717 ( 
.A(n_5458),
.B(n_5006),
.Y(n_5717)
);

NOR2xp33_ASAP7_75t_L g5718 ( 
.A(n_5352),
.B(n_4994),
.Y(n_5718)
);

INVx2_ASAP7_75t_L g5719 ( 
.A(n_5134),
.Y(n_5719)
);

INVx1_ASAP7_75t_L g5720 ( 
.A(n_5271),
.Y(n_5720)
);

INVx2_ASAP7_75t_SL g5721 ( 
.A(n_5142),
.Y(n_5721)
);

BUFx2_ASAP7_75t_L g5722 ( 
.A(n_5604),
.Y(n_5722)
);

AND2x4_ASAP7_75t_L g5723 ( 
.A(n_5470),
.B(n_4992),
.Y(n_5723)
);

NOR2xp33_ASAP7_75t_L g5724 ( 
.A(n_5168),
.B(n_5449),
.Y(n_5724)
);

INVx1_ASAP7_75t_L g5725 ( 
.A(n_5281),
.Y(n_5725)
);

NOR2xp33_ASAP7_75t_L g5726 ( 
.A(n_5256),
.B(n_4993),
.Y(n_5726)
);

AND2x6_ASAP7_75t_L g5727 ( 
.A(n_5369),
.B(n_5003),
.Y(n_5727)
);

INVx1_ASAP7_75t_L g5728 ( 
.A(n_5283),
.Y(n_5728)
);

NAND2xp5_ASAP7_75t_SL g5729 ( 
.A(n_5514),
.B(n_4913),
.Y(n_5729)
);

NOR2xp33_ASAP7_75t_L g5730 ( 
.A(n_5133),
.B(n_5022),
.Y(n_5730)
);

BUFx6f_ASAP7_75t_L g5731 ( 
.A(n_5242),
.Y(n_5731)
);

INVx1_ASAP7_75t_L g5732 ( 
.A(n_5285),
.Y(n_5732)
);

INVxp67_ASAP7_75t_SL g5733 ( 
.A(n_5441),
.Y(n_5733)
);

NAND2xp5_ASAP7_75t_L g5734 ( 
.A(n_5374),
.B(n_4815),
.Y(n_5734)
);

AND2x2_ASAP7_75t_L g5735 ( 
.A(n_5382),
.B(n_5245),
.Y(n_5735)
);

HB1xp67_ASAP7_75t_L g5736 ( 
.A(n_5522),
.Y(n_5736)
);

BUFx2_ASAP7_75t_L g5737 ( 
.A(n_5487),
.Y(n_5737)
);

BUFx3_ASAP7_75t_L g5738 ( 
.A(n_5368),
.Y(n_5738)
);

BUFx2_ASAP7_75t_L g5739 ( 
.A(n_5491),
.Y(n_5739)
);

NAND2xp5_ASAP7_75t_L g5740 ( 
.A(n_5383),
.B(n_4815),
.Y(n_5740)
);

INVx8_ASAP7_75t_L g5741 ( 
.A(n_5293),
.Y(n_5741)
);

INVx2_ASAP7_75t_L g5742 ( 
.A(n_5144),
.Y(n_5742)
);

NOR2xp33_ASAP7_75t_L g5743 ( 
.A(n_5652),
.B(n_5004),
.Y(n_5743)
);

INVx2_ASAP7_75t_L g5744 ( 
.A(n_5148),
.Y(n_5744)
);

NAND2x1p5_ASAP7_75t_L g5745 ( 
.A(n_5392),
.B(n_4703),
.Y(n_5745)
);

INVx1_ASAP7_75t_L g5746 ( 
.A(n_5286),
.Y(n_5746)
);

NOR2xp33_ASAP7_75t_L g5747 ( 
.A(n_5118),
.B(n_4622),
.Y(n_5747)
);

INVx1_ASAP7_75t_L g5748 ( 
.A(n_5301),
.Y(n_5748)
);

CKINVDCx20_ASAP7_75t_R g5749 ( 
.A(n_5507),
.Y(n_5749)
);

AOI22xp5_ASAP7_75t_L g5750 ( 
.A1(n_5259),
.A2(n_5011),
.B1(n_5021),
.B2(n_4906),
.Y(n_5750)
);

INVx2_ASAP7_75t_L g5751 ( 
.A(n_5149),
.Y(n_5751)
);

BUFx6f_ASAP7_75t_L g5752 ( 
.A(n_5268),
.Y(n_5752)
);

INVx1_ASAP7_75t_L g5753 ( 
.A(n_5311),
.Y(n_5753)
);

INVx1_ASAP7_75t_L g5754 ( 
.A(n_5317),
.Y(n_5754)
);

BUFx10_ASAP7_75t_L g5755 ( 
.A(n_5527),
.Y(n_5755)
);

INVx1_ASAP7_75t_L g5756 ( 
.A(n_5320),
.Y(n_5756)
);

INVx1_ASAP7_75t_L g5757 ( 
.A(n_5321),
.Y(n_5757)
);

BUFx3_ASAP7_75t_L g5758 ( 
.A(n_5268),
.Y(n_5758)
);

INVx2_ASAP7_75t_L g5759 ( 
.A(n_5153),
.Y(n_5759)
);

INVx1_ASAP7_75t_L g5760 ( 
.A(n_5330),
.Y(n_5760)
);

NAND2xp5_ASAP7_75t_L g5761 ( 
.A(n_5325),
.B(n_2561),
.Y(n_5761)
);

NAND2xp5_ASAP7_75t_SL g5762 ( 
.A(n_5517),
.B(n_4627),
.Y(n_5762)
);

NAND2xp5_ASAP7_75t_L g5763 ( 
.A(n_5476),
.B(n_2562),
.Y(n_5763)
);

NAND2xp5_ASAP7_75t_SL g5764 ( 
.A(n_5530),
.B(n_4633),
.Y(n_5764)
);

NAND2xp5_ASAP7_75t_SL g5765 ( 
.A(n_5635),
.B(n_4996),
.Y(n_5765)
);

INVx2_ASAP7_75t_L g5766 ( 
.A(n_5158),
.Y(n_5766)
);

BUFx6f_ASAP7_75t_L g5767 ( 
.A(n_5345),
.Y(n_5767)
);

INVx5_ASAP7_75t_L g5768 ( 
.A(n_5658),
.Y(n_5768)
);

NAND3xp33_ASAP7_75t_L g5769 ( 
.A(n_5370),
.B(n_5001),
.C(n_4795),
.Y(n_5769)
);

INVx2_ASAP7_75t_L g5770 ( 
.A(n_5164),
.Y(n_5770)
);

INVx1_ASAP7_75t_L g5771 ( 
.A(n_5331),
.Y(n_5771)
);

INVx2_ASAP7_75t_L g5772 ( 
.A(n_5177),
.Y(n_5772)
);

INVx2_ASAP7_75t_L g5773 ( 
.A(n_5179),
.Y(n_5773)
);

AND2x4_ASAP7_75t_L g5774 ( 
.A(n_5483),
.B(n_5028),
.Y(n_5774)
);

NAND2xp33_ASAP7_75t_L g5775 ( 
.A(n_5174),
.B(n_5227),
.Y(n_5775)
);

INVx2_ASAP7_75t_L g5776 ( 
.A(n_5180),
.Y(n_5776)
);

INVx2_ASAP7_75t_L g5777 ( 
.A(n_5184),
.Y(n_5777)
);

AND2x4_ASAP7_75t_L g5778 ( 
.A(n_5489),
.B(n_5020),
.Y(n_5778)
);

INVx1_ASAP7_75t_L g5779 ( 
.A(n_5335),
.Y(n_5779)
);

AOI22xp33_ASAP7_75t_L g5780 ( 
.A1(n_5354),
.A2(n_3080),
.B1(n_3085),
.B2(n_3071),
.Y(n_5780)
);

AND2x4_ASAP7_75t_L g5781 ( 
.A(n_5337),
.B(n_4628),
.Y(n_5781)
);

NAND2xp5_ASAP7_75t_L g5782 ( 
.A(n_5356),
.B(n_2564),
.Y(n_5782)
);

INVx2_ASAP7_75t_L g5783 ( 
.A(n_5186),
.Y(n_5783)
);

AND2x6_ASAP7_75t_L g5784 ( 
.A(n_5411),
.B(n_4990),
.Y(n_5784)
);

BUFx3_ASAP7_75t_L g5785 ( 
.A(n_5345),
.Y(n_5785)
);

AND2x4_ASAP7_75t_L g5786 ( 
.A(n_5346),
.B(n_5029),
.Y(n_5786)
);

NOR2xp33_ASAP7_75t_L g5787 ( 
.A(n_5414),
.B(n_5425),
.Y(n_5787)
);

NAND2xp5_ASAP7_75t_L g5788 ( 
.A(n_5357),
.B(n_2565),
.Y(n_5788)
);

NOR2xp33_ASAP7_75t_L g5789 ( 
.A(n_5255),
.B(n_4664),
.Y(n_5789)
);

INVx2_ASAP7_75t_L g5790 ( 
.A(n_5187),
.Y(n_5790)
);

BUFx3_ASAP7_75t_L g5791 ( 
.A(n_5435),
.Y(n_5791)
);

AND2x4_ASAP7_75t_L g5792 ( 
.A(n_5365),
.B(n_5019),
.Y(n_5792)
);

BUFx3_ASAP7_75t_L g5793 ( 
.A(n_5435),
.Y(n_5793)
);

AND2x4_ASAP7_75t_L g5794 ( 
.A(n_5377),
.B(n_4579),
.Y(n_5794)
);

OAI22xp33_ASAP7_75t_L g5795 ( 
.A1(n_5191),
.A2(n_3074),
.B1(n_3086),
.B2(n_3065),
.Y(n_5795)
);

INVx4_ASAP7_75t_SL g5796 ( 
.A(n_5504),
.Y(n_5796)
);

NAND2xp5_ASAP7_75t_L g5797 ( 
.A(n_5360),
.B(n_2570),
.Y(n_5797)
);

INVx8_ASAP7_75t_L g5798 ( 
.A(n_5293),
.Y(n_5798)
);

AND2x4_ASAP7_75t_L g5799 ( 
.A(n_5433),
.B(n_5142),
.Y(n_5799)
);

AND2x2_ASAP7_75t_L g5800 ( 
.A(n_5154),
.B(n_4577),
.Y(n_5800)
);

AND2x4_ASAP7_75t_L g5801 ( 
.A(n_5125),
.B(n_4591),
.Y(n_5801)
);

NAND2xp5_ASAP7_75t_SL g5802 ( 
.A(n_5198),
.B(n_4857),
.Y(n_5802)
);

NAND2xp5_ASAP7_75t_L g5803 ( 
.A(n_5361),
.B(n_2574),
.Y(n_5803)
);

INVx1_ASAP7_75t_L g5804 ( 
.A(n_5336),
.Y(n_5804)
);

BUFx6f_ASAP7_75t_L g5805 ( 
.A(n_5497),
.Y(n_5805)
);

INVx1_ASAP7_75t_L g5806 ( 
.A(n_5350),
.Y(n_5806)
);

CKINVDCx16_ASAP7_75t_R g5807 ( 
.A(n_5117),
.Y(n_5807)
);

INVx1_ASAP7_75t_L g5808 ( 
.A(n_5396),
.Y(n_5808)
);

INVx2_ASAP7_75t_L g5809 ( 
.A(n_5188),
.Y(n_5809)
);

INVx1_ASAP7_75t_L g5810 ( 
.A(n_5401),
.Y(n_5810)
);

INVx4_ASAP7_75t_L g5811 ( 
.A(n_5624),
.Y(n_5811)
);

OAI22xp33_ASAP7_75t_L g5812 ( 
.A1(n_5225),
.A2(n_5228),
.B1(n_5250),
.B2(n_5328),
.Y(n_5812)
);

INVx2_ASAP7_75t_L g5813 ( 
.A(n_5197),
.Y(n_5813)
);

AND2x4_ASAP7_75t_L g5814 ( 
.A(n_5208),
.B(n_4936),
.Y(n_5814)
);

CKINVDCx5p33_ASAP7_75t_R g5815 ( 
.A(n_5196),
.Y(n_5815)
);

NAND2xp5_ASAP7_75t_L g5816 ( 
.A(n_5579),
.B(n_2575),
.Y(n_5816)
);

INVx1_ASAP7_75t_L g5817 ( 
.A(n_5332),
.Y(n_5817)
);

OAI22xp33_ASAP7_75t_SL g5818 ( 
.A1(n_5130),
.A2(n_3089),
.B1(n_3097),
.B2(n_3090),
.Y(n_5818)
);

BUFx2_ASAP7_75t_L g5819 ( 
.A(n_5367),
.Y(n_5819)
);

INVx1_ASAP7_75t_L g5820 ( 
.A(n_5342),
.Y(n_5820)
);

BUFx3_ASAP7_75t_L g5821 ( 
.A(n_5497),
.Y(n_5821)
);

INVx2_ASAP7_75t_L g5822 ( 
.A(n_5200),
.Y(n_5822)
);

INVx2_ASAP7_75t_L g5823 ( 
.A(n_5203),
.Y(n_5823)
);

INVx2_ASAP7_75t_L g5824 ( 
.A(n_5205),
.Y(n_5824)
);

INVx1_ASAP7_75t_L g5825 ( 
.A(n_5353),
.Y(n_5825)
);

NAND2xp5_ASAP7_75t_L g5826 ( 
.A(n_5580),
.B(n_2576),
.Y(n_5826)
);

INVx1_ASAP7_75t_L g5827 ( 
.A(n_5172),
.Y(n_5827)
);

INVx1_ASAP7_75t_L g5828 ( 
.A(n_5190),
.Y(n_5828)
);

INVx2_ASAP7_75t_L g5829 ( 
.A(n_5207),
.Y(n_5829)
);

INVx2_ASAP7_75t_L g5830 ( 
.A(n_5210),
.Y(n_5830)
);

INVx2_ASAP7_75t_SL g5831 ( 
.A(n_5209),
.Y(n_5831)
);

OAI22xp5_ASAP7_75t_SL g5832 ( 
.A1(n_5334),
.A2(n_3105),
.B1(n_3111),
.B2(n_3102),
.Y(n_5832)
);

INVx1_ASAP7_75t_L g5833 ( 
.A(n_5202),
.Y(n_5833)
);

AND2x4_ASAP7_75t_L g5834 ( 
.A(n_5363),
.B(n_3087),
.Y(n_5834)
);

INVx8_ASAP7_75t_L g5835 ( 
.A(n_5624),
.Y(n_5835)
);

INVx1_ASAP7_75t_L g5836 ( 
.A(n_5206),
.Y(n_5836)
);

INVx2_ASAP7_75t_L g5837 ( 
.A(n_5213),
.Y(n_5837)
);

NOR2xp33_ASAP7_75t_L g5838 ( 
.A(n_5139),
.B(n_2577),
.Y(n_5838)
);

BUFx6f_ASAP7_75t_L g5839 ( 
.A(n_5511),
.Y(n_5839)
);

NOR2xp33_ASAP7_75t_L g5840 ( 
.A(n_5230),
.B(n_2578),
.Y(n_5840)
);

BUFx6f_ASAP7_75t_L g5841 ( 
.A(n_5558),
.Y(n_5841)
);

INVx2_ASAP7_75t_L g5842 ( 
.A(n_5214),
.Y(n_5842)
);

INVx2_ASAP7_75t_L g5843 ( 
.A(n_5235),
.Y(n_5843)
);

AND2x4_ASAP7_75t_L g5844 ( 
.A(n_5547),
.B(n_3092),
.Y(n_5844)
);

AND2x2_ASAP7_75t_L g5845 ( 
.A(n_5480),
.B(n_3119),
.Y(n_5845)
);

AO21x2_ASAP7_75t_L g5846 ( 
.A1(n_5467),
.A2(n_5469),
.B(n_5413),
.Y(n_5846)
);

INVx1_ASAP7_75t_L g5847 ( 
.A(n_5218),
.Y(n_5847)
);

INVx2_ASAP7_75t_L g5848 ( 
.A(n_5236),
.Y(n_5848)
);

BUFx3_ASAP7_75t_L g5849 ( 
.A(n_5569),
.Y(n_5849)
);

NAND2xp5_ASAP7_75t_SL g5850 ( 
.A(n_5171),
.B(n_4920),
.Y(n_5850)
);

INVx3_ASAP7_75t_L g5851 ( 
.A(n_5170),
.Y(n_5851)
);

AND2x4_ASAP7_75t_L g5852 ( 
.A(n_5248),
.B(n_3101),
.Y(n_5852)
);

AND2x2_ASAP7_75t_L g5853 ( 
.A(n_5562),
.B(n_3123),
.Y(n_5853)
);

INVx2_ASAP7_75t_L g5854 ( 
.A(n_5237),
.Y(n_5854)
);

INVx1_ASAP7_75t_L g5855 ( 
.A(n_5220),
.Y(n_5855)
);

INVx1_ASAP7_75t_L g5856 ( 
.A(n_5226),
.Y(n_5856)
);

AND2x2_ASAP7_75t_SL g5857 ( 
.A(n_5537),
.B(n_3110),
.Y(n_5857)
);

BUFx6f_ASAP7_75t_L g5858 ( 
.A(n_5591),
.Y(n_5858)
);

INVx2_ASAP7_75t_L g5859 ( 
.A(n_5238),
.Y(n_5859)
);

INVx4_ASAP7_75t_L g5860 ( 
.A(n_5298),
.Y(n_5860)
);

INVx4_ASAP7_75t_L g5861 ( 
.A(n_5324),
.Y(n_5861)
);

AND2x2_ASAP7_75t_L g5862 ( 
.A(n_5572),
.B(n_3128),
.Y(n_5862)
);

INVxp67_ASAP7_75t_L g5863 ( 
.A(n_5559),
.Y(n_5863)
);

BUFx6f_ASAP7_75t_L g5864 ( 
.A(n_5601),
.Y(n_5864)
);

INVx1_ASAP7_75t_L g5865 ( 
.A(n_5233),
.Y(n_5865)
);

NAND2xp5_ASAP7_75t_L g5866 ( 
.A(n_5456),
.B(n_2585),
.Y(n_5866)
);

NAND2xp33_ASAP7_75t_L g5867 ( 
.A(n_5174),
.B(n_3129),
.Y(n_5867)
);

AND2x4_ASAP7_75t_L g5868 ( 
.A(n_5534),
.B(n_3124),
.Y(n_5868)
);

NOR2xp33_ASAP7_75t_L g5869 ( 
.A(n_5216),
.B(n_2591),
.Y(n_5869)
);

NOR2xp33_ASAP7_75t_SL g5870 ( 
.A(n_5141),
.B(n_5305),
.Y(n_5870)
);

XNOR2xp5_ASAP7_75t_L g5871 ( 
.A(n_5262),
.B(n_4610),
.Y(n_5871)
);

BUFx3_ASAP7_75t_L g5872 ( 
.A(n_5138),
.Y(n_5872)
);

INVx1_ASAP7_75t_SL g5873 ( 
.A(n_5182),
.Y(n_5873)
);

AND2x4_ASAP7_75t_L g5874 ( 
.A(n_5395),
.B(n_5313),
.Y(n_5874)
);

INVx1_ASAP7_75t_L g5875 ( 
.A(n_5249),
.Y(n_5875)
);

NOR2xp33_ASAP7_75t_L g5876 ( 
.A(n_5223),
.B(n_5625),
.Y(n_5876)
);

AND2x4_ASAP7_75t_L g5877 ( 
.A(n_5419),
.B(n_3130),
.Y(n_5877)
);

INVx1_ASAP7_75t_SL g5878 ( 
.A(n_5241),
.Y(n_5878)
);

INVx1_ASAP7_75t_L g5879 ( 
.A(n_5239),
.Y(n_5879)
);

BUFx6f_ASAP7_75t_L g5880 ( 
.A(n_5308),
.Y(n_5880)
);

BUFx6f_ASAP7_75t_L g5881 ( 
.A(n_5341),
.Y(n_5881)
);

NAND2xp5_ASAP7_75t_SL g5882 ( 
.A(n_5340),
.B(n_4923),
.Y(n_5882)
);

INVx1_ASAP7_75t_L g5883 ( 
.A(n_5240),
.Y(n_5883)
);

NAND2xp5_ASAP7_75t_L g5884 ( 
.A(n_5445),
.B(n_5452),
.Y(n_5884)
);

INVx1_ASAP7_75t_L g5885 ( 
.A(n_5246),
.Y(n_5885)
);

AND2x4_ASAP7_75t_L g5886 ( 
.A(n_5459),
.B(n_3133),
.Y(n_5886)
);

NOR2xp33_ASAP7_75t_L g5887 ( 
.A(n_5461),
.B(n_2592),
.Y(n_5887)
);

INVx1_ASAP7_75t_L g5888 ( 
.A(n_5252),
.Y(n_5888)
);

AO21x2_ASAP7_75t_L g5889 ( 
.A1(n_5424),
.A2(n_3142),
.B(n_3141),
.Y(n_5889)
);

INVx1_ASAP7_75t_L g5890 ( 
.A(n_5253),
.Y(n_5890)
);

AOI22xp5_ASAP7_75t_L g5891 ( 
.A1(n_5372),
.A2(n_5169),
.B1(n_5227),
.B2(n_5174),
.Y(n_5891)
);

INVx3_ASAP7_75t_L g5892 ( 
.A(n_5112),
.Y(n_5892)
);

INVx4_ASAP7_75t_SL g5893 ( 
.A(n_5504),
.Y(n_5893)
);

AND2x2_ASAP7_75t_L g5894 ( 
.A(n_5585),
.B(n_3138),
.Y(n_5894)
);

INVx1_ASAP7_75t_L g5895 ( 
.A(n_5260),
.Y(n_5895)
);

NAND3xp33_ASAP7_75t_L g5896 ( 
.A(n_5421),
.B(n_2594),
.C(n_2593),
.Y(n_5896)
);

INVx4_ASAP7_75t_L g5897 ( 
.A(n_5431),
.Y(n_5897)
);

OR2x6_ASAP7_75t_L g5898 ( 
.A(n_5630),
.B(n_3145),
.Y(n_5898)
);

AO22x2_ASAP7_75t_L g5899 ( 
.A1(n_5152),
.A2(n_5306),
.B1(n_5300),
.B2(n_5162),
.Y(n_5899)
);

AND2x4_ASAP7_75t_L g5900 ( 
.A(n_5309),
.B(n_3198),
.Y(n_5900)
);

NOR2x1p5_ASAP7_75t_L g5901 ( 
.A(n_5274),
.B(n_3144),
.Y(n_5901)
);

INVx4_ASAP7_75t_SL g5902 ( 
.A(n_5504),
.Y(n_5902)
);

INVx2_ASAP7_75t_L g5903 ( 
.A(n_5263),
.Y(n_5903)
);

BUFx6f_ASAP7_75t_L g5904 ( 
.A(n_5115),
.Y(n_5904)
);

AND2x2_ASAP7_75t_L g5905 ( 
.A(n_5621),
.B(n_3149),
.Y(n_5905)
);

NOR2xp33_ASAP7_75t_L g5906 ( 
.A(n_5593),
.B(n_2595),
.Y(n_5906)
);

INVx1_ASAP7_75t_SL g5907 ( 
.A(n_5423),
.Y(n_5907)
);

NAND2xp5_ASAP7_75t_L g5908 ( 
.A(n_5454),
.B(n_2597),
.Y(n_5908)
);

AND2x4_ASAP7_75t_L g5909 ( 
.A(n_5655),
.B(n_3201),
.Y(n_5909)
);

INVx1_ASAP7_75t_L g5910 ( 
.A(n_5265),
.Y(n_5910)
);

INVx2_ASAP7_75t_SL g5911 ( 
.A(n_5302),
.Y(n_5911)
);

NAND2xp5_ASAP7_75t_SL g5912 ( 
.A(n_5222),
.B(n_2600),
.Y(n_5912)
);

INVx2_ASAP7_75t_L g5913 ( 
.A(n_5273),
.Y(n_5913)
);

AO22x2_ASAP7_75t_L g5914 ( 
.A1(n_5645),
.A2(n_3227),
.B1(n_3241),
.B2(n_3232),
.Y(n_5914)
);

INVx1_ASAP7_75t_L g5915 ( 
.A(n_5275),
.Y(n_5915)
);

INVx1_ASAP7_75t_L g5916 ( 
.A(n_5277),
.Y(n_5916)
);

AND2x4_ASAP7_75t_L g5917 ( 
.A(n_5656),
.B(n_3247),
.Y(n_5917)
);

INVx1_ASAP7_75t_L g5918 ( 
.A(n_5278),
.Y(n_5918)
);

AND2x4_ASAP7_75t_L g5919 ( 
.A(n_5657),
.B(n_3260),
.Y(n_5919)
);

INVx3_ASAP7_75t_L g5920 ( 
.A(n_5120),
.Y(n_5920)
);

INVx4_ASAP7_75t_L g5921 ( 
.A(n_5329),
.Y(n_5921)
);

INVx2_ASAP7_75t_L g5922 ( 
.A(n_5282),
.Y(n_5922)
);

AO21x2_ASAP7_75t_L g5923 ( 
.A1(n_5427),
.A2(n_3289),
.B(n_3277),
.Y(n_5923)
);

INVx1_ASAP7_75t_L g5924 ( 
.A(n_5284),
.Y(n_5924)
);

NAND2xp5_ASAP7_75t_L g5925 ( 
.A(n_5359),
.B(n_2613),
.Y(n_5925)
);

INVx1_ASAP7_75t_L g5926 ( 
.A(n_5287),
.Y(n_5926)
);

INVx2_ASAP7_75t_L g5927 ( 
.A(n_5290),
.Y(n_5927)
);

INVx2_ASAP7_75t_L g5928 ( 
.A(n_5297),
.Y(n_5928)
);

NOR2xp33_ASAP7_75t_L g5929 ( 
.A(n_5532),
.B(n_2617),
.Y(n_5929)
);

INVx1_ASAP7_75t_L g5930 ( 
.A(n_5299),
.Y(n_5930)
);

INVx2_ASAP7_75t_L g5931 ( 
.A(n_5304),
.Y(n_5931)
);

NAND2xp5_ASAP7_75t_SL g5932 ( 
.A(n_5506),
.B(n_2618),
.Y(n_5932)
);

BUFx3_ASAP7_75t_L g5933 ( 
.A(n_5128),
.Y(n_5933)
);

INVx2_ASAP7_75t_L g5934 ( 
.A(n_5310),
.Y(n_5934)
);

BUFx6f_ASAP7_75t_L g5935 ( 
.A(n_5131),
.Y(n_5935)
);

INVx1_ASAP7_75t_L g5936 ( 
.A(n_5312),
.Y(n_5936)
);

INVx2_ASAP7_75t_SL g5937 ( 
.A(n_5358),
.Y(n_5937)
);

OAI22xp33_ASAP7_75t_L g5938 ( 
.A1(n_5264),
.A2(n_5151),
.B1(n_5588),
.B2(n_5584),
.Y(n_5938)
);

OAI221xp5_ASAP7_75t_L g5939 ( 
.A1(n_5373),
.A2(n_3323),
.B1(n_3324),
.B2(n_3318),
.C(n_3302),
.Y(n_5939)
);

INVxp33_ASAP7_75t_L g5940 ( 
.A(n_5529),
.Y(n_5940)
);

NAND2x1p5_ASAP7_75t_L g5941 ( 
.A(n_5610),
.B(n_5147),
.Y(n_5941)
);

BUFx10_ASAP7_75t_L g5942 ( 
.A(n_5348),
.Y(n_5942)
);

NOR2x1p5_ASAP7_75t_L g5943 ( 
.A(n_5403),
.B(n_3157),
.Y(n_5943)
);

BUFx6f_ASAP7_75t_SL g5944 ( 
.A(n_5355),
.Y(n_5944)
);

INVx5_ASAP7_75t_L g5945 ( 
.A(n_5503),
.Y(n_5945)
);

INVx1_ASAP7_75t_L g5946 ( 
.A(n_5314),
.Y(n_5946)
);

AND2x6_ASAP7_75t_L g5947 ( 
.A(n_5643),
.B(n_3341),
.Y(n_5947)
);

BUFx3_ASAP7_75t_L g5948 ( 
.A(n_5155),
.Y(n_5948)
);

AND2x2_ASAP7_75t_L g5949 ( 
.A(n_5499),
.B(n_3158),
.Y(n_5949)
);

INVx1_ASAP7_75t_L g5950 ( 
.A(n_5319),
.Y(n_5950)
);

INVx1_ASAP7_75t_L g5951 ( 
.A(n_5326),
.Y(n_5951)
);

INVx3_ASAP7_75t_L g5952 ( 
.A(n_5156),
.Y(n_5952)
);

INVx1_ASAP7_75t_L g5953 ( 
.A(n_5327),
.Y(n_5953)
);

NAND2xp33_ASAP7_75t_L g5954 ( 
.A(n_5227),
.B(n_5457),
.Y(n_5954)
);

HB1xp67_ASAP7_75t_L g5955 ( 
.A(n_5623),
.Y(n_5955)
);

INVx1_ASAP7_75t_L g5956 ( 
.A(n_5316),
.Y(n_5956)
);

AND2x2_ASAP7_75t_L g5957 ( 
.A(n_5500),
.B(n_5509),
.Y(n_5957)
);

NAND2xp5_ASAP7_75t_L g5958 ( 
.A(n_5371),
.B(n_2620),
.Y(n_5958)
);

NOR2xp33_ASAP7_75t_L g5959 ( 
.A(n_5617),
.B(n_2622),
.Y(n_5959)
);

OAI22xp5_ASAP7_75t_L g5960 ( 
.A1(n_5173),
.A2(n_2626),
.B1(n_2631),
.B2(n_2624),
.Y(n_5960)
);

AND2x4_ASAP7_75t_L g5961 ( 
.A(n_5462),
.B(n_3345),
.Y(n_5961)
);

NOR2xp33_ASAP7_75t_L g5962 ( 
.A(n_5626),
.B(n_2634),
.Y(n_5962)
);

INVx1_ASAP7_75t_L g5963 ( 
.A(n_5318),
.Y(n_5963)
);

INVx2_ASAP7_75t_L g5964 ( 
.A(n_5366),
.Y(n_5964)
);

INVx2_ASAP7_75t_SL g5965 ( 
.A(n_5622),
.Y(n_5965)
);

BUFx6f_ASAP7_75t_L g5966 ( 
.A(n_5175),
.Y(n_5966)
);

INVx1_ASAP7_75t_L g5967 ( 
.A(n_5376),
.Y(n_5967)
);

INVx4_ASAP7_75t_L g5968 ( 
.A(n_5426),
.Y(n_5968)
);

INVx8_ASAP7_75t_L g5969 ( 
.A(n_5457),
.Y(n_5969)
);

INVx1_ASAP7_75t_L g5970 ( 
.A(n_5381),
.Y(n_5970)
);

BUFx3_ASAP7_75t_L g5971 ( 
.A(n_5178),
.Y(n_5971)
);

BUFx2_ASAP7_75t_L g5972 ( 
.A(n_5457),
.Y(n_5972)
);

BUFx6f_ASAP7_75t_L g5973 ( 
.A(n_5201),
.Y(n_5973)
);

AO22x2_ASAP7_75t_L g5974 ( 
.A1(n_5642),
.A2(n_3348),
.B1(n_3359),
.B2(n_3353),
.Y(n_5974)
);

INVx1_ASAP7_75t_L g5975 ( 
.A(n_5409),
.Y(n_5975)
);

BUFx2_ASAP7_75t_L g5976 ( 
.A(n_5176),
.Y(n_5976)
);

INVx1_ASAP7_75t_L g5977 ( 
.A(n_5412),
.Y(n_5977)
);

AOI22xp33_ASAP7_75t_L g5978 ( 
.A1(n_5244),
.A2(n_3371),
.B1(n_3373),
.B2(n_3369),
.Y(n_5978)
);

INVx1_ASAP7_75t_L g5979 ( 
.A(n_5185),
.Y(n_5979)
);

INVx4_ASAP7_75t_L g5980 ( 
.A(n_5477),
.Y(n_5980)
);

INVx2_ASAP7_75t_L g5981 ( 
.A(n_5405),
.Y(n_5981)
);

INVx1_ASAP7_75t_L g5982 ( 
.A(n_5189),
.Y(n_5982)
);

INVx1_ASAP7_75t_L g5983 ( 
.A(n_5404),
.Y(n_5983)
);

NAND2xp5_ASAP7_75t_L g5984 ( 
.A(n_5157),
.B(n_2638),
.Y(n_5984)
);

AND2x4_ASAP7_75t_L g5985 ( 
.A(n_5474),
.B(n_5485),
.Y(n_5985)
);

INVx1_ASAP7_75t_L g5986 ( 
.A(n_5416),
.Y(n_5986)
);

AO21x2_ASAP7_75t_L g5987 ( 
.A1(n_5387),
.A2(n_3384),
.B(n_3382),
.Y(n_5987)
);

INVx1_ASAP7_75t_SL g5988 ( 
.A(n_5561),
.Y(n_5988)
);

INVx1_ASAP7_75t_L g5989 ( 
.A(n_5417),
.Y(n_5989)
);

NAND2xp5_ASAP7_75t_SL g5990 ( 
.A(n_5612),
.B(n_2644),
.Y(n_5990)
);

INVx1_ASAP7_75t_L g5991 ( 
.A(n_5420),
.Y(n_5991)
);

NOR3xp33_ASAP7_75t_SL g5992 ( 
.A(n_5339),
.B(n_3160),
.C(n_3159),
.Y(n_5992)
);

INVx1_ASAP7_75t_L g5993 ( 
.A(n_5429),
.Y(n_5993)
);

INVx2_ASAP7_75t_L g5994 ( 
.A(n_5406),
.Y(n_5994)
);

NOR2xp33_ASAP7_75t_SL g5995 ( 
.A(n_5574),
.B(n_5503),
.Y(n_5995)
);

CKINVDCx5p33_ASAP7_75t_R g5996 ( 
.A(n_5453),
.Y(n_5996)
);

AOI22xp33_ASAP7_75t_L g5997 ( 
.A1(n_5519),
.A2(n_3390),
.B1(n_3401),
.B2(n_3385),
.Y(n_5997)
);

INVx1_ASAP7_75t_L g5998 ( 
.A(n_5430),
.Y(n_5998)
);

INVx1_ASAP7_75t_L g5999 ( 
.A(n_5434),
.Y(n_5999)
);

INVx1_ASAP7_75t_L g6000 ( 
.A(n_5439),
.Y(n_6000)
);

AND2x4_ASAP7_75t_L g6001 ( 
.A(n_5651),
.B(n_3415),
.Y(n_6001)
);

INVx4_ASAP7_75t_L g6002 ( 
.A(n_5232),
.Y(n_6002)
);

INVx1_ASAP7_75t_L g6003 ( 
.A(n_5440),
.Y(n_6003)
);

NAND3xp33_ASAP7_75t_L g6004 ( 
.A(n_5204),
.B(n_2648),
.C(n_2646),
.Y(n_6004)
);

INVx2_ASAP7_75t_L g6005 ( 
.A(n_5408),
.Y(n_6005)
);

INVx1_ASAP7_75t_L g6006 ( 
.A(n_5442),
.Y(n_6006)
);

INVx4_ASAP7_75t_L g6007 ( 
.A(n_5257),
.Y(n_6007)
);

INVx1_ASAP7_75t_L g6008 ( 
.A(n_5444),
.Y(n_6008)
);

NOR2xp33_ASAP7_75t_L g6009 ( 
.A(n_5418),
.B(n_2650),
.Y(n_6009)
);

INVx4_ASAP7_75t_L g6010 ( 
.A(n_5266),
.Y(n_6010)
);

CKINVDCx14_ASAP7_75t_R g6011 ( 
.A(n_5280),
.Y(n_6011)
);

AO22x2_ASAP7_75t_L g6012 ( 
.A1(n_5267),
.A2(n_3418),
.B1(n_3429),
.B2(n_3424),
.Y(n_6012)
);

INVx1_ASAP7_75t_L g6013 ( 
.A(n_5447),
.Y(n_6013)
);

AND2x4_ASAP7_75t_L g6014 ( 
.A(n_5641),
.B(n_5648),
.Y(n_6014)
);

INVx3_ASAP7_75t_L g6015 ( 
.A(n_5279),
.Y(n_6015)
);

AND2x6_ASAP7_75t_L g6016 ( 
.A(n_5629),
.B(n_3430),
.Y(n_6016)
);

INVx1_ASAP7_75t_L g6017 ( 
.A(n_5448),
.Y(n_6017)
);

AND2x2_ASAP7_75t_L g6018 ( 
.A(n_5528),
.B(n_3163),
.Y(n_6018)
);

AND2x2_ASAP7_75t_L g6019 ( 
.A(n_5443),
.B(n_3173),
.Y(n_6019)
);

AOI22xp33_ASAP7_75t_L g6020 ( 
.A1(n_5515),
.A2(n_3437),
.B1(n_3440),
.B2(n_3434),
.Y(n_6020)
);

AOI21x1_ASAP7_75t_L g6021 ( 
.A1(n_5181),
.A2(n_3448),
.B(n_3442),
.Y(n_6021)
);

OR2x6_ASAP7_75t_L g6022 ( 
.A(n_5630),
.B(n_3450),
.Y(n_6022)
);

INVx2_ASAP7_75t_L g6023 ( 
.A(n_5475),
.Y(n_6023)
);

NAND3xp33_ASAP7_75t_L g6024 ( 
.A(n_5465),
.B(n_2654),
.C(n_2651),
.Y(n_6024)
);

INVx2_ASAP7_75t_SL g6025 ( 
.A(n_5495),
.Y(n_6025)
);

CKINVDCx5p33_ASAP7_75t_R g6026 ( 
.A(n_5586),
.Y(n_6026)
);

AND2x6_ASAP7_75t_L g6027 ( 
.A(n_5647),
.B(n_5478),
.Y(n_6027)
);

AND2x4_ASAP7_75t_L g6028 ( 
.A(n_5294),
.B(n_3457),
.Y(n_6028)
);

INVx2_ASAP7_75t_L g6029 ( 
.A(n_5486),
.Y(n_6029)
);

INVx1_ASAP7_75t_L g6030 ( 
.A(n_5490),
.Y(n_6030)
);

INVx2_ASAP7_75t_L g6031 ( 
.A(n_5493),
.Y(n_6031)
);

BUFx3_ASAP7_75t_L g6032 ( 
.A(n_5343),
.Y(n_6032)
);

INVx4_ASAP7_75t_L g6033 ( 
.A(n_5349),
.Y(n_6033)
);

AND2x4_ASAP7_75t_L g6034 ( 
.A(n_5364),
.B(n_3464),
.Y(n_6034)
);

NOR2xp33_ASAP7_75t_L g6035 ( 
.A(n_5472),
.B(n_2658),
.Y(n_6035)
);

NAND2xp5_ASAP7_75t_L g6036 ( 
.A(n_5385),
.B(n_2661),
.Y(n_6036)
);

NOR2xp33_ASAP7_75t_L g6037 ( 
.A(n_5473),
.B(n_2666),
.Y(n_6037)
);

AND2x2_ASAP7_75t_L g6038 ( 
.A(n_5571),
.B(n_3181),
.Y(n_6038)
);

BUFx3_ASAP7_75t_L g6039 ( 
.A(n_5393),
.Y(n_6039)
);

AND2x2_ASAP7_75t_L g6040 ( 
.A(n_5270),
.B(n_3188),
.Y(n_6040)
);

INVx1_ASAP7_75t_L g6041 ( 
.A(n_5496),
.Y(n_6041)
);

OR2x2_ASAP7_75t_L g6042 ( 
.A(n_5344),
.B(n_3192),
.Y(n_6042)
);

INVx4_ASAP7_75t_L g6043 ( 
.A(n_5410),
.Y(n_6043)
);

INVx5_ASAP7_75t_L g6044 ( 
.A(n_5135),
.Y(n_6044)
);

AND2x2_ASAP7_75t_L g6045 ( 
.A(n_5272),
.B(n_3195),
.Y(n_6045)
);

NAND2xp5_ASAP7_75t_L g6046 ( 
.A(n_5386),
.B(n_2673),
.Y(n_6046)
);

BUFx2_ASAP7_75t_L g6047 ( 
.A(n_5451),
.Y(n_6047)
);

BUFx6f_ASAP7_75t_L g6048 ( 
.A(n_5446),
.Y(n_6048)
);

BUFx6f_ASAP7_75t_L g6049 ( 
.A(n_5450),
.Y(n_6049)
);

INVx2_ASAP7_75t_L g6050 ( 
.A(n_5498),
.Y(n_6050)
);

CKINVDCx5p33_ASAP7_75t_R g6051 ( 
.A(n_5614),
.Y(n_6051)
);

INVx1_ASAP7_75t_L g6052 ( 
.A(n_5512),
.Y(n_6052)
);

NOR2x1p5_ASAP7_75t_L g6053 ( 
.A(n_5650),
.B(n_5492),
.Y(n_6053)
);

OR2x2_ASAP7_75t_L g6054 ( 
.A(n_5291),
.B(n_3204),
.Y(n_6054)
);

INVx1_ASAP7_75t_L g6055 ( 
.A(n_5516),
.Y(n_6055)
);

BUFx2_ASAP7_75t_L g6056 ( 
.A(n_5523),
.Y(n_6056)
);

INVx2_ASAP7_75t_SL g6057 ( 
.A(n_5482),
.Y(n_6057)
);

INVx1_ASAP7_75t_L g6058 ( 
.A(n_5548),
.Y(n_6058)
);

AND2x4_ASAP7_75t_L g6059 ( 
.A(n_5484),
.B(n_5510),
.Y(n_6059)
);

NAND2xp5_ASAP7_75t_SL g6060 ( 
.A(n_5502),
.B(n_2677),
.Y(n_6060)
);

INVx4_ASAP7_75t_SL g6061 ( 
.A(n_5135),
.Y(n_6061)
);

AND2x2_ASAP7_75t_L g6062 ( 
.A(n_5546),
.B(n_5407),
.Y(n_6062)
);

INVx3_ASAP7_75t_L g6063 ( 
.A(n_5539),
.Y(n_6063)
);

INVx1_ASAP7_75t_L g6064 ( 
.A(n_5552),
.Y(n_6064)
);

INVx1_ASAP7_75t_L g6065 ( 
.A(n_5553),
.Y(n_6065)
);

BUFx2_ASAP7_75t_L g6066 ( 
.A(n_5541),
.Y(n_6066)
);

INVx1_ASAP7_75t_L g6067 ( 
.A(n_5557),
.Y(n_6067)
);

INVx2_ASAP7_75t_L g6068 ( 
.A(n_5513),
.Y(n_6068)
);

OR2x6_ASAP7_75t_L g6069 ( 
.A(n_5276),
.B(n_3475),
.Y(n_6069)
);

AOI22xp5_ASAP7_75t_L g6070 ( 
.A1(n_5362),
.A2(n_5471),
.B1(n_5520),
.B2(n_5518),
.Y(n_6070)
);

INVx1_ASAP7_75t_L g6071 ( 
.A(n_5521),
.Y(n_6071)
);

INVx1_ASAP7_75t_L g6072 ( 
.A(n_5560),
.Y(n_6072)
);

INVx1_ASAP7_75t_L g6073 ( 
.A(n_5563),
.Y(n_6073)
);

INVx1_ASAP7_75t_L g6074 ( 
.A(n_5570),
.Y(n_6074)
);

BUFx2_ASAP7_75t_L g6075 ( 
.A(n_5575),
.Y(n_6075)
);

AND2x4_ASAP7_75t_L g6076 ( 
.A(n_5581),
.B(n_3487),
.Y(n_6076)
);

INVx2_ASAP7_75t_L g6077 ( 
.A(n_5538),
.Y(n_6077)
);

INVx4_ASAP7_75t_L g6078 ( 
.A(n_5587),
.Y(n_6078)
);

INVx1_ASAP7_75t_L g6079 ( 
.A(n_5573),
.Y(n_6079)
);

BUFx6f_ASAP7_75t_L g6080 ( 
.A(n_5598),
.Y(n_6080)
);

INVx1_ASAP7_75t_L g6081 ( 
.A(n_5576),
.Y(n_6081)
);

NAND2xp5_ASAP7_75t_L g6082 ( 
.A(n_5390),
.B(n_2679),
.Y(n_6082)
);

NAND2x1p5_ASAP7_75t_L g6083 ( 
.A(n_5620),
.B(n_3493),
.Y(n_6083)
);

BUFx6f_ASAP7_75t_L g6084 ( 
.A(n_5632),
.Y(n_6084)
);

INVx8_ASAP7_75t_L g6085 ( 
.A(n_5276),
.Y(n_6085)
);

INVx1_ASAP7_75t_L g6086 ( 
.A(n_5582),
.Y(n_6086)
);

INVx2_ASAP7_75t_L g6087 ( 
.A(n_5542),
.Y(n_6087)
);

INVx2_ASAP7_75t_L g6088 ( 
.A(n_5549),
.Y(n_6088)
);

BUFx6f_ASAP7_75t_L g6089 ( 
.A(n_5633),
.Y(n_6089)
);

BUFx3_ASAP7_75t_L g6090 ( 
.A(n_5627),
.Y(n_6090)
);

AND2x6_ASAP7_75t_L g6091 ( 
.A(n_5589),
.B(n_3495),
.Y(n_6091)
);

NOR2xp33_ASAP7_75t_L g6092 ( 
.A(n_5231),
.B(n_2685),
.Y(n_6092)
);

NAND2xp5_ASAP7_75t_L g6093 ( 
.A(n_5556),
.B(n_2688),
.Y(n_6093)
);

INVx4_ASAP7_75t_L g6094 ( 
.A(n_5428),
.Y(n_6094)
);

INVx2_ASAP7_75t_L g6095 ( 
.A(n_5555),
.Y(n_6095)
);

INVx5_ASAP7_75t_L g6096 ( 
.A(n_5428),
.Y(n_6096)
);

INVx1_ASAP7_75t_L g6097 ( 
.A(n_5590),
.Y(n_6097)
);

AND2x4_ASAP7_75t_L g6098 ( 
.A(n_5583),
.B(n_3501),
.Y(n_6098)
);

INVx1_ASAP7_75t_L g6099 ( 
.A(n_5592),
.Y(n_6099)
);

INVx1_ASAP7_75t_SL g6100 ( 
.A(n_5619),
.Y(n_6100)
);

INVx1_ASAP7_75t_L g6101 ( 
.A(n_5595),
.Y(n_6101)
);

NAND2xp5_ASAP7_75t_L g6102 ( 
.A(n_5566),
.B(n_2700),
.Y(n_6102)
);

O2A1O1Ixp33_ASAP7_75t_L g6103 ( 
.A1(n_5211),
.A2(n_5243),
.B(n_5351),
.C(n_5347),
.Y(n_6103)
);

INVxp67_ASAP7_75t_SL g6104 ( 
.A(n_5464),
.Y(n_6104)
);

NAND2xp5_ASAP7_75t_SL g6105 ( 
.A(n_5578),
.B(n_5505),
.Y(n_6105)
);

INVx3_ASAP7_75t_L g6106 ( 
.A(n_5525),
.Y(n_6106)
);

AO22x2_ASAP7_75t_L g6107 ( 
.A1(n_5599),
.A2(n_3511),
.B1(n_3524),
.B2(n_3522),
.Y(n_6107)
);

INVxp67_ASAP7_75t_L g6108 ( 
.A(n_5397),
.Y(n_6108)
);

NOR2xp33_ASAP7_75t_L g6109 ( 
.A(n_5649),
.B(n_2701),
.Y(n_6109)
);

INVx1_ASAP7_75t_L g6110 ( 
.A(n_5597),
.Y(n_6110)
);

NAND2xp5_ASAP7_75t_L g6111 ( 
.A(n_5199),
.B(n_5212),
.Y(n_6111)
);

NAND3x1_ASAP7_75t_L g6112 ( 
.A(n_5378),
.B(n_3536),
.C(n_3530),
.Y(n_6112)
);

INVx1_ASAP7_75t_L g6113 ( 
.A(n_5564),
.Y(n_6113)
);

INVx3_ASAP7_75t_L g6114 ( 
.A(n_5531),
.Y(n_6114)
);

INVx1_ASAP7_75t_L g6115 ( 
.A(n_5565),
.Y(n_6115)
);

NAND2xp5_ASAP7_75t_L g6116 ( 
.A(n_5646),
.B(n_2702),
.Y(n_6116)
);

NAND2xp5_ASAP7_75t_SL g6117 ( 
.A(n_5288),
.B(n_2704),
.Y(n_6117)
);

INVx1_ASAP7_75t_L g6118 ( 
.A(n_5568),
.Y(n_6118)
);

BUFx6f_ASAP7_75t_L g6119 ( 
.A(n_5653),
.Y(n_6119)
);

BUFx6f_ASAP7_75t_L g6120 ( 
.A(n_5600),
.Y(n_6120)
);

INVx4_ASAP7_75t_SL g6121 ( 
.A(n_5631),
.Y(n_6121)
);

INVx3_ASAP7_75t_L g6122 ( 
.A(n_5533),
.Y(n_6122)
);

AND2x4_ASAP7_75t_L g6123 ( 
.A(n_5602),
.B(n_3538),
.Y(n_6123)
);

INVx1_ASAP7_75t_L g6124 ( 
.A(n_5577),
.Y(n_6124)
);

NAND2xp5_ASAP7_75t_L g6125 ( 
.A(n_5323),
.B(n_2705),
.Y(n_6125)
);

BUFx3_ASAP7_75t_L g6126 ( 
.A(n_5637),
.Y(n_6126)
);

INVx2_ASAP7_75t_SL g6127 ( 
.A(n_5605),
.Y(n_6127)
);

INVx2_ASAP7_75t_L g6128 ( 
.A(n_5606),
.Y(n_6128)
);

NAND3x1_ASAP7_75t_L g6129 ( 
.A(n_5550),
.B(n_3559),
.C(n_3557),
.Y(n_6129)
);

AOI22xp5_ASAP7_75t_L g6130 ( 
.A1(n_5468),
.A2(n_2707),
.B1(n_2710),
.B2(n_2706),
.Y(n_6130)
);

OAI22xp5_ASAP7_75t_SL g6131 ( 
.A1(n_5544),
.A2(n_3208),
.B1(n_3210),
.B2(n_3206),
.Y(n_6131)
);

INVx1_ASAP7_75t_L g6132 ( 
.A(n_5607),
.Y(n_6132)
);

INVx4_ASAP7_75t_L g6133 ( 
.A(n_5479),
.Y(n_6133)
);

INVx1_ASAP7_75t_L g6134 ( 
.A(n_5608),
.Y(n_6134)
);

INVx2_ASAP7_75t_L g6135 ( 
.A(n_5609),
.Y(n_6135)
);

INVx2_ASAP7_75t_SL g6136 ( 
.A(n_5611),
.Y(n_6136)
);

INVx1_ASAP7_75t_L g6137 ( 
.A(n_5615),
.Y(n_6137)
);

NAND2xp5_ASAP7_75t_L g6138 ( 
.A(n_5455),
.B(n_2715),
.Y(n_6138)
);

BUFx6f_ASAP7_75t_L g6139 ( 
.A(n_5618),
.Y(n_6139)
);

INVx1_ASAP7_75t_L g6140 ( 
.A(n_5251),
.Y(n_6140)
);

BUFx6f_ASAP7_75t_L g6141 ( 
.A(n_5638),
.Y(n_6141)
);

AND2x4_ASAP7_75t_L g6142 ( 
.A(n_5258),
.B(n_5639),
.Y(n_6142)
);

INVx2_ASAP7_75t_L g6143 ( 
.A(n_5535),
.Y(n_6143)
);

AND2x4_ASAP7_75t_L g6144 ( 
.A(n_5536),
.B(n_3560),
.Y(n_6144)
);

NAND2xp5_ASAP7_75t_SL g6145 ( 
.A(n_5391),
.B(n_2716),
.Y(n_6145)
);

INVx1_ASAP7_75t_L g6146 ( 
.A(n_5540),
.Y(n_6146)
);

AND2x4_ASAP7_75t_L g6147 ( 
.A(n_5545),
.B(n_3566),
.Y(n_6147)
);

OR2x2_ASAP7_75t_L g6148 ( 
.A(n_5567),
.B(n_3225),
.Y(n_6148)
);

INVx2_ASAP7_75t_L g6149 ( 
.A(n_5289),
.Y(n_6149)
);

BUFx6f_ASAP7_75t_L g6150 ( 
.A(n_5613),
.Y(n_6150)
);

INVx2_ASAP7_75t_SL g6151 ( 
.A(n_5261),
.Y(n_6151)
);

AND2x6_ASAP7_75t_L g6152 ( 
.A(n_5654),
.B(n_3568),
.Y(n_6152)
);

NAND2xp5_ASAP7_75t_L g6153 ( 
.A(n_5554),
.B(n_5399),
.Y(n_6153)
);

INVx1_ASAP7_75t_L g6154 ( 
.A(n_5460),
.Y(n_6154)
);

NAND2xp5_ASAP7_75t_L g6155 ( 
.A(n_5524),
.B(n_2723),
.Y(n_6155)
);

INVxp67_ASAP7_75t_L g6156 ( 
.A(n_5634),
.Y(n_6156)
);

INVxp33_ASAP7_75t_L g6157 ( 
.A(n_5463),
.Y(n_6157)
);

AND2x4_ASAP7_75t_L g6158 ( 
.A(n_5292),
.B(n_3588),
.Y(n_6158)
);

AND2x4_ASAP7_75t_L g6159 ( 
.A(n_5526),
.B(n_3596),
.Y(n_6159)
);

NAND2x1p5_ASAP7_75t_L g6160 ( 
.A(n_5315),
.B(n_3612),
.Y(n_6160)
);

INVx2_ASAP7_75t_L g6161 ( 
.A(n_5215),
.Y(n_6161)
);

INVx1_ASAP7_75t_L g6162 ( 
.A(n_5338),
.Y(n_6162)
);

BUFx6f_ASAP7_75t_L g6163 ( 
.A(n_5166),
.Y(n_6163)
);

INVx2_ASAP7_75t_L g6164 ( 
.A(n_5422),
.Y(n_6164)
);

INVx1_ASAP7_75t_L g6165 ( 
.A(n_5432),
.Y(n_6165)
);

INVx1_ASAP7_75t_L g6166 ( 
.A(n_5438),
.Y(n_6166)
);

HB1xp67_ASAP7_75t_L g6167 ( 
.A(n_5466),
.Y(n_6167)
);

INVx1_ASAP7_75t_L g6168 ( 
.A(n_5488),
.Y(n_6168)
);

NAND2xp5_ASAP7_75t_L g6169 ( 
.A(n_5375),
.B(n_2735),
.Y(n_6169)
);

BUFx3_ASAP7_75t_L g6170 ( 
.A(n_5616),
.Y(n_6170)
);

INVx4_ASAP7_75t_L g6171 ( 
.A(n_5269),
.Y(n_6171)
);

AOI22xp5_ASAP7_75t_L g6172 ( 
.A1(n_5494),
.A2(n_5636),
.B1(n_5415),
.B2(n_5254),
.Y(n_6172)
);

AND2x2_ASAP7_75t_SL g6173 ( 
.A(n_5596),
.B(n_3614),
.Y(n_6173)
);

INVx1_ASAP7_75t_L g6174 ( 
.A(n_5379),
.Y(n_6174)
);

INVx1_ASAP7_75t_L g6175 ( 
.A(n_5384),
.Y(n_6175)
);

AND2x2_ASAP7_75t_L g6176 ( 
.A(n_5628),
.B(n_3237),
.Y(n_6176)
);

AO22x2_ASAP7_75t_L g6177 ( 
.A1(n_5551),
.A2(n_3616),
.B1(n_3623),
.B2(n_5167),
.Y(n_6177)
);

BUFx3_ASAP7_75t_L g6178 ( 
.A(n_5389),
.Y(n_6178)
);

OR2x6_ASAP7_75t_L g6179 ( 
.A(n_5594),
.B(n_3196),
.Y(n_6179)
);

INVx4_ASAP7_75t_L g6180 ( 
.A(n_5603),
.Y(n_6180)
);

AND2x2_ASAP7_75t_L g6181 ( 
.A(n_5543),
.B(n_3238),
.Y(n_6181)
);

INVx2_ASAP7_75t_L g6182 ( 
.A(n_5437),
.Y(n_6182)
);

AND2x4_ASAP7_75t_L g6183 ( 
.A(n_5501),
.B(n_3245),
.Y(n_6183)
);

BUFx6f_ASAP7_75t_L g6184 ( 
.A(n_5644),
.Y(n_6184)
);

AND2x4_ASAP7_75t_L g6185 ( 
.A(n_5458),
.B(n_3251),
.Y(n_6185)
);

CKINVDCx5p33_ASAP7_75t_R g6186 ( 
.A(n_5137),
.Y(n_6186)
);

NAND2xp5_ASAP7_75t_SL g6187 ( 
.A(n_5193),
.B(n_2737),
.Y(n_6187)
);

AO22x2_ASAP7_75t_L g6188 ( 
.A1(n_5152),
.A2(n_4),
.B1(n_2),
.B2(n_3),
.Y(n_6188)
);

NOR2x1p5_ASAP7_75t_L g6189 ( 
.A(n_5872),
.B(n_3255),
.Y(n_6189)
);

INVx1_ASAP7_75t_L g6190 ( 
.A(n_5660),
.Y(n_6190)
);

AO221x1_ASAP7_75t_L g6191 ( 
.A1(n_6188),
.A2(n_3265),
.B1(n_3274),
.B2(n_3261),
.C(n_3256),
.Y(n_6191)
);

OAI22xp5_ASAP7_75t_L g6192 ( 
.A1(n_5669),
.A2(n_2740),
.B1(n_2741),
.B2(n_2738),
.Y(n_6192)
);

INVx1_ASAP7_75t_L g6193 ( 
.A(n_5662),
.Y(n_6193)
);

INVx2_ASAP7_75t_SL g6194 ( 
.A(n_5675),
.Y(n_6194)
);

NAND2xp5_ASAP7_75t_L g6195 ( 
.A(n_5957),
.B(n_2742),
.Y(n_6195)
);

INVx1_ASAP7_75t_L g6196 ( 
.A(n_5663),
.Y(n_6196)
);

NAND2xp5_ASAP7_75t_L g6197 ( 
.A(n_5661),
.B(n_2744),
.Y(n_6197)
);

NAND2xp5_ASAP7_75t_L g6198 ( 
.A(n_5812),
.B(n_2746),
.Y(n_6198)
);

INVx2_ASAP7_75t_SL g6199 ( 
.A(n_5675),
.Y(n_6199)
);

NAND2xp5_ASAP7_75t_L g6200 ( 
.A(n_5735),
.B(n_2748),
.Y(n_6200)
);

INVx2_ASAP7_75t_L g6201 ( 
.A(n_5703),
.Y(n_6201)
);

NAND2xp5_ASAP7_75t_L g6202 ( 
.A(n_5697),
.B(n_2749),
.Y(n_6202)
);

NOR2xp33_ASAP7_75t_L g6203 ( 
.A(n_5863),
.B(n_2752),
.Y(n_6203)
);

AOI22xp33_ASAP7_75t_L g6204 ( 
.A1(n_6182),
.A2(n_2755),
.B1(n_2760),
.B2(n_2753),
.Y(n_6204)
);

OAI21xp5_ASAP7_75t_L g6205 ( 
.A1(n_5668),
.A2(n_2767),
.B(n_2765),
.Y(n_6205)
);

NAND2xp5_ASAP7_75t_SL g6206 ( 
.A(n_5724),
.B(n_2769),
.Y(n_6206)
);

NOR2xp33_ASAP7_75t_L g6207 ( 
.A(n_6009),
.B(n_2775),
.Y(n_6207)
);

NAND2xp5_ASAP7_75t_L g6208 ( 
.A(n_5869),
.B(n_2777),
.Y(n_6208)
);

INVx2_ASAP7_75t_L g6209 ( 
.A(n_5710),
.Y(n_6209)
);

NAND2xp5_ASAP7_75t_L g6210 ( 
.A(n_6035),
.B(n_2780),
.Y(n_6210)
);

BUFx6f_ASAP7_75t_SL g6211 ( 
.A(n_5717),
.Y(n_6211)
);

INVx1_ASAP7_75t_L g6212 ( 
.A(n_5666),
.Y(n_6212)
);

NAND2xp5_ASAP7_75t_L g6213 ( 
.A(n_6037),
.B(n_2793),
.Y(n_6213)
);

NAND2xp5_ASAP7_75t_L g6214 ( 
.A(n_5763),
.B(n_2795),
.Y(n_6214)
);

NOR2xp33_ASAP7_75t_L g6215 ( 
.A(n_5730),
.B(n_2801),
.Y(n_6215)
);

INVx2_ASAP7_75t_L g6216 ( 
.A(n_5712),
.Y(n_6216)
);

NOR2xp67_ASAP7_75t_L g6217 ( 
.A(n_5897),
.B(n_3275),
.Y(n_6217)
);

NAND2xp5_ASAP7_75t_SL g6218 ( 
.A(n_5938),
.B(n_2803),
.Y(n_6218)
);

NAND2xp5_ASAP7_75t_L g6219 ( 
.A(n_5761),
.B(n_2805),
.Y(n_6219)
);

NAND2xp5_ASAP7_75t_SL g6220 ( 
.A(n_5787),
.B(n_6100),
.Y(n_6220)
);

HB1xp67_ASAP7_75t_L g6221 ( 
.A(n_5678),
.Y(n_6221)
);

NAND2xp5_ASAP7_75t_L g6222 ( 
.A(n_5876),
.B(n_2811),
.Y(n_6222)
);

INVx4_ASAP7_75t_L g6223 ( 
.A(n_5768),
.Y(n_6223)
);

NAND2xp5_ASAP7_75t_SL g6224 ( 
.A(n_5684),
.B(n_2816),
.Y(n_6224)
);

INVx2_ASAP7_75t_L g6225 ( 
.A(n_5719),
.Y(n_6225)
);

OR2x6_ASAP7_75t_L g6226 ( 
.A(n_5741),
.B(n_5798),
.Y(n_6226)
);

OR2x6_ASAP7_75t_L g6227 ( 
.A(n_5835),
.B(n_1047),
.Y(n_6227)
);

NOR2xp33_ASAP7_75t_L g6228 ( 
.A(n_5683),
.B(n_2822),
.Y(n_6228)
);

OAI22xp5_ASAP7_75t_L g6229 ( 
.A1(n_6111),
.A2(n_2830),
.B1(n_2831),
.B2(n_2827),
.Y(n_6229)
);

A2O1A1Ixp33_ASAP7_75t_L g6230 ( 
.A1(n_6103),
.A2(n_5838),
.B(n_5840),
.C(n_5959),
.Y(n_6230)
);

NAND2xp5_ASAP7_75t_L g6231 ( 
.A(n_5853),
.B(n_2833),
.Y(n_6231)
);

NAND2xp5_ASAP7_75t_L g6232 ( 
.A(n_5862),
.B(n_5894),
.Y(n_6232)
);

NAND2xp5_ASAP7_75t_L g6233 ( 
.A(n_5905),
.B(n_5949),
.Y(n_6233)
);

INVx1_ASAP7_75t_L g6234 ( 
.A(n_5667),
.Y(n_6234)
);

INVx1_ASAP7_75t_L g6235 ( 
.A(n_5672),
.Y(n_6235)
);

INVx1_ASAP7_75t_L g6236 ( 
.A(n_5674),
.Y(n_6236)
);

INVx2_ASAP7_75t_SL g6237 ( 
.A(n_5768),
.Y(n_6237)
);

AND2x4_ASAP7_75t_L g6238 ( 
.A(n_5799),
.B(n_3276),
.Y(n_6238)
);

AOI22x1_ASAP7_75t_L g6239 ( 
.A1(n_5899),
.A2(n_3280),
.B1(n_3283),
.B2(n_3279),
.Y(n_6239)
);

AOI22xp5_ASAP7_75t_L g6240 ( 
.A1(n_6062),
.A2(n_2836),
.B1(n_2839),
.B2(n_2834),
.Y(n_6240)
);

OR2x2_ASAP7_75t_L g6241 ( 
.A(n_5698),
.B(n_3284),
.Y(n_6241)
);

INVx5_ASAP7_75t_L g6242 ( 
.A(n_6184),
.Y(n_6242)
);

O2A1O1Ixp5_ASAP7_75t_L g6243 ( 
.A1(n_6105),
.A2(n_3291),
.B(n_3298),
.C(n_3290),
.Y(n_6243)
);

AOI22xp5_ASAP7_75t_L g6244 ( 
.A1(n_5691),
.A2(n_2859),
.B1(n_2860),
.B2(n_2857),
.Y(n_6244)
);

INVx1_ASAP7_75t_L g6245 ( 
.A(n_5676),
.Y(n_6245)
);

AOI22xp33_ASAP7_75t_L g6246 ( 
.A1(n_6173),
.A2(n_2868),
.B1(n_2878),
.B2(n_2864),
.Y(n_6246)
);

NAND2xp5_ASAP7_75t_SL g6247 ( 
.A(n_5696),
.B(n_2880),
.Y(n_6247)
);

NAND2xp5_ASAP7_75t_L g6248 ( 
.A(n_6018),
.B(n_2881),
.Y(n_6248)
);

OR2x6_ASAP7_75t_L g6249 ( 
.A(n_6085),
.B(n_1047),
.Y(n_6249)
);

NAND2xp5_ASAP7_75t_L g6250 ( 
.A(n_6019),
.B(n_2886),
.Y(n_6250)
);

INVx1_ASAP7_75t_L g6251 ( 
.A(n_5679),
.Y(n_6251)
);

O2A1O1Ixp33_ASAP7_75t_L g6252 ( 
.A1(n_6187),
.A2(n_5706),
.B(n_5818),
.C(n_6167),
.Y(n_6252)
);

OAI22xp5_ASAP7_75t_L g6253 ( 
.A1(n_6171),
.A2(n_2895),
.B1(n_2901),
.B2(n_2887),
.Y(n_6253)
);

NAND2xp5_ASAP7_75t_L g6254 ( 
.A(n_5866),
.B(n_5681),
.Y(n_6254)
);

AOI22xp33_ASAP7_75t_L g6255 ( 
.A1(n_6181),
.A2(n_2905),
.B1(n_2906),
.B2(n_2903),
.Y(n_6255)
);

NAND2xp5_ASAP7_75t_L g6256 ( 
.A(n_5686),
.B(n_2908),
.Y(n_6256)
);

NAND2xp5_ASAP7_75t_L g6257 ( 
.A(n_5687),
.B(n_2910),
.Y(n_6257)
);

OR2x2_ASAP7_75t_L g6258 ( 
.A(n_5699),
.B(n_3306),
.Y(n_6258)
);

INVx1_ASAP7_75t_L g6259 ( 
.A(n_5702),
.Y(n_6259)
);

NAND2x1_ASAP7_75t_L g6260 ( 
.A(n_5851),
.B(n_1048),
.Y(n_6260)
);

NOR2xp33_ASAP7_75t_L g6261 ( 
.A(n_5705),
.B(n_2918),
.Y(n_6261)
);

OR2x2_ASAP7_75t_L g6262 ( 
.A(n_5736),
.B(n_3312),
.Y(n_6262)
);

INVx1_ASAP7_75t_L g6263 ( 
.A(n_5704),
.Y(n_6263)
);

NAND2xp5_ASAP7_75t_L g6264 ( 
.A(n_5707),
.B(n_2921),
.Y(n_6264)
);

INVx2_ASAP7_75t_SL g6265 ( 
.A(n_6184),
.Y(n_6265)
);

NAND2xp5_ASAP7_75t_L g6266 ( 
.A(n_5714),
.B(n_2923),
.Y(n_6266)
);

INVx2_ASAP7_75t_L g6267 ( 
.A(n_5742),
.Y(n_6267)
);

NAND3xp33_ASAP7_75t_SL g6268 ( 
.A(n_5996),
.B(n_3319),
.C(n_3313),
.Y(n_6268)
);

A2O1A1Ixp33_ASAP7_75t_L g6269 ( 
.A1(n_6092),
.A2(n_3340),
.B(n_3343),
.C(n_3328),
.Y(n_6269)
);

INVx2_ASAP7_75t_L g6270 ( 
.A(n_5744),
.Y(n_6270)
);

NOR2xp33_ASAP7_75t_L g6271 ( 
.A(n_5711),
.B(n_2924),
.Y(n_6271)
);

INVx2_ASAP7_75t_L g6272 ( 
.A(n_5751),
.Y(n_6272)
);

INVx1_ASAP7_75t_L g6273 ( 
.A(n_5720),
.Y(n_6273)
);

NAND2xp5_ASAP7_75t_SL g6274 ( 
.A(n_5695),
.B(n_2925),
.Y(n_6274)
);

NAND2xp5_ASAP7_75t_SL g6275 ( 
.A(n_5734),
.B(n_2928),
.Y(n_6275)
);

INVxp67_ASAP7_75t_SL g6276 ( 
.A(n_5955),
.Y(n_6276)
);

NOR2x1p5_ASAP7_75t_L g6277 ( 
.A(n_5694),
.B(n_3344),
.Y(n_6277)
);

INVx2_ASAP7_75t_SL g6278 ( 
.A(n_5685),
.Y(n_6278)
);

BUFx6f_ASAP7_75t_L g6279 ( 
.A(n_5670),
.Y(n_6279)
);

INVx1_ASAP7_75t_L g6280 ( 
.A(n_5725),
.Y(n_6280)
);

NAND2xp5_ASAP7_75t_L g6281 ( 
.A(n_5728),
.B(n_2930),
.Y(n_6281)
);

NOR2xp33_ASAP7_75t_L g6282 ( 
.A(n_6026),
.B(n_2931),
.Y(n_6282)
);

AOI21xp5_ASAP7_75t_L g6283 ( 
.A1(n_6149),
.A2(n_2936),
.B(n_2933),
.Y(n_6283)
);

BUFx3_ASAP7_75t_L g6284 ( 
.A(n_5839),
.Y(n_6284)
);

AND2x4_ASAP7_75t_L g6285 ( 
.A(n_5700),
.B(n_3346),
.Y(n_6285)
);

NAND2xp5_ASAP7_75t_L g6286 ( 
.A(n_5732),
.B(n_2938),
.Y(n_6286)
);

A2O1A1Ixp33_ASAP7_75t_SL g6287 ( 
.A1(n_6109),
.A2(n_5743),
.B(n_5690),
.C(n_6011),
.Y(n_6287)
);

NOR2xp33_ASAP7_75t_L g6288 ( 
.A(n_5988),
.B(n_2940),
.Y(n_6288)
);

NAND2xp5_ASAP7_75t_L g6289 ( 
.A(n_5746),
.B(n_2945),
.Y(n_6289)
);

INVx2_ASAP7_75t_SL g6290 ( 
.A(n_5758),
.Y(n_6290)
);

BUFx3_ASAP7_75t_L g6291 ( 
.A(n_5688),
.Y(n_6291)
);

NOR2xp33_ASAP7_75t_L g6292 ( 
.A(n_5740),
.B(n_2948),
.Y(n_6292)
);

NAND2xp5_ASAP7_75t_L g6293 ( 
.A(n_5748),
.B(n_2949),
.Y(n_6293)
);

INVx2_ASAP7_75t_L g6294 ( 
.A(n_5759),
.Y(n_6294)
);

O2A1O1Ixp5_ASAP7_75t_L g6295 ( 
.A1(n_6154),
.A2(n_3354),
.B(n_3356),
.C(n_3349),
.Y(n_6295)
);

NAND2xp5_ASAP7_75t_L g6296 ( 
.A(n_5753),
.B(n_5754),
.Y(n_6296)
);

NOR2xp33_ASAP7_75t_L g6297 ( 
.A(n_5925),
.B(n_2956),
.Y(n_6297)
);

NAND2xp5_ASAP7_75t_L g6298 ( 
.A(n_5756),
.B(n_2958),
.Y(n_6298)
);

NAND2xp5_ASAP7_75t_SL g6299 ( 
.A(n_6180),
.B(n_2959),
.Y(n_6299)
);

INVx1_ASAP7_75t_L g6300 ( 
.A(n_5757),
.Y(n_6300)
);

NAND2xp5_ASAP7_75t_L g6301 ( 
.A(n_5760),
.B(n_2964),
.Y(n_6301)
);

INVx4_ASAP7_75t_L g6302 ( 
.A(n_5880),
.Y(n_6302)
);

NAND2xp5_ASAP7_75t_L g6303 ( 
.A(n_5771),
.B(n_2967),
.Y(n_6303)
);

CKINVDCx5p33_ASAP7_75t_R g6304 ( 
.A(n_5673),
.Y(n_6304)
);

NAND2xp5_ASAP7_75t_L g6305 ( 
.A(n_5779),
.B(n_2969),
.Y(n_6305)
);

INVxp67_ASAP7_75t_L g6306 ( 
.A(n_5737),
.Y(n_6306)
);

INVx1_ASAP7_75t_L g6307 ( 
.A(n_5804),
.Y(n_6307)
);

OAI22xp33_ASAP7_75t_L g6308 ( 
.A1(n_5750),
.A2(n_3364),
.B1(n_3365),
.B2(n_3361),
.Y(n_6308)
);

AND2x4_ASAP7_75t_L g6309 ( 
.A(n_5738),
.B(n_3370),
.Y(n_6309)
);

NAND2xp5_ASAP7_75t_SL g6310 ( 
.A(n_5870),
.B(n_2972),
.Y(n_6310)
);

NAND2xp5_ASAP7_75t_L g6311 ( 
.A(n_5806),
.B(n_2974),
.Y(n_6311)
);

INVx2_ASAP7_75t_L g6312 ( 
.A(n_5766),
.Y(n_6312)
);

AOI22xp5_ASAP7_75t_L g6313 ( 
.A1(n_6151),
.A2(n_2977),
.B1(n_2981),
.B2(n_2976),
.Y(n_6313)
);

AOI221xp5_ASAP7_75t_L g6314 ( 
.A1(n_5795),
.A2(n_3387),
.B1(n_3393),
.B2(n_3380),
.C(n_3374),
.Y(n_6314)
);

INVx2_ASAP7_75t_L g6315 ( 
.A(n_5770),
.Y(n_6315)
);

INVx1_ASAP7_75t_L g6316 ( 
.A(n_5808),
.Y(n_6316)
);

AOI22xp33_ASAP7_75t_L g6317 ( 
.A1(n_5896),
.A2(n_2987),
.B1(n_2991),
.B2(n_2984),
.Y(n_6317)
);

INVx1_ASAP7_75t_L g6318 ( 
.A(n_5810),
.Y(n_6318)
);

NOR2xp67_ASAP7_75t_L g6319 ( 
.A(n_5921),
.B(n_3394),
.Y(n_6319)
);

BUFx3_ASAP7_75t_L g6320 ( 
.A(n_5709),
.Y(n_6320)
);

AOI22xp33_ASAP7_75t_L g6321 ( 
.A1(n_6183),
.A2(n_3008),
.B1(n_3012),
.B2(n_2998),
.Y(n_6321)
);

AOI22xp5_ASAP7_75t_L g6322 ( 
.A1(n_6108),
.A2(n_6156),
.B1(n_5664),
.B2(n_6104),
.Y(n_6322)
);

HB1xp67_ASAP7_75t_L g6323 ( 
.A(n_5739),
.Y(n_6323)
);

INVx5_ASAP7_75t_L g6324 ( 
.A(n_5755),
.Y(n_6324)
);

NAND2xp5_ASAP7_75t_L g6325 ( 
.A(n_5958),
.B(n_3015),
.Y(n_6325)
);

INVx2_ASAP7_75t_SL g6326 ( 
.A(n_5785),
.Y(n_6326)
);

INVx5_ASAP7_75t_L g6327 ( 
.A(n_5713),
.Y(n_6327)
);

INVx1_ASAP7_75t_L g6328 ( 
.A(n_5975),
.Y(n_6328)
);

AOI22xp33_ASAP7_75t_L g6329 ( 
.A1(n_5659),
.A2(n_5677),
.B1(n_5693),
.B2(n_5680),
.Y(n_6329)
);

OAI22xp5_ASAP7_75t_L g6330 ( 
.A1(n_5682),
.A2(n_3018),
.B1(n_3022),
.B2(n_3017),
.Y(n_6330)
);

NAND2xp5_ASAP7_75t_SL g6331 ( 
.A(n_6139),
.B(n_3023),
.Y(n_6331)
);

AND2x2_ASAP7_75t_L g6332 ( 
.A(n_5845),
.B(n_3395),
.Y(n_6332)
);

NAND2xp5_ASAP7_75t_L g6333 ( 
.A(n_6036),
.B(n_3024),
.Y(n_6333)
);

NAND2xp5_ASAP7_75t_L g6334 ( 
.A(n_6046),
.B(n_3026),
.Y(n_6334)
);

INVx2_ASAP7_75t_SL g6335 ( 
.A(n_5791),
.Y(n_6335)
);

INVx1_ASAP7_75t_L g6336 ( 
.A(n_5977),
.Y(n_6336)
);

CKINVDCx5p33_ASAP7_75t_R g6337 ( 
.A(n_5815),
.Y(n_6337)
);

NOR2xp33_ASAP7_75t_L g6338 ( 
.A(n_5906),
.B(n_3027),
.Y(n_6338)
);

INVx2_ASAP7_75t_L g6339 ( 
.A(n_5772),
.Y(n_6339)
);

NAND2xp5_ASAP7_75t_L g6340 ( 
.A(n_6082),
.B(n_6093),
.Y(n_6340)
);

NAND2xp5_ASAP7_75t_L g6341 ( 
.A(n_6102),
.B(n_3031),
.Y(n_6341)
);

NAND2xp5_ASAP7_75t_SL g6342 ( 
.A(n_6139),
.B(n_3034),
.Y(n_6342)
);

NAND2xp5_ASAP7_75t_SL g6343 ( 
.A(n_5665),
.B(n_3037),
.Y(n_6343)
);

NAND2xp5_ASAP7_75t_L g6344 ( 
.A(n_5817),
.B(n_3041),
.Y(n_6344)
);

NAND2xp5_ASAP7_75t_SL g6345 ( 
.A(n_6172),
.B(n_3044),
.Y(n_6345)
);

NAND2xp5_ASAP7_75t_L g6346 ( 
.A(n_5820),
.B(n_3046),
.Y(n_6346)
);

NAND2xp5_ASAP7_75t_L g6347 ( 
.A(n_5825),
.B(n_3049),
.Y(n_6347)
);

NOR2xp33_ASAP7_75t_L g6348 ( 
.A(n_5887),
.B(n_3054),
.Y(n_6348)
);

AOI22xp33_ASAP7_75t_L g6349 ( 
.A1(n_5913),
.A2(n_3058),
.B1(n_3061),
.B2(n_3056),
.Y(n_6349)
);

O2A1O1Ixp33_ASAP7_75t_L g6350 ( 
.A1(n_5912),
.A2(n_3402),
.B(n_3427),
.C(n_3398),
.Y(n_6350)
);

OR2x6_ASAP7_75t_L g6351 ( 
.A(n_5881),
.B(n_1048),
.Y(n_6351)
);

NOR3xp33_ASAP7_75t_L g6352 ( 
.A(n_6004),
.B(n_3070),
.C(n_3062),
.Y(n_6352)
);

AND2x4_ASAP7_75t_L g6353 ( 
.A(n_5814),
.B(n_3428),
.Y(n_6353)
);

INVx2_ASAP7_75t_L g6354 ( 
.A(n_5773),
.Y(n_6354)
);

CKINVDCx5p33_ASAP7_75t_R g6355 ( 
.A(n_6186),
.Y(n_6355)
);

INVx4_ASAP7_75t_L g6356 ( 
.A(n_5864),
.Y(n_6356)
);

INVx4_ASAP7_75t_L g6357 ( 
.A(n_5715),
.Y(n_6357)
);

NAND2xp5_ASAP7_75t_SL g6358 ( 
.A(n_6163),
.B(n_3076),
.Y(n_6358)
);

INVx2_ASAP7_75t_SL g6359 ( 
.A(n_5793),
.Y(n_6359)
);

AOI21xp5_ASAP7_75t_L g6360 ( 
.A1(n_5733),
.A2(n_3078),
.B(n_3077),
.Y(n_6360)
);

AND2x4_ASAP7_75t_SL g6361 ( 
.A(n_5942),
.B(n_3431),
.Y(n_6361)
);

AOI22xp33_ASAP7_75t_L g6362 ( 
.A1(n_5922),
.A2(n_3088),
.B1(n_3091),
.B2(n_3083),
.Y(n_6362)
);

NAND2xp5_ASAP7_75t_SL g6363 ( 
.A(n_6163),
.B(n_3094),
.Y(n_6363)
);

INVx2_ASAP7_75t_L g6364 ( 
.A(n_5776),
.Y(n_6364)
);

NAND2xp5_ASAP7_75t_L g6365 ( 
.A(n_5986),
.B(n_3100),
.Y(n_6365)
);

AOI21xp5_ASAP7_75t_L g6366 ( 
.A1(n_6161),
.A2(n_3107),
.B(n_3103),
.Y(n_6366)
);

NAND2xp5_ASAP7_75t_L g6367 ( 
.A(n_5989),
.B(n_3115),
.Y(n_6367)
);

HB1xp67_ASAP7_75t_L g6368 ( 
.A(n_5821),
.Y(n_6368)
);

NAND2xp5_ASAP7_75t_L g6369 ( 
.A(n_5991),
.B(n_3116),
.Y(n_6369)
);

AOI22xp5_ASAP7_75t_L g6370 ( 
.A1(n_5664),
.A2(n_3121),
.B1(n_3125),
.B2(n_3118),
.Y(n_6370)
);

NAND2xp5_ASAP7_75t_SL g6371 ( 
.A(n_6056),
.B(n_3131),
.Y(n_6371)
);

NAND2xp5_ASAP7_75t_L g6372 ( 
.A(n_5993),
.B(n_3134),
.Y(n_6372)
);

AOI22xp5_ASAP7_75t_L g6373 ( 
.A1(n_6176),
.A2(n_6165),
.B1(n_6168),
.B2(n_6166),
.Y(n_6373)
);

NOR2xp33_ASAP7_75t_SL g6374 ( 
.A(n_5968),
.B(n_5980),
.Y(n_6374)
);

NAND2xp5_ASAP7_75t_L g6375 ( 
.A(n_5998),
.B(n_3136),
.Y(n_6375)
);

NAND2xp5_ASAP7_75t_L g6376 ( 
.A(n_5999),
.B(n_6000),
.Y(n_6376)
);

NAND2xp5_ASAP7_75t_L g6377 ( 
.A(n_6003),
.B(n_3139),
.Y(n_6377)
);

A2O1A1Ixp33_ASAP7_75t_L g6378 ( 
.A1(n_6153),
.A2(n_3452),
.B(n_3454),
.C(n_3438),
.Y(n_6378)
);

NAND2xp5_ASAP7_75t_L g6379 ( 
.A(n_6006),
.B(n_3140),
.Y(n_6379)
);

NOR2xp33_ASAP7_75t_L g6380 ( 
.A(n_5873),
.B(n_3148),
.Y(n_6380)
);

AND2x6_ASAP7_75t_SL g6381 ( 
.A(n_5789),
.B(n_3455),
.Y(n_6381)
);

NOR2xp33_ASAP7_75t_L g6382 ( 
.A(n_5878),
.B(n_3153),
.Y(n_6382)
);

NAND2xp5_ASAP7_75t_L g6383 ( 
.A(n_6008),
.B(n_3154),
.Y(n_6383)
);

INVx1_ASAP7_75t_L g6384 ( 
.A(n_6013),
.Y(n_6384)
);

NAND2xp5_ASAP7_75t_SL g6385 ( 
.A(n_6017),
.B(n_3162),
.Y(n_6385)
);

NAND2xp5_ASAP7_75t_L g6386 ( 
.A(n_6030),
.B(n_3169),
.Y(n_6386)
);

BUFx3_ASAP7_75t_L g6387 ( 
.A(n_5731),
.Y(n_6387)
);

INVx2_ASAP7_75t_SL g6388 ( 
.A(n_5752),
.Y(n_6388)
);

NOR2xp33_ASAP7_75t_L g6389 ( 
.A(n_5907),
.B(n_3174),
.Y(n_6389)
);

INVxp67_ASAP7_75t_L g6390 ( 
.A(n_5718),
.Y(n_6390)
);

OAI22xp5_ASAP7_75t_L g6391 ( 
.A1(n_6041),
.A2(n_6052),
.B1(n_6058),
.B2(n_6055),
.Y(n_6391)
);

O2A1O1Ixp5_ASAP7_75t_L g6392 ( 
.A1(n_6162),
.A2(n_3461),
.B(n_3462),
.C(n_3459),
.Y(n_6392)
);

AND2x6_ASAP7_75t_SL g6393 ( 
.A(n_5747),
.B(n_3463),
.Y(n_6393)
);

INVx1_ASAP7_75t_L g6394 ( 
.A(n_6064),
.Y(n_6394)
);

NOR3xp33_ASAP7_75t_SL g6395 ( 
.A(n_5769),
.B(n_3481),
.C(n_3467),
.Y(n_6395)
);

NAND2xp5_ASAP7_75t_L g6396 ( 
.A(n_6065),
.B(n_6067),
.Y(n_6396)
);

INVxp33_ASAP7_75t_L g6397 ( 
.A(n_5722),
.Y(n_6397)
);

NOR2xp33_ASAP7_75t_L g6398 ( 
.A(n_6169),
.B(n_3176),
.Y(n_6398)
);

NAND2xp5_ASAP7_75t_L g6399 ( 
.A(n_5816),
.B(n_3177),
.Y(n_6399)
);

INVx2_ASAP7_75t_L g6400 ( 
.A(n_5777),
.Y(n_6400)
);

NOR2xp33_ASAP7_75t_L g6401 ( 
.A(n_5800),
.B(n_3178),
.Y(n_6401)
);

NAND2xp5_ASAP7_75t_L g6402 ( 
.A(n_5826),
.B(n_3180),
.Y(n_6402)
);

INVx2_ASAP7_75t_L g6403 ( 
.A(n_5783),
.Y(n_6403)
);

INVx1_ASAP7_75t_L g6404 ( 
.A(n_6072),
.Y(n_6404)
);

HB1xp67_ASAP7_75t_L g6405 ( 
.A(n_5767),
.Y(n_6405)
);

INVx1_ASAP7_75t_L g6406 ( 
.A(n_6073),
.Y(n_6406)
);

NAND2xp5_ASAP7_75t_L g6407 ( 
.A(n_5915),
.B(n_3182),
.Y(n_6407)
);

NAND2xp5_ASAP7_75t_L g6408 ( 
.A(n_5916),
.B(n_3183),
.Y(n_6408)
);

NAND2x1_ASAP7_75t_L g6409 ( 
.A(n_5790),
.B(n_1049),
.Y(n_6409)
);

NAND2xp5_ASAP7_75t_L g6410 ( 
.A(n_5918),
.B(n_3186),
.Y(n_6410)
);

INVx2_ASAP7_75t_L g6411 ( 
.A(n_5809),
.Y(n_6411)
);

AOI22xp33_ASAP7_75t_L g6412 ( 
.A1(n_5927),
.A2(n_3190),
.B1(n_3200),
.B2(n_3189),
.Y(n_6412)
);

INVx2_ASAP7_75t_L g6413 ( 
.A(n_5813),
.Y(n_6413)
);

BUFx3_ASAP7_75t_L g6414 ( 
.A(n_5805),
.Y(n_6414)
);

INVx1_ASAP7_75t_L g6415 ( 
.A(n_6074),
.Y(n_6415)
);

NOR2xp33_ASAP7_75t_L g6416 ( 
.A(n_5976),
.B(n_3203),
.Y(n_6416)
);

NAND2xp5_ASAP7_75t_L g6417 ( 
.A(n_5924),
.B(n_3207),
.Y(n_6417)
);

OAI22xp33_ASAP7_75t_L g6418 ( 
.A1(n_6157),
.A2(n_3488),
.B1(n_3492),
.B2(n_3483),
.Y(n_6418)
);

INVx1_ASAP7_75t_L g6419 ( 
.A(n_6079),
.Y(n_6419)
);

BUFx6f_ASAP7_75t_SL g6420 ( 
.A(n_5858),
.Y(n_6420)
);

INVx3_ASAP7_75t_L g6421 ( 
.A(n_5811),
.Y(n_6421)
);

NAND2xp5_ASAP7_75t_L g6422 ( 
.A(n_5926),
.B(n_3211),
.Y(n_6422)
);

INVx2_ASAP7_75t_L g6423 ( 
.A(n_5822),
.Y(n_6423)
);

INVx1_ASAP7_75t_L g6424 ( 
.A(n_6081),
.Y(n_6424)
);

NAND2xp33_ASAP7_75t_SL g6425 ( 
.A(n_5992),
.B(n_3497),
.Y(n_6425)
);

NAND2xp5_ASAP7_75t_L g6426 ( 
.A(n_5930),
.B(n_3212),
.Y(n_6426)
);

BUFx2_ASAP7_75t_L g6427 ( 
.A(n_5819),
.Y(n_6427)
);

NAND2x1_ASAP7_75t_L g6428 ( 
.A(n_5823),
.B(n_1049),
.Y(n_6428)
);

NAND2xp5_ASAP7_75t_L g6429 ( 
.A(n_5936),
.B(n_3213),
.Y(n_6429)
);

AOI22xp5_ASAP7_75t_L g6430 ( 
.A1(n_6164),
.A2(n_3216),
.B1(n_3218),
.B2(n_3214),
.Y(n_6430)
);

O2A1O1Ixp33_ASAP7_75t_L g6431 ( 
.A1(n_5932),
.A2(n_6117),
.B(n_5782),
.C(n_5797),
.Y(n_6431)
);

BUFx3_ASAP7_75t_L g6432 ( 
.A(n_5841),
.Y(n_6432)
);

NAND2x1_ASAP7_75t_L g6433 ( 
.A(n_5824),
.B(n_1050),
.Y(n_6433)
);

AND2x2_ASAP7_75t_L g6434 ( 
.A(n_6038),
.B(n_3509),
.Y(n_6434)
);

INVx4_ASAP7_75t_L g6435 ( 
.A(n_5841),
.Y(n_6435)
);

NOR2xp67_ASAP7_75t_L g6436 ( 
.A(n_5945),
.B(n_3516),
.Y(n_6436)
);

NAND2xp5_ASAP7_75t_L g6437 ( 
.A(n_5946),
.B(n_3219),
.Y(n_6437)
);

INVx1_ASAP7_75t_L g6438 ( 
.A(n_6086),
.Y(n_6438)
);

O2A1O1Ixp33_ASAP7_75t_L g6439 ( 
.A1(n_5788),
.A2(n_3537),
.B(n_3541),
.C(n_3526),
.Y(n_6439)
);

NAND2xp5_ASAP7_75t_L g6440 ( 
.A(n_5950),
.B(n_3221),
.Y(n_6440)
);

NAND2xp5_ASAP7_75t_L g6441 ( 
.A(n_5951),
.B(n_3224),
.Y(n_6441)
);

NAND2xp5_ASAP7_75t_L g6442 ( 
.A(n_5953),
.B(n_3226),
.Y(n_6442)
);

INVx2_ASAP7_75t_SL g6443 ( 
.A(n_6044),
.Y(n_6443)
);

NAND2xp5_ASAP7_75t_L g6444 ( 
.A(n_5827),
.B(n_3230),
.Y(n_6444)
);

NAND2xp5_ASAP7_75t_L g6445 ( 
.A(n_5828),
.B(n_3231),
.Y(n_6445)
);

INVx2_ASAP7_75t_SL g6446 ( 
.A(n_6044),
.Y(n_6446)
);

NAND2xp5_ASAP7_75t_L g6447 ( 
.A(n_5833),
.B(n_5836),
.Y(n_6447)
);

INVx1_ASAP7_75t_L g6448 ( 
.A(n_6097),
.Y(n_6448)
);

INVxp67_ASAP7_75t_SL g6449 ( 
.A(n_5692),
.Y(n_6449)
);

AND2x2_ASAP7_75t_L g6450 ( 
.A(n_6040),
.B(n_3550),
.Y(n_6450)
);

AOI22xp33_ASAP7_75t_L g6451 ( 
.A1(n_5928),
.A2(n_3240),
.B1(n_3242),
.B2(n_3236),
.Y(n_6451)
);

NAND2xp5_ASAP7_75t_L g6452 ( 
.A(n_5847),
.B(n_3243),
.Y(n_6452)
);

NAND2xp5_ASAP7_75t_L g6453 ( 
.A(n_5855),
.B(n_3246),
.Y(n_6453)
);

INVx2_ASAP7_75t_L g6454 ( 
.A(n_5829),
.Y(n_6454)
);

INVx1_ASAP7_75t_L g6455 ( 
.A(n_6099),
.Y(n_6455)
);

NAND2xp5_ASAP7_75t_L g6456 ( 
.A(n_5856),
.B(n_3248),
.Y(n_6456)
);

NOR2xp33_ASAP7_75t_L g6457 ( 
.A(n_6042),
.B(n_6047),
.Y(n_6457)
);

INVx5_ASAP7_75t_L g6458 ( 
.A(n_5858),
.Y(n_6458)
);

AOI22xp33_ASAP7_75t_L g6459 ( 
.A1(n_5931),
.A2(n_3250),
.B1(n_3259),
.B2(n_3249),
.Y(n_6459)
);

NAND2xp5_ASAP7_75t_L g6460 ( 
.A(n_5865),
.B(n_5875),
.Y(n_6460)
);

NAND2xp5_ASAP7_75t_L g6461 ( 
.A(n_5934),
.B(n_5879),
.Y(n_6461)
);

AOI22xp5_ASAP7_75t_L g6462 ( 
.A1(n_6174),
.A2(n_3266),
.B1(n_3268),
.B2(n_3262),
.Y(n_6462)
);

NAND2xp5_ASAP7_75t_L g6463 ( 
.A(n_5883),
.B(n_3269),
.Y(n_6463)
);

OAI22xp5_ASAP7_75t_L g6464 ( 
.A1(n_6070),
.A2(n_3278),
.B1(n_3281),
.B2(n_3273),
.Y(n_6464)
);

NAND2xp5_ASAP7_75t_L g6465 ( 
.A(n_5885),
.B(n_3282),
.Y(n_6465)
);

NOR2x1p5_ASAP7_75t_L g6466 ( 
.A(n_6094),
.B(n_3556),
.Y(n_6466)
);

NAND2xp5_ASAP7_75t_L g6467 ( 
.A(n_5888),
.B(n_3285),
.Y(n_6467)
);

AND2x6_ASAP7_75t_SL g6468 ( 
.A(n_5898),
.B(n_3564),
.Y(n_6468)
);

NAND2xp5_ASAP7_75t_L g6469 ( 
.A(n_5890),
.B(n_3287),
.Y(n_6469)
);

NOR2xp33_ASAP7_75t_L g6470 ( 
.A(n_6054),
.B(n_3295),
.Y(n_6470)
);

INVx1_ASAP7_75t_L g6471 ( 
.A(n_6101),
.Y(n_6471)
);

INVx1_ASAP7_75t_L g6472 ( 
.A(n_6110),
.Y(n_6472)
);

OR2x2_ASAP7_75t_L g6473 ( 
.A(n_5803),
.B(n_3572),
.Y(n_6473)
);

NAND2xp5_ASAP7_75t_SL g6474 ( 
.A(n_6120),
.B(n_3296),
.Y(n_6474)
);

NAND2xp5_ASAP7_75t_L g6475 ( 
.A(n_5895),
.B(n_3300),
.Y(n_6475)
);

NAND2xp5_ASAP7_75t_L g6476 ( 
.A(n_5910),
.B(n_3303),
.Y(n_6476)
);

CKINVDCx20_ASAP7_75t_R g6477 ( 
.A(n_5749),
.Y(n_6477)
);

INVx3_ASAP7_75t_L g6478 ( 
.A(n_5860),
.Y(n_6478)
);

O2A1O1Ixp5_ASAP7_75t_L g6479 ( 
.A1(n_6021),
.A2(n_3582),
.B(n_3583),
.C(n_3573),
.Y(n_6479)
);

INVx2_ASAP7_75t_L g6480 ( 
.A(n_5830),
.Y(n_6480)
);

INVxp33_ASAP7_75t_SL g6481 ( 
.A(n_5871),
.Y(n_6481)
);

INVx1_ASAP7_75t_L g6482 ( 
.A(n_5979),
.Y(n_6482)
);

INVx2_ASAP7_75t_L g6483 ( 
.A(n_5837),
.Y(n_6483)
);

NOR2xp33_ASAP7_75t_L g6484 ( 
.A(n_5940),
.B(n_3308),
.Y(n_6484)
);

O2A1O1Ixp33_ASAP7_75t_L g6485 ( 
.A1(n_6145),
.A2(n_3594),
.B(n_3598),
.C(n_3590),
.Y(n_6485)
);

AOI21xp5_ASAP7_75t_L g6486 ( 
.A1(n_5884),
.A2(n_3314),
.B(n_3310),
.Y(n_6486)
);

BUFx6f_ASAP7_75t_L g6487 ( 
.A(n_6119),
.Y(n_6487)
);

NAND2xp5_ASAP7_75t_L g6488 ( 
.A(n_5967),
.B(n_3315),
.Y(n_6488)
);

NAND2x1_ASAP7_75t_L g6489 ( 
.A(n_5842),
.B(n_1051),
.Y(n_6489)
);

NAND2xp5_ASAP7_75t_SL g6490 ( 
.A(n_6116),
.B(n_3316),
.Y(n_6490)
);

NAND2xp5_ASAP7_75t_L g6491 ( 
.A(n_5970),
.B(n_3317),
.Y(n_6491)
);

INVx4_ASAP7_75t_L g6492 ( 
.A(n_5945),
.Y(n_6492)
);

NOR2x1p5_ASAP7_75t_L g6493 ( 
.A(n_6051),
.B(n_3602),
.Y(n_6493)
);

NAND2xp5_ASAP7_75t_L g6494 ( 
.A(n_5956),
.B(n_3320),
.Y(n_6494)
);

AOI22xp5_ASAP7_75t_L g6495 ( 
.A1(n_6175),
.A2(n_3326),
.B1(n_3329),
.B2(n_3322),
.Y(n_6495)
);

INVxp67_ASAP7_75t_L g6496 ( 
.A(n_6119),
.Y(n_6496)
);

NAND2xp5_ASAP7_75t_L g6497 ( 
.A(n_5963),
.B(n_3331),
.Y(n_6497)
);

AOI22xp5_ASAP7_75t_L g6498 ( 
.A1(n_6024),
.A2(n_3333),
.B1(n_3335),
.B2(n_3332),
.Y(n_6498)
);

NAND2xp5_ASAP7_75t_SL g6499 ( 
.A(n_6096),
.B(n_3336),
.Y(n_6499)
);

INVx1_ASAP7_75t_L g6500 ( 
.A(n_5982),
.Y(n_6500)
);

AND2x4_ASAP7_75t_L g6501 ( 
.A(n_5723),
.B(n_3606),
.Y(n_6501)
);

INVx4_ASAP7_75t_L g6502 ( 
.A(n_5861),
.Y(n_6502)
);

NAND2xp5_ASAP7_75t_L g6503 ( 
.A(n_5843),
.B(n_3337),
.Y(n_6503)
);

INVx2_ASAP7_75t_L g6504 ( 
.A(n_5848),
.Y(n_6504)
);

AOI22xp33_ASAP7_75t_L g6505 ( 
.A1(n_6023),
.A2(n_3339),
.B1(n_3350),
.B2(n_3338),
.Y(n_6505)
);

NAND2xp5_ASAP7_75t_L g6506 ( 
.A(n_5854),
.B(n_3351),
.Y(n_6506)
);

INVx5_ASAP7_75t_L g6507 ( 
.A(n_5784),
.Y(n_6507)
);

NAND2xp5_ASAP7_75t_L g6508 ( 
.A(n_5859),
.B(n_3352),
.Y(n_6508)
);

NAND2xp5_ASAP7_75t_L g6509 ( 
.A(n_5903),
.B(n_3357),
.Y(n_6509)
);

NAND2xp5_ASAP7_75t_L g6510 ( 
.A(n_5964),
.B(n_6016),
.Y(n_6510)
);

AND2x2_ASAP7_75t_L g6511 ( 
.A(n_6045),
.B(n_3607),
.Y(n_6511)
);

NAND2xp5_ASAP7_75t_L g6512 ( 
.A(n_6016),
.B(n_3360),
.Y(n_6512)
);

INVx1_ASAP7_75t_L g6513 ( 
.A(n_5983),
.Y(n_6513)
);

AOI22xp33_ASAP7_75t_L g6514 ( 
.A1(n_6029),
.A2(n_3363),
.B1(n_3367),
.B2(n_3362),
.Y(n_6514)
);

INVx2_ASAP7_75t_SL g6515 ( 
.A(n_6096),
.Y(n_6515)
);

NOR2xp33_ASAP7_75t_L g6516 ( 
.A(n_5962),
.B(n_3368),
.Y(n_6516)
);

NAND2xp5_ASAP7_75t_L g6517 ( 
.A(n_6071),
.B(n_3372),
.Y(n_6517)
);

NAND2xp5_ASAP7_75t_SL g6518 ( 
.A(n_6031),
.B(n_3377),
.Y(n_6518)
);

NAND2xp5_ASAP7_75t_L g6519 ( 
.A(n_6050),
.B(n_3378),
.Y(n_6519)
);

NAND2xp5_ASAP7_75t_L g6520 ( 
.A(n_6068),
.B(n_5981),
.Y(n_6520)
);

INVx1_ASAP7_75t_L g6521 ( 
.A(n_5994),
.Y(n_6521)
);

INVx1_ASAP7_75t_L g6522 ( 
.A(n_6005),
.Y(n_6522)
);

NAND2xp5_ASAP7_75t_SL g6523 ( 
.A(n_6127),
.B(n_3392),
.Y(n_6523)
);

OAI22xp5_ASAP7_75t_L g6524 ( 
.A1(n_5891),
.A2(n_3397),
.B1(n_3399),
.B2(n_3396),
.Y(n_6524)
);

INVx1_ASAP7_75t_L g6525 ( 
.A(n_6132),
.Y(n_6525)
);

INVx1_ASAP7_75t_L g6526 ( 
.A(n_6134),
.Y(n_6526)
);

NAND2xp5_ASAP7_75t_L g6527 ( 
.A(n_6027),
.B(n_3404),
.Y(n_6527)
);

OAI21xp5_ASAP7_75t_L g6528 ( 
.A1(n_5908),
.A2(n_3408),
.B(n_3405),
.Y(n_6528)
);

NAND2xp5_ASAP7_75t_L g6529 ( 
.A(n_6027),
.B(n_3410),
.Y(n_6529)
);

CKINVDCx20_ASAP7_75t_R g6530 ( 
.A(n_5807),
.Y(n_6530)
);

NAND2xp5_ASAP7_75t_SL g6531 ( 
.A(n_6136),
.B(n_3420),
.Y(n_6531)
);

INVx4_ASAP7_75t_L g6532 ( 
.A(n_5849),
.Y(n_6532)
);

NAND2xp5_ASAP7_75t_L g6533 ( 
.A(n_6077),
.B(n_3421),
.Y(n_6533)
);

NAND2xp5_ASAP7_75t_L g6534 ( 
.A(n_6087),
.B(n_3422),
.Y(n_6534)
);

NAND2xp5_ASAP7_75t_L g6535 ( 
.A(n_6088),
.B(n_3426),
.Y(n_6535)
);

INVx1_ASAP7_75t_L g6536 ( 
.A(n_6137),
.Y(n_6536)
);

AOI221xp5_ASAP7_75t_L g6537 ( 
.A1(n_5832),
.A2(n_3435),
.B1(n_3436),
.B2(n_3433),
.C(n_3432),
.Y(n_6537)
);

NOR2xp33_ASAP7_75t_L g6538 ( 
.A(n_5929),
.B(n_3447),
.Y(n_6538)
);

NAND2xp5_ASAP7_75t_SL g6539 ( 
.A(n_5972),
.B(n_3451),
.Y(n_6539)
);

A2O1A1Ixp33_ASAP7_75t_L g6540 ( 
.A1(n_5984),
.A2(n_3456),
.B(n_3458),
.C(n_3453),
.Y(n_6540)
);

NAND2xp5_ASAP7_75t_L g6541 ( 
.A(n_6095),
.B(n_3465),
.Y(n_6541)
);

NAND2xp5_ASAP7_75t_L g6542 ( 
.A(n_6113),
.B(n_3470),
.Y(n_6542)
);

NOR2xp33_ASAP7_75t_L g6543 ( 
.A(n_6148),
.B(n_3476),
.Y(n_6543)
);

INVx1_ASAP7_75t_L g6544 ( 
.A(n_6115),
.Y(n_6544)
);

INVxp67_ASAP7_75t_L g6545 ( 
.A(n_6066),
.Y(n_6545)
);

NAND2xp5_ASAP7_75t_L g6546 ( 
.A(n_6118),
.B(n_6124),
.Y(n_6546)
);

NOR2xp33_ASAP7_75t_L g6547 ( 
.A(n_5726),
.B(n_3485),
.Y(n_6547)
);

AOI22xp5_ASAP7_75t_L g6548 ( 
.A1(n_5671),
.A2(n_5727),
.B1(n_6177),
.B2(n_6060),
.Y(n_6548)
);

NOR2xp33_ASAP7_75t_L g6549 ( 
.A(n_6143),
.B(n_3489),
.Y(n_6549)
);

INVx2_ASAP7_75t_L g6550 ( 
.A(n_5846),
.Y(n_6550)
);

NAND2xp5_ASAP7_75t_L g6551 ( 
.A(n_5978),
.B(n_3490),
.Y(n_6551)
);

HB1xp67_ASAP7_75t_L g6552 ( 
.A(n_5701),
.Y(n_6552)
);

NAND2xp5_ASAP7_75t_SL g6553 ( 
.A(n_5857),
.B(n_3491),
.Y(n_6553)
);

AOI22xp33_ASAP7_75t_L g6554 ( 
.A1(n_6012),
.A2(n_3504),
.B1(n_3505),
.B2(n_3496),
.Y(n_6554)
);

INVx2_ASAP7_75t_SL g6555 ( 
.A(n_5904),
.Y(n_6555)
);

OAI22xp5_ASAP7_75t_L g6556 ( 
.A1(n_6140),
.A2(n_3510),
.B1(n_3512),
.B2(n_3507),
.Y(n_6556)
);

INVx2_ASAP7_75t_L g6557 ( 
.A(n_6128),
.Y(n_6557)
);

NOR2xp33_ASAP7_75t_L g6558 ( 
.A(n_6146),
.B(n_6178),
.Y(n_6558)
);

INVx2_ASAP7_75t_SL g6559 ( 
.A(n_5904),
.Y(n_6559)
);

AOI22xp5_ASAP7_75t_L g6560 ( 
.A1(n_5727),
.A2(n_3519),
.B1(n_3525),
.B2(n_3515),
.Y(n_6560)
);

NAND2xp5_ASAP7_75t_L g6561 ( 
.A(n_6135),
.B(n_3528),
.Y(n_6561)
);

NOR2xp33_ASAP7_75t_L g6562 ( 
.A(n_6125),
.B(n_3534),
.Y(n_6562)
);

INVx1_ASAP7_75t_L g6563 ( 
.A(n_6001),
.Y(n_6563)
);

INVx2_ASAP7_75t_L g6564 ( 
.A(n_6106),
.Y(n_6564)
);

NOR2xp33_ASAP7_75t_L g6565 ( 
.A(n_5708),
.B(n_3535),
.Y(n_6565)
);

NAND2xp5_ASAP7_75t_L g6566 ( 
.A(n_5997),
.B(n_3539),
.Y(n_6566)
);

OR2x6_ASAP7_75t_L g6567 ( 
.A(n_5969),
.B(n_1052),
.Y(n_6567)
);

OR2x2_ASAP7_75t_L g6568 ( 
.A(n_6138),
.B(n_3543),
.Y(n_6568)
);

INVx2_ASAP7_75t_L g6569 ( 
.A(n_6114),
.Y(n_6569)
);

NAND2xp5_ASAP7_75t_L g6570 ( 
.A(n_6020),
.B(n_3546),
.Y(n_6570)
);

AND2x2_ASAP7_75t_L g6571 ( 
.A(n_5877),
.B(n_3551),
.Y(n_6571)
);

NAND2xp5_ASAP7_75t_L g6572 ( 
.A(n_6122),
.B(n_3552),
.Y(n_6572)
);

NOR2xp67_ASAP7_75t_L g6573 ( 
.A(n_6002),
.B(n_6007),
.Y(n_6573)
);

NAND2xp5_ASAP7_75t_L g6574 ( 
.A(n_6091),
.B(n_3554),
.Y(n_6574)
);

AND2x2_ASAP7_75t_L g6575 ( 
.A(n_5886),
.B(n_3558),
.Y(n_6575)
);

OAI21xp5_ASAP7_75t_L g6576 ( 
.A1(n_6155),
.A2(n_3565),
.B(n_3561),
.Y(n_6576)
);

NAND2xp5_ASAP7_75t_SL g6577 ( 
.A(n_5985),
.B(n_3576),
.Y(n_6577)
);

INVx3_ASAP7_75t_L g6578 ( 
.A(n_6010),
.Y(n_6578)
);

OAI22xp5_ASAP7_75t_L g6579 ( 
.A1(n_5965),
.A2(n_3579),
.B1(n_3581),
.B2(n_3577),
.Y(n_6579)
);

NAND2xp5_ASAP7_75t_L g6580 ( 
.A(n_6091),
.B(n_3584),
.Y(n_6580)
);

INVx2_ASAP7_75t_SL g6581 ( 
.A(n_5966),
.Y(n_6581)
);

NAND2xp5_ASAP7_75t_SL g6582 ( 
.A(n_6141),
.B(n_3586),
.Y(n_6582)
);

NAND2xp5_ASAP7_75t_L g6583 ( 
.A(n_6098),
.B(n_3592),
.Y(n_6583)
);

NAND2xp5_ASAP7_75t_L g6584 ( 
.A(n_6123),
.B(n_3593),
.Y(n_6584)
);

AOI22xp33_ASAP7_75t_L g6585 ( 
.A1(n_5947),
.A2(n_3604),
.B1(n_3609),
.B2(n_3601),
.Y(n_6585)
);

CKINVDCx5p33_ASAP7_75t_R g6586 ( 
.A(n_5944),
.Y(n_6586)
);

AOI22xp33_ASAP7_75t_L g6587 ( 
.A1(n_5947),
.A2(n_3615),
.B1(n_3617),
.B2(n_3611),
.Y(n_6587)
);

OR2x2_ASAP7_75t_L g6588 ( 
.A(n_5831),
.B(n_3619),
.Y(n_6588)
);

INVx2_ASAP7_75t_L g6589 ( 
.A(n_5987),
.Y(n_6589)
);

NAND2xp5_ASAP7_75t_L g6590 ( 
.A(n_5961),
.B(n_3624),
.Y(n_6590)
);

NOR2xp33_ASAP7_75t_L g6591 ( 
.A(n_5765),
.B(n_5990),
.Y(n_6591)
);

NAND2xp5_ASAP7_75t_SL g6592 ( 
.A(n_6141),
.B(n_3625),
.Y(n_6592)
);

NAND2xp5_ASAP7_75t_SL g6593 ( 
.A(n_6142),
.B(n_3628),
.Y(n_6593)
);

AOI22xp5_ASAP7_75t_L g6594 ( 
.A1(n_5775),
.A2(n_1054),
.B1(n_1055),
.B2(n_1053),
.Y(n_6594)
);

INVx1_ASAP7_75t_L g6595 ( 
.A(n_6144),
.Y(n_6595)
);

NAND2xp5_ASAP7_75t_SL g6596 ( 
.A(n_5874),
.B(n_6084),
.Y(n_6596)
);

NAND2xp5_ASAP7_75t_L g6597 ( 
.A(n_6152),
.B(n_2),
.Y(n_6597)
);

NOR2xp33_ASAP7_75t_L g6598 ( 
.A(n_5995),
.B(n_1054),
.Y(n_6598)
);

INVx1_ASAP7_75t_L g6599 ( 
.A(n_6147),
.Y(n_6599)
);

NAND2xp5_ASAP7_75t_SL g6600 ( 
.A(n_6089),
.B(n_1055),
.Y(n_6600)
);

AO22x1_ASAP7_75t_L g6601 ( 
.A1(n_5784),
.A2(n_5),
.B1(n_2),
.B2(n_3),
.Y(n_6601)
);

AOI22xp33_ASAP7_75t_L g6602 ( 
.A1(n_6107),
.A2(n_1057),
.B1(n_1058),
.B2(n_1056),
.Y(n_6602)
);

NOR2xp33_ASAP7_75t_L g6603 ( 
.A(n_6033),
.B(n_6043),
.Y(n_6603)
);

AOI21xp5_ASAP7_75t_L g6604 ( 
.A1(n_5954),
.A2(n_1059),
.B(n_1056),
.Y(n_6604)
);

NAND2xp5_ASAP7_75t_L g6605 ( 
.A(n_6152),
.B(n_3),
.Y(n_6605)
);

NAND2xp5_ASAP7_75t_L g6606 ( 
.A(n_5780),
.B(n_5),
.Y(n_6606)
);

NAND2xp5_ASAP7_75t_L g6607 ( 
.A(n_5909),
.B(n_6),
.Y(n_6607)
);

INVx2_ASAP7_75t_L g6608 ( 
.A(n_5917),
.Y(n_6608)
);

NAND2x1_ASAP7_75t_L g6609 ( 
.A(n_6078),
.B(n_1060),
.Y(n_6609)
);

NAND2xp5_ASAP7_75t_L g6610 ( 
.A(n_5919),
.B(n_6160),
.Y(n_6610)
);

NAND2xp5_ASAP7_75t_L g6611 ( 
.A(n_5900),
.B(n_6),
.Y(n_6611)
);

INVx1_ASAP7_75t_L g6612 ( 
.A(n_5889),
.Y(n_6612)
);

AND2x6_ASAP7_75t_SL g6613 ( 
.A(n_6022),
.B(n_6),
.Y(n_6613)
);

NOR2xp33_ASAP7_75t_SL g6614 ( 
.A(n_5778),
.B(n_5774),
.Y(n_6614)
);

NAND2xp5_ASAP7_75t_SL g6615 ( 
.A(n_6150),
.B(n_1060),
.Y(n_6615)
);

INVxp67_ASAP7_75t_L g6616 ( 
.A(n_6075),
.Y(n_6616)
);

AND2x2_ASAP7_75t_L g6617 ( 
.A(n_5868),
.B(n_1061),
.Y(n_6617)
);

BUFx2_ASAP7_75t_L g6618 ( 
.A(n_6170),
.Y(n_6618)
);

NAND2xp5_ASAP7_75t_L g6619 ( 
.A(n_5923),
.B(n_7),
.Y(n_6619)
);

INVx1_ASAP7_75t_L g6620 ( 
.A(n_6126),
.Y(n_6620)
);

OAI221xp5_ASAP7_75t_L g6621 ( 
.A1(n_6131),
.A2(n_9),
.B1(n_7),
.B2(n_8),
.C(n_10),
.Y(n_6621)
);

NAND2xp5_ASAP7_75t_SL g6622 ( 
.A(n_6014),
.B(n_1062),
.Y(n_6622)
);

NOR2xp33_ASAP7_75t_L g6623 ( 
.A(n_6090),
.B(n_1063),
.Y(n_6623)
);

BUFx6f_ASAP7_75t_L g6624 ( 
.A(n_5935),
.Y(n_6624)
);

NOR2xp33_ASAP7_75t_L g6625 ( 
.A(n_5716),
.B(n_1063),
.Y(n_6625)
);

NAND2xp5_ASAP7_75t_L g6626 ( 
.A(n_5960),
.B(n_7),
.Y(n_6626)
);

INVx1_ASAP7_75t_L g6627 ( 
.A(n_6028),
.Y(n_6627)
);

NAND2xp5_ASAP7_75t_L g6628 ( 
.A(n_5867),
.B(n_8),
.Y(n_6628)
);

INVx1_ASAP7_75t_L g6629 ( 
.A(n_6034),
.Y(n_6629)
);

OR2x2_ASAP7_75t_L g6630 ( 
.A(n_5911),
.B(n_1064),
.Y(n_6630)
);

INVx2_ASAP7_75t_L g6631 ( 
.A(n_5892),
.Y(n_6631)
);

AOI22xp33_ASAP7_75t_L g6632 ( 
.A1(n_6076),
.A2(n_1066),
.B1(n_1067),
.B2(n_1065),
.Y(n_6632)
);

INVx2_ASAP7_75t_L g6633 ( 
.A(n_5920),
.Y(n_6633)
);

AOI22xp33_ASAP7_75t_L g6634 ( 
.A1(n_5834),
.A2(n_1068),
.B1(n_1069),
.B2(n_1066),
.Y(n_6634)
);

NOR2xp33_ASAP7_75t_L g6635 ( 
.A(n_5762),
.B(n_1068),
.Y(n_6635)
);

NAND2xp5_ASAP7_75t_SL g6636 ( 
.A(n_5801),
.B(n_1069),
.Y(n_6636)
);

NOR2xp33_ASAP7_75t_L g6637 ( 
.A(n_5729),
.B(n_1070),
.Y(n_6637)
);

AND2x2_ASAP7_75t_L g6638 ( 
.A(n_5914),
.B(n_1070),
.Y(n_6638)
);

NAND2xp5_ASAP7_75t_SL g6639 ( 
.A(n_5937),
.B(n_1071),
.Y(n_6639)
);

NOR2x2_ASAP7_75t_L g6640 ( 
.A(n_6179),
.B(n_9),
.Y(n_6640)
);

INVx2_ASAP7_75t_L g6641 ( 
.A(n_5952),
.Y(n_6641)
);

INVx1_ASAP7_75t_L g6642 ( 
.A(n_6015),
.Y(n_6642)
);

NOR2xp33_ASAP7_75t_L g6643 ( 
.A(n_6063),
.B(n_1071),
.Y(n_6643)
);

BUFx8_ASAP7_75t_L g6644 ( 
.A(n_5781),
.Y(n_6644)
);

NAND2xp5_ASAP7_75t_SL g6645 ( 
.A(n_6025),
.B(n_1072),
.Y(n_6645)
);

NAND2xp5_ASAP7_75t_L g6646 ( 
.A(n_5974),
.B(n_9),
.Y(n_6646)
);

INVx3_ASAP7_75t_L g6647 ( 
.A(n_5966),
.Y(n_6647)
);

AOI22xp5_ASAP7_75t_L g6648 ( 
.A1(n_6112),
.A2(n_1074),
.B1(n_1075),
.B2(n_1073),
.Y(n_6648)
);

BUFx6f_ASAP7_75t_L g6649 ( 
.A(n_5973),
.Y(n_6649)
);

NAND2xp5_ASAP7_75t_L g6650 ( 
.A(n_6130),
.B(n_10),
.Y(n_6650)
);

AND2x2_ASAP7_75t_L g6651 ( 
.A(n_5852),
.B(n_1073),
.Y(n_6651)
);

NAND2xp5_ASAP7_75t_L g6652 ( 
.A(n_6053),
.B(n_11),
.Y(n_6652)
);

INVx1_ASAP7_75t_L g6653 ( 
.A(n_5844),
.Y(n_6653)
);

INVx1_ASAP7_75t_L g6654 ( 
.A(n_6057),
.Y(n_6654)
);

AOI22xp33_ASAP7_75t_L g6655 ( 
.A1(n_5792),
.A2(n_1076),
.B1(n_1077),
.B2(n_1074),
.Y(n_6655)
);

NAND2xp5_ASAP7_75t_L g6656 ( 
.A(n_5941),
.B(n_11),
.Y(n_6656)
);

NAND2xp5_ASAP7_75t_L g6657 ( 
.A(n_6129),
.B(n_11),
.Y(n_6657)
);

INVx4_ASAP7_75t_L g6658 ( 
.A(n_6048),
.Y(n_6658)
);

NOR2xp33_ASAP7_75t_SL g6659 ( 
.A(n_5786),
.B(n_12),
.Y(n_6659)
);

NAND2xp5_ASAP7_75t_L g6660 ( 
.A(n_6059),
.B(n_12),
.Y(n_6660)
);

BUFx4f_ASAP7_75t_SL g6661 ( 
.A(n_6477),
.Y(n_6661)
);

INVx5_ASAP7_75t_L g6662 ( 
.A(n_6223),
.Y(n_6662)
);

INVx2_ASAP7_75t_L g6663 ( 
.A(n_6190),
.Y(n_6663)
);

INVx1_ASAP7_75t_L g6664 ( 
.A(n_6193),
.Y(n_6664)
);

CKINVDCx5p33_ASAP7_75t_R g6665 ( 
.A(n_6304),
.Y(n_6665)
);

AND2x4_ASAP7_75t_L g6666 ( 
.A(n_6432),
.B(n_6356),
.Y(n_6666)
);

NAND2xp5_ASAP7_75t_SL g6667 ( 
.A(n_6457),
.B(n_6061),
.Y(n_6667)
);

INVx3_ASAP7_75t_L g6668 ( 
.A(n_6532),
.Y(n_6668)
);

INVx2_ASAP7_75t_L g6669 ( 
.A(n_6196),
.Y(n_6669)
);

INVx2_ASAP7_75t_L g6670 ( 
.A(n_6212),
.Y(n_6670)
);

INVx5_ASAP7_75t_L g6671 ( 
.A(n_6226),
.Y(n_6671)
);

OR2x6_ASAP7_75t_L g6672 ( 
.A(n_6226),
.B(n_6302),
.Y(n_6672)
);

INVx2_ASAP7_75t_L g6673 ( 
.A(n_6234),
.Y(n_6673)
);

NOR2xp33_ASAP7_75t_SL g6674 ( 
.A(n_6337),
.B(n_5721),
.Y(n_6674)
);

INVx1_ASAP7_75t_L g6675 ( 
.A(n_6235),
.Y(n_6675)
);

OR2x6_ASAP7_75t_L g6676 ( 
.A(n_6194),
.B(n_5745),
.Y(n_6676)
);

INVx1_ASAP7_75t_L g6677 ( 
.A(n_6236),
.Y(n_6677)
);

INVx1_ASAP7_75t_L g6678 ( 
.A(n_6245),
.Y(n_6678)
);

NOR2xp33_ASAP7_75t_L g6679 ( 
.A(n_6207),
.B(n_5802),
.Y(n_6679)
);

HB1xp67_ASAP7_75t_L g6680 ( 
.A(n_6323),
.Y(n_6680)
);

INVx1_ASAP7_75t_L g6681 ( 
.A(n_6251),
.Y(n_6681)
);

AND2x6_ASAP7_75t_L g6682 ( 
.A(n_6594),
.B(n_6159),
.Y(n_6682)
);

BUFx2_ASAP7_75t_L g6683 ( 
.A(n_6427),
.Y(n_6683)
);

HB1xp67_ASAP7_75t_L g6684 ( 
.A(n_6221),
.Y(n_6684)
);

INVx1_ASAP7_75t_L g6685 ( 
.A(n_6259),
.Y(n_6685)
);

BUFx6f_ASAP7_75t_L g6686 ( 
.A(n_6487),
.Y(n_6686)
);

NAND2xp5_ASAP7_75t_L g6687 ( 
.A(n_6340),
.B(n_5796),
.Y(n_6687)
);

NAND2xp5_ASAP7_75t_L g6688 ( 
.A(n_6232),
.B(n_5893),
.Y(n_6688)
);

INVx2_ASAP7_75t_L g6689 ( 
.A(n_6263),
.Y(n_6689)
);

INVx1_ASAP7_75t_L g6690 ( 
.A(n_6273),
.Y(n_6690)
);

INVx1_ASAP7_75t_L g6691 ( 
.A(n_6280),
.Y(n_6691)
);

AOI22xp5_ASAP7_75t_L g6692 ( 
.A1(n_6516),
.A2(n_5943),
.B1(n_5882),
.B2(n_6185),
.Y(n_6692)
);

BUFx4f_ASAP7_75t_L g6693 ( 
.A(n_6487),
.Y(n_6693)
);

BUFx2_ASAP7_75t_L g6694 ( 
.A(n_6306),
.Y(n_6694)
);

NOR2xp33_ASAP7_75t_L g6695 ( 
.A(n_6220),
.B(n_5764),
.Y(n_6695)
);

INVx1_ASAP7_75t_L g6696 ( 
.A(n_6300),
.Y(n_6696)
);

INVx2_ASAP7_75t_L g6697 ( 
.A(n_6307),
.Y(n_6697)
);

BUFx3_ASAP7_75t_L g6698 ( 
.A(n_6327),
.Y(n_6698)
);

NAND2xp5_ASAP7_75t_L g6699 ( 
.A(n_6233),
.B(n_5902),
.Y(n_6699)
);

INVx1_ASAP7_75t_L g6700 ( 
.A(n_6316),
.Y(n_6700)
);

BUFx6f_ASAP7_75t_L g6701 ( 
.A(n_6279),
.Y(n_6701)
);

O2A1O1Ixp33_ASAP7_75t_L g6702 ( 
.A1(n_6215),
.A2(n_5939),
.B(n_5850),
.C(n_6158),
.Y(n_6702)
);

CKINVDCx8_ASAP7_75t_R g6703 ( 
.A(n_6458),
.Y(n_6703)
);

AOI22xp33_ASAP7_75t_L g6704 ( 
.A1(n_6538),
.A2(n_5933),
.B1(n_5971),
.B2(n_5948),
.Y(n_6704)
);

INVx2_ASAP7_75t_SL g6705 ( 
.A(n_6327),
.Y(n_6705)
);

NOR2xp33_ASAP7_75t_L g6706 ( 
.A(n_6390),
.B(n_6049),
.Y(n_6706)
);

AOI22xp33_ASAP7_75t_L g6707 ( 
.A1(n_6338),
.A2(n_6032),
.B1(n_6039),
.B2(n_6080),
.Y(n_6707)
);

INVx2_ASAP7_75t_L g6708 ( 
.A(n_6318),
.Y(n_6708)
);

INVx1_ASAP7_75t_L g6709 ( 
.A(n_6328),
.Y(n_6709)
);

INVx1_ASAP7_75t_L g6710 ( 
.A(n_6336),
.Y(n_6710)
);

INVx1_ASAP7_75t_L g6711 ( 
.A(n_6384),
.Y(n_6711)
);

A2O1A1Ixp33_ASAP7_75t_L g6712 ( 
.A1(n_6230),
.A2(n_5794),
.B(n_5901),
.C(n_6121),
.Y(n_6712)
);

NAND2xp5_ASAP7_75t_L g6713 ( 
.A(n_6202),
.B(n_6254),
.Y(n_6713)
);

AOI22xp33_ASAP7_75t_L g6714 ( 
.A1(n_6348),
.A2(n_6069),
.B1(n_6083),
.B2(n_6133),
.Y(n_6714)
);

INVx3_ASAP7_75t_L g6715 ( 
.A(n_6502),
.Y(n_6715)
);

NAND2xp5_ASAP7_75t_SL g6716 ( 
.A(n_6322),
.B(n_5689),
.Y(n_6716)
);

NAND2x1p5_ASAP7_75t_L g6717 ( 
.A(n_6242),
.B(n_1076),
.Y(n_6717)
);

INVx3_ASAP7_75t_L g6718 ( 
.A(n_6435),
.Y(n_6718)
);

INVx1_ASAP7_75t_L g6719 ( 
.A(n_6394),
.Y(n_6719)
);

INVx1_ASAP7_75t_L g6720 ( 
.A(n_6404),
.Y(n_6720)
);

INVx1_ASAP7_75t_L g6721 ( 
.A(n_6406),
.Y(n_6721)
);

AOI22xp5_ASAP7_75t_L g6722 ( 
.A1(n_6484),
.A2(n_1078),
.B1(n_1079),
.B2(n_1077),
.Y(n_6722)
);

AND2x4_ASAP7_75t_L g6723 ( 
.A(n_6658),
.B(n_1078),
.Y(n_6723)
);

AND2x2_ASAP7_75t_L g6724 ( 
.A(n_6450),
.B(n_1079),
.Y(n_6724)
);

BUFx6f_ASAP7_75t_L g6725 ( 
.A(n_6279),
.Y(n_6725)
);

AOI22xp33_ASAP7_75t_L g6726 ( 
.A1(n_6218),
.A2(n_16),
.B1(n_13),
.B2(n_15),
.Y(n_6726)
);

INVx2_ASAP7_75t_L g6727 ( 
.A(n_6415),
.Y(n_6727)
);

INVx3_ASAP7_75t_L g6728 ( 
.A(n_6284),
.Y(n_6728)
);

INVx1_ASAP7_75t_L g6729 ( 
.A(n_6419),
.Y(n_6729)
);

AOI22xp5_ASAP7_75t_L g6730 ( 
.A1(n_6282),
.A2(n_1082),
.B1(n_1083),
.B2(n_1081),
.Y(n_6730)
);

NAND2xp5_ASAP7_75t_SL g6731 ( 
.A(n_6558),
.B(n_1084),
.Y(n_6731)
);

BUFx6f_ASAP7_75t_L g6732 ( 
.A(n_6242),
.Y(n_6732)
);

AOI22xp33_ASAP7_75t_L g6733 ( 
.A1(n_6239),
.A2(n_16),
.B1(n_13),
.B2(n_15),
.Y(n_6733)
);

INVx1_ASAP7_75t_L g6734 ( 
.A(n_6424),
.Y(n_6734)
);

BUFx2_ASAP7_75t_L g6735 ( 
.A(n_6291),
.Y(n_6735)
);

AOI22xp33_ASAP7_75t_L g6736 ( 
.A1(n_6470),
.A2(n_6543),
.B1(n_6398),
.B2(n_6191),
.Y(n_6736)
);

NAND2xp5_ASAP7_75t_L g6737 ( 
.A(n_6297),
.B(n_15),
.Y(n_6737)
);

BUFx2_ASAP7_75t_L g6738 ( 
.A(n_6320),
.Y(n_6738)
);

INVx1_ASAP7_75t_L g6739 ( 
.A(n_6438),
.Y(n_6739)
);

BUFx6f_ASAP7_75t_L g6740 ( 
.A(n_6242),
.Y(n_6740)
);

NAND2xp5_ASAP7_75t_SL g6741 ( 
.A(n_6614),
.B(n_1085),
.Y(n_6741)
);

INVx2_ASAP7_75t_L g6742 ( 
.A(n_6448),
.Y(n_6742)
);

INVx4_ASAP7_75t_L g6743 ( 
.A(n_6327),
.Y(n_6743)
);

BUFx2_ASAP7_75t_SL g6744 ( 
.A(n_6458),
.Y(n_6744)
);

BUFx12f_ASAP7_75t_SL g6745 ( 
.A(n_6492),
.Y(n_6745)
);

INVx3_ASAP7_75t_L g6746 ( 
.A(n_6624),
.Y(n_6746)
);

INVx5_ASAP7_75t_L g6747 ( 
.A(n_6624),
.Y(n_6747)
);

INVx2_ASAP7_75t_L g6748 ( 
.A(n_6455),
.Y(n_6748)
);

OR2x6_ASAP7_75t_L g6749 ( 
.A(n_6199),
.B(n_6237),
.Y(n_6749)
);

NAND2xp5_ASAP7_75t_L g6750 ( 
.A(n_6208),
.B(n_17),
.Y(n_6750)
);

INVx1_ASAP7_75t_L g6751 ( 
.A(n_6471),
.Y(n_6751)
);

INVx2_ASAP7_75t_L g6752 ( 
.A(n_6472),
.Y(n_6752)
);

NAND2x1p5_ASAP7_75t_L g6753 ( 
.A(n_6458),
.B(n_1086),
.Y(n_6753)
);

INVx2_ASAP7_75t_L g6754 ( 
.A(n_6482),
.Y(n_6754)
);

NAND2xp5_ASAP7_75t_L g6755 ( 
.A(n_6210),
.B(n_18),
.Y(n_6755)
);

AND2x6_ASAP7_75t_L g6756 ( 
.A(n_6373),
.B(n_19),
.Y(n_6756)
);

INVx1_ASAP7_75t_SL g6757 ( 
.A(n_6355),
.Y(n_6757)
);

INVx2_ASAP7_75t_L g6758 ( 
.A(n_6500),
.Y(n_6758)
);

AOI22xp5_ASAP7_75t_L g6759 ( 
.A1(n_6228),
.A2(n_1087),
.B1(n_1089),
.B2(n_1086),
.Y(n_6759)
);

INVx2_ASAP7_75t_L g6760 ( 
.A(n_6513),
.Y(n_6760)
);

INVx1_ASAP7_75t_L g6761 ( 
.A(n_6296),
.Y(n_6761)
);

BUFx12f_ASAP7_75t_L g6762 ( 
.A(n_6644),
.Y(n_6762)
);

INVx1_ASAP7_75t_L g6763 ( 
.A(n_6376),
.Y(n_6763)
);

AND2x4_ASAP7_75t_L g6764 ( 
.A(n_6387),
.B(n_1089),
.Y(n_6764)
);

BUFx4f_ASAP7_75t_SL g6765 ( 
.A(n_6530),
.Y(n_6765)
);

HB1xp67_ASAP7_75t_L g6766 ( 
.A(n_6368),
.Y(n_6766)
);

HB1xp67_ASAP7_75t_L g6767 ( 
.A(n_6276),
.Y(n_6767)
);

BUFx3_ASAP7_75t_L g6768 ( 
.A(n_6414),
.Y(n_6768)
);

INVx2_ASAP7_75t_SL g6769 ( 
.A(n_6649),
.Y(n_6769)
);

AND2x4_ASAP7_75t_L g6770 ( 
.A(n_6443),
.B(n_1090),
.Y(n_6770)
);

NAND2xp5_ASAP7_75t_L g6771 ( 
.A(n_6213),
.B(n_6222),
.Y(n_6771)
);

OR2x4_ASAP7_75t_L g6772 ( 
.A(n_6268),
.B(n_19),
.Y(n_6772)
);

INVx1_ASAP7_75t_L g6773 ( 
.A(n_6396),
.Y(n_6773)
);

AND3x1_ASAP7_75t_SL g6774 ( 
.A(n_6621),
.B(n_19),
.C(n_20),
.Y(n_6774)
);

INVx2_ASAP7_75t_L g6775 ( 
.A(n_6525),
.Y(n_6775)
);

AND2x2_ASAP7_75t_L g6776 ( 
.A(n_6511),
.B(n_1090),
.Y(n_6776)
);

INVx1_ASAP7_75t_L g6777 ( 
.A(n_6447),
.Y(n_6777)
);

CKINVDCx5p33_ASAP7_75t_R g6778 ( 
.A(n_6420),
.Y(n_6778)
);

INVx1_ASAP7_75t_L g6779 ( 
.A(n_6460),
.Y(n_6779)
);

INVx1_ASAP7_75t_L g6780 ( 
.A(n_6526),
.Y(n_6780)
);

INVx1_ASAP7_75t_L g6781 ( 
.A(n_6536),
.Y(n_6781)
);

BUFx6f_ASAP7_75t_L g6782 ( 
.A(n_6649),
.Y(n_6782)
);

INVx1_ASAP7_75t_L g6783 ( 
.A(n_6546),
.Y(n_6783)
);

NAND2xp5_ASAP7_75t_SL g6784 ( 
.A(n_6374),
.B(n_1091),
.Y(n_6784)
);

NAND2xp5_ASAP7_75t_L g6785 ( 
.A(n_6562),
.B(n_20),
.Y(n_6785)
);

INVxp67_ASAP7_75t_L g6786 ( 
.A(n_6405),
.Y(n_6786)
);

INVx2_ASAP7_75t_L g6787 ( 
.A(n_6544),
.Y(n_6787)
);

BUFx6f_ASAP7_75t_L g6788 ( 
.A(n_6357),
.Y(n_6788)
);

INVx1_ASAP7_75t_L g6789 ( 
.A(n_6391),
.Y(n_6789)
);

INVx2_ASAP7_75t_L g6790 ( 
.A(n_6557),
.Y(n_6790)
);

BUFx6f_ASAP7_75t_L g6791 ( 
.A(n_6265),
.Y(n_6791)
);

NAND2x1p5_ASAP7_75t_L g6792 ( 
.A(n_6478),
.B(n_1092),
.Y(n_6792)
);

BUFx6f_ASAP7_75t_L g6793 ( 
.A(n_6446),
.Y(n_6793)
);

AND2x2_ASAP7_75t_L g6794 ( 
.A(n_6434),
.B(n_1093),
.Y(n_6794)
);

AOI22xp33_ASAP7_75t_L g6795 ( 
.A1(n_6626),
.A2(n_22),
.B1(n_20),
.B2(n_21),
.Y(n_6795)
);

NAND2xp5_ASAP7_75t_L g6796 ( 
.A(n_6547),
.B(n_21),
.Y(n_6796)
);

INVx1_ASAP7_75t_L g6797 ( 
.A(n_6461),
.Y(n_6797)
);

INVx1_ASAP7_75t_L g6798 ( 
.A(n_6520),
.Y(n_6798)
);

NOR2xp33_ASAP7_75t_L g6799 ( 
.A(n_6219),
.B(n_1093),
.Y(n_6799)
);

INVx2_ASAP7_75t_L g6800 ( 
.A(n_6201),
.Y(n_6800)
);

AOI22xp5_ASAP7_75t_L g6801 ( 
.A1(n_6591),
.A2(n_1095),
.B1(n_1096),
.B2(n_1094),
.Y(n_6801)
);

NAND2xp5_ASAP7_75t_L g6802 ( 
.A(n_6214),
.B(n_6401),
.Y(n_6802)
);

NAND2xp5_ASAP7_75t_SL g6803 ( 
.A(n_6288),
.B(n_1094),
.Y(n_6803)
);

INVx6_ASAP7_75t_L g6804 ( 
.A(n_6324),
.Y(n_6804)
);

BUFx4f_ASAP7_75t_L g6805 ( 
.A(n_6515),
.Y(n_6805)
);

INVx5_ASAP7_75t_L g6806 ( 
.A(n_6324),
.Y(n_6806)
);

CKINVDCx5p33_ASAP7_75t_R g6807 ( 
.A(n_6586),
.Y(n_6807)
);

INVx2_ASAP7_75t_L g6808 ( 
.A(n_6209),
.Y(n_6808)
);

INVx1_ASAP7_75t_L g6809 ( 
.A(n_6521),
.Y(n_6809)
);

INVx4_ASAP7_75t_L g6810 ( 
.A(n_6507),
.Y(n_6810)
);

INVx2_ASAP7_75t_SL g6811 ( 
.A(n_6388),
.Y(n_6811)
);

INVx1_ASAP7_75t_L g6812 ( 
.A(n_6522),
.Y(n_6812)
);

AOI22xp33_ASAP7_75t_SL g6813 ( 
.A1(n_6659),
.A2(n_1099),
.B1(n_1100),
.B2(n_1097),
.Y(n_6813)
);

BUFx2_ASAP7_75t_L g6814 ( 
.A(n_6618),
.Y(n_6814)
);

BUFx6f_ASAP7_75t_L g6815 ( 
.A(n_6324),
.Y(n_6815)
);

INVx3_ASAP7_75t_SL g6816 ( 
.A(n_6640),
.Y(n_6816)
);

NAND2xp5_ASAP7_75t_L g6817 ( 
.A(n_6195),
.B(n_21),
.Y(n_6817)
);

INVx1_ASAP7_75t_SL g6818 ( 
.A(n_6241),
.Y(n_6818)
);

INVxp67_ASAP7_75t_L g6819 ( 
.A(n_6258),
.Y(n_6819)
);

INVx4_ASAP7_75t_L g6820 ( 
.A(n_6507),
.Y(n_6820)
);

INVx4_ASAP7_75t_L g6821 ( 
.A(n_6507),
.Y(n_6821)
);

BUFx3_ASAP7_75t_L g6822 ( 
.A(n_6647),
.Y(n_6822)
);

HB1xp67_ASAP7_75t_L g6823 ( 
.A(n_6545),
.Y(n_6823)
);

AND2x4_ASAP7_75t_L g6824 ( 
.A(n_6496),
.B(n_1097),
.Y(n_6824)
);

BUFx8_ASAP7_75t_L g6825 ( 
.A(n_6211),
.Y(n_6825)
);

INVx1_ASAP7_75t_L g6826 ( 
.A(n_6216),
.Y(n_6826)
);

INVx2_ASAP7_75t_L g6827 ( 
.A(n_6225),
.Y(n_6827)
);

NAND2xp5_ASAP7_75t_SL g6828 ( 
.A(n_6416),
.B(n_6620),
.Y(n_6828)
);

NAND2xp5_ASAP7_75t_SL g6829 ( 
.A(n_6252),
.B(n_1099),
.Y(n_6829)
);

NOR2xp67_ASAP7_75t_L g6830 ( 
.A(n_6421),
.B(n_22),
.Y(n_6830)
);

NOR2x1_ASAP7_75t_R g6831 ( 
.A(n_6636),
.B(n_1100),
.Y(n_6831)
);

BUFx4f_ASAP7_75t_L g6832 ( 
.A(n_6351),
.Y(n_6832)
);

NAND2xp5_ASAP7_75t_SL g6833 ( 
.A(n_6610),
.B(n_1101),
.Y(n_6833)
);

AOI22xp5_ASAP7_75t_L g6834 ( 
.A1(n_6261),
.A2(n_1102),
.B1(n_1103),
.B2(n_1101),
.Y(n_6834)
);

INVx1_ASAP7_75t_L g6835 ( 
.A(n_6267),
.Y(n_6835)
);

INVx2_ASAP7_75t_L g6836 ( 
.A(n_6270),
.Y(n_6836)
);

INVx1_ASAP7_75t_L g6837 ( 
.A(n_6272),
.Y(n_6837)
);

AND2x2_ASAP7_75t_L g6838 ( 
.A(n_6332),
.B(n_1102),
.Y(n_6838)
);

AND2x4_ASAP7_75t_L g6839 ( 
.A(n_6555),
.B(n_1104),
.Y(n_6839)
);

INVx5_ASAP7_75t_L g6840 ( 
.A(n_6227),
.Y(n_6840)
);

OR2x6_ASAP7_75t_L g6841 ( 
.A(n_6573),
.B(n_1108),
.Y(n_6841)
);

BUFx2_ASAP7_75t_L g6842 ( 
.A(n_6616),
.Y(n_6842)
);

BUFx4f_ASAP7_75t_L g6843 ( 
.A(n_6351),
.Y(n_6843)
);

BUFx3_ASAP7_75t_L g6844 ( 
.A(n_6278),
.Y(n_6844)
);

NOR2xp33_ASAP7_75t_L g6845 ( 
.A(n_6341),
.B(n_1108),
.Y(n_6845)
);

CKINVDCx8_ASAP7_75t_R g6846 ( 
.A(n_6468),
.Y(n_6846)
);

AOI22xp33_ASAP7_75t_L g6847 ( 
.A1(n_6537),
.A2(n_24),
.B1(n_22),
.B2(n_23),
.Y(n_6847)
);

INVx1_ASAP7_75t_SL g6848 ( 
.A(n_6397),
.Y(n_6848)
);

NAND2xp5_ASAP7_75t_L g6849 ( 
.A(n_6197),
.B(n_23),
.Y(n_6849)
);

INVx2_ASAP7_75t_L g6850 ( 
.A(n_6294),
.Y(n_6850)
);

INVxp67_ASAP7_75t_L g6851 ( 
.A(n_6552),
.Y(n_6851)
);

NOR2x1p5_ASAP7_75t_L g6852 ( 
.A(n_6653),
.B(n_6574),
.Y(n_6852)
);

INVx1_ASAP7_75t_L g6853 ( 
.A(n_6312),
.Y(n_6853)
);

HB1xp67_ASAP7_75t_L g6854 ( 
.A(n_6290),
.Y(n_6854)
);

AND2x4_ASAP7_75t_SL g6855 ( 
.A(n_6578),
.B(n_1109),
.Y(n_6855)
);

BUFx3_ASAP7_75t_L g6856 ( 
.A(n_6326),
.Y(n_6856)
);

NAND2xp5_ASAP7_75t_SL g6857 ( 
.A(n_6431),
.B(n_1109),
.Y(n_6857)
);

INVxp67_ASAP7_75t_SL g6858 ( 
.A(n_6449),
.Y(n_6858)
);

BUFx6f_ASAP7_75t_L g6859 ( 
.A(n_6335),
.Y(n_6859)
);

INVx1_ASAP7_75t_L g6860 ( 
.A(n_6315),
.Y(n_6860)
);

INVx1_ASAP7_75t_L g6861 ( 
.A(n_6339),
.Y(n_6861)
);

INVx2_ASAP7_75t_SL g6862 ( 
.A(n_6359),
.Y(n_6862)
);

INVx3_ASAP7_75t_L g6863 ( 
.A(n_6559),
.Y(n_6863)
);

AOI22xp5_ASAP7_75t_L g6864 ( 
.A1(n_6371),
.A2(n_1111),
.B1(n_1112),
.B2(n_1110),
.Y(n_6864)
);

BUFx2_ASAP7_75t_L g6865 ( 
.A(n_6285),
.Y(n_6865)
);

INVx1_ASAP7_75t_L g6866 ( 
.A(n_6354),
.Y(n_6866)
);

NAND2xp5_ASAP7_75t_L g6867 ( 
.A(n_6292),
.B(n_23),
.Y(n_6867)
);

BUFx3_ASAP7_75t_L g6868 ( 
.A(n_6581),
.Y(n_6868)
);

BUFx3_ASAP7_75t_L g6869 ( 
.A(n_6353),
.Y(n_6869)
);

AND2x4_ASAP7_75t_L g6870 ( 
.A(n_6595),
.B(n_1113),
.Y(n_6870)
);

INVx1_ASAP7_75t_L g6871 ( 
.A(n_6364),
.Y(n_6871)
);

HB1xp67_ASAP7_75t_L g6872 ( 
.A(n_6608),
.Y(n_6872)
);

BUFx3_ASAP7_75t_L g6873 ( 
.A(n_6309),
.Y(n_6873)
);

INVx1_ASAP7_75t_L g6874 ( 
.A(n_6400),
.Y(n_6874)
);

AOI22xp33_ASAP7_75t_L g6875 ( 
.A1(n_6650),
.A2(n_26),
.B1(n_24),
.B2(n_25),
.Y(n_6875)
);

NAND2xp5_ASAP7_75t_L g6876 ( 
.A(n_6271),
.B(n_24),
.Y(n_6876)
);

NAND2xp5_ASAP7_75t_L g6877 ( 
.A(n_6333),
.B(n_25),
.Y(n_6877)
);

INVx2_ASAP7_75t_L g6878 ( 
.A(n_6403),
.Y(n_6878)
);

INVx2_ASAP7_75t_L g6879 ( 
.A(n_6411),
.Y(n_6879)
);

NOR2xp33_ASAP7_75t_L g6880 ( 
.A(n_6334),
.B(n_1114),
.Y(n_6880)
);

INVx1_ASAP7_75t_L g6881 ( 
.A(n_6413),
.Y(n_6881)
);

AOI22xp33_ASAP7_75t_L g6882 ( 
.A1(n_6198),
.A2(n_27),
.B1(n_25),
.B2(n_26),
.Y(n_6882)
);

BUFx2_ASAP7_75t_R g6883 ( 
.A(n_6499),
.Y(n_6883)
);

NOR2xp33_ASAP7_75t_L g6884 ( 
.A(n_6203),
.B(n_1114),
.Y(n_6884)
);

AOI21xp5_ASAP7_75t_L g6885 ( 
.A1(n_6247),
.A2(n_1116),
.B(n_1115),
.Y(n_6885)
);

INVx1_ASAP7_75t_L g6886 ( 
.A(n_6423),
.Y(n_6886)
);

HB1xp67_ASAP7_75t_L g6887 ( 
.A(n_6563),
.Y(n_6887)
);

INVx1_ASAP7_75t_L g6888 ( 
.A(n_6454),
.Y(n_6888)
);

AND2x4_ASAP7_75t_SL g6889 ( 
.A(n_6603),
.B(n_1116),
.Y(n_6889)
);

INVx2_ASAP7_75t_L g6890 ( 
.A(n_6480),
.Y(n_6890)
);

AOI22xp33_ASAP7_75t_L g6891 ( 
.A1(n_6345),
.A2(n_28),
.B1(n_26),
.B2(n_27),
.Y(n_6891)
);

INVx2_ASAP7_75t_L g6892 ( 
.A(n_6483),
.Y(n_6892)
);

OAI22xp5_ASAP7_75t_L g6893 ( 
.A1(n_6329),
.A2(n_1118),
.B1(n_1119),
.B2(n_1117),
.Y(n_6893)
);

AOI22xp33_ASAP7_75t_L g6894 ( 
.A1(n_6343),
.A2(n_29),
.B1(n_27),
.B2(n_28),
.Y(n_6894)
);

NAND2xp5_ASAP7_75t_SL g6895 ( 
.A(n_6548),
.B(n_1117),
.Y(n_6895)
);

INVx5_ASAP7_75t_L g6896 ( 
.A(n_6227),
.Y(n_6896)
);

INVx3_ASAP7_75t_L g6897 ( 
.A(n_6631),
.Y(n_6897)
);

INVx1_ASAP7_75t_L g6898 ( 
.A(n_6504),
.Y(n_6898)
);

NOR2xp33_ASAP7_75t_L g6899 ( 
.A(n_6325),
.B(n_1118),
.Y(n_6899)
);

NAND2xp5_ASAP7_75t_L g6900 ( 
.A(n_6231),
.B(n_28),
.Y(n_6900)
);

INVx4_ASAP7_75t_L g6901 ( 
.A(n_6249),
.Y(n_6901)
);

BUFx6f_ASAP7_75t_L g6902 ( 
.A(n_6596),
.Y(n_6902)
);

NAND2xp5_ASAP7_75t_L g6903 ( 
.A(n_6248),
.B(n_30),
.Y(n_6903)
);

OAI22xp5_ASAP7_75t_SL g6904 ( 
.A1(n_6321),
.A2(n_32),
.B1(n_30),
.B2(n_31),
.Y(n_6904)
);

INVx1_ASAP7_75t_L g6905 ( 
.A(n_6564),
.Y(n_6905)
);

AND2x4_ASAP7_75t_SL g6906 ( 
.A(n_6599),
.B(n_6627),
.Y(n_6906)
);

BUFx3_ASAP7_75t_L g6907 ( 
.A(n_6654),
.Y(n_6907)
);

CKINVDCx20_ASAP7_75t_R g6908 ( 
.A(n_6425),
.Y(n_6908)
);

NAND2xp5_ASAP7_75t_L g6909 ( 
.A(n_6250),
.B(n_30),
.Y(n_6909)
);

AND2x4_ASAP7_75t_L g6910 ( 
.A(n_6629),
.B(n_1119),
.Y(n_6910)
);

INVx2_ASAP7_75t_L g6911 ( 
.A(n_6550),
.Y(n_6911)
);

INVx1_ASAP7_75t_L g6912 ( 
.A(n_6569),
.Y(n_6912)
);

INVx1_ASAP7_75t_SL g6913 ( 
.A(n_6588),
.Y(n_6913)
);

INVx2_ASAP7_75t_L g6914 ( 
.A(n_6589),
.Y(n_6914)
);

INVx5_ASAP7_75t_L g6915 ( 
.A(n_6249),
.Y(n_6915)
);

INVx1_ASAP7_75t_L g6916 ( 
.A(n_6612),
.Y(n_6916)
);

INVx5_ASAP7_75t_L g6917 ( 
.A(n_6567),
.Y(n_6917)
);

INVx2_ASAP7_75t_L g6918 ( 
.A(n_6633),
.Y(n_6918)
);

INVx4_ASAP7_75t_L g6919 ( 
.A(n_6238),
.Y(n_6919)
);

INVx2_ASAP7_75t_SL g6920 ( 
.A(n_6466),
.Y(n_6920)
);

NAND2xp5_ASAP7_75t_L g6921 ( 
.A(n_6399),
.B(n_31),
.Y(n_6921)
);

NAND2xp33_ASAP7_75t_SL g6922 ( 
.A(n_6395),
.B(n_1120),
.Y(n_6922)
);

NAND2xp5_ASAP7_75t_SL g6923 ( 
.A(n_6380),
.B(n_6382),
.Y(n_6923)
);

INVx2_ASAP7_75t_SL g6924 ( 
.A(n_6277),
.Y(n_6924)
);

INVx2_ASAP7_75t_L g6925 ( 
.A(n_6641),
.Y(n_6925)
);

INVx1_ASAP7_75t_SL g6926 ( 
.A(n_6262),
.Y(n_6926)
);

AOI221xp5_ASAP7_75t_SL g6927 ( 
.A1(n_6308),
.A2(n_6269),
.B1(n_6314),
.B2(n_6524),
.C(n_6246),
.Y(n_6927)
);

INVx1_ASAP7_75t_L g6928 ( 
.A(n_6503),
.Y(n_6928)
);

CKINVDCx5p33_ASAP7_75t_R g6929 ( 
.A(n_6481),
.Y(n_6929)
);

INVx1_ASAP7_75t_L g6930 ( 
.A(n_6506),
.Y(n_6930)
);

BUFx6f_ASAP7_75t_L g6931 ( 
.A(n_6501),
.Y(n_6931)
);

CKINVDCx5p33_ASAP7_75t_R g6932 ( 
.A(n_6393),
.Y(n_6932)
);

BUFx8_ASAP7_75t_L g6933 ( 
.A(n_6617),
.Y(n_6933)
);

CKINVDCx8_ASAP7_75t_R g6934 ( 
.A(n_6381),
.Y(n_6934)
);

AND2x2_ASAP7_75t_L g6935 ( 
.A(n_6571),
.B(n_1121),
.Y(n_6935)
);

NAND2x1p5_ASAP7_75t_L g6936 ( 
.A(n_6642),
.B(n_1121),
.Y(n_6936)
);

AND2x2_ASAP7_75t_L g6937 ( 
.A(n_6575),
.B(n_1122),
.Y(n_6937)
);

OAI22xp5_ASAP7_75t_L g6938 ( 
.A1(n_6402),
.A2(n_1123),
.B1(n_1124),
.B2(n_1122),
.Y(n_6938)
);

INVx2_ASAP7_75t_L g6939 ( 
.A(n_6508),
.Y(n_6939)
);

AOI22xp5_ASAP7_75t_L g6940 ( 
.A1(n_6352),
.A2(n_1125),
.B1(n_1126),
.B2(n_1124),
.Y(n_6940)
);

OR2x2_ASAP7_75t_L g6941 ( 
.A(n_6200),
.B(n_32),
.Y(n_6941)
);

AND2x4_ASAP7_75t_L g6942 ( 
.A(n_6358),
.B(n_1127),
.Y(n_6942)
);

NAND2xp5_ASAP7_75t_L g6943 ( 
.A(n_6287),
.B(n_33),
.Y(n_6943)
);

BUFx6f_ASAP7_75t_L g6944 ( 
.A(n_6660),
.Y(n_6944)
);

NAND2xp5_ASAP7_75t_L g6945 ( 
.A(n_6205),
.B(n_33),
.Y(n_6945)
);

NAND2xp5_ASAP7_75t_L g6946 ( 
.A(n_6473),
.B(n_33),
.Y(n_6946)
);

INVx2_ASAP7_75t_L g6947 ( 
.A(n_6509),
.Y(n_6947)
);

CKINVDCx5p33_ASAP7_75t_R g6948 ( 
.A(n_6613),
.Y(n_6948)
);

INVx1_ASAP7_75t_L g6949 ( 
.A(n_6533),
.Y(n_6949)
);

NOR2xp33_ASAP7_75t_L g6950 ( 
.A(n_6206),
.B(n_1128),
.Y(n_6950)
);

AND2x4_ASAP7_75t_L g6951 ( 
.A(n_6363),
.B(n_1128),
.Y(n_6951)
);

INVxp67_ASAP7_75t_L g6952 ( 
.A(n_6389),
.Y(n_6952)
);

NAND2xp5_ASAP7_75t_SL g6953 ( 
.A(n_6510),
.B(n_1129),
.Y(n_6953)
);

BUFx2_ASAP7_75t_L g6954 ( 
.A(n_6630),
.Y(n_6954)
);

INVx1_ASAP7_75t_L g6955 ( 
.A(n_6534),
.Y(n_6955)
);

INVx1_ASAP7_75t_L g6956 ( 
.A(n_6535),
.Y(n_6956)
);

INVx1_ASAP7_75t_L g6957 ( 
.A(n_6541),
.Y(n_6957)
);

BUFx2_ASAP7_75t_L g6958 ( 
.A(n_6656),
.Y(n_6958)
);

INVx1_ASAP7_75t_L g6959 ( 
.A(n_6519),
.Y(n_6959)
);

AOI22xp5_ASAP7_75t_L g6960 ( 
.A1(n_6565),
.A2(n_1130),
.B1(n_1131),
.B2(n_1129),
.Y(n_6960)
);

NAND2xp5_ASAP7_75t_L g6961 ( 
.A(n_6549),
.B(n_34),
.Y(n_6961)
);

INVx2_ASAP7_75t_SL g6962 ( 
.A(n_6361),
.Y(n_6962)
);

INVx1_ASAP7_75t_L g6963 ( 
.A(n_6561),
.Y(n_6963)
);

INVx2_ASAP7_75t_L g6964 ( 
.A(n_6463),
.Y(n_6964)
);

INVx2_ASAP7_75t_L g6965 ( 
.A(n_6465),
.Y(n_6965)
);

BUFx8_ASAP7_75t_L g6966 ( 
.A(n_6638),
.Y(n_6966)
);

INVx1_ASAP7_75t_L g6967 ( 
.A(n_6467),
.Y(n_6967)
);

NAND2xp5_ASAP7_75t_L g6968 ( 
.A(n_6256),
.B(n_34),
.Y(n_6968)
);

INVx5_ASAP7_75t_L g6969 ( 
.A(n_6567),
.Y(n_6969)
);

INVx4_ASAP7_75t_L g6970 ( 
.A(n_6651),
.Y(n_6970)
);

AOI22xp5_ASAP7_75t_L g6971 ( 
.A1(n_6299),
.A2(n_1132),
.B1(n_1133),
.B2(n_1130),
.Y(n_6971)
);

CKINVDCx5p33_ASAP7_75t_R g6972 ( 
.A(n_6493),
.Y(n_6972)
);

INVx1_ASAP7_75t_L g6973 ( 
.A(n_6469),
.Y(n_6973)
);

OR2x6_ASAP7_75t_L g6974 ( 
.A(n_6260),
.B(n_1132),
.Y(n_6974)
);

NOR2xp33_ASAP7_75t_L g6975 ( 
.A(n_6553),
.B(n_1134),
.Y(n_6975)
);

AND2x4_ASAP7_75t_L g6976 ( 
.A(n_6582),
.B(n_1134),
.Y(n_6976)
);

INVx5_ASAP7_75t_L g6977 ( 
.A(n_6189),
.Y(n_6977)
);

INVx2_ASAP7_75t_L g6978 ( 
.A(n_6475),
.Y(n_6978)
);

INVx2_ASAP7_75t_SL g6979 ( 
.A(n_6474),
.Y(n_6979)
);

INVx1_ASAP7_75t_L g6980 ( 
.A(n_6476),
.Y(n_6980)
);

AOI22xp33_ASAP7_75t_L g6981 ( 
.A1(n_6628),
.A2(n_37),
.B1(n_35),
.B2(n_36),
.Y(n_6981)
);

INVx1_ASAP7_75t_L g6982 ( 
.A(n_6488),
.Y(n_6982)
);

INVx2_ASAP7_75t_SL g6983 ( 
.A(n_6577),
.Y(n_6983)
);

HB1xp67_ASAP7_75t_L g6984 ( 
.A(n_6409),
.Y(n_6984)
);

CKINVDCx5p33_ASAP7_75t_R g6985 ( 
.A(n_6310),
.Y(n_6985)
);

INVx1_ASAP7_75t_L g6986 ( 
.A(n_6491),
.Y(n_6986)
);

NAND3xp33_ASAP7_75t_SL g6987 ( 
.A(n_6255),
.B(n_35),
.C(n_36),
.Y(n_6987)
);

NAND2xp5_ASAP7_75t_L g6988 ( 
.A(n_6257),
.B(n_36),
.Y(n_6988)
);

INVx3_ASAP7_75t_L g6989 ( 
.A(n_6609),
.Y(n_6989)
);

INVx2_ASAP7_75t_L g6990 ( 
.A(n_6494),
.Y(n_6990)
);

BUFx6f_ASAP7_75t_L g6991 ( 
.A(n_6428),
.Y(n_6991)
);

NOR2xp33_ASAP7_75t_L g6992 ( 
.A(n_6490),
.B(n_1135),
.Y(n_6992)
);

NOR2xp33_ASAP7_75t_L g6993 ( 
.A(n_6568),
.B(n_1135),
.Y(n_6993)
);

BUFx3_ASAP7_75t_L g6994 ( 
.A(n_6623),
.Y(n_6994)
);

INVx1_ASAP7_75t_L g6995 ( 
.A(n_6497),
.Y(n_6995)
);

INVx1_ASAP7_75t_L g6996 ( 
.A(n_6542),
.Y(n_6996)
);

AND2x2_ASAP7_75t_L g6997 ( 
.A(n_6576),
.B(n_6240),
.Y(n_6997)
);

BUFx2_ASAP7_75t_L g6998 ( 
.A(n_6611),
.Y(n_6998)
);

INVx2_ASAP7_75t_L g6999 ( 
.A(n_6344),
.Y(n_6999)
);

BUFx6f_ASAP7_75t_L g7000 ( 
.A(n_6433),
.Y(n_7000)
);

AND2x4_ASAP7_75t_L g7001 ( 
.A(n_6592),
.B(n_1137),
.Y(n_7001)
);

NOR2xp33_ASAP7_75t_R g7002 ( 
.A(n_6527),
.B(n_1137),
.Y(n_7002)
);

BUFx3_ASAP7_75t_L g7003 ( 
.A(n_6652),
.Y(n_7003)
);

CKINVDCx5p33_ASAP7_75t_R g7004 ( 
.A(n_6637),
.Y(n_7004)
);

INVx1_ASAP7_75t_L g7005 ( 
.A(n_6346),
.Y(n_7005)
);

INVx1_ASAP7_75t_L g7006 ( 
.A(n_6347),
.Y(n_7006)
);

INVx1_ASAP7_75t_L g7007 ( 
.A(n_6407),
.Y(n_7007)
);

NOR2xp33_ASAP7_75t_R g7008 ( 
.A(n_6529),
.B(n_1138),
.Y(n_7008)
);

OR2x2_ASAP7_75t_L g7009 ( 
.A(n_6264),
.B(n_37),
.Y(n_7009)
);

BUFx2_ASAP7_75t_L g7010 ( 
.A(n_6607),
.Y(n_7010)
);

NAND2xp5_ASAP7_75t_L g7011 ( 
.A(n_6266),
.B(n_37),
.Y(n_7011)
);

BUFx3_ASAP7_75t_L g7012 ( 
.A(n_6625),
.Y(n_7012)
);

NAND2xp5_ASAP7_75t_L g7013 ( 
.A(n_6281),
.B(n_38),
.Y(n_7013)
);

INVx2_ASAP7_75t_SL g7014 ( 
.A(n_6331),
.Y(n_7014)
);

NAND2x1p5_ASAP7_75t_L g7015 ( 
.A(n_6489),
.B(n_1138),
.Y(n_7015)
);

CKINVDCx5p33_ASAP7_75t_R g7016 ( 
.A(n_6598),
.Y(n_7016)
);

BUFx12f_ASAP7_75t_L g7017 ( 
.A(n_6436),
.Y(n_7017)
);

OR2x6_ASAP7_75t_L g7018 ( 
.A(n_6601),
.B(n_1139),
.Y(n_7018)
);

INVx2_ASAP7_75t_L g7019 ( 
.A(n_6408),
.Y(n_7019)
);

OR2x2_ASAP7_75t_L g7020 ( 
.A(n_6286),
.B(n_38),
.Y(n_7020)
);

INVx1_ASAP7_75t_L g7021 ( 
.A(n_6410),
.Y(n_7021)
);

OR2x6_ASAP7_75t_L g7022 ( 
.A(n_6604),
.B(n_1139),
.Y(n_7022)
);

BUFx3_ASAP7_75t_L g7023 ( 
.A(n_6635),
.Y(n_7023)
);

INVx1_ASAP7_75t_SL g7024 ( 
.A(n_6572),
.Y(n_7024)
);

BUFx3_ASAP7_75t_L g7025 ( 
.A(n_6643),
.Y(n_7025)
);

BUFx5_ASAP7_75t_L g7026 ( 
.A(n_6479),
.Y(n_7026)
);

INVx3_ASAP7_75t_L g7027 ( 
.A(n_6580),
.Y(n_7027)
);

NOR2xp33_ASAP7_75t_L g7028 ( 
.A(n_6385),
.B(n_1140),
.Y(n_7028)
);

AND2x4_ASAP7_75t_L g7029 ( 
.A(n_6342),
.B(n_1140),
.Y(n_7029)
);

AND2x4_ASAP7_75t_L g7030 ( 
.A(n_6593),
.B(n_1141),
.Y(n_7030)
);

INVxp67_ASAP7_75t_SL g7031 ( 
.A(n_6417),
.Y(n_7031)
);

INVx1_ASAP7_75t_L g7032 ( 
.A(n_6422),
.Y(n_7032)
);

INVx1_ASAP7_75t_L g7033 ( 
.A(n_6426),
.Y(n_7033)
);

HB1xp67_ASAP7_75t_L g7034 ( 
.A(n_6622),
.Y(n_7034)
);

INVx1_ASAP7_75t_L g7035 ( 
.A(n_6429),
.Y(n_7035)
);

NAND2xp5_ASAP7_75t_L g7036 ( 
.A(n_6289),
.B(n_39),
.Y(n_7036)
);

NAND2xp5_ASAP7_75t_L g7037 ( 
.A(n_6293),
.B(n_39),
.Y(n_7037)
);

NAND2xp5_ASAP7_75t_SL g7038 ( 
.A(n_6319),
.B(n_1141),
.Y(n_7038)
);

INVx3_ASAP7_75t_L g7039 ( 
.A(n_6512),
.Y(n_7039)
);

NAND2xp5_ASAP7_75t_L g7040 ( 
.A(n_6298),
.B(n_6301),
.Y(n_7040)
);

INVx1_ASAP7_75t_L g7041 ( 
.A(n_6437),
.Y(n_7041)
);

INVx2_ASAP7_75t_L g7042 ( 
.A(n_6440),
.Y(n_7042)
);

INVx2_ASAP7_75t_L g7043 ( 
.A(n_6441),
.Y(n_7043)
);

INVx1_ASAP7_75t_L g7044 ( 
.A(n_6442),
.Y(n_7044)
);

NOR2xp33_ASAP7_75t_L g7045 ( 
.A(n_6275),
.B(n_1142),
.Y(n_7045)
);

INVx1_ASAP7_75t_L g7046 ( 
.A(n_6517),
.Y(n_7046)
);

NAND2xp5_ASAP7_75t_L g7047 ( 
.A(n_6303),
.B(n_6305),
.Y(n_7047)
);

INVx5_ASAP7_75t_L g7048 ( 
.A(n_6539),
.Y(n_7048)
);

INVx4_ASAP7_75t_L g7049 ( 
.A(n_6615),
.Y(n_7049)
);

INVx5_ASAP7_75t_L g7050 ( 
.A(n_6600),
.Y(n_7050)
);

INVx1_ASAP7_75t_L g7051 ( 
.A(n_6619),
.Y(n_7051)
);

INVx3_ASAP7_75t_L g7052 ( 
.A(n_6583),
.Y(n_7052)
);

INVx2_ASAP7_75t_SL g7053 ( 
.A(n_6274),
.Y(n_7053)
);

BUFx2_ASAP7_75t_L g7054 ( 
.A(n_6584),
.Y(n_7054)
);

BUFx3_ASAP7_75t_L g7055 ( 
.A(n_6590),
.Y(n_7055)
);

A2O1A1Ixp33_ASAP7_75t_L g7056 ( 
.A1(n_6439),
.A2(n_41),
.B(n_39),
.C(n_40),
.Y(n_7056)
);

BUFx6f_ASAP7_75t_L g7057 ( 
.A(n_6657),
.Y(n_7057)
);

NOR2x1_ASAP7_75t_L g7058 ( 
.A(n_6224),
.B(n_1142),
.Y(n_7058)
);

HB1xp67_ASAP7_75t_L g7059 ( 
.A(n_6639),
.Y(n_7059)
);

NAND2xp5_ASAP7_75t_SL g7060 ( 
.A(n_6350),
.B(n_6418),
.Y(n_7060)
);

INVx4_ASAP7_75t_L g7061 ( 
.A(n_6243),
.Y(n_7061)
);

INVx2_ASAP7_75t_SL g7062 ( 
.A(n_6523),
.Y(n_7062)
);

CKINVDCx20_ASAP7_75t_R g7063 ( 
.A(n_6531),
.Y(n_7063)
);

NOR2x1p5_ASAP7_75t_L g7064 ( 
.A(n_6606),
.B(n_1143),
.Y(n_7064)
);

NOR2xp67_ASAP7_75t_L g7065 ( 
.A(n_6444),
.B(n_40),
.Y(n_7065)
);

BUFx6f_ASAP7_75t_L g7066 ( 
.A(n_6646),
.Y(n_7066)
);

INVx1_ASAP7_75t_L g7067 ( 
.A(n_6311),
.Y(n_7067)
);

INVx2_ASAP7_75t_L g7068 ( 
.A(n_6445),
.Y(n_7068)
);

INVx1_ASAP7_75t_L g7069 ( 
.A(n_6365),
.Y(n_7069)
);

AOI22xp33_ASAP7_75t_L g7070 ( 
.A1(n_6204),
.A2(n_6655),
.B1(n_6645),
.B2(n_6566),
.Y(n_7070)
);

NOR2xp33_ASAP7_75t_L g7071 ( 
.A(n_6253),
.B(n_1143),
.Y(n_7071)
);

AND2x2_ASAP7_75t_L g7072 ( 
.A(n_6528),
.B(n_1144),
.Y(n_7072)
);

INVx5_ASAP7_75t_L g7073 ( 
.A(n_6217),
.Y(n_7073)
);

OAI21xp5_ASAP7_75t_L g7074 ( 
.A1(n_6378),
.A2(n_6392),
.B(n_6295),
.Y(n_7074)
);

NAND2xp5_ASAP7_75t_L g7075 ( 
.A(n_6367),
.B(n_40),
.Y(n_7075)
);

AND2x4_ASAP7_75t_L g7076 ( 
.A(n_6518),
.B(n_1144),
.Y(n_7076)
);

NAND2xp5_ASAP7_75t_L g7077 ( 
.A(n_6369),
.B(n_41),
.Y(n_7077)
);

INVx1_ASAP7_75t_L g7078 ( 
.A(n_6372),
.Y(n_7078)
);

INVx1_ASAP7_75t_L g7079 ( 
.A(n_6375),
.Y(n_7079)
);

CKINVDCx20_ASAP7_75t_R g7080 ( 
.A(n_6648),
.Y(n_7080)
);

NAND2xp5_ASAP7_75t_L g7081 ( 
.A(n_6377),
.B(n_41),
.Y(n_7081)
);

NAND2xp5_ASAP7_75t_L g7082 ( 
.A(n_6379),
.B(n_42),
.Y(n_7082)
);

INVx1_ASAP7_75t_L g7083 ( 
.A(n_6383),
.Y(n_7083)
);

INVx1_ASAP7_75t_L g7084 ( 
.A(n_6386),
.Y(n_7084)
);

BUFx8_ASAP7_75t_L g7085 ( 
.A(n_6597),
.Y(n_7085)
);

NAND2xp5_ASAP7_75t_L g7086 ( 
.A(n_6452),
.B(n_42),
.Y(n_7086)
);

INVx4_ASAP7_75t_L g7087 ( 
.A(n_6366),
.Y(n_7087)
);

OR2x2_ASAP7_75t_L g7088 ( 
.A(n_6453),
.B(n_42),
.Y(n_7088)
);

INVx2_ASAP7_75t_L g7089 ( 
.A(n_6456),
.Y(n_7089)
);

INVx1_ASAP7_75t_L g7090 ( 
.A(n_6551),
.Y(n_7090)
);

NAND2xp5_ASAP7_75t_L g7091 ( 
.A(n_6192),
.B(n_43),
.Y(n_7091)
);

INVxp67_ASAP7_75t_L g7092 ( 
.A(n_6605),
.Y(n_7092)
);

INVx5_ASAP7_75t_L g7093 ( 
.A(n_6634),
.Y(n_7093)
);

INVx2_ASAP7_75t_SL g7094 ( 
.A(n_6579),
.Y(n_7094)
);

INVx4_ASAP7_75t_SL g7095 ( 
.A(n_6632),
.Y(n_7095)
);

CKINVDCx8_ASAP7_75t_R g7096 ( 
.A(n_6540),
.Y(n_7096)
);

INVx1_ASAP7_75t_L g7097 ( 
.A(n_6570),
.Y(n_7097)
);

INVx2_ASAP7_75t_L g7098 ( 
.A(n_6229),
.Y(n_7098)
);

NAND2xp5_ASAP7_75t_SL g7099 ( 
.A(n_6313),
.B(n_1145),
.Y(n_7099)
);

NAND2xp5_ASAP7_75t_L g7100 ( 
.A(n_6486),
.B(n_43),
.Y(n_7100)
);

INVx3_ASAP7_75t_L g7101 ( 
.A(n_6485),
.Y(n_7101)
);

BUFx2_ASAP7_75t_L g7102 ( 
.A(n_6370),
.Y(n_7102)
);

OAI22xp5_ASAP7_75t_L g7103 ( 
.A1(n_6736),
.A2(n_6554),
.B1(n_6244),
.B2(n_6317),
.Y(n_7103)
);

NAND2xp5_ASAP7_75t_L g7104 ( 
.A(n_6713),
.B(n_6602),
.Y(n_7104)
);

BUFx3_ASAP7_75t_L g7105 ( 
.A(n_6747),
.Y(n_7105)
);

INVx1_ASAP7_75t_L g7106 ( 
.A(n_6663),
.Y(n_7106)
);

AOI21xp5_ASAP7_75t_L g7107 ( 
.A1(n_6771),
.A2(n_6283),
.B(n_6360),
.Y(n_7107)
);

AOI21xp5_ASAP7_75t_L g7108 ( 
.A1(n_6802),
.A2(n_6464),
.B(n_6330),
.Y(n_7108)
);

CKINVDCx5p33_ASAP7_75t_R g7109 ( 
.A(n_6665),
.Y(n_7109)
);

O2A1O1Ixp33_ASAP7_75t_L g7110 ( 
.A1(n_6884),
.A2(n_6556),
.B(n_6587),
.C(n_6585),
.Y(n_7110)
);

NOR2xp33_ASAP7_75t_L g7111 ( 
.A(n_7004),
.B(n_6498),
.Y(n_7111)
);

INVx2_ASAP7_75t_L g7112 ( 
.A(n_6669),
.Y(n_7112)
);

AOI21xp5_ASAP7_75t_L g7113 ( 
.A1(n_7040),
.A2(n_6495),
.B(n_6462),
.Y(n_7113)
);

NAND2xp33_ASAP7_75t_L g7114 ( 
.A(n_6796),
.B(n_6349),
.Y(n_7114)
);

AOI21xp5_ASAP7_75t_L g7115 ( 
.A1(n_7047),
.A2(n_7031),
.B(n_6997),
.Y(n_7115)
);

INVx1_ASAP7_75t_L g7116 ( 
.A(n_6670),
.Y(n_7116)
);

OR2x6_ASAP7_75t_L g7117 ( 
.A(n_6744),
.B(n_6560),
.Y(n_7117)
);

NAND2xp5_ASAP7_75t_L g7118 ( 
.A(n_6761),
.B(n_6362),
.Y(n_7118)
);

NAND2xp5_ASAP7_75t_L g7119 ( 
.A(n_6763),
.B(n_6412),
.Y(n_7119)
);

AND2x2_ASAP7_75t_L g7120 ( 
.A(n_7023),
.B(n_6430),
.Y(n_7120)
);

INVx1_ASAP7_75t_L g7121 ( 
.A(n_6673),
.Y(n_7121)
);

NAND2x1p5_ASAP7_75t_L g7122 ( 
.A(n_6806),
.B(n_6451),
.Y(n_7122)
);

INVx4_ASAP7_75t_L g7123 ( 
.A(n_6747),
.Y(n_7123)
);

A2O1A1Ixp33_ASAP7_75t_L g7124 ( 
.A1(n_6679),
.A2(n_6505),
.B(n_6514),
.C(n_6459),
.Y(n_7124)
);

INVxp67_ASAP7_75t_L g7125 ( 
.A(n_6680),
.Y(n_7125)
);

AOI21xp5_ASAP7_75t_L g7126 ( 
.A1(n_6857),
.A2(n_1146),
.B(n_1145),
.Y(n_7126)
);

INVx3_ASAP7_75t_L g7127 ( 
.A(n_6703),
.Y(n_7127)
);

AOI21xp5_ASAP7_75t_L g7128 ( 
.A1(n_7074),
.A2(n_1147),
.B(n_1146),
.Y(n_7128)
);

NOR2xp33_ASAP7_75t_L g7129 ( 
.A(n_6952),
.B(n_1147),
.Y(n_7129)
);

INVx1_ASAP7_75t_SL g7130 ( 
.A(n_6848),
.Y(n_7130)
);

AOI21xp5_ASAP7_75t_L g7131 ( 
.A1(n_6716),
.A2(n_1149),
.B(n_1148),
.Y(n_7131)
);

AND2x2_ASAP7_75t_L g7132 ( 
.A(n_6724),
.B(n_6776),
.Y(n_7132)
);

BUFx2_ASAP7_75t_L g7133 ( 
.A(n_6683),
.Y(n_7133)
);

INVx1_ASAP7_75t_L g7134 ( 
.A(n_6689),
.Y(n_7134)
);

INVx3_ASAP7_75t_L g7135 ( 
.A(n_6666),
.Y(n_7135)
);

INVx1_ASAP7_75t_L g7136 ( 
.A(n_6697),
.Y(n_7136)
);

INVx2_ASAP7_75t_L g7137 ( 
.A(n_6708),
.Y(n_7137)
);

O2A1O1Ixp33_ASAP7_75t_L g7138 ( 
.A1(n_6785),
.A2(n_46),
.B(n_44),
.C(n_45),
.Y(n_7138)
);

INVx2_ASAP7_75t_L g7139 ( 
.A(n_6727),
.Y(n_7139)
);

NOR2xp33_ASAP7_75t_L g7140 ( 
.A(n_6923),
.B(n_7016),
.Y(n_7140)
);

NAND2xp5_ASAP7_75t_SL g7141 ( 
.A(n_6994),
.B(n_1148),
.Y(n_7141)
);

AOI21x1_ASAP7_75t_L g7142 ( 
.A1(n_6829),
.A2(n_44),
.B(n_45),
.Y(n_7142)
);

NOR2xp33_ASAP7_75t_L g7143 ( 
.A(n_7025),
.B(n_1149),
.Y(n_7143)
);

BUFx2_ASAP7_75t_L g7144 ( 
.A(n_6814),
.Y(n_7144)
);

AND2x2_ASAP7_75t_L g7145 ( 
.A(n_6794),
.B(n_44),
.Y(n_7145)
);

INVx1_ASAP7_75t_L g7146 ( 
.A(n_6742),
.Y(n_7146)
);

AOI22xp33_ASAP7_75t_L g7147 ( 
.A1(n_7072),
.A2(n_47),
.B1(n_45),
.B2(n_46),
.Y(n_7147)
);

NOR2xp33_ASAP7_75t_L g7148 ( 
.A(n_7012),
.B(n_1150),
.Y(n_7148)
);

OAI21xp5_ASAP7_75t_L g7149 ( 
.A1(n_6737),
.A2(n_46),
.B(n_47),
.Y(n_7149)
);

NOR2xp33_ASAP7_75t_L g7150 ( 
.A(n_7024),
.B(n_7102),
.Y(n_7150)
);

NAND2xp5_ASAP7_75t_L g7151 ( 
.A(n_6773),
.B(n_47),
.Y(n_7151)
);

A2O1A1Ixp33_ASAP7_75t_L g7152 ( 
.A1(n_6702),
.A2(n_50),
.B(n_48),
.C(n_49),
.Y(n_7152)
);

NOR2xp67_ASAP7_75t_SL g7153 ( 
.A(n_6934),
.B(n_48),
.Y(n_7153)
);

AOI22xp33_ASAP7_75t_L g7154 ( 
.A1(n_6987),
.A2(n_50),
.B1(n_48),
.B2(n_49),
.Y(n_7154)
);

AOI22xp5_ASAP7_75t_L g7155 ( 
.A1(n_6993),
.A2(n_51),
.B1(n_49),
.B2(n_50),
.Y(n_7155)
);

NOR2xp33_ASAP7_75t_L g7156 ( 
.A(n_7067),
.B(n_1150),
.Y(n_7156)
);

OR2x6_ASAP7_75t_L g7157 ( 
.A(n_6672),
.B(n_1151),
.Y(n_7157)
);

NAND2xp5_ASAP7_75t_L g7158 ( 
.A(n_6777),
.B(n_52),
.Y(n_7158)
);

NAND2xp5_ASAP7_75t_L g7159 ( 
.A(n_6779),
.B(n_52),
.Y(n_7159)
);

AOI21xp5_ASAP7_75t_L g7160 ( 
.A1(n_7060),
.A2(n_1152),
.B(n_1151),
.Y(n_7160)
);

AO21x2_ASAP7_75t_L g7161 ( 
.A1(n_6916),
.A2(n_53),
.B(n_54),
.Y(n_7161)
);

INVx1_ASAP7_75t_L g7162 ( 
.A(n_6748),
.Y(n_7162)
);

AND2x4_ASAP7_75t_L g7163 ( 
.A(n_6768),
.B(n_1155),
.Y(n_7163)
);

AND2x2_ASAP7_75t_L g7164 ( 
.A(n_6838),
.B(n_53),
.Y(n_7164)
);

AOI21x1_ASAP7_75t_L g7165 ( 
.A1(n_6943),
.A2(n_53),
.B(n_54),
.Y(n_7165)
);

NAND2xp5_ASAP7_75t_SL g7166 ( 
.A(n_7050),
.B(n_1155),
.Y(n_7166)
);

NAND2xp5_ASAP7_75t_L g7167 ( 
.A(n_6783),
.B(n_54),
.Y(n_7167)
);

AOI21xp5_ASAP7_75t_L g7168 ( 
.A1(n_7087),
.A2(n_1157),
.B(n_1156),
.Y(n_7168)
);

BUFx8_ASAP7_75t_SL g7169 ( 
.A(n_6762),
.Y(n_7169)
);

INVx1_ASAP7_75t_L g7170 ( 
.A(n_6752),
.Y(n_7170)
);

INVx5_ASAP7_75t_L g7171 ( 
.A(n_6732),
.Y(n_7171)
);

INVx1_ASAP7_75t_L g7172 ( 
.A(n_6754),
.Y(n_7172)
);

INVx1_ASAP7_75t_L g7173 ( 
.A(n_6758),
.Y(n_7173)
);

OAI21xp33_ASAP7_75t_L g7174 ( 
.A1(n_6961),
.A2(n_55),
.B(n_56),
.Y(n_7174)
);

OAI22xp5_ASAP7_75t_L g7175 ( 
.A1(n_7093),
.A2(n_57),
.B1(n_55),
.B2(n_56),
.Y(n_7175)
);

BUFx3_ASAP7_75t_L g7176 ( 
.A(n_6693),
.Y(n_7176)
);

OAI21xp33_ASAP7_75t_L g7177 ( 
.A1(n_6845),
.A2(n_57),
.B(n_58),
.Y(n_7177)
);

NAND2xp5_ASAP7_75t_L g7178 ( 
.A(n_6797),
.B(n_58),
.Y(n_7178)
);

INVx4_ASAP7_75t_L g7179 ( 
.A(n_6732),
.Y(n_7179)
);

INVx4_ASAP7_75t_L g7180 ( 
.A(n_6740),
.Y(n_7180)
);

AOI21xp5_ASAP7_75t_L g7181 ( 
.A1(n_6967),
.A2(n_1157),
.B(n_1156),
.Y(n_7181)
);

OAI21x1_ASAP7_75t_SL g7182 ( 
.A1(n_6945),
.A2(n_59),
.B(n_60),
.Y(n_7182)
);

NAND2xp5_ASAP7_75t_L g7183 ( 
.A(n_7069),
.B(n_59),
.Y(n_7183)
);

O2A1O1Ixp33_ASAP7_75t_L g7184 ( 
.A1(n_6803),
.A2(n_62),
.B(n_60),
.C(n_61),
.Y(n_7184)
);

HB1xp67_ASAP7_75t_L g7185 ( 
.A(n_6684),
.Y(n_7185)
);

NAND2xp5_ASAP7_75t_L g7186 ( 
.A(n_7078),
.B(n_60),
.Y(n_7186)
);

OAI22xp5_ASAP7_75t_L g7187 ( 
.A1(n_7093),
.A2(n_63),
.B1(n_61),
.B2(n_62),
.Y(n_7187)
);

AOI21xp5_ASAP7_75t_L g7188 ( 
.A1(n_6973),
.A2(n_1159),
.B(n_1158),
.Y(n_7188)
);

CKINVDCx5p33_ASAP7_75t_R g7189 ( 
.A(n_6661),
.Y(n_7189)
);

AND2x4_ASAP7_75t_L g7190 ( 
.A(n_6671),
.B(n_1159),
.Y(n_7190)
);

NAND2xp5_ASAP7_75t_L g7191 ( 
.A(n_7079),
.B(n_7083),
.Y(n_7191)
);

NAND2xp5_ASAP7_75t_L g7192 ( 
.A(n_7084),
.B(n_62),
.Y(n_7192)
);

AOI21xp5_ASAP7_75t_L g7193 ( 
.A1(n_6980),
.A2(n_1162),
.B(n_1161),
.Y(n_7193)
);

AOI21xp5_ASAP7_75t_L g7194 ( 
.A1(n_6982),
.A2(n_1162),
.B(n_1161),
.Y(n_7194)
);

CKINVDCx5p33_ASAP7_75t_R g7195 ( 
.A(n_6807),
.Y(n_7195)
);

O2A1O1Ixp33_ASAP7_75t_L g7196 ( 
.A1(n_6876),
.A2(n_6867),
.B(n_7099),
.C(n_6731),
.Y(n_7196)
);

INVx1_ASAP7_75t_L g7197 ( 
.A(n_6760),
.Y(n_7197)
);

NAND2xp5_ASAP7_75t_L g7198 ( 
.A(n_7051),
.B(n_63),
.Y(n_7198)
);

INVx1_ASAP7_75t_L g7199 ( 
.A(n_6664),
.Y(n_7199)
);

NAND2xp5_ASAP7_75t_L g7200 ( 
.A(n_7068),
.B(n_63),
.Y(n_7200)
);

NAND2xp5_ASAP7_75t_L g7201 ( 
.A(n_7089),
.B(n_64),
.Y(n_7201)
);

INVx1_ASAP7_75t_L g7202 ( 
.A(n_6675),
.Y(n_7202)
);

NAND2xp5_ASAP7_75t_L g7203 ( 
.A(n_6986),
.B(n_64),
.Y(n_7203)
);

BUFx4f_ASAP7_75t_L g7204 ( 
.A(n_6740),
.Y(n_7204)
);

NAND3xp33_ASAP7_75t_L g7205 ( 
.A(n_6799),
.B(n_64),
.C(n_65),
.Y(n_7205)
);

O2A1O1Ixp33_ASAP7_75t_SL g7206 ( 
.A1(n_6712),
.A2(n_1165),
.B(n_1166),
.C(n_1164),
.Y(n_7206)
);

O2A1O1Ixp33_ASAP7_75t_L g7207 ( 
.A1(n_6895),
.A2(n_67),
.B(n_65),
.C(n_66),
.Y(n_7207)
);

OAI21xp33_ASAP7_75t_L g7208 ( 
.A1(n_6880),
.A2(n_65),
.B(n_66),
.Y(n_7208)
);

O2A1O1Ixp33_ASAP7_75t_L g7209 ( 
.A1(n_7071),
.A2(n_68),
.B(n_66),
.C(n_67),
.Y(n_7209)
);

NAND2xp5_ASAP7_75t_L g7210 ( 
.A(n_6995),
.B(n_67),
.Y(n_7210)
);

NAND2xp5_ASAP7_75t_L g7211 ( 
.A(n_6996),
.B(n_68),
.Y(n_7211)
);

O2A1O1Ixp33_ASAP7_75t_L g7212 ( 
.A1(n_6899),
.A2(n_71),
.B(n_69),
.C(n_70),
.Y(n_7212)
);

AO21x2_ASAP7_75t_L g7213 ( 
.A1(n_6789),
.A2(n_69),
.B(n_71),
.Y(n_7213)
);

BUFx2_ASAP7_75t_L g7214 ( 
.A(n_6735),
.Y(n_7214)
);

NOR2xp33_ASAP7_75t_L g7215 ( 
.A(n_7005),
.B(n_1164),
.Y(n_7215)
);

OAI21xp5_ASAP7_75t_L g7216 ( 
.A1(n_7006),
.A2(n_71),
.B(n_72),
.Y(n_7216)
);

NAND2xp5_ASAP7_75t_SL g7217 ( 
.A(n_7050),
.B(n_1165),
.Y(n_7217)
);

BUFx4f_ASAP7_75t_L g7218 ( 
.A(n_6701),
.Y(n_7218)
);

NOR2xp33_ASAP7_75t_L g7219 ( 
.A(n_7007),
.B(n_1166),
.Y(n_7219)
);

OAI22xp5_ASAP7_75t_L g7220 ( 
.A1(n_7070),
.A2(n_74),
.B1(n_72),
.B2(n_73),
.Y(n_7220)
);

AND2x4_ASAP7_75t_L g7221 ( 
.A(n_6671),
.B(n_1168),
.Y(n_7221)
);

NAND2xp5_ASAP7_75t_L g7222 ( 
.A(n_7021),
.B(n_72),
.Y(n_7222)
);

A2O1A1Ixp33_ASAP7_75t_SL g7223 ( 
.A1(n_7101),
.A2(n_6992),
.B(n_6950),
.C(n_7045),
.Y(n_7223)
);

O2A1O1Ixp33_ASAP7_75t_L g7224 ( 
.A1(n_7056),
.A2(n_75),
.B(n_73),
.C(n_74),
.Y(n_7224)
);

INVx2_ASAP7_75t_L g7225 ( 
.A(n_6775),
.Y(n_7225)
);

NOR2xp33_ASAP7_75t_L g7226 ( 
.A(n_7032),
.B(n_1168),
.Y(n_7226)
);

AOI21xp5_ASAP7_75t_L g7227 ( 
.A1(n_7033),
.A2(n_1170),
.B(n_1169),
.Y(n_7227)
);

BUFx2_ASAP7_75t_L g7228 ( 
.A(n_6738),
.Y(n_7228)
);

NAND2xp5_ASAP7_75t_L g7229 ( 
.A(n_7035),
.B(n_73),
.Y(n_7229)
);

NAND2xp5_ASAP7_75t_L g7230 ( 
.A(n_7041),
.B(n_74),
.Y(n_7230)
);

INVx5_ASAP7_75t_L g7231 ( 
.A(n_6701),
.Y(n_7231)
);

CKINVDCx20_ASAP7_75t_R g7232 ( 
.A(n_6765),
.Y(n_7232)
);

BUFx12f_ASAP7_75t_L g7233 ( 
.A(n_6778),
.Y(n_7233)
);

INVx1_ASAP7_75t_L g7234 ( 
.A(n_6677),
.Y(n_7234)
);

A2O1A1Ixp33_ASAP7_75t_L g7235 ( 
.A1(n_6927),
.A2(n_77),
.B(n_75),
.C(n_76),
.Y(n_7235)
);

AND2x2_ASAP7_75t_L g7236 ( 
.A(n_7066),
.B(n_75),
.Y(n_7236)
);

AOI21xp5_ASAP7_75t_L g7237 ( 
.A1(n_7044),
.A2(n_1170),
.B(n_1169),
.Y(n_7237)
);

NAND2xp5_ASAP7_75t_L g7238 ( 
.A(n_7046),
.B(n_76),
.Y(n_7238)
);

NOR2xp33_ASAP7_75t_R g7239 ( 
.A(n_6929),
.B(n_1171),
.Y(n_7239)
);

BUFx8_ASAP7_75t_L g7240 ( 
.A(n_6782),
.Y(n_7240)
);

NAND2xp5_ASAP7_75t_L g7241 ( 
.A(n_6964),
.B(n_77),
.Y(n_7241)
);

OAI22xp5_ASAP7_75t_L g7242 ( 
.A1(n_6913),
.A2(n_80),
.B1(n_78),
.B2(n_79),
.Y(n_7242)
);

NOR2xp33_ASAP7_75t_L g7243 ( 
.A(n_6818),
.B(n_1171),
.Y(n_7243)
);

INVx4_ASAP7_75t_L g7244 ( 
.A(n_6662),
.Y(n_7244)
);

NAND2xp5_ASAP7_75t_L g7245 ( 
.A(n_6965),
.B(n_78),
.Y(n_7245)
);

NAND2xp5_ASAP7_75t_SL g7246 ( 
.A(n_7057),
.B(n_1172),
.Y(n_7246)
);

AOI21x1_ASAP7_75t_L g7247 ( 
.A1(n_7098),
.A2(n_79),
.B(n_80),
.Y(n_7247)
);

CKINVDCx5p33_ASAP7_75t_R g7248 ( 
.A(n_6825),
.Y(n_7248)
);

AOI21xp5_ASAP7_75t_L g7249 ( 
.A1(n_6928),
.A2(n_1173),
.B(n_1172),
.Y(n_7249)
);

AND2x2_ASAP7_75t_L g7250 ( 
.A(n_7066),
.B(n_79),
.Y(n_7250)
);

CKINVDCx5p33_ASAP7_75t_R g7251 ( 
.A(n_6757),
.Y(n_7251)
);

AOI21xp5_ASAP7_75t_L g7252 ( 
.A1(n_6930),
.A2(n_1175),
.B(n_1174),
.Y(n_7252)
);

INVx1_ASAP7_75t_L g7253 ( 
.A(n_6678),
.Y(n_7253)
);

AOI22xp33_ASAP7_75t_L g7254 ( 
.A1(n_7080),
.A2(n_82),
.B1(n_80),
.B2(n_81),
.Y(n_7254)
);

AOI22xp33_ASAP7_75t_L g7255 ( 
.A1(n_6756),
.A2(n_83),
.B1(n_81),
.B2(n_82),
.Y(n_7255)
);

NOR2xp67_ASAP7_75t_SL g7256 ( 
.A(n_6846),
.B(n_81),
.Y(n_7256)
);

A2O1A1Ixp33_ASAP7_75t_SL g7257 ( 
.A1(n_6975),
.A2(n_85),
.B(n_82),
.C(n_84),
.Y(n_7257)
);

AOI21xp5_ASAP7_75t_L g7258 ( 
.A1(n_6949),
.A2(n_1176),
.B(n_1175),
.Y(n_7258)
);

NOR2xp33_ASAP7_75t_L g7259 ( 
.A(n_7003),
.B(n_1178),
.Y(n_7259)
);

INVx2_ASAP7_75t_L g7260 ( 
.A(n_6787),
.Y(n_7260)
);

INVx1_ASAP7_75t_L g7261 ( 
.A(n_6681),
.Y(n_7261)
);

INVx1_ASAP7_75t_L g7262 ( 
.A(n_6685),
.Y(n_7262)
);

OAI22xp5_ASAP7_75t_L g7263 ( 
.A1(n_6819),
.A2(n_87),
.B1(n_85),
.B2(n_86),
.Y(n_7263)
);

INVx1_ASAP7_75t_L g7264 ( 
.A(n_6690),
.Y(n_7264)
);

AND2x2_ASAP7_75t_L g7265 ( 
.A(n_6998),
.B(n_85),
.Y(n_7265)
);

INVxp67_ASAP7_75t_SL g7266 ( 
.A(n_6767),
.Y(n_7266)
);

NOR2xp33_ASAP7_75t_L g7267 ( 
.A(n_6978),
.B(n_1180),
.Y(n_7267)
);

NAND2xp5_ASAP7_75t_L g7268 ( 
.A(n_6990),
.B(n_86),
.Y(n_7268)
);

AOI22xp33_ASAP7_75t_SL g7269 ( 
.A1(n_6756),
.A2(n_1181),
.B1(n_1182),
.B2(n_1180),
.Y(n_7269)
);

NAND2xp5_ASAP7_75t_L g7270 ( 
.A(n_6999),
.B(n_86),
.Y(n_7270)
);

AOI21x1_ASAP7_75t_L g7271 ( 
.A1(n_6984),
.A2(n_87),
.B(n_88),
.Y(n_7271)
);

INVx1_ASAP7_75t_L g7272 ( 
.A(n_6691),
.Y(n_7272)
);

OR2x6_ASAP7_75t_L g7273 ( 
.A(n_6788),
.B(n_1181),
.Y(n_7273)
);

OAI22xp5_ASAP7_75t_L g7274 ( 
.A1(n_6926),
.A2(n_90),
.B1(n_88),
.B2(n_89),
.Y(n_7274)
);

OAI21x1_ASAP7_75t_L g7275 ( 
.A1(n_6914),
.A2(n_88),
.B(n_89),
.Y(n_7275)
);

OR2x2_ASAP7_75t_L g7276 ( 
.A(n_6849),
.B(n_1182),
.Y(n_7276)
);

NAND2xp5_ASAP7_75t_SL g7277 ( 
.A(n_7057),
.B(n_1183),
.Y(n_7277)
);

INVx1_ASAP7_75t_L g7278 ( 
.A(n_6696),
.Y(n_7278)
);

NAND2xp5_ASAP7_75t_SL g7279 ( 
.A(n_7049),
.B(n_1183),
.Y(n_7279)
);

INVx2_ASAP7_75t_L g7280 ( 
.A(n_6790),
.Y(n_7280)
);

NOR2xp33_ASAP7_75t_L g7281 ( 
.A(n_7019),
.B(n_1184),
.Y(n_7281)
);

BUFx12f_ASAP7_75t_L g7282 ( 
.A(n_6788),
.Y(n_7282)
);

AOI21xp5_ASAP7_75t_L g7283 ( 
.A1(n_6955),
.A2(n_1186),
.B(n_1184),
.Y(n_7283)
);

AOI21xp5_ASAP7_75t_L g7284 ( 
.A1(n_6956),
.A2(n_1188),
.B(n_1187),
.Y(n_7284)
);

NAND2xp5_ASAP7_75t_L g7285 ( 
.A(n_7042),
.B(n_89),
.Y(n_7285)
);

NOR2xp67_ASAP7_75t_SL g7286 ( 
.A(n_6806),
.B(n_90),
.Y(n_7286)
);

O2A1O1Ixp5_ASAP7_75t_L g7287 ( 
.A1(n_7061),
.A2(n_92),
.B(n_90),
.C(n_91),
.Y(n_7287)
);

INVx2_ASAP7_75t_L g7288 ( 
.A(n_6800),
.Y(n_7288)
);

INVx1_ASAP7_75t_SL g7289 ( 
.A(n_6694),
.Y(n_7289)
);

INVx2_ASAP7_75t_L g7290 ( 
.A(n_6808),
.Y(n_7290)
);

OAI22xp5_ASAP7_75t_L g7291 ( 
.A1(n_6958),
.A2(n_93),
.B1(n_91),
.B2(n_92),
.Y(n_7291)
);

NAND2xp5_ASAP7_75t_L g7292 ( 
.A(n_7043),
.B(n_92),
.Y(n_7292)
);

O2A1O1Ixp33_ASAP7_75t_L g7293 ( 
.A1(n_7091),
.A2(n_95),
.B(n_93),
.C(n_94),
.Y(n_7293)
);

AOI21xp5_ASAP7_75t_L g7294 ( 
.A1(n_6957),
.A2(n_1188),
.B(n_1187),
.Y(n_7294)
);

INVx2_ASAP7_75t_L g7295 ( 
.A(n_6827),
.Y(n_7295)
);

NAND2xp5_ASAP7_75t_L g7296 ( 
.A(n_6959),
.B(n_93),
.Y(n_7296)
);

NAND2xp5_ASAP7_75t_L g7297 ( 
.A(n_6963),
.B(n_94),
.Y(n_7297)
);

NOR3xp33_ASAP7_75t_L g7298 ( 
.A(n_6904),
.B(n_94),
.C(n_95),
.Y(n_7298)
);

NAND2xp5_ASAP7_75t_L g7299 ( 
.A(n_6939),
.B(n_95),
.Y(n_7299)
);

O2A1O1Ixp33_ASAP7_75t_L g7300 ( 
.A1(n_7038),
.A2(n_98),
.B(n_96),
.C(n_97),
.Y(n_7300)
);

OR2x6_ASAP7_75t_SL g7301 ( 
.A(n_6985),
.B(n_6932),
.Y(n_7301)
);

BUFx6f_ASAP7_75t_L g7302 ( 
.A(n_6725),
.Y(n_7302)
);

AND2x2_ASAP7_75t_SL g7303 ( 
.A(n_6832),
.B(n_1189),
.Y(n_7303)
);

NAND2xp5_ASAP7_75t_L g7304 ( 
.A(n_6947),
.B(n_6798),
.Y(n_7304)
);

AOI21xp5_ASAP7_75t_L g7305 ( 
.A1(n_7090),
.A2(n_7097),
.B(n_6687),
.Y(n_7305)
);

AND2x2_ASAP7_75t_L g7306 ( 
.A(n_7010),
.B(n_96),
.Y(n_7306)
);

OAI22xp5_ASAP7_75t_SL g7307 ( 
.A1(n_6813),
.A2(n_7063),
.B1(n_7018),
.B2(n_6714),
.Y(n_7307)
);

BUFx3_ASAP7_75t_L g7308 ( 
.A(n_6782),
.Y(n_7308)
);

INVx1_ASAP7_75t_L g7309 ( 
.A(n_6700),
.Y(n_7309)
);

BUFx2_ASAP7_75t_L g7310 ( 
.A(n_6842),
.Y(n_7310)
);

AO32x2_ASAP7_75t_L g7311 ( 
.A1(n_6938),
.A2(n_98),
.A3(n_96),
.B1(n_97),
.B2(n_99),
.Y(n_7311)
);

A2O1A1Ixp33_ASAP7_75t_L g7312 ( 
.A1(n_6750),
.A2(n_101),
.B(n_99),
.C(n_100),
.Y(n_7312)
);

INVx2_ASAP7_75t_L g7313 ( 
.A(n_6836),
.Y(n_7313)
);

INVx2_ASAP7_75t_L g7314 ( 
.A(n_6850),
.Y(n_7314)
);

INVx1_ASAP7_75t_L g7315 ( 
.A(n_6709),
.Y(n_7315)
);

HB1xp67_ASAP7_75t_L g7316 ( 
.A(n_6823),
.Y(n_7316)
);

OAI21x1_ASAP7_75t_L g7317 ( 
.A1(n_6911),
.A2(n_99),
.B(n_100),
.Y(n_7317)
);

AOI21x1_ASAP7_75t_L g7318 ( 
.A1(n_6817),
.A2(n_100),
.B(n_101),
.Y(n_7318)
);

INVx3_ASAP7_75t_L g7319 ( 
.A(n_6743),
.Y(n_7319)
);

AOI21xp5_ASAP7_75t_L g7320 ( 
.A1(n_7022),
.A2(n_1190),
.B(n_1189),
.Y(n_7320)
);

AOI21xp5_ASAP7_75t_L g7321 ( 
.A1(n_6755),
.A2(n_1191),
.B(n_1190),
.Y(n_7321)
);

AOI33xp33_ASAP7_75t_L g7322 ( 
.A1(n_6795),
.A2(n_103),
.A3(n_105),
.B1(n_101),
.B2(n_102),
.B3(n_104),
.Y(n_7322)
);

NAND2xp5_ASAP7_75t_L g7323 ( 
.A(n_7054),
.B(n_102),
.Y(n_7323)
);

OAI21xp5_ASAP7_75t_L g7324 ( 
.A1(n_6877),
.A2(n_102),
.B(n_103),
.Y(n_7324)
);

NAND2xp5_ASAP7_75t_SL g7325 ( 
.A(n_7048),
.B(n_1191),
.Y(n_7325)
);

OAI22xp5_ASAP7_75t_L g7326 ( 
.A1(n_7092),
.A2(n_6704),
.B1(n_6695),
.B2(n_6692),
.Y(n_7326)
);

O2A1O1Ixp33_ASAP7_75t_L g7327 ( 
.A1(n_7028),
.A2(n_6828),
.B(n_6741),
.C(n_6833),
.Y(n_7327)
);

AND2x4_ASAP7_75t_L g7328 ( 
.A(n_6728),
.B(n_1192),
.Y(n_7328)
);

AOI22xp5_ASAP7_75t_L g7329 ( 
.A1(n_6682),
.A2(n_105),
.B1(n_103),
.B2(n_104),
.Y(n_7329)
);

AOI21xp5_ASAP7_75t_L g7330 ( 
.A1(n_6921),
.A2(n_1194),
.B(n_1193),
.Y(n_7330)
);

AOI21xp5_ASAP7_75t_L g7331 ( 
.A1(n_7094),
.A2(n_1194),
.B(n_1193),
.Y(n_7331)
);

AOI21xp5_ASAP7_75t_L g7332 ( 
.A1(n_6858),
.A2(n_1196),
.B(n_1195),
.Y(n_7332)
);

NAND2xp5_ASAP7_75t_SL g7333 ( 
.A(n_7048),
.B(n_6944),
.Y(n_7333)
);

NOR2xp67_ASAP7_75t_L g7334 ( 
.A(n_6715),
.B(n_104),
.Y(n_7334)
);

NAND2xp5_ASAP7_75t_L g7335 ( 
.A(n_7052),
.B(n_105),
.Y(n_7335)
);

O2A1O1Ixp33_ASAP7_75t_L g7336 ( 
.A1(n_6784),
.A2(n_108),
.B(n_106),
.C(n_107),
.Y(n_7336)
);

AOI21xp33_ASAP7_75t_L g7337 ( 
.A1(n_7100),
.A2(n_106),
.B(n_107),
.Y(n_7337)
);

NAND2xp5_ASAP7_75t_SL g7338 ( 
.A(n_6944),
.B(n_1196),
.Y(n_7338)
);

AOI21xp5_ASAP7_75t_L g7339 ( 
.A1(n_6688),
.A2(n_1198),
.B(n_1197),
.Y(n_7339)
);

NAND2xp5_ASAP7_75t_SL g7340 ( 
.A(n_7055),
.B(n_1197),
.Y(n_7340)
);

INVx1_ASAP7_75t_L g7341 ( 
.A(n_6710),
.Y(n_7341)
);

AOI22xp33_ASAP7_75t_L g7342 ( 
.A1(n_6756),
.A2(n_108),
.B1(n_106),
.B2(n_107),
.Y(n_7342)
);

INVx1_ASAP7_75t_L g7343 ( 
.A(n_6711),
.Y(n_7343)
);

OAI22xp5_ASAP7_75t_L g7344 ( 
.A1(n_7034),
.A2(n_111),
.B1(n_109),
.B2(n_110),
.Y(n_7344)
);

NOR2xp33_ASAP7_75t_L g7345 ( 
.A(n_6970),
.B(n_1198),
.Y(n_7345)
);

BUFx2_ASAP7_75t_L g7346 ( 
.A(n_6854),
.Y(n_7346)
);

OAI22xp5_ASAP7_75t_SL g7347 ( 
.A1(n_6772),
.A2(n_111),
.B1(n_109),
.B2(n_110),
.Y(n_7347)
);

BUFx6f_ASAP7_75t_L g7348 ( 
.A(n_6725),
.Y(n_7348)
);

INVx1_ASAP7_75t_L g7349 ( 
.A(n_6719),
.Y(n_7349)
);

A2O1A1Ixp33_ASAP7_75t_L g7350 ( 
.A1(n_6900),
.A2(n_112),
.B(n_109),
.C(n_110),
.Y(n_7350)
);

NAND2xp5_ASAP7_75t_SL g7351 ( 
.A(n_7062),
.B(n_1199),
.Y(n_7351)
);

NAND2xp33_ASAP7_75t_SL g7352 ( 
.A(n_6815),
.B(n_1200),
.Y(n_7352)
);

AOI21xp5_ASAP7_75t_L g7353 ( 
.A1(n_6699),
.A2(n_1203),
.B(n_1201),
.Y(n_7353)
);

OAI22xp33_ASAP7_75t_L g7354 ( 
.A1(n_6730),
.A2(n_115),
.B1(n_113),
.B2(n_114),
.Y(n_7354)
);

INVxp67_ASAP7_75t_L g7355 ( 
.A(n_6766),
.Y(n_7355)
);

NOR2xp33_ASAP7_75t_L g7356 ( 
.A(n_6816),
.B(n_1204),
.Y(n_7356)
);

OAI22xp5_ASAP7_75t_L g7357 ( 
.A1(n_7053),
.A2(n_116),
.B1(n_113),
.B2(n_114),
.Y(n_7357)
);

INVx2_ASAP7_75t_L g7358 ( 
.A(n_6878),
.Y(n_7358)
);

O2A1O1Ixp33_ASAP7_75t_L g7359 ( 
.A1(n_6946),
.A2(n_116),
.B(n_113),
.C(n_114),
.Y(n_7359)
);

BUFx3_ASAP7_75t_L g7360 ( 
.A(n_6686),
.Y(n_7360)
);

INVx1_ASAP7_75t_L g7361 ( 
.A(n_6720),
.Y(n_7361)
);

NAND2xp5_ASAP7_75t_SL g7362 ( 
.A(n_7014),
.B(n_1205),
.Y(n_7362)
);

OAI21xp5_ASAP7_75t_L g7363 ( 
.A1(n_6903),
.A2(n_117),
.B(n_118),
.Y(n_7363)
);

CKINVDCx14_ASAP7_75t_R g7364 ( 
.A(n_6843),
.Y(n_7364)
);

NAND2xp5_ASAP7_75t_SL g7365 ( 
.A(n_7027),
.B(n_1205),
.Y(n_7365)
);

INVx2_ASAP7_75t_L g7366 ( 
.A(n_6879),
.Y(n_7366)
);

AOI21xp5_ASAP7_75t_L g7367 ( 
.A1(n_6989),
.A2(n_1207),
.B(n_1206),
.Y(n_7367)
);

AOI21xp5_ASAP7_75t_L g7368 ( 
.A1(n_6909),
.A2(n_1207),
.B(n_1206),
.Y(n_7368)
);

OAI22xp5_ASAP7_75t_L g7369 ( 
.A1(n_7059),
.A2(n_120),
.B1(n_118),
.B2(n_119),
.Y(n_7369)
);

OR2x6_ASAP7_75t_L g7370 ( 
.A(n_6962),
.B(n_6919),
.Y(n_7370)
);

BUFx6f_ASAP7_75t_L g7371 ( 
.A(n_6686),
.Y(n_7371)
);

NOR3xp33_ASAP7_75t_L g7372 ( 
.A(n_6831),
.B(n_119),
.C(n_120),
.Y(n_7372)
);

BUFx3_ASAP7_75t_L g7373 ( 
.A(n_6698),
.Y(n_7373)
);

NAND2xp5_ASAP7_75t_SL g7374 ( 
.A(n_7039),
.B(n_1208),
.Y(n_7374)
);

NAND2xp5_ASAP7_75t_L g7375 ( 
.A(n_7095),
.B(n_119),
.Y(n_7375)
);

O2A1O1Ixp33_ASAP7_75t_L g7376 ( 
.A1(n_6953),
.A2(n_6988),
.B(n_7011),
.C(n_6968),
.Y(n_7376)
);

NAND2xp5_ASAP7_75t_L g7377 ( 
.A(n_7013),
.B(n_120),
.Y(n_7377)
);

AND2x2_ASAP7_75t_L g7378 ( 
.A(n_6935),
.B(n_121),
.Y(n_7378)
);

HB1xp67_ASAP7_75t_L g7379 ( 
.A(n_6872),
.Y(n_7379)
);

HB1xp67_ASAP7_75t_L g7380 ( 
.A(n_6786),
.Y(n_7380)
);

NOR2xp33_ASAP7_75t_L g7381 ( 
.A(n_6706),
.B(n_1208),
.Y(n_7381)
);

NOR2xp33_ASAP7_75t_L g7382 ( 
.A(n_7096),
.B(n_1209),
.Y(n_7382)
);

AOI21xp5_ASAP7_75t_L g7383 ( 
.A1(n_7036),
.A2(n_1210),
.B(n_1209),
.Y(n_7383)
);

NOR2xp33_ASAP7_75t_L g7384 ( 
.A(n_6667),
.B(n_1211),
.Y(n_7384)
);

CKINVDCx5p33_ASAP7_75t_R g7385 ( 
.A(n_6972),
.Y(n_7385)
);

INVx2_ASAP7_75t_L g7386 ( 
.A(n_6890),
.Y(n_7386)
);

NOR2xp33_ASAP7_75t_L g7387 ( 
.A(n_6983),
.B(n_1211),
.Y(n_7387)
);

NOR3xp33_ASAP7_75t_L g7388 ( 
.A(n_6922),
.B(n_121),
.C(n_122),
.Y(n_7388)
);

HB1xp67_ASAP7_75t_L g7389 ( 
.A(n_6887),
.Y(n_7389)
);

BUFx6f_ASAP7_75t_L g7390 ( 
.A(n_6815),
.Y(n_7390)
);

OAI21x1_ASAP7_75t_L g7391 ( 
.A1(n_6809),
.A2(n_122),
.B(n_123),
.Y(n_7391)
);

NAND2xp5_ASAP7_75t_SL g7392 ( 
.A(n_6979),
.B(n_1212),
.Y(n_7392)
);

O2A1O1Ixp33_ASAP7_75t_L g7393 ( 
.A1(n_7037),
.A2(n_125),
.B(n_123),
.C(n_124),
.Y(n_7393)
);

CKINVDCx5p33_ASAP7_75t_R g7394 ( 
.A(n_7017),
.Y(n_7394)
);

A2O1A1Ixp33_ASAP7_75t_L g7395 ( 
.A1(n_7075),
.A2(n_125),
.B(n_123),
.C(n_124),
.Y(n_7395)
);

INVx2_ASAP7_75t_L g7396 ( 
.A(n_6892),
.Y(n_7396)
);

INVx1_ASAP7_75t_L g7397 ( 
.A(n_6721),
.Y(n_7397)
);

O2A1O1Ixp33_ASAP7_75t_L g7398 ( 
.A1(n_7077),
.A2(n_127),
.B(n_125),
.C(n_126),
.Y(n_7398)
);

NOR2xp33_ASAP7_75t_L g7399 ( 
.A(n_6851),
.B(n_1212),
.Y(n_7399)
);

INVx1_ASAP7_75t_L g7400 ( 
.A(n_6729),
.Y(n_7400)
);

AND3x1_ASAP7_75t_SL g7401 ( 
.A(n_7064),
.B(n_126),
.C(n_127),
.Y(n_7401)
);

AOI22x1_ASAP7_75t_L g7402 ( 
.A1(n_6885),
.A2(n_6852),
.B1(n_7000),
.B2(n_6991),
.Y(n_7402)
);

O2A1O1Ixp33_ASAP7_75t_L g7403 ( 
.A1(n_7081),
.A2(n_7086),
.B(n_7082),
.C(n_6893),
.Y(n_7403)
);

A2O1A1Ixp33_ASAP7_75t_L g7404 ( 
.A1(n_6940),
.A2(n_128),
.B(n_126),
.C(n_127),
.Y(n_7404)
);

INVx1_ASAP7_75t_L g7405 ( 
.A(n_6734),
.Y(n_7405)
);

AOI21xp5_ASAP7_75t_L g7406 ( 
.A1(n_6991),
.A2(n_1214),
.B(n_1213),
.Y(n_7406)
);

AOI21xp5_ASAP7_75t_L g7407 ( 
.A1(n_7000),
.A2(n_1215),
.B(n_1214),
.Y(n_7407)
);

AOI21xp5_ASAP7_75t_L g7408 ( 
.A1(n_6739),
.A2(n_1216),
.B(n_1215),
.Y(n_7408)
);

INVx2_ASAP7_75t_L g7409 ( 
.A(n_6751),
.Y(n_7409)
);

BUFx6f_ASAP7_75t_L g7410 ( 
.A(n_6859),
.Y(n_7410)
);

OAI22xp5_ASAP7_75t_L g7411 ( 
.A1(n_6707),
.A2(n_130),
.B1(n_128),
.B2(n_129),
.Y(n_7411)
);

AOI21x1_ASAP7_75t_L g7412 ( 
.A1(n_6812),
.A2(n_129),
.B(n_130),
.Y(n_7412)
);

BUFx6f_ASAP7_75t_L g7413 ( 
.A(n_6859),
.Y(n_7413)
);

BUFx3_ASAP7_75t_L g7414 ( 
.A(n_6746),
.Y(n_7414)
);

AOI21xp5_ASAP7_75t_L g7415 ( 
.A1(n_6780),
.A2(n_1217),
.B(n_1216),
.Y(n_7415)
);

AOI21xp5_ASAP7_75t_L g7416 ( 
.A1(n_6781),
.A2(n_1218),
.B(n_1217),
.Y(n_7416)
);

NOR2x1_ASAP7_75t_L g7417 ( 
.A(n_6810),
.B(n_1218),
.Y(n_7417)
);

AND2x2_ASAP7_75t_L g7418 ( 
.A(n_6937),
.B(n_129),
.Y(n_7418)
);

OAI21xp33_ASAP7_75t_L g7419 ( 
.A1(n_6847),
.A2(n_130),
.B(n_131),
.Y(n_7419)
);

BUFx4f_ASAP7_75t_L g7420 ( 
.A(n_6931),
.Y(n_7420)
);

NOR3xp33_ASAP7_75t_SL g7421 ( 
.A(n_6948),
.B(n_131),
.C(n_132),
.Y(n_7421)
);

INVx1_ASAP7_75t_L g7422 ( 
.A(n_6826),
.Y(n_7422)
);

AOI21xp5_ASAP7_75t_L g7423 ( 
.A1(n_6733),
.A2(n_1221),
.B(n_1220),
.Y(n_7423)
);

AOI21xp5_ASAP7_75t_L g7424 ( 
.A1(n_7015),
.A2(n_1221),
.B(n_1220),
.Y(n_7424)
);

AOI21xp5_ASAP7_75t_L g7425 ( 
.A1(n_6835),
.A2(n_1223),
.B(n_1222),
.Y(n_7425)
);

OAI21xp5_ASAP7_75t_L g7426 ( 
.A1(n_6726),
.A2(n_132),
.B(n_133),
.Y(n_7426)
);

NAND2xp5_ASAP7_75t_SL g7427 ( 
.A(n_6915),
.B(n_1223),
.Y(n_7427)
);

HB1xp67_ASAP7_75t_L g7428 ( 
.A(n_6954),
.Y(n_7428)
);

AOI21xp5_ASAP7_75t_L g7429 ( 
.A1(n_6837),
.A2(n_1225),
.B(n_1224),
.Y(n_7429)
);

INVxp33_ASAP7_75t_SL g7430 ( 
.A(n_6674),
.Y(n_7430)
);

OR2x2_ASAP7_75t_L g7431 ( 
.A(n_6941),
.B(n_1226),
.Y(n_7431)
);

INVx1_ASAP7_75t_L g7432 ( 
.A(n_6853),
.Y(n_7432)
);

OAI22xp5_ASAP7_75t_L g7433 ( 
.A1(n_6907),
.A2(n_134),
.B1(n_132),
.B2(n_133),
.Y(n_7433)
);

NAND2xp5_ASAP7_75t_SL g7434 ( 
.A(n_6915),
.B(n_1227),
.Y(n_7434)
);

AOI21xp5_ASAP7_75t_L g7435 ( 
.A1(n_6860),
.A2(n_1228),
.B(n_1227),
.Y(n_7435)
);

NAND2x1p5_ASAP7_75t_L g7436 ( 
.A(n_6820),
.B(n_1228),
.Y(n_7436)
);

BUFx6f_ASAP7_75t_L g7437 ( 
.A(n_6791),
.Y(n_7437)
);

AOI21xp5_ASAP7_75t_L g7438 ( 
.A1(n_6861),
.A2(n_1230),
.B(n_1229),
.Y(n_7438)
);

AOI21xp5_ASAP7_75t_L g7439 ( 
.A1(n_6866),
.A2(n_1231),
.B(n_1230),
.Y(n_7439)
);

NAND2xp5_ASAP7_75t_L g7440 ( 
.A(n_6682),
.B(n_133),
.Y(n_7440)
);

CKINVDCx14_ASAP7_75t_R g7441 ( 
.A(n_6745),
.Y(n_7441)
);

NAND2xp5_ASAP7_75t_L g7442 ( 
.A(n_6682),
.B(n_134),
.Y(n_7442)
);

INVx1_ASAP7_75t_L g7443 ( 
.A(n_6871),
.Y(n_7443)
);

NAND2xp5_ASAP7_75t_L g7444 ( 
.A(n_7009),
.B(n_135),
.Y(n_7444)
);

INVx1_ASAP7_75t_L g7445 ( 
.A(n_6874),
.Y(n_7445)
);

INVx1_ASAP7_75t_L g7446 ( 
.A(n_6881),
.Y(n_7446)
);

OAI21xp5_ASAP7_75t_L g7447 ( 
.A1(n_6894),
.A2(n_135),
.B(n_136),
.Y(n_7447)
);

NOR2xp33_ASAP7_75t_R g7448 ( 
.A(n_6908),
.B(n_1231),
.Y(n_7448)
);

NAND2xp5_ASAP7_75t_L g7449 ( 
.A(n_7020),
.B(n_7088),
.Y(n_7449)
);

AND2x4_ASAP7_75t_L g7450 ( 
.A(n_6822),
.B(n_1232),
.Y(n_7450)
);

NAND2x1p5_ASAP7_75t_L g7451 ( 
.A(n_6821),
.B(n_1233),
.Y(n_7451)
);

AOI21xp5_ASAP7_75t_L g7452 ( 
.A1(n_6886),
.A2(n_1234),
.B(n_1233),
.Y(n_7452)
);

NAND2xp5_ASAP7_75t_SL g7453 ( 
.A(n_6902),
.B(n_1234),
.Y(n_7453)
);

AND2x4_ASAP7_75t_L g7454 ( 
.A(n_6873),
.B(n_1235),
.Y(n_7454)
);

OAI22x1_ASAP7_75t_L g7455 ( 
.A1(n_6801),
.A2(n_137),
.B1(n_135),
.B2(n_136),
.Y(n_7455)
);

BUFx6f_ASAP7_75t_L g7456 ( 
.A(n_6791),
.Y(n_7456)
);

INVx1_ASAP7_75t_L g7457 ( 
.A(n_6888),
.Y(n_7457)
);

INVx2_ASAP7_75t_L g7458 ( 
.A(n_6898),
.Y(n_7458)
);

NAND2xp5_ASAP7_75t_SL g7459 ( 
.A(n_6902),
.B(n_1236),
.Y(n_7459)
);

OAI22xp5_ASAP7_75t_L g7460 ( 
.A1(n_6917),
.A2(n_139),
.B1(n_136),
.B2(n_138),
.Y(n_7460)
);

INVx1_ASAP7_75t_L g7461 ( 
.A(n_6905),
.Y(n_7461)
);

AOI33xp33_ASAP7_75t_L g7462 ( 
.A1(n_6875),
.A2(n_140),
.A3(n_142),
.B1(n_138),
.B2(n_139),
.B3(n_141),
.Y(n_7462)
);

OAI22xp5_ASAP7_75t_L g7463 ( 
.A1(n_6917),
.A2(n_141),
.B1(n_139),
.B2(n_140),
.Y(n_7463)
);

AOI21xp33_ASAP7_75t_L g7464 ( 
.A1(n_6882),
.A2(n_142),
.B(n_143),
.Y(n_7464)
);

AOI21xp5_ASAP7_75t_L g7465 ( 
.A1(n_6974),
.A2(n_1237),
.B(n_1236),
.Y(n_7465)
);

BUFx6f_ASAP7_75t_L g7466 ( 
.A(n_6805),
.Y(n_7466)
);

O2A1O1Ixp33_ASAP7_75t_L g7467 ( 
.A1(n_6936),
.A2(n_144),
.B(n_142),
.C(n_143),
.Y(n_7467)
);

A2O1A1Ixp33_ASAP7_75t_L g7468 ( 
.A1(n_7058),
.A2(n_146),
.B(n_144),
.C(n_145),
.Y(n_7468)
);

NAND2xp5_ASAP7_75t_SL g7469 ( 
.A(n_6969),
.B(n_1237),
.Y(n_7469)
);

BUFx6f_ASAP7_75t_L g7470 ( 
.A(n_6662),
.Y(n_7470)
);

NAND2xp5_ASAP7_75t_L g7471 ( 
.A(n_6906),
.B(n_145),
.Y(n_7471)
);

AOI21xp5_ASAP7_75t_L g7472 ( 
.A1(n_7026),
.A2(n_1240),
.B(n_1239),
.Y(n_7472)
);

INVxp67_ASAP7_75t_L g7473 ( 
.A(n_6811),
.Y(n_7473)
);

O2A1O1Ixp5_ASAP7_75t_L g7474 ( 
.A1(n_7076),
.A2(n_148),
.B(n_146),
.C(n_147),
.Y(n_7474)
);

NAND2xp5_ASAP7_75t_L g7475 ( 
.A(n_7030),
.B(n_147),
.Y(n_7475)
);

INVx1_ASAP7_75t_L g7476 ( 
.A(n_6912),
.Y(n_7476)
);

INVx1_ASAP7_75t_L g7477 ( 
.A(n_6918),
.Y(n_7477)
);

NAND2xp5_ASAP7_75t_L g7478 ( 
.A(n_6981),
.B(n_147),
.Y(n_7478)
);

HB1xp67_ASAP7_75t_L g7479 ( 
.A(n_6844),
.Y(n_7479)
);

NAND2xp5_ASAP7_75t_L g7480 ( 
.A(n_7065),
.B(n_148),
.Y(n_7480)
);

INVx2_ASAP7_75t_L g7481 ( 
.A(n_6925),
.Y(n_7481)
);

NOR3xp33_ASAP7_75t_SL g7482 ( 
.A(n_6774),
.B(n_149),
.C(n_150),
.Y(n_7482)
);

OAI21xp5_ASAP7_75t_L g7483 ( 
.A1(n_6891),
.A2(n_149),
.B(n_150),
.Y(n_7483)
);

NOR2xp33_ASAP7_75t_R g7484 ( 
.A(n_6668),
.B(n_1240),
.Y(n_7484)
);

OAI21xp33_ASAP7_75t_L g7485 ( 
.A1(n_6759),
.A2(n_149),
.B(n_150),
.Y(n_7485)
);

NAND2xp5_ASAP7_75t_L g7486 ( 
.A(n_6976),
.B(n_151),
.Y(n_7486)
);

AOI21xp5_ASAP7_75t_L g7487 ( 
.A1(n_7026),
.A2(n_1242),
.B(n_1241),
.Y(n_7487)
);

AND2x4_ASAP7_75t_L g7488 ( 
.A(n_6856),
.B(n_1241),
.Y(n_7488)
);

AOI22xp5_ASAP7_75t_L g7489 ( 
.A1(n_6942),
.A2(n_6951),
.B1(n_6920),
.B2(n_7029),
.Y(n_7489)
);

INVx2_ASAP7_75t_L g7490 ( 
.A(n_6897),
.Y(n_7490)
);

BUFx6f_ASAP7_75t_L g7491 ( 
.A(n_6804),
.Y(n_7491)
);

INVx3_ASAP7_75t_L g7492 ( 
.A(n_6718),
.Y(n_7492)
);

AOI21xp5_ASAP7_75t_L g7493 ( 
.A1(n_7026),
.A2(n_1243),
.B(n_1242),
.Y(n_7493)
);

AOI21xp5_ASAP7_75t_L g7494 ( 
.A1(n_6830),
.A2(n_1244),
.B(n_1243),
.Y(n_7494)
);

A2O1A1Ixp33_ASAP7_75t_L g7495 ( 
.A1(n_6960),
.A2(n_153),
.B(n_151),
.C(n_152),
.Y(n_7495)
);

AOI21xp5_ASAP7_75t_L g7496 ( 
.A1(n_6889),
.A2(n_1246),
.B(n_1245),
.Y(n_7496)
);

NAND2xp5_ASAP7_75t_L g7497 ( 
.A(n_7001),
.B(n_152),
.Y(n_7497)
);

A2O1A1Ixp33_ASAP7_75t_L g7498 ( 
.A1(n_6722),
.A2(n_155),
.B(n_153),
.C(n_154),
.Y(n_7498)
);

INVx1_ASAP7_75t_L g7499 ( 
.A(n_6971),
.Y(n_7499)
);

NAND2xp5_ASAP7_75t_L g7500 ( 
.A(n_6870),
.B(n_154),
.Y(n_7500)
);

OAI21xp33_ASAP7_75t_L g7501 ( 
.A1(n_6834),
.A2(n_154),
.B(n_155),
.Y(n_7501)
);

OAI22x1_ASAP7_75t_L g7502 ( 
.A1(n_6864),
.A2(n_158),
.B1(n_156),
.B2(n_157),
.Y(n_7502)
);

OAI21xp33_ASAP7_75t_SL g7503 ( 
.A1(n_6841),
.A2(n_6676),
.B(n_6901),
.Y(n_7503)
);

OAI21x1_ASAP7_75t_L g7504 ( 
.A1(n_6792),
.A2(n_6717),
.B(n_6753),
.Y(n_7504)
);

NOR2xp33_ASAP7_75t_L g7505 ( 
.A(n_6883),
.B(n_1245),
.Y(n_7505)
);

BUFx6f_ASAP7_75t_L g7506 ( 
.A(n_6793),
.Y(n_7506)
);

AND2x4_ASAP7_75t_L g7507 ( 
.A(n_6769),
.B(n_1246),
.Y(n_7507)
);

OAI21xp5_ASAP7_75t_L g7508 ( 
.A1(n_7073),
.A2(n_6924),
.B(n_6910),
.Y(n_7508)
);

NAND2xp5_ASAP7_75t_L g7509 ( 
.A(n_6862),
.B(n_6931),
.Y(n_7509)
);

AOI21xp5_ASAP7_75t_L g7510 ( 
.A1(n_7073),
.A2(n_1249),
.B(n_1248),
.Y(n_7510)
);

NAND2xp5_ASAP7_75t_SL g7511 ( 
.A(n_6969),
.B(n_1249),
.Y(n_7511)
);

INVx1_ASAP7_75t_L g7512 ( 
.A(n_6839),
.Y(n_7512)
);

CKINVDCx5p33_ASAP7_75t_R g7513 ( 
.A(n_7085),
.Y(n_7513)
);

NAND2xp5_ASAP7_75t_L g7514 ( 
.A(n_6865),
.B(n_156),
.Y(n_7514)
);

BUFx6f_ASAP7_75t_L g7515 ( 
.A(n_6793),
.Y(n_7515)
);

INVx3_ASAP7_75t_L g7516 ( 
.A(n_6868),
.Y(n_7516)
);

OAI22xp5_ASAP7_75t_L g7517 ( 
.A1(n_6840),
.A2(n_159),
.B1(n_156),
.B2(n_157),
.Y(n_7517)
);

NAND2xp5_ASAP7_75t_L g7518 ( 
.A(n_6863),
.B(n_157),
.Y(n_7518)
);

NAND2xp5_ASAP7_75t_L g7519 ( 
.A(n_6824),
.B(n_159),
.Y(n_7519)
);

AOI21xp5_ASAP7_75t_L g7520 ( 
.A1(n_6855),
.A2(n_6896),
.B(n_6840),
.Y(n_7520)
);

NAND2xp5_ASAP7_75t_L g7521 ( 
.A(n_6869),
.B(n_160),
.Y(n_7521)
);

AND2x2_ASAP7_75t_L g7522 ( 
.A(n_6770),
.B(n_160),
.Y(n_7522)
);

NOR2xp67_ASAP7_75t_L g7523 ( 
.A(n_6977),
.B(n_6896),
.Y(n_7523)
);

INVx1_ASAP7_75t_L g7524 ( 
.A(n_6705),
.Y(n_7524)
);

NAND2xp5_ASAP7_75t_L g7525 ( 
.A(n_6933),
.B(n_161),
.Y(n_7525)
);

BUFx8_ASAP7_75t_L g7526 ( 
.A(n_6764),
.Y(n_7526)
);

CKINVDCx10_ASAP7_75t_R g7527 ( 
.A(n_6749),
.Y(n_7527)
);

AOI21xp5_ASAP7_75t_L g7528 ( 
.A1(n_6977),
.A2(n_1251),
.B(n_1250),
.Y(n_7528)
);

A2O1A1Ixp33_ASAP7_75t_L g7529 ( 
.A1(n_6723),
.A2(n_163),
.B(n_161),
.C(n_162),
.Y(n_7529)
);

AND2x2_ASAP7_75t_L g7530 ( 
.A(n_7008),
.B(n_161),
.Y(n_7530)
);

NOR2xp33_ASAP7_75t_L g7531 ( 
.A(n_6966),
.B(n_1250),
.Y(n_7531)
);

AOI22xp33_ASAP7_75t_L g7532 ( 
.A1(n_7002),
.A2(n_164),
.B1(n_162),
.B2(n_163),
.Y(n_7532)
);

INVx2_ASAP7_75t_L g7533 ( 
.A(n_6663),
.Y(n_7533)
);

INVx1_ASAP7_75t_L g7534 ( 
.A(n_6663),
.Y(n_7534)
);

OAI22xp5_ASAP7_75t_L g7535 ( 
.A1(n_6736),
.A2(n_165),
.B1(n_163),
.B2(n_164),
.Y(n_7535)
);

INVx1_ASAP7_75t_L g7536 ( 
.A(n_7199),
.Y(n_7536)
);

INVx2_ASAP7_75t_L g7537 ( 
.A(n_7112),
.Y(n_7537)
);

BUFx6f_ASAP7_75t_L g7538 ( 
.A(n_7218),
.Y(n_7538)
);

AOI22xp33_ASAP7_75t_L g7539 ( 
.A1(n_7298),
.A2(n_167),
.B1(n_165),
.B2(n_166),
.Y(n_7539)
);

NAND2xp5_ASAP7_75t_L g7540 ( 
.A(n_7115),
.B(n_1251),
.Y(n_7540)
);

INVx1_ASAP7_75t_L g7541 ( 
.A(n_7202),
.Y(n_7541)
);

BUFx6f_ASAP7_75t_L g7542 ( 
.A(n_7176),
.Y(n_7542)
);

INVx1_ASAP7_75t_L g7543 ( 
.A(n_7234),
.Y(n_7543)
);

INVx1_ASAP7_75t_L g7544 ( 
.A(n_7253),
.Y(n_7544)
);

NAND2x1p5_ASAP7_75t_L g7545 ( 
.A(n_7171),
.B(n_1252),
.Y(n_7545)
);

NAND2xp33_ASAP7_75t_L g7546 ( 
.A(n_7501),
.B(n_166),
.Y(n_7546)
);

OAI22xp33_ASAP7_75t_L g7547 ( 
.A1(n_7329),
.A2(n_1253),
.B1(n_1254),
.B2(n_1252),
.Y(n_7547)
);

INVx3_ASAP7_75t_L g7548 ( 
.A(n_7437),
.Y(n_7548)
);

AOI22xp33_ASAP7_75t_L g7549 ( 
.A1(n_7103),
.A2(n_168),
.B1(n_166),
.B2(n_167),
.Y(n_7549)
);

INVx2_ASAP7_75t_L g7550 ( 
.A(n_7137),
.Y(n_7550)
);

HB1xp67_ASAP7_75t_L g7551 ( 
.A(n_7389),
.Y(n_7551)
);

AOI21xp5_ASAP7_75t_L g7552 ( 
.A1(n_7107),
.A2(n_1254),
.B(n_1253),
.Y(n_7552)
);

AOI22xp33_ASAP7_75t_L g7553 ( 
.A1(n_7485),
.A2(n_169),
.B1(n_167),
.B2(n_168),
.Y(n_7553)
);

BUFx6f_ASAP7_75t_L g7554 ( 
.A(n_7466),
.Y(n_7554)
);

INVxp67_ASAP7_75t_SL g7555 ( 
.A(n_7266),
.Y(n_7555)
);

INVx1_ASAP7_75t_L g7556 ( 
.A(n_7261),
.Y(n_7556)
);

INVx1_ASAP7_75t_L g7557 ( 
.A(n_7262),
.Y(n_7557)
);

NAND2xp5_ASAP7_75t_L g7558 ( 
.A(n_7191),
.B(n_1255),
.Y(n_7558)
);

INVx3_ASAP7_75t_L g7559 ( 
.A(n_7437),
.Y(n_7559)
);

INVx2_ASAP7_75t_SL g7560 ( 
.A(n_7420),
.Y(n_7560)
);

INVx1_ASAP7_75t_L g7561 ( 
.A(n_7264),
.Y(n_7561)
);

AND2x4_ASAP7_75t_L g7562 ( 
.A(n_7214),
.B(n_1255),
.Y(n_7562)
);

OAI21x1_ASAP7_75t_L g7563 ( 
.A1(n_7275),
.A2(n_168),
.B(n_169),
.Y(n_7563)
);

AND2x4_ASAP7_75t_L g7564 ( 
.A(n_7228),
.B(n_1256),
.Y(n_7564)
);

INVx1_ASAP7_75t_SL g7565 ( 
.A(n_7130),
.Y(n_7565)
);

HB1xp67_ASAP7_75t_L g7566 ( 
.A(n_7185),
.Y(n_7566)
);

BUFx6f_ASAP7_75t_L g7567 ( 
.A(n_7466),
.Y(n_7567)
);

INVx2_ASAP7_75t_SL g7568 ( 
.A(n_7231),
.Y(n_7568)
);

INVx2_ASAP7_75t_L g7569 ( 
.A(n_7139),
.Y(n_7569)
);

INVx2_ASAP7_75t_L g7570 ( 
.A(n_7225),
.Y(n_7570)
);

AND3x1_ASAP7_75t_SL g7571 ( 
.A(n_7524),
.B(n_169),
.C(n_170),
.Y(n_7571)
);

INVx3_ASAP7_75t_L g7572 ( 
.A(n_7456),
.Y(n_7572)
);

INVx6_ASAP7_75t_L g7573 ( 
.A(n_7240),
.Y(n_7573)
);

BUFx6f_ASAP7_75t_L g7574 ( 
.A(n_7302),
.Y(n_7574)
);

INVx2_ASAP7_75t_SL g7575 ( 
.A(n_7231),
.Y(n_7575)
);

INVx1_ASAP7_75t_L g7576 ( 
.A(n_7272),
.Y(n_7576)
);

OAI22xp5_ASAP7_75t_L g7577 ( 
.A1(n_7111),
.A2(n_172),
.B1(n_170),
.B2(n_171),
.Y(n_7577)
);

BUFx6f_ASAP7_75t_L g7578 ( 
.A(n_7302),
.Y(n_7578)
);

INVx3_ASAP7_75t_L g7579 ( 
.A(n_7456),
.Y(n_7579)
);

INVx2_ASAP7_75t_L g7580 ( 
.A(n_7260),
.Y(n_7580)
);

INVx1_ASAP7_75t_L g7581 ( 
.A(n_7278),
.Y(n_7581)
);

AOI21xp5_ASAP7_75t_L g7582 ( 
.A1(n_7108),
.A2(n_1257),
.B(n_1256),
.Y(n_7582)
);

AND2x4_ASAP7_75t_L g7583 ( 
.A(n_7310),
.B(n_1257),
.Y(n_7583)
);

NAND2xp5_ASAP7_75t_L g7584 ( 
.A(n_7304),
.B(n_1258),
.Y(n_7584)
);

INVx2_ASAP7_75t_L g7585 ( 
.A(n_7533),
.Y(n_7585)
);

CKINVDCx8_ASAP7_75t_R g7586 ( 
.A(n_7527),
.Y(n_7586)
);

INVx1_ASAP7_75t_L g7587 ( 
.A(n_7309),
.Y(n_7587)
);

INVx3_ASAP7_75t_L g7588 ( 
.A(n_7410),
.Y(n_7588)
);

BUFx12f_ASAP7_75t_L g7589 ( 
.A(n_7248),
.Y(n_7589)
);

INVx2_ASAP7_75t_L g7590 ( 
.A(n_7409),
.Y(n_7590)
);

AND2x4_ASAP7_75t_L g7591 ( 
.A(n_7133),
.B(n_1258),
.Y(n_7591)
);

INVx5_ASAP7_75t_L g7592 ( 
.A(n_7282),
.Y(n_7592)
);

INVx1_ASAP7_75t_L g7593 ( 
.A(n_7315),
.Y(n_7593)
);

BUFx6f_ASAP7_75t_L g7594 ( 
.A(n_7348),
.Y(n_7594)
);

A2O1A1Ixp33_ASAP7_75t_L g7595 ( 
.A1(n_7110),
.A2(n_1261),
.B(n_1262),
.C(n_1259),
.Y(n_7595)
);

BUFx8_ASAP7_75t_L g7596 ( 
.A(n_7233),
.Y(n_7596)
);

OAI21xp33_ASAP7_75t_SL g7597 ( 
.A1(n_7447),
.A2(n_1262),
.B(n_1261),
.Y(n_7597)
);

A2O1A1Ixp33_ASAP7_75t_SL g7598 ( 
.A1(n_7128),
.A2(n_173),
.B(n_171),
.C(n_172),
.Y(n_7598)
);

OAI22xp5_ASAP7_75t_L g7599 ( 
.A1(n_7124),
.A2(n_7150),
.B1(n_7140),
.B2(n_7307),
.Y(n_7599)
);

NAND2xp5_ASAP7_75t_L g7600 ( 
.A(n_7104),
.B(n_1263),
.Y(n_7600)
);

OR2x6_ASAP7_75t_L g7601 ( 
.A(n_7520),
.B(n_1264),
.Y(n_7601)
);

AOI22xp33_ASAP7_75t_L g7602 ( 
.A1(n_7177),
.A2(n_175),
.B1(n_172),
.B2(n_174),
.Y(n_7602)
);

INVx4_ASAP7_75t_L g7603 ( 
.A(n_7231),
.Y(n_7603)
);

NAND2xp5_ASAP7_75t_L g7604 ( 
.A(n_7223),
.B(n_1264),
.Y(n_7604)
);

O2A1O1Ixp33_ASAP7_75t_L g7605 ( 
.A1(n_7152),
.A2(n_176),
.B(n_174),
.C(n_175),
.Y(n_7605)
);

INVx4_ASAP7_75t_L g7606 ( 
.A(n_7171),
.Y(n_7606)
);

CKINVDCx5p33_ASAP7_75t_R g7607 ( 
.A(n_7109),
.Y(n_7607)
);

NAND2xp5_ASAP7_75t_SL g7608 ( 
.A(n_7326),
.B(n_1265),
.Y(n_7608)
);

BUFx6f_ASAP7_75t_L g7609 ( 
.A(n_7348),
.Y(n_7609)
);

BUFx2_ASAP7_75t_L g7610 ( 
.A(n_7144),
.Y(n_7610)
);

BUFx6f_ASAP7_75t_L g7611 ( 
.A(n_7204),
.Y(n_7611)
);

AND2x4_ASAP7_75t_L g7612 ( 
.A(n_7370),
.B(n_1265),
.Y(n_7612)
);

NAND2xp5_ASAP7_75t_L g7613 ( 
.A(n_7316),
.B(n_1266),
.Y(n_7613)
);

INVxp67_ASAP7_75t_SL g7614 ( 
.A(n_7379),
.Y(n_7614)
);

NAND2xp5_ASAP7_75t_L g7615 ( 
.A(n_7305),
.B(n_1266),
.Y(n_7615)
);

INVx1_ASAP7_75t_L g7616 ( 
.A(n_7341),
.Y(n_7616)
);

OAI22xp5_ASAP7_75t_L g7617 ( 
.A1(n_7489),
.A2(n_176),
.B1(n_174),
.B2(n_175),
.Y(n_7617)
);

BUFx2_ASAP7_75t_L g7618 ( 
.A(n_7428),
.Y(n_7618)
);

BUFx2_ASAP7_75t_L g7619 ( 
.A(n_7346),
.Y(n_7619)
);

AOI22xp33_ASAP7_75t_L g7620 ( 
.A1(n_7208),
.A2(n_179),
.B1(n_177),
.B2(n_178),
.Y(n_7620)
);

OR2x2_ASAP7_75t_L g7621 ( 
.A(n_7449),
.B(n_7289),
.Y(n_7621)
);

NAND2x1p5_ASAP7_75t_L g7622 ( 
.A(n_7171),
.B(n_1267),
.Y(n_7622)
);

BUFx2_ASAP7_75t_SL g7623 ( 
.A(n_7523),
.Y(n_7623)
);

INVx1_ASAP7_75t_L g7624 ( 
.A(n_7343),
.Y(n_7624)
);

INVx5_ASAP7_75t_L g7625 ( 
.A(n_7470),
.Y(n_7625)
);

INVx8_ASAP7_75t_L g7626 ( 
.A(n_7470),
.Y(n_7626)
);

HB1xp67_ASAP7_75t_L g7627 ( 
.A(n_7355),
.Y(n_7627)
);

INVx2_ASAP7_75t_SL g7628 ( 
.A(n_7506),
.Y(n_7628)
);

INVx1_ASAP7_75t_L g7629 ( 
.A(n_7349),
.Y(n_7629)
);

INVx1_ASAP7_75t_L g7630 ( 
.A(n_7361),
.Y(n_7630)
);

AND2x2_ASAP7_75t_L g7631 ( 
.A(n_7132),
.B(n_1267),
.Y(n_7631)
);

BUFx6f_ASAP7_75t_L g7632 ( 
.A(n_7506),
.Y(n_7632)
);

INVxp67_ASAP7_75t_L g7633 ( 
.A(n_7380),
.Y(n_7633)
);

BUFx6f_ASAP7_75t_L g7634 ( 
.A(n_7515),
.Y(n_7634)
);

HB1xp67_ASAP7_75t_L g7635 ( 
.A(n_7125),
.Y(n_7635)
);

INVx1_ASAP7_75t_L g7636 ( 
.A(n_7397),
.Y(n_7636)
);

NOR2xp33_ASAP7_75t_SL g7637 ( 
.A(n_7430),
.B(n_177),
.Y(n_7637)
);

BUFx2_ASAP7_75t_L g7638 ( 
.A(n_7503),
.Y(n_7638)
);

NAND2xp5_ASAP7_75t_L g7639 ( 
.A(n_7118),
.B(n_7119),
.Y(n_7639)
);

INVx2_ASAP7_75t_L g7640 ( 
.A(n_7481),
.Y(n_7640)
);

INVx2_ASAP7_75t_L g7641 ( 
.A(n_7280),
.Y(n_7641)
);

INVx1_ASAP7_75t_L g7642 ( 
.A(n_7400),
.Y(n_7642)
);

OAI22xp5_ASAP7_75t_L g7643 ( 
.A1(n_7255),
.A2(n_181),
.B1(n_179),
.B2(n_180),
.Y(n_7643)
);

INVx2_ASAP7_75t_L g7644 ( 
.A(n_7288),
.Y(n_7644)
);

INVx4_ASAP7_75t_L g7645 ( 
.A(n_7123),
.Y(n_7645)
);

NOR2xp33_ASAP7_75t_L g7646 ( 
.A(n_7251),
.B(n_1268),
.Y(n_7646)
);

INVxp67_ASAP7_75t_SL g7647 ( 
.A(n_7458),
.Y(n_7647)
);

AOI21xp5_ASAP7_75t_L g7648 ( 
.A1(n_7113),
.A2(n_1270),
.B(n_1269),
.Y(n_7648)
);

INVx3_ASAP7_75t_L g7649 ( 
.A(n_7410),
.Y(n_7649)
);

AND2x2_ASAP7_75t_L g7650 ( 
.A(n_7236),
.B(n_1271),
.Y(n_7650)
);

AOI22xp5_ASAP7_75t_L g7651 ( 
.A1(n_7114),
.A2(n_182),
.B1(n_180),
.B2(n_181),
.Y(n_7651)
);

AND3x2_ASAP7_75t_L g7652 ( 
.A(n_7372),
.B(n_180),
.C(n_181),
.Y(n_7652)
);

BUFx12f_ASAP7_75t_L g7653 ( 
.A(n_7189),
.Y(n_7653)
);

A2O1A1Ixp33_ASAP7_75t_L g7654 ( 
.A1(n_7196),
.A2(n_1272),
.B(n_1274),
.C(n_1271),
.Y(n_7654)
);

INVx3_ASAP7_75t_L g7655 ( 
.A(n_7413),
.Y(n_7655)
);

AOI22xp33_ASAP7_75t_L g7656 ( 
.A1(n_7419),
.A2(n_184),
.B1(n_182),
.B2(n_183),
.Y(n_7656)
);

INVx2_ASAP7_75t_SL g7657 ( 
.A(n_7515),
.Y(n_7657)
);

INVx2_ASAP7_75t_L g7658 ( 
.A(n_7290),
.Y(n_7658)
);

OR2x6_ASAP7_75t_L g7659 ( 
.A(n_7370),
.B(n_1272),
.Y(n_7659)
);

NAND2x1p5_ASAP7_75t_L g7660 ( 
.A(n_7333),
.B(n_1274),
.Y(n_7660)
);

NAND2xp5_ASAP7_75t_L g7661 ( 
.A(n_7376),
.B(n_1275),
.Y(n_7661)
);

INVx1_ASAP7_75t_L g7662 ( 
.A(n_7405),
.Y(n_7662)
);

AOI22xp5_ASAP7_75t_L g7663 ( 
.A1(n_7382),
.A2(n_184),
.B1(n_182),
.B2(n_183),
.Y(n_7663)
);

OR2x6_ASAP7_75t_L g7664 ( 
.A(n_7508),
.B(n_1275),
.Y(n_7664)
);

NAND3xp33_ASAP7_75t_L g7665 ( 
.A(n_7149),
.B(n_184),
.C(n_185),
.Y(n_7665)
);

INVx1_ASAP7_75t_L g7666 ( 
.A(n_7422),
.Y(n_7666)
);

OAI22xp5_ASAP7_75t_L g7667 ( 
.A1(n_7342),
.A2(n_187),
.B1(n_185),
.B2(n_186),
.Y(n_7667)
);

INVx2_ASAP7_75t_L g7668 ( 
.A(n_7295),
.Y(n_7668)
);

NAND2xp5_ASAP7_75t_L g7669 ( 
.A(n_7327),
.B(n_1276),
.Y(n_7669)
);

INVx1_ASAP7_75t_SL g7670 ( 
.A(n_7479),
.Y(n_7670)
);

NAND2xp5_ASAP7_75t_L g7671 ( 
.A(n_7324),
.B(n_1277),
.Y(n_7671)
);

INVx5_ASAP7_75t_L g7672 ( 
.A(n_7169),
.Y(n_7672)
);

INVxp67_ASAP7_75t_L g7673 ( 
.A(n_7509),
.Y(n_7673)
);

NAND2x1p5_ASAP7_75t_L g7674 ( 
.A(n_7105),
.B(n_1277),
.Y(n_7674)
);

CKINVDCx11_ASAP7_75t_R g7675 ( 
.A(n_7232),
.Y(n_7675)
);

OR2x6_ASAP7_75t_L g7676 ( 
.A(n_7273),
.B(n_1278),
.Y(n_7676)
);

BUFx6f_ASAP7_75t_L g7677 ( 
.A(n_7371),
.Y(n_7677)
);

HB1xp67_ASAP7_75t_L g7678 ( 
.A(n_7106),
.Y(n_7678)
);

AND2x4_ASAP7_75t_L g7679 ( 
.A(n_7135),
.B(n_1279),
.Y(n_7679)
);

INVxp67_ASAP7_75t_SL g7680 ( 
.A(n_7116),
.Y(n_7680)
);

INVx5_ASAP7_75t_L g7681 ( 
.A(n_7371),
.Y(n_7681)
);

INVx2_ASAP7_75t_SL g7682 ( 
.A(n_7413),
.Y(n_7682)
);

INVx1_ASAP7_75t_L g7683 ( 
.A(n_7432),
.Y(n_7683)
);

BUFx2_ASAP7_75t_L g7684 ( 
.A(n_7516),
.Y(n_7684)
);

INVx5_ASAP7_75t_L g7685 ( 
.A(n_7491),
.Y(n_7685)
);

NOR2xp33_ASAP7_75t_L g7686 ( 
.A(n_7120),
.B(n_1280),
.Y(n_7686)
);

INVxp67_ASAP7_75t_L g7687 ( 
.A(n_7414),
.Y(n_7687)
);

INVx2_ASAP7_75t_SL g7688 ( 
.A(n_7308),
.Y(n_7688)
);

INVx3_ASAP7_75t_L g7689 ( 
.A(n_7491),
.Y(n_7689)
);

INVx1_ASAP7_75t_SL g7690 ( 
.A(n_7360),
.Y(n_7690)
);

INVx2_ASAP7_75t_L g7691 ( 
.A(n_7313),
.Y(n_7691)
);

OAI22xp5_ASAP7_75t_L g7692 ( 
.A1(n_7154),
.A2(n_187),
.B1(n_185),
.B2(n_186),
.Y(n_7692)
);

HB1xp67_ASAP7_75t_L g7693 ( 
.A(n_7121),
.Y(n_7693)
);

OAI22xp5_ASAP7_75t_L g7694 ( 
.A1(n_7269),
.A2(n_189),
.B1(n_187),
.B2(n_188),
.Y(n_7694)
);

BUFx4f_ASAP7_75t_L g7695 ( 
.A(n_7390),
.Y(n_7695)
);

AND2x4_ASAP7_75t_L g7696 ( 
.A(n_7373),
.B(n_1280),
.Y(n_7696)
);

OAI21x1_ASAP7_75t_SL g7697 ( 
.A1(n_7247),
.A2(n_188),
.B(n_189),
.Y(n_7697)
);

INVx1_ASAP7_75t_L g7698 ( 
.A(n_7443),
.Y(n_7698)
);

NAND2xp5_ASAP7_75t_SL g7699 ( 
.A(n_7402),
.B(n_1281),
.Y(n_7699)
);

INVx1_ASAP7_75t_L g7700 ( 
.A(n_7445),
.Y(n_7700)
);

HB1xp67_ASAP7_75t_L g7701 ( 
.A(n_7134),
.Y(n_7701)
);

AOI221x1_ASAP7_75t_L g7702 ( 
.A1(n_7160),
.A2(n_1285),
.B1(n_1286),
.B2(n_1283),
.C(n_1282),
.Y(n_7702)
);

BUFx2_ASAP7_75t_L g7703 ( 
.A(n_7117),
.Y(n_7703)
);

CKINVDCx6p67_ASAP7_75t_R g7704 ( 
.A(n_7273),
.Y(n_7704)
);

BUFx2_ASAP7_75t_L g7705 ( 
.A(n_7117),
.Y(n_7705)
);

NAND2xp33_ASAP7_75t_L g7706 ( 
.A(n_7495),
.B(n_189),
.Y(n_7706)
);

INVx1_ASAP7_75t_L g7707 ( 
.A(n_7446),
.Y(n_7707)
);

INVx3_ASAP7_75t_L g7708 ( 
.A(n_7390),
.Y(n_7708)
);

INVx4_ASAP7_75t_L g7709 ( 
.A(n_7195),
.Y(n_7709)
);

BUFx3_ASAP7_75t_L g7710 ( 
.A(n_7526),
.Y(n_7710)
);

AOI21x1_ASAP7_75t_L g7711 ( 
.A1(n_7142),
.A2(n_7165),
.B(n_7271),
.Y(n_7711)
);

BUFx2_ASAP7_75t_L g7712 ( 
.A(n_7122),
.Y(n_7712)
);

INVx2_ASAP7_75t_L g7713 ( 
.A(n_7314),
.Y(n_7713)
);

BUFx2_ASAP7_75t_SL g7714 ( 
.A(n_7244),
.Y(n_7714)
);

AND2x4_ASAP7_75t_L g7715 ( 
.A(n_7512),
.B(n_1283),
.Y(n_7715)
);

NAND2xp5_ASAP7_75t_L g7716 ( 
.A(n_7363),
.B(n_1286),
.Y(n_7716)
);

CKINVDCx5p33_ASAP7_75t_R g7717 ( 
.A(n_7385),
.Y(n_7717)
);

OR2x6_ASAP7_75t_L g7718 ( 
.A(n_7157),
.B(n_1287),
.Y(n_7718)
);

INVx4_ASAP7_75t_L g7719 ( 
.A(n_7179),
.Y(n_7719)
);

INVx3_ASAP7_75t_L g7720 ( 
.A(n_7180),
.Y(n_7720)
);

BUFx3_ASAP7_75t_L g7721 ( 
.A(n_7127),
.Y(n_7721)
);

A2O1A1Ixp33_ASAP7_75t_L g7722 ( 
.A1(n_7403),
.A2(n_1289),
.B(n_1290),
.C(n_1288),
.Y(n_7722)
);

AOI22xp33_ASAP7_75t_L g7723 ( 
.A1(n_7499),
.A2(n_7205),
.B1(n_7388),
.B2(n_7535),
.Y(n_7723)
);

CKINVDCx6p67_ASAP7_75t_R g7724 ( 
.A(n_7301),
.Y(n_7724)
);

BUFx3_ASAP7_75t_L g7725 ( 
.A(n_7492),
.Y(n_7725)
);

INVx1_ASAP7_75t_L g7726 ( 
.A(n_7457),
.Y(n_7726)
);

INVx1_ASAP7_75t_L g7727 ( 
.A(n_7534),
.Y(n_7727)
);

INVx3_ASAP7_75t_L g7728 ( 
.A(n_7319),
.Y(n_7728)
);

CKINVDCx11_ASAP7_75t_R g7729 ( 
.A(n_7157),
.Y(n_7729)
);

BUFx2_ASAP7_75t_L g7730 ( 
.A(n_7473),
.Y(n_7730)
);

BUFx6f_ASAP7_75t_L g7731 ( 
.A(n_7454),
.Y(n_7731)
);

INVx1_ASAP7_75t_L g7732 ( 
.A(n_7136),
.Y(n_7732)
);

AOI22xp33_ASAP7_75t_L g7733 ( 
.A1(n_7483),
.A2(n_192),
.B1(n_190),
.B2(n_191),
.Y(n_7733)
);

NAND2x1p5_ASAP7_75t_L g7734 ( 
.A(n_7504),
.B(n_7286),
.Y(n_7734)
);

AOI221x1_ASAP7_75t_L g7735 ( 
.A1(n_7502),
.A2(n_1290),
.B1(n_1291),
.B2(n_1289),
.C(n_1288),
.Y(n_7735)
);

AND2x2_ASAP7_75t_L g7736 ( 
.A(n_7250),
.B(n_1292),
.Y(n_7736)
);

AND2x4_ASAP7_75t_L g7737 ( 
.A(n_7490),
.B(n_1292),
.Y(n_7737)
);

INVx1_ASAP7_75t_L g7738 ( 
.A(n_7146),
.Y(n_7738)
);

INVx4_ASAP7_75t_L g7739 ( 
.A(n_7394),
.Y(n_7739)
);

INVx2_ASAP7_75t_L g7740 ( 
.A(n_7358),
.Y(n_7740)
);

AOI22xp33_ASAP7_75t_L g7741 ( 
.A1(n_7426),
.A2(n_192),
.B1(n_190),
.B2(n_191),
.Y(n_7741)
);

OR2x6_ASAP7_75t_L g7742 ( 
.A(n_7163),
.B(n_1293),
.Y(n_7742)
);

OR2x6_ASAP7_75t_L g7743 ( 
.A(n_7488),
.B(n_1294),
.Y(n_7743)
);

BUFx6f_ASAP7_75t_L g7744 ( 
.A(n_7450),
.Y(n_7744)
);

INVx3_ASAP7_75t_L g7745 ( 
.A(n_7366),
.Y(n_7745)
);

OR2x6_ASAP7_75t_L g7746 ( 
.A(n_7328),
.B(n_1294),
.Y(n_7746)
);

INVx2_ASAP7_75t_L g7747 ( 
.A(n_7386),
.Y(n_7747)
);

NAND2xp5_ASAP7_75t_L g7748 ( 
.A(n_7174),
.B(n_1297),
.Y(n_7748)
);

BUFx2_ASAP7_75t_L g7749 ( 
.A(n_7162),
.Y(n_7749)
);

BUFx2_ASAP7_75t_L g7750 ( 
.A(n_7170),
.Y(n_7750)
);

CKINVDCx20_ASAP7_75t_R g7751 ( 
.A(n_7441),
.Y(n_7751)
);

CKINVDCx11_ASAP7_75t_R g7752 ( 
.A(n_7190),
.Y(n_7752)
);

AOI22xp33_ASAP7_75t_L g7753 ( 
.A1(n_7354),
.A2(n_193),
.B1(n_190),
.B2(n_191),
.Y(n_7753)
);

INVx3_ASAP7_75t_L g7754 ( 
.A(n_7396),
.Y(n_7754)
);

AOI221x1_ASAP7_75t_L g7755 ( 
.A1(n_7472),
.A2(n_1299),
.B1(n_1301),
.B2(n_1298),
.C(n_1297),
.Y(n_7755)
);

OR2x2_ASAP7_75t_L g7756 ( 
.A(n_7276),
.B(n_1302),
.Y(n_7756)
);

HB1xp67_ASAP7_75t_L g7757 ( 
.A(n_7172),
.Y(n_7757)
);

AOI22xp33_ASAP7_75t_L g7758 ( 
.A1(n_7220),
.A2(n_195),
.B1(n_193),
.B2(n_194),
.Y(n_7758)
);

O2A1O1Ixp33_ASAP7_75t_L g7759 ( 
.A1(n_7404),
.A2(n_195),
.B(n_193),
.C(n_194),
.Y(n_7759)
);

INVx1_ASAP7_75t_L g7760 ( 
.A(n_7173),
.Y(n_7760)
);

INVx1_ASAP7_75t_L g7761 ( 
.A(n_7197),
.Y(n_7761)
);

BUFx2_ASAP7_75t_L g7762 ( 
.A(n_7477),
.Y(n_7762)
);

AOI21xp5_ASAP7_75t_L g7763 ( 
.A1(n_7235),
.A2(n_1305),
.B(n_1303),
.Y(n_7763)
);

BUFx6f_ASAP7_75t_L g7764 ( 
.A(n_7507),
.Y(n_7764)
);

OR2x2_ASAP7_75t_L g7765 ( 
.A(n_7323),
.B(n_7444),
.Y(n_7765)
);

BUFx6f_ASAP7_75t_L g7766 ( 
.A(n_7221),
.Y(n_7766)
);

INVx2_ASAP7_75t_L g7767 ( 
.A(n_7461),
.Y(n_7767)
);

INVx3_ASAP7_75t_L g7768 ( 
.A(n_7476),
.Y(n_7768)
);

INVx1_ASAP7_75t_L g7769 ( 
.A(n_7317),
.Y(n_7769)
);

AND2x2_ASAP7_75t_L g7770 ( 
.A(n_7145),
.B(n_1303),
.Y(n_7770)
);

INVx1_ASAP7_75t_L g7771 ( 
.A(n_7161),
.Y(n_7771)
);

NOR2x1p5_ASAP7_75t_L g7772 ( 
.A(n_7440),
.B(n_194),
.Y(n_7772)
);

NAND2xp5_ASAP7_75t_L g7773 ( 
.A(n_7322),
.B(n_1305),
.Y(n_7773)
);

INVx2_ASAP7_75t_L g7774 ( 
.A(n_7391),
.Y(n_7774)
);

BUFx4_ASAP7_75t_SL g7775 ( 
.A(n_7513),
.Y(n_7775)
);

AOI21xp5_ASAP7_75t_L g7776 ( 
.A1(n_7487),
.A2(n_1307),
.B(n_1306),
.Y(n_7776)
);

AND2x2_ASAP7_75t_L g7777 ( 
.A(n_7164),
.B(n_1306),
.Y(n_7777)
);

CKINVDCx20_ASAP7_75t_R g7778 ( 
.A(n_7364),
.Y(n_7778)
);

INVx1_ASAP7_75t_L g7779 ( 
.A(n_7412),
.Y(n_7779)
);

INVx1_ASAP7_75t_SL g7780 ( 
.A(n_7265),
.Y(n_7780)
);

NOR2xp33_ASAP7_75t_L g7781 ( 
.A(n_7375),
.B(n_1307),
.Y(n_7781)
);

AOI22xp33_ASAP7_75t_L g7782 ( 
.A1(n_7464),
.A2(n_197),
.B1(n_195),
.B2(n_196),
.Y(n_7782)
);

INVx4_ASAP7_75t_L g7783 ( 
.A(n_7306),
.Y(n_7783)
);

OR2x6_ASAP7_75t_L g7784 ( 
.A(n_7406),
.B(n_1309),
.Y(n_7784)
);

AOI22xp33_ASAP7_75t_L g7785 ( 
.A1(n_7216),
.A2(n_198),
.B1(n_196),
.B2(n_197),
.Y(n_7785)
);

INVx3_ASAP7_75t_L g7786 ( 
.A(n_7436),
.Y(n_7786)
);

INVx3_ASAP7_75t_L g7787 ( 
.A(n_7451),
.Y(n_7787)
);

INVx5_ASAP7_75t_L g7788 ( 
.A(n_7522),
.Y(n_7788)
);

NAND2xp5_ASAP7_75t_L g7789 ( 
.A(n_7462),
.B(n_1310),
.Y(n_7789)
);

INVx3_ASAP7_75t_L g7790 ( 
.A(n_7318),
.Y(n_7790)
);

NAND2xp5_ASAP7_75t_L g7791 ( 
.A(n_7198),
.B(n_1310),
.Y(n_7791)
);

NAND2xp5_ASAP7_75t_L g7792 ( 
.A(n_7151),
.B(n_1311),
.Y(n_7792)
);

NAND2xp5_ASAP7_75t_L g7793 ( 
.A(n_7158),
.B(n_1311),
.Y(n_7793)
);

INVx5_ASAP7_75t_L g7794 ( 
.A(n_7378),
.Y(n_7794)
);

AOI22xp33_ASAP7_75t_L g7795 ( 
.A1(n_7337),
.A2(n_199),
.B1(n_197),
.B2(n_198),
.Y(n_7795)
);

HB1xp67_ASAP7_75t_L g7796 ( 
.A(n_7442),
.Y(n_7796)
);

NOR2xp33_ASAP7_75t_R g7797 ( 
.A(n_7352),
.B(n_199),
.Y(n_7797)
);

INVx3_ASAP7_75t_L g7798 ( 
.A(n_7431),
.Y(n_7798)
);

INVx1_ASAP7_75t_L g7799 ( 
.A(n_7213),
.Y(n_7799)
);

INVx3_ASAP7_75t_L g7800 ( 
.A(n_7471),
.Y(n_7800)
);

AOI21xp33_ASAP7_75t_L g7801 ( 
.A1(n_7224),
.A2(n_199),
.B(n_200),
.Y(n_7801)
);

NOR2xp33_ASAP7_75t_L g7802 ( 
.A(n_7141),
.B(n_7340),
.Y(n_7802)
);

NAND2xp5_ASAP7_75t_L g7803 ( 
.A(n_7159),
.B(n_1312),
.Y(n_7803)
);

OAI21xp33_ASAP7_75t_L g7804 ( 
.A1(n_7155),
.A2(n_200),
.B(n_201),
.Y(n_7804)
);

NOR2xp33_ASAP7_75t_L g7805 ( 
.A(n_7279),
.B(n_1313),
.Y(n_7805)
);

AOI21xp5_ASAP7_75t_L g7806 ( 
.A1(n_7493),
.A2(n_1314),
.B(n_1313),
.Y(n_7806)
);

NOR2xp33_ASAP7_75t_L g7807 ( 
.A(n_7303),
.B(n_1314),
.Y(n_7807)
);

AOI221xp5_ASAP7_75t_L g7808 ( 
.A1(n_7212),
.A2(n_202),
.B1(n_200),
.B2(n_201),
.C(n_203),
.Y(n_7808)
);

AND2x2_ASAP7_75t_L g7809 ( 
.A(n_7418),
.B(n_1315),
.Y(n_7809)
);

NAND2xp5_ASAP7_75t_L g7810 ( 
.A(n_7167),
.B(n_1315),
.Y(n_7810)
);

INVx4_ASAP7_75t_L g7811 ( 
.A(n_7530),
.Y(n_7811)
);

INVx2_ASAP7_75t_L g7812 ( 
.A(n_7178),
.Y(n_7812)
);

INVxp67_ASAP7_75t_SL g7813 ( 
.A(n_7299),
.Y(n_7813)
);

BUFx2_ASAP7_75t_L g7814 ( 
.A(n_7484),
.Y(n_7814)
);

NAND2xp5_ASAP7_75t_L g7815 ( 
.A(n_7156),
.B(n_1316),
.Y(n_7815)
);

AND2x4_ASAP7_75t_L g7816 ( 
.A(n_7334),
.B(n_1316),
.Y(n_7816)
);

NAND2xp5_ASAP7_75t_L g7817 ( 
.A(n_7215),
.B(n_1318),
.Y(n_7817)
);

INVx1_ASAP7_75t_L g7818 ( 
.A(n_7200),
.Y(n_7818)
);

AOI22xp33_ASAP7_75t_L g7819 ( 
.A1(n_7455),
.A2(n_204),
.B1(n_202),
.B2(n_203),
.Y(n_7819)
);

INVx2_ASAP7_75t_L g7820 ( 
.A(n_7201),
.Y(n_7820)
);

BUFx2_ASAP7_75t_L g7821 ( 
.A(n_7335),
.Y(n_7821)
);

A2O1A1Ixp33_ASAP7_75t_L g7822 ( 
.A1(n_7423),
.A2(n_7209),
.B(n_7207),
.C(n_7126),
.Y(n_7822)
);

BUFx6f_ASAP7_75t_L g7823 ( 
.A(n_7514),
.Y(n_7823)
);

NOR2xp67_ASAP7_75t_L g7824 ( 
.A(n_7241),
.B(n_202),
.Y(n_7824)
);

AOI22xp5_ASAP7_75t_L g7825 ( 
.A1(n_7219),
.A2(n_206),
.B1(n_204),
.B2(n_205),
.Y(n_7825)
);

INVx1_ASAP7_75t_L g7826 ( 
.A(n_7245),
.Y(n_7826)
);

INVx1_ASAP7_75t_L g7827 ( 
.A(n_7268),
.Y(n_7827)
);

AOI21xp33_ASAP7_75t_L g7828 ( 
.A1(n_7257),
.A2(n_204),
.B(n_205),
.Y(n_7828)
);

INVx1_ASAP7_75t_L g7829 ( 
.A(n_7270),
.Y(n_7829)
);

AOI22xp5_ASAP7_75t_L g7830 ( 
.A1(n_7226),
.A2(n_209),
.B1(n_206),
.B2(n_207),
.Y(n_7830)
);

AOI22xp5_ASAP7_75t_L g7831 ( 
.A1(n_7351),
.A2(n_209),
.B1(n_206),
.B2(n_207),
.Y(n_7831)
);

NAND2xp5_ASAP7_75t_L g7832 ( 
.A(n_7183),
.B(n_1318),
.Y(n_7832)
);

NOR2xp33_ASAP7_75t_L g7833 ( 
.A(n_7325),
.B(n_1319),
.Y(n_7833)
);

NAND2xp5_ASAP7_75t_L g7834 ( 
.A(n_7186),
.B(n_1319),
.Y(n_7834)
);

INVx1_ASAP7_75t_L g7835 ( 
.A(n_7285),
.Y(n_7835)
);

INVx3_ASAP7_75t_L g7836 ( 
.A(n_7518),
.Y(n_7836)
);

CKINVDCx8_ASAP7_75t_R g7837 ( 
.A(n_7143),
.Y(n_7837)
);

AOI22xp33_ASAP7_75t_L g7838 ( 
.A1(n_7320),
.A2(n_210),
.B1(n_207),
.B2(n_209),
.Y(n_7838)
);

AOI22xp5_ASAP7_75t_L g7839 ( 
.A1(n_7362),
.A2(n_212),
.B1(n_210),
.B2(n_211),
.Y(n_7839)
);

INVx1_ASAP7_75t_L g7840 ( 
.A(n_7292),
.Y(n_7840)
);

AOI22xp5_ASAP7_75t_L g7841 ( 
.A1(n_7392),
.A2(n_212),
.B1(n_210),
.B2(n_211),
.Y(n_7841)
);

BUFx6f_ASAP7_75t_L g7842 ( 
.A(n_7521),
.Y(n_7842)
);

INVx1_ASAP7_75t_L g7843 ( 
.A(n_7296),
.Y(n_7843)
);

AOI22xp33_ASAP7_75t_L g7844 ( 
.A1(n_7532),
.A2(n_215),
.B1(n_213),
.B2(n_214),
.Y(n_7844)
);

NAND3xp33_ASAP7_75t_L g7845 ( 
.A(n_7321),
.B(n_213),
.C(n_214),
.Y(n_7845)
);

AOI22xp33_ASAP7_75t_L g7846 ( 
.A1(n_7424),
.A2(n_215),
.B1(n_213),
.B2(n_214),
.Y(n_7846)
);

OAI22xp33_ASAP7_75t_L g7847 ( 
.A1(n_7465),
.A2(n_1321),
.B1(n_1322),
.B2(n_1320),
.Y(n_7847)
);

OR2x2_ASAP7_75t_L g7848 ( 
.A(n_7297),
.B(n_1320),
.Y(n_7848)
);

NAND2xp5_ASAP7_75t_L g7849 ( 
.A(n_7192),
.B(n_1321),
.Y(n_7849)
);

BUFx12f_ASAP7_75t_L g7850 ( 
.A(n_7153),
.Y(n_7850)
);

A2O1A1Ixp33_ASAP7_75t_L g7851 ( 
.A1(n_7131),
.A2(n_1324),
.B(n_1325),
.C(n_1323),
.Y(n_7851)
);

OR2x6_ASAP7_75t_L g7852 ( 
.A(n_7407),
.B(n_1325),
.Y(n_7852)
);

CKINVDCx20_ASAP7_75t_R g7853 ( 
.A(n_7448),
.Y(n_7853)
);

INVx3_ASAP7_75t_SL g7854 ( 
.A(n_7338),
.Y(n_7854)
);

AOI21xp33_ASAP7_75t_L g7855 ( 
.A1(n_7138),
.A2(n_215),
.B(n_216),
.Y(n_7855)
);

AOI22xp33_ASAP7_75t_L g7856 ( 
.A1(n_7478),
.A2(n_218),
.B1(n_216),
.B2(n_217),
.Y(n_7856)
);

NOR2x1_ASAP7_75t_L g7857 ( 
.A(n_7365),
.B(n_1326),
.Y(n_7857)
);

BUFx2_ASAP7_75t_L g7858 ( 
.A(n_7239),
.Y(n_7858)
);

OAI22xp5_ASAP7_75t_L g7859 ( 
.A1(n_7498),
.A2(n_219),
.B1(n_217),
.B2(n_218),
.Y(n_7859)
);

INVx2_ASAP7_75t_L g7860 ( 
.A(n_7203),
.Y(n_7860)
);

AOI222xp33_ASAP7_75t_L g7861 ( 
.A1(n_7347),
.A2(n_7254),
.B1(n_7256),
.B2(n_7274),
.C1(n_7242),
.C2(n_7147),
.Y(n_7861)
);

NOR2x1_ASAP7_75t_SL g7862 ( 
.A(n_7374),
.B(n_1326),
.Y(n_7862)
);

CKINVDCx5p33_ASAP7_75t_R g7863 ( 
.A(n_7421),
.Y(n_7863)
);

BUFx6f_ASAP7_75t_L g7864 ( 
.A(n_7500),
.Y(n_7864)
);

NAND2xp5_ASAP7_75t_L g7865 ( 
.A(n_7210),
.B(n_1328),
.Y(n_7865)
);

INVx2_ASAP7_75t_L g7866 ( 
.A(n_7211),
.Y(n_7866)
);

INVx1_ASAP7_75t_L g7867 ( 
.A(n_7222),
.Y(n_7867)
);

INVx1_ASAP7_75t_L g7868 ( 
.A(n_7229),
.Y(n_7868)
);

BUFx6f_ASAP7_75t_L g7869 ( 
.A(n_7519),
.Y(n_7869)
);

NAND2xp5_ASAP7_75t_L g7870 ( 
.A(n_7230),
.B(n_1328),
.Y(n_7870)
);

AOI22xp33_ASAP7_75t_SL g7871 ( 
.A1(n_7175),
.A2(n_220),
.B1(n_217),
.B2(n_219),
.Y(n_7871)
);

INVx1_ASAP7_75t_SL g7872 ( 
.A(n_7238),
.Y(n_7872)
);

BUFx2_ASAP7_75t_L g7873 ( 
.A(n_7417),
.Y(n_7873)
);

BUFx2_ASAP7_75t_L g7874 ( 
.A(n_7377),
.Y(n_7874)
);

INVx1_ASAP7_75t_SL g7875 ( 
.A(n_7475),
.Y(n_7875)
);

OAI21x1_ASAP7_75t_L g7876 ( 
.A1(n_7168),
.A2(n_219),
.B(n_220),
.Y(n_7876)
);

AND2x6_ASAP7_75t_L g7877 ( 
.A(n_7384),
.B(n_1330),
.Y(n_7877)
);

NAND2xp5_ASAP7_75t_L g7878 ( 
.A(n_7267),
.B(n_1330),
.Y(n_7878)
);

NAND2xp5_ASAP7_75t_L g7879 ( 
.A(n_7281),
.B(n_1331),
.Y(n_7879)
);

NOR2xp33_ASAP7_75t_L g7880 ( 
.A(n_7246),
.B(n_1332),
.Y(n_7880)
);

AOI21xp5_ASAP7_75t_L g7881 ( 
.A1(n_7206),
.A2(n_1333),
.B(n_1332),
.Y(n_7881)
);

BUFx3_ASAP7_75t_L g7882 ( 
.A(n_7148),
.Y(n_7882)
);

INVx1_ASAP7_75t_L g7883 ( 
.A(n_7287),
.Y(n_7883)
);

INVx2_ASAP7_75t_L g7884 ( 
.A(n_7182),
.Y(n_7884)
);

NAND2xp5_ASAP7_75t_L g7885 ( 
.A(n_7482),
.B(n_1333),
.Y(n_7885)
);

NOR2xp33_ASAP7_75t_R g7886 ( 
.A(n_7345),
.B(n_7486),
.Y(n_7886)
);

INVx2_ASAP7_75t_L g7887 ( 
.A(n_7474),
.Y(n_7887)
);

BUFx2_ASAP7_75t_L g7888 ( 
.A(n_7497),
.Y(n_7888)
);

INVx1_ASAP7_75t_L g7889 ( 
.A(n_7311),
.Y(n_7889)
);

NAND2xp5_ASAP7_75t_L g7890 ( 
.A(n_7395),
.B(n_1334),
.Y(n_7890)
);

INVx3_ASAP7_75t_L g7891 ( 
.A(n_7480),
.Y(n_7891)
);

BUFx6f_ASAP7_75t_L g7892 ( 
.A(n_7277),
.Y(n_7892)
);

INVx2_ASAP7_75t_SL g7893 ( 
.A(n_7166),
.Y(n_7893)
);

BUFx6f_ASAP7_75t_L g7894 ( 
.A(n_7217),
.Y(n_7894)
);

NOR2x1_ASAP7_75t_SL g7895 ( 
.A(n_7453),
.B(n_1334),
.Y(n_7895)
);

CKINVDCx6p67_ASAP7_75t_R g7896 ( 
.A(n_7525),
.Y(n_7896)
);

AOI22xp33_ASAP7_75t_L g7897 ( 
.A1(n_7383),
.A2(n_222),
.B1(n_220),
.B2(n_221),
.Y(n_7897)
);

OAI22xp5_ASAP7_75t_SL g7898 ( 
.A1(n_7505),
.A2(n_223),
.B1(n_221),
.B2(n_222),
.Y(n_7898)
);

AOI22xp33_ASAP7_75t_L g7899 ( 
.A1(n_7330),
.A2(n_224),
.B1(n_222),
.B2(n_223),
.Y(n_7899)
);

INVx3_ASAP7_75t_L g7900 ( 
.A(n_7401),
.Y(n_7900)
);

CKINVDCx20_ASAP7_75t_R g7901 ( 
.A(n_7381),
.Y(n_7901)
);

INVx1_ASAP7_75t_SL g7902 ( 
.A(n_7259),
.Y(n_7902)
);

INVx1_ASAP7_75t_L g7903 ( 
.A(n_7311),
.Y(n_7903)
);

BUFx6f_ASAP7_75t_L g7904 ( 
.A(n_7459),
.Y(n_7904)
);

AND2x4_ASAP7_75t_L g7905 ( 
.A(n_7427),
.B(n_1335),
.Y(n_7905)
);

NAND2xp5_ASAP7_75t_L g7906 ( 
.A(n_7350),
.B(n_1335),
.Y(n_7906)
);

OAI21xp5_ASAP7_75t_L g7907 ( 
.A1(n_7368),
.A2(n_224),
.B(n_226),
.Y(n_7907)
);

BUFx3_ASAP7_75t_L g7908 ( 
.A(n_7243),
.Y(n_7908)
);

INVx3_ASAP7_75t_L g7909 ( 
.A(n_7434),
.Y(n_7909)
);

AO21x2_ASAP7_75t_L g7910 ( 
.A1(n_7332),
.A2(n_224),
.B(n_226),
.Y(n_7910)
);

AOI22xp33_ASAP7_75t_L g7911 ( 
.A1(n_7187),
.A2(n_228),
.B1(n_226),
.B2(n_227),
.Y(n_7911)
);

BUFx3_ASAP7_75t_L g7912 ( 
.A(n_7399),
.Y(n_7912)
);

INVx1_ASAP7_75t_L g7913 ( 
.A(n_7393),
.Y(n_7913)
);

INVx4_ASAP7_75t_L g7914 ( 
.A(n_7469),
.Y(n_7914)
);

HB1xp67_ASAP7_75t_L g7915 ( 
.A(n_7387),
.Y(n_7915)
);

BUFx4f_ASAP7_75t_SL g7916 ( 
.A(n_7511),
.Y(n_7916)
);

INVx1_ASAP7_75t_L g7917 ( 
.A(n_7398),
.Y(n_7917)
);

AND2x2_ASAP7_75t_L g7918 ( 
.A(n_7339),
.B(n_1336),
.Y(n_7918)
);

INVx2_ASAP7_75t_L g7919 ( 
.A(n_7357),
.Y(n_7919)
);

BUFx2_ASAP7_75t_SL g7920 ( 
.A(n_7496),
.Y(n_7920)
);

AOI21xp5_ASAP7_75t_L g7921 ( 
.A1(n_7552),
.A2(n_7188),
.B(n_7181),
.Y(n_7921)
);

OAI22x1_ASAP7_75t_L g7922 ( 
.A1(n_7807),
.A2(n_7531),
.B1(n_7356),
.B2(n_7129),
.Y(n_7922)
);

INVx1_ASAP7_75t_L g7923 ( 
.A(n_7536),
.Y(n_7923)
);

O2A1O1Ixp33_ASAP7_75t_SL g7924 ( 
.A1(n_7595),
.A2(n_7468),
.B(n_7529),
.C(n_7312),
.Y(n_7924)
);

AO31x2_ASAP7_75t_L g7925 ( 
.A1(n_7771),
.A2(n_7415),
.A3(n_7416),
.B(n_7408),
.Y(n_7925)
);

AO31x2_ASAP7_75t_L g7926 ( 
.A1(n_7799),
.A2(n_7252),
.A3(n_7258),
.B(n_7249),
.Y(n_7926)
);

OAI21x1_ASAP7_75t_L g7927 ( 
.A1(n_7774),
.A2(n_7429),
.B(n_7425),
.Y(n_7927)
);

AOI21xp5_ASAP7_75t_L g7928 ( 
.A1(n_7546),
.A2(n_7194),
.B(n_7193),
.Y(n_7928)
);

OAI22xp5_ASAP7_75t_L g7929 ( 
.A1(n_7599),
.A2(n_7467),
.B1(n_7411),
.B2(n_7184),
.Y(n_7929)
);

AOI21xp5_ASAP7_75t_L g7930 ( 
.A1(n_7582),
.A2(n_7237),
.B(n_7227),
.Y(n_7930)
);

INVx5_ASAP7_75t_L g7931 ( 
.A(n_7601),
.Y(n_7931)
);

NOR2xp67_ASAP7_75t_L g7932 ( 
.A(n_7728),
.B(n_7353),
.Y(n_7932)
);

BUFx2_ASAP7_75t_L g7933 ( 
.A(n_7619),
.Y(n_7933)
);

OAI21xp5_ASAP7_75t_L g7934 ( 
.A1(n_7648),
.A2(n_7284),
.B(n_7283),
.Y(n_7934)
);

INVx1_ASAP7_75t_L g7935 ( 
.A(n_7541),
.Y(n_7935)
);

OAI21xp5_ASAP7_75t_L g7936 ( 
.A1(n_7776),
.A2(n_7294),
.B(n_7331),
.Y(n_7936)
);

OAI21xp5_ASAP7_75t_L g7937 ( 
.A1(n_7806),
.A2(n_7293),
.B(n_7359),
.Y(n_7937)
);

O2A1O1Ixp33_ASAP7_75t_SL g7938 ( 
.A1(n_7654),
.A2(n_7463),
.B(n_7517),
.C(n_7460),
.Y(n_7938)
);

NAND2xp5_ASAP7_75t_L g7939 ( 
.A(n_7639),
.B(n_7813),
.Y(n_7939)
);

O2A1O1Ixp33_ASAP7_75t_L g7940 ( 
.A1(n_7822),
.A2(n_7300),
.B(n_7336),
.C(n_7263),
.Y(n_7940)
);

INVx1_ASAP7_75t_L g7941 ( 
.A(n_7543),
.Y(n_7941)
);

AO32x2_ASAP7_75t_L g7942 ( 
.A1(n_7898),
.A2(n_7291),
.A3(n_7369),
.B1(n_7344),
.B2(n_7433),
.Y(n_7942)
);

INVx8_ASAP7_75t_L g7943 ( 
.A(n_7626),
.Y(n_7943)
);

NAND2xp5_ASAP7_75t_L g7944 ( 
.A(n_7566),
.B(n_7435),
.Y(n_7944)
);

A2O1A1Ixp33_ASAP7_75t_L g7945 ( 
.A1(n_7605),
.A2(n_7528),
.B(n_7494),
.C(n_7510),
.Y(n_7945)
);

INVx1_ASAP7_75t_L g7946 ( 
.A(n_7544),
.Y(n_7946)
);

INVx1_ASAP7_75t_L g7947 ( 
.A(n_7556),
.Y(n_7947)
);

NAND2xp5_ASAP7_75t_L g7948 ( 
.A(n_7551),
.B(n_7438),
.Y(n_7948)
);

AND2x2_ASAP7_75t_L g7949 ( 
.A(n_7796),
.B(n_7367),
.Y(n_7949)
);

AO31x2_ASAP7_75t_L g7950 ( 
.A1(n_7779),
.A2(n_7452),
.A3(n_7439),
.B(n_229),
.Y(n_7950)
);

OAI21x1_ASAP7_75t_L g7951 ( 
.A1(n_7711),
.A2(n_227),
.B(n_228),
.Y(n_7951)
);

INVx1_ASAP7_75t_L g7952 ( 
.A(n_7557),
.Y(n_7952)
);

AOI21xp5_ASAP7_75t_L g7953 ( 
.A1(n_7699),
.A2(n_227),
.B(n_228),
.Y(n_7953)
);

AO31x2_ASAP7_75t_L g7954 ( 
.A1(n_7755),
.A2(n_231),
.A3(n_229),
.B(n_230),
.Y(n_7954)
);

OAI21xp5_ASAP7_75t_L g7955 ( 
.A1(n_7722),
.A2(n_229),
.B(n_230),
.Y(n_7955)
);

OAI21xp5_ASAP7_75t_L g7956 ( 
.A1(n_7665),
.A2(n_230),
.B(n_231),
.Y(n_7956)
);

AOI22xp33_ASAP7_75t_L g7957 ( 
.A1(n_7608),
.A2(n_233),
.B1(n_231),
.B2(n_232),
.Y(n_7957)
);

OAI21xp33_ASAP7_75t_SL g7958 ( 
.A1(n_7907),
.A2(n_1337),
.B(n_1336),
.Y(n_7958)
);

INVx1_ASAP7_75t_L g7959 ( 
.A(n_7561),
.Y(n_7959)
);

BUFx2_ASAP7_75t_L g7960 ( 
.A(n_7703),
.Y(n_7960)
);

A2O1A1Ixp33_ASAP7_75t_L g7961 ( 
.A1(n_7759),
.A2(n_1338),
.B(n_1340),
.C(n_1337),
.Y(n_7961)
);

OR2x2_ASAP7_75t_L g7962 ( 
.A(n_7614),
.B(n_1341),
.Y(n_7962)
);

A2O1A1Ixp33_ASAP7_75t_L g7963 ( 
.A1(n_7804),
.A2(n_1342),
.B(n_1343),
.C(n_1341),
.Y(n_7963)
);

INVx1_ASAP7_75t_L g7964 ( 
.A(n_7576),
.Y(n_7964)
);

AOI22xp33_ASAP7_75t_L g7965 ( 
.A1(n_7877),
.A2(n_234),
.B1(n_232),
.B2(n_233),
.Y(n_7965)
);

NAND2x1p5_ASAP7_75t_L g7966 ( 
.A(n_7606),
.B(n_1343),
.Y(n_7966)
);

AOI21xp5_ASAP7_75t_L g7967 ( 
.A1(n_7540),
.A2(n_232),
.B(n_233),
.Y(n_7967)
);

HB1xp67_ASAP7_75t_L g7968 ( 
.A(n_7749),
.Y(n_7968)
);

AOI21x1_ASAP7_75t_L g7969 ( 
.A1(n_7604),
.A2(n_234),
.B(n_235),
.Y(n_7969)
);

O2A1O1Ixp33_ASAP7_75t_SL g7970 ( 
.A1(n_7851),
.A2(n_237),
.B(n_235),
.C(n_236),
.Y(n_7970)
);

A2O1A1Ixp33_ASAP7_75t_L g7971 ( 
.A1(n_7763),
.A2(n_1345),
.B(n_1346),
.C(n_1344),
.Y(n_7971)
);

CKINVDCx6p67_ASAP7_75t_R g7972 ( 
.A(n_7672),
.Y(n_7972)
);

NAND2xp5_ASAP7_75t_SL g7973 ( 
.A(n_7638),
.B(n_1346),
.Y(n_7973)
);

OAI21xp5_ASAP7_75t_L g7974 ( 
.A1(n_7845),
.A2(n_236),
.B(n_237),
.Y(n_7974)
);

INVx2_ASAP7_75t_L g7975 ( 
.A(n_7590),
.Y(n_7975)
);

O2A1O1Ixp33_ASAP7_75t_L g7976 ( 
.A1(n_7706),
.A2(n_7598),
.B(n_7801),
.C(n_7669),
.Y(n_7976)
);

AO32x2_ASAP7_75t_L g7977 ( 
.A1(n_7577),
.A2(n_7617),
.A3(n_7859),
.B1(n_7694),
.B2(n_7893),
.Y(n_7977)
);

INVx2_ASAP7_75t_L g7978 ( 
.A(n_7768),
.Y(n_7978)
);

OAI22xp5_ASAP7_75t_L g7979 ( 
.A1(n_7539),
.A2(n_239),
.B1(n_236),
.B2(n_238),
.Y(n_7979)
);

NAND2xp33_ASAP7_75t_SL g7980 ( 
.A(n_7797),
.B(n_1348),
.Y(n_7980)
);

INVx1_ASAP7_75t_SL g7981 ( 
.A(n_7565),
.Y(n_7981)
);

BUFx12f_ASAP7_75t_L g7982 ( 
.A(n_7675),
.Y(n_7982)
);

NAND2xp5_ASAP7_75t_SL g7983 ( 
.A(n_7892),
.B(n_1348),
.Y(n_7983)
);

AOI221x1_ASAP7_75t_L g7984 ( 
.A1(n_7881),
.A2(n_240),
.B1(n_238),
.B2(n_239),
.C(n_241),
.Y(n_7984)
);

OR2x2_ASAP7_75t_L g7985 ( 
.A(n_7555),
.B(n_1349),
.Y(n_7985)
);

INVx1_ASAP7_75t_L g7986 ( 
.A(n_7581),
.Y(n_7986)
);

BUFx10_ASAP7_75t_L g7987 ( 
.A(n_7611),
.Y(n_7987)
);

INVx3_ASAP7_75t_L g7988 ( 
.A(n_7574),
.Y(n_7988)
);

INVx4_ASAP7_75t_SL g7989 ( 
.A(n_7573),
.Y(n_7989)
);

INVx1_ASAP7_75t_L g7990 ( 
.A(n_7587),
.Y(n_7990)
);

A2O1A1Ixp33_ASAP7_75t_L g7991 ( 
.A1(n_7597),
.A2(n_1350),
.B(n_1352),
.C(n_1349),
.Y(n_7991)
);

INVx1_ASAP7_75t_L g7992 ( 
.A(n_7593),
.Y(n_7992)
);

INVx4_ASAP7_75t_L g7993 ( 
.A(n_7611),
.Y(n_7993)
);

INVx1_ASAP7_75t_L g7994 ( 
.A(n_7616),
.Y(n_7994)
);

A2O1A1Ixp33_ASAP7_75t_L g7995 ( 
.A1(n_7808),
.A2(n_1354),
.B(n_1355),
.C(n_1350),
.Y(n_7995)
);

OAI21xp5_ASAP7_75t_L g7996 ( 
.A1(n_7661),
.A2(n_239),
.B(n_240),
.Y(n_7996)
);

A2O1A1Ixp33_ASAP7_75t_L g7997 ( 
.A1(n_7802),
.A2(n_1358),
.B(n_1359),
.C(n_1356),
.Y(n_7997)
);

AOI221x1_ASAP7_75t_L g7998 ( 
.A1(n_7855),
.A2(n_243),
.B1(n_241),
.B2(n_242),
.C(n_244),
.Y(n_7998)
);

NOR2xp33_ASAP7_75t_L g7999 ( 
.A(n_7837),
.B(n_1356),
.Y(n_7999)
);

O2A1O1Ixp33_ASAP7_75t_L g8000 ( 
.A1(n_7671),
.A2(n_243),
.B(n_241),
.C(n_242),
.Y(n_8000)
);

AO31x2_ASAP7_75t_L g8001 ( 
.A1(n_7883),
.A2(n_7702),
.A3(n_7769),
.B(n_7887),
.Y(n_8001)
);

NAND2xp5_ASAP7_75t_L g8002 ( 
.A(n_7647),
.B(n_1358),
.Y(n_8002)
);

OAI22xp5_ASAP7_75t_L g8003 ( 
.A1(n_7723),
.A2(n_245),
.B1(n_243),
.B2(n_244),
.Y(n_8003)
);

INVx1_ASAP7_75t_L g8004 ( 
.A(n_7624),
.Y(n_8004)
);

INVx1_ASAP7_75t_L g8005 ( 
.A(n_7629),
.Y(n_8005)
);

O2A1O1Ixp33_ASAP7_75t_SL g8006 ( 
.A1(n_7716),
.A2(n_246),
.B(n_244),
.C(n_245),
.Y(n_8006)
);

A2O1A1Ixp33_ASAP7_75t_L g8007 ( 
.A1(n_7913),
.A2(n_1360),
.B(n_1361),
.C(n_1359),
.Y(n_8007)
);

AO31x2_ASAP7_75t_L g8008 ( 
.A1(n_7735),
.A2(n_248),
.A3(n_245),
.B(n_247),
.Y(n_8008)
);

AOI221x1_ASAP7_75t_L g8009 ( 
.A1(n_7828),
.A2(n_249),
.B1(n_247),
.B2(n_248),
.C(n_250),
.Y(n_8009)
);

AND2x2_ASAP7_75t_L g8010 ( 
.A(n_7750),
.B(n_1360),
.Y(n_8010)
);

INVx1_ASAP7_75t_L g8011 ( 
.A(n_7630),
.Y(n_8011)
);

A2O1A1Ixp33_ASAP7_75t_L g8012 ( 
.A1(n_7917),
.A2(n_1362),
.B(n_1363),
.C(n_1361),
.Y(n_8012)
);

AOI21xp5_ASAP7_75t_L g8013 ( 
.A1(n_7615),
.A2(n_7680),
.B(n_7733),
.Y(n_8013)
);

O2A1O1Ixp33_ASAP7_75t_SL g8014 ( 
.A1(n_7847),
.A2(n_249),
.B(n_247),
.C(n_248),
.Y(n_8014)
);

AO32x2_ASAP7_75t_L g8015 ( 
.A1(n_7914),
.A2(n_251),
.A3(n_249),
.B1(n_250),
.B2(n_252),
.Y(n_8015)
);

INVx1_ASAP7_75t_L g8016 ( 
.A(n_7636),
.Y(n_8016)
);

NAND2xp5_ASAP7_75t_L g8017 ( 
.A(n_7872),
.B(n_1362),
.Y(n_8017)
);

NAND2xp5_ASAP7_75t_L g8018 ( 
.A(n_7618),
.B(n_1364),
.Y(n_8018)
);

INVx1_ASAP7_75t_L g8019 ( 
.A(n_7642),
.Y(n_8019)
);

BUFx2_ASAP7_75t_L g8020 ( 
.A(n_7705),
.Y(n_8020)
);

OAI22x1_ASAP7_75t_L g8021 ( 
.A1(n_7663),
.A2(n_7854),
.B1(n_7873),
.B2(n_7830),
.Y(n_8021)
);

AOI22xp33_ASAP7_75t_L g8022 ( 
.A1(n_7877),
.A2(n_252),
.B1(n_250),
.B2(n_251),
.Y(n_8022)
);

BUFx10_ASAP7_75t_L g8023 ( 
.A(n_7538),
.Y(n_8023)
);

INVx1_ASAP7_75t_L g8024 ( 
.A(n_7662),
.Y(n_8024)
);

AOI21xp5_ASAP7_75t_L g8025 ( 
.A1(n_7741),
.A2(n_253),
.B(n_254),
.Y(n_8025)
);

OR2x2_ASAP7_75t_L g8026 ( 
.A(n_7621),
.B(n_1364),
.Y(n_8026)
);

O2A1O1Ixp33_ASAP7_75t_SL g8027 ( 
.A1(n_7547),
.A2(n_7890),
.B(n_7906),
.C(n_7885),
.Y(n_8027)
);

OAI22x1_ASAP7_75t_L g8028 ( 
.A1(n_7825),
.A2(n_255),
.B1(n_253),
.B2(n_254),
.Y(n_8028)
);

AOI22xp5_ASAP7_75t_L g8029 ( 
.A1(n_7877),
.A2(n_255),
.B1(n_253),
.B2(n_254),
.Y(n_8029)
);

AO31x2_ASAP7_75t_L g8030 ( 
.A1(n_7884),
.A2(n_257),
.A3(n_255),
.B(n_256),
.Y(n_8030)
);

AOI21xp5_ASAP7_75t_L g8031 ( 
.A1(n_7785),
.A2(n_256),
.B(n_257),
.Y(n_8031)
);

NAND2xp5_ASAP7_75t_L g8032 ( 
.A(n_7820),
.B(n_1365),
.Y(n_8032)
);

INVx3_ASAP7_75t_L g8033 ( 
.A(n_7574),
.Y(n_8033)
);

AOI21xp5_ASAP7_75t_L g8034 ( 
.A1(n_7734),
.A2(n_258),
.B(n_259),
.Y(n_8034)
);

AOI22xp33_ASAP7_75t_SL g8035 ( 
.A1(n_7637),
.A2(n_260),
.B1(n_258),
.B2(n_259),
.Y(n_8035)
);

CKINVDCx20_ASAP7_75t_R g8036 ( 
.A(n_7778),
.Y(n_8036)
);

NOR2xp33_ASAP7_75t_SL g8037 ( 
.A(n_7586),
.B(n_258),
.Y(n_8037)
);

BUFx8_ASAP7_75t_SL g8038 ( 
.A(n_7589),
.Y(n_8038)
);

O2A1O1Ixp33_ASAP7_75t_L g8039 ( 
.A1(n_7773),
.A2(n_7789),
.B(n_7817),
.C(n_7815),
.Y(n_8039)
);

NOR2xp67_ASAP7_75t_SL g8040 ( 
.A(n_7672),
.B(n_260),
.Y(n_8040)
);

AOI21xp5_ASAP7_75t_L g8041 ( 
.A1(n_7910),
.A2(n_261),
.B(n_262),
.Y(n_8041)
);

O2A1O1Ixp33_ASAP7_75t_SL g8042 ( 
.A1(n_7748),
.A2(n_7878),
.B(n_7879),
.C(n_7651),
.Y(n_8042)
);

INVx5_ASAP7_75t_L g8043 ( 
.A(n_7538),
.Y(n_8043)
);

INVxp67_ASAP7_75t_L g8044 ( 
.A(n_7730),
.Y(n_8044)
);

INVx1_ASAP7_75t_L g8045 ( 
.A(n_7666),
.Y(n_8045)
);

INVx2_ASAP7_75t_L g8046 ( 
.A(n_7767),
.Y(n_8046)
);

AOI21xp33_ASAP7_75t_L g8047 ( 
.A1(n_7549),
.A2(n_261),
.B(n_262),
.Y(n_8047)
);

INVx3_ASAP7_75t_SL g8048 ( 
.A(n_7607),
.Y(n_8048)
);

AOI222xp33_ASAP7_75t_L g8049 ( 
.A1(n_7553),
.A2(n_264),
.B1(n_267),
.B2(n_262),
.C1(n_263),
.C2(n_266),
.Y(n_8049)
);

NOR2xp33_ASAP7_75t_L g8050 ( 
.A(n_7902),
.B(n_1365),
.Y(n_8050)
);

AOI22xp5_ASAP7_75t_L g8051 ( 
.A1(n_7805),
.A2(n_266),
.B1(n_263),
.B2(n_264),
.Y(n_8051)
);

NAND2xp5_ASAP7_75t_L g8052 ( 
.A(n_7821),
.B(n_7812),
.Y(n_8052)
);

INVx1_ASAP7_75t_L g8053 ( 
.A(n_7683),
.Y(n_8053)
);

INVx3_ASAP7_75t_L g8054 ( 
.A(n_7578),
.Y(n_8054)
);

AOI21xp5_ASAP7_75t_L g8055 ( 
.A1(n_7876),
.A2(n_266),
.B(n_267),
.Y(n_8055)
);

INVx1_ASAP7_75t_L g8056 ( 
.A(n_7698),
.Y(n_8056)
);

AND2x2_ASAP7_75t_L g8057 ( 
.A(n_7762),
.B(n_1366),
.Y(n_8057)
);

INVx1_ASAP7_75t_L g8058 ( 
.A(n_7700),
.Y(n_8058)
);

NAND2xp5_ASAP7_75t_L g8059 ( 
.A(n_7860),
.B(n_1368),
.Y(n_8059)
);

OAI21xp5_ASAP7_75t_L g8060 ( 
.A1(n_7897),
.A2(n_7899),
.B(n_7846),
.Y(n_8060)
);

OAI22xp33_ASAP7_75t_L g8061 ( 
.A1(n_7664),
.A2(n_269),
.B1(n_267),
.B2(n_268),
.Y(n_8061)
);

INVx1_ASAP7_75t_L g8062 ( 
.A(n_7707),
.Y(n_8062)
);

OA21x2_ASAP7_75t_L g8063 ( 
.A1(n_7563),
.A2(n_268),
.B(n_269),
.Y(n_8063)
);

AOI21xp5_ASAP7_75t_L g8064 ( 
.A1(n_7784),
.A2(n_269),
.B(n_270),
.Y(n_8064)
);

AOI22xp33_ASAP7_75t_L g8065 ( 
.A1(n_7861),
.A2(n_272),
.B1(n_270),
.B2(n_271),
.Y(n_8065)
);

AOI21xp5_ASAP7_75t_L g8066 ( 
.A1(n_7852),
.A2(n_7826),
.B(n_7818),
.Y(n_8066)
);

NAND2xp5_ASAP7_75t_L g8067 ( 
.A(n_7866),
.B(n_1368),
.Y(n_8067)
);

AO21x1_ASAP7_75t_L g8068 ( 
.A1(n_7880),
.A2(n_270),
.B(n_271),
.Y(n_8068)
);

INVx2_ASAP7_75t_SL g8069 ( 
.A(n_7625),
.Y(n_8069)
);

NAND2xp5_ASAP7_75t_L g8070 ( 
.A(n_7678),
.B(n_1369),
.Y(n_8070)
);

NAND2xp5_ASAP7_75t_L g8071 ( 
.A(n_7693),
.B(n_1369),
.Y(n_8071)
);

INVx1_ASAP7_75t_L g8072 ( 
.A(n_7726),
.Y(n_8072)
);

INVx2_ASAP7_75t_L g8073 ( 
.A(n_7727),
.Y(n_8073)
);

O2A1O1Ixp33_ASAP7_75t_L g8074 ( 
.A1(n_7833),
.A2(n_274),
.B(n_272),
.C(n_273),
.Y(n_8074)
);

BUFx10_ASAP7_75t_L g8075 ( 
.A(n_7717),
.Y(n_8075)
);

OAI21xp5_ASAP7_75t_L g8076 ( 
.A1(n_7782),
.A2(n_273),
.B(n_274),
.Y(n_8076)
);

INVx1_ASAP7_75t_SL g8077 ( 
.A(n_7684),
.Y(n_8077)
);

A2O1A1Ixp33_ASAP7_75t_L g8078 ( 
.A1(n_7602),
.A2(n_1371),
.B(n_1372),
.C(n_1370),
.Y(n_8078)
);

AOI21xp33_ASAP7_75t_L g8079 ( 
.A1(n_7600),
.A2(n_273),
.B(n_274),
.Y(n_8079)
);

OR2x6_ASAP7_75t_L g8080 ( 
.A(n_7920),
.B(n_1370),
.Y(n_8080)
);

INVx2_ASAP7_75t_L g8081 ( 
.A(n_7732),
.Y(n_8081)
);

INVx1_ASAP7_75t_L g8082 ( 
.A(n_7701),
.Y(n_8082)
);

AOI22xp33_ASAP7_75t_L g8083 ( 
.A1(n_7900),
.A2(n_277),
.B1(n_275),
.B2(n_276),
.Y(n_8083)
);

INVx1_ASAP7_75t_L g8084 ( 
.A(n_7757),
.Y(n_8084)
);

INVx1_ASAP7_75t_L g8085 ( 
.A(n_7738),
.Y(n_8085)
);

INVx1_ASAP7_75t_L g8086 ( 
.A(n_7760),
.Y(n_8086)
);

AOI222xp33_ASAP7_75t_L g8087 ( 
.A1(n_7692),
.A2(n_278),
.B1(n_280),
.B2(n_276),
.C1(n_277),
.C2(n_279),
.Y(n_8087)
);

HB1xp67_ASAP7_75t_L g8088 ( 
.A(n_7610),
.Y(n_8088)
);

NAND2xp5_ASAP7_75t_L g8089 ( 
.A(n_7633),
.B(n_1372),
.Y(n_8089)
);

INVx1_ASAP7_75t_L g8090 ( 
.A(n_7761),
.Y(n_8090)
);

OAI21xp5_ASAP7_75t_L g8091 ( 
.A1(n_7620),
.A2(n_277),
.B(n_278),
.Y(n_8091)
);

NAND2xp5_ASAP7_75t_L g8092 ( 
.A(n_7874),
.B(n_1373),
.Y(n_8092)
);

O2A1O1Ixp33_ASAP7_75t_L g8093 ( 
.A1(n_7643),
.A2(n_280),
.B(n_278),
.C(n_279),
.Y(n_8093)
);

AOI21xp5_ASAP7_75t_L g8094 ( 
.A1(n_7827),
.A2(n_279),
.B(n_280),
.Y(n_8094)
);

AOI21xp5_ASAP7_75t_L g8095 ( 
.A1(n_7829),
.A2(n_281),
.B(n_282),
.Y(n_8095)
);

NAND2xp5_ASAP7_75t_L g8096 ( 
.A(n_7835),
.B(n_1374),
.Y(n_8096)
);

INVx1_ASAP7_75t_L g8097 ( 
.A(n_7537),
.Y(n_8097)
);

NOR2xp33_ASAP7_75t_L g8098 ( 
.A(n_7811),
.B(n_1375),
.Y(n_8098)
);

NAND2x1p5_ASAP7_75t_L g8099 ( 
.A(n_7670),
.B(n_1375),
.Y(n_8099)
);

OAI21x1_ASAP7_75t_L g8100 ( 
.A1(n_7790),
.A2(n_281),
.B(n_282),
.Y(n_8100)
);

AOI21xp5_ASAP7_75t_L g8101 ( 
.A1(n_7840),
.A2(n_281),
.B(n_282),
.Y(n_8101)
);

INVx2_ASAP7_75t_L g8102 ( 
.A(n_7550),
.Y(n_8102)
);

INVx3_ASAP7_75t_L g8103 ( 
.A(n_7578),
.Y(n_8103)
);

INVx2_ASAP7_75t_L g8104 ( 
.A(n_7569),
.Y(n_8104)
);

AOI21xp5_ASAP7_75t_L g8105 ( 
.A1(n_7656),
.A2(n_283),
.B(n_284),
.Y(n_8105)
);

OAI21xp5_ASAP7_75t_L g8106 ( 
.A1(n_7838),
.A2(n_283),
.B(n_284),
.Y(n_8106)
);

NAND2xp5_ASAP7_75t_SL g8107 ( 
.A(n_7892),
.B(n_1376),
.Y(n_8107)
);

BUFx12f_ASAP7_75t_L g8108 ( 
.A(n_7596),
.Y(n_8108)
);

INVx2_ASAP7_75t_L g8109 ( 
.A(n_7570),
.Y(n_8109)
);

OAI211xp5_ASAP7_75t_SL g8110 ( 
.A1(n_7791),
.A2(n_286),
.B(n_284),
.C(n_285),
.Y(n_8110)
);

OAI22xp5_ASAP7_75t_L g8111 ( 
.A1(n_7916),
.A2(n_287),
.B1(n_285),
.B2(n_286),
.Y(n_8111)
);

NAND2xp5_ASAP7_75t_L g8112 ( 
.A(n_7843),
.B(n_1376),
.Y(n_8112)
);

A2O1A1Ixp33_ASAP7_75t_L g8113 ( 
.A1(n_7831),
.A2(n_1378),
.B(n_1379),
.C(n_1377),
.Y(n_8113)
);

AO31x2_ASAP7_75t_L g8114 ( 
.A1(n_7889),
.A2(n_287),
.A3(n_285),
.B(n_286),
.Y(n_8114)
);

AO31x2_ASAP7_75t_L g8115 ( 
.A1(n_7903),
.A2(n_289),
.A3(n_287),
.B(n_288),
.Y(n_8115)
);

A2O1A1Ixp33_ASAP7_75t_L g8116 ( 
.A1(n_7839),
.A2(n_1379),
.B(n_1380),
.C(n_1377),
.Y(n_8116)
);

AOI22xp33_ASAP7_75t_L g8117 ( 
.A1(n_7908),
.A2(n_290),
.B1(n_288),
.B2(n_289),
.Y(n_8117)
);

A2O1A1Ixp33_ASAP7_75t_L g8118 ( 
.A1(n_7841),
.A2(n_1382),
.B(n_1384),
.C(n_1381),
.Y(n_8118)
);

AND2x2_ASAP7_75t_L g8119 ( 
.A(n_7798),
.B(n_1381),
.Y(n_8119)
);

CKINVDCx5p33_ASAP7_75t_R g8120 ( 
.A(n_7775),
.Y(n_8120)
);

BUFx3_ASAP7_75t_L g8121 ( 
.A(n_7632),
.Y(n_8121)
);

NAND2xp5_ASAP7_75t_L g8122 ( 
.A(n_7867),
.B(n_1384),
.Y(n_8122)
);

NOR2xp33_ASAP7_75t_L g8123 ( 
.A(n_7882),
.B(n_1387),
.Y(n_8123)
);

A2O1A1Ixp33_ASAP7_75t_L g8124 ( 
.A1(n_7753),
.A2(n_1389),
.B(n_1390),
.C(n_1388),
.Y(n_8124)
);

CKINVDCx11_ASAP7_75t_R g8125 ( 
.A(n_7751),
.Y(n_8125)
);

INVx1_ASAP7_75t_L g8126 ( 
.A(n_7580),
.Y(n_8126)
);

OAI21xp5_ASAP7_75t_L g8127 ( 
.A1(n_7795),
.A2(n_288),
.B(n_290),
.Y(n_8127)
);

AO32x2_ASAP7_75t_L g8128 ( 
.A1(n_7667),
.A2(n_293),
.A3(n_291),
.B1(n_292),
.B2(n_294),
.Y(n_8128)
);

NOR2xp33_ASAP7_75t_L g8129 ( 
.A(n_7783),
.B(n_1388),
.Y(n_8129)
);

A2O1A1Ixp33_ASAP7_75t_L g8130 ( 
.A1(n_7844),
.A2(n_1390),
.B(n_1392),
.C(n_1389),
.Y(n_8130)
);

AOI22xp33_ASAP7_75t_SL g8131 ( 
.A1(n_7862),
.A2(n_293),
.B1(n_291),
.B2(n_292),
.Y(n_8131)
);

OAI22xp33_ASAP7_75t_L g8132 ( 
.A1(n_7794),
.A2(n_7676),
.B1(n_7718),
.B2(n_7901),
.Y(n_8132)
);

O2A1O1Ixp33_ASAP7_75t_L g8133 ( 
.A1(n_7909),
.A2(n_296),
.B(n_292),
.C(n_295),
.Y(n_8133)
);

OAI21xp5_ASAP7_75t_L g8134 ( 
.A1(n_7857),
.A2(n_296),
.B(n_297),
.Y(n_8134)
);

INVx2_ASAP7_75t_L g8135 ( 
.A(n_7585),
.Y(n_8135)
);

NOR2xp33_ASAP7_75t_L g8136 ( 
.A(n_7673),
.B(n_1393),
.Y(n_8136)
);

A2O1A1Ixp33_ASAP7_75t_L g8137 ( 
.A1(n_7824),
.A2(n_7686),
.B(n_7758),
.C(n_7819),
.Y(n_8137)
);

INVx2_ASAP7_75t_L g8138 ( 
.A(n_7640),
.Y(n_8138)
);

NOR2xp33_ASAP7_75t_L g8139 ( 
.A(n_7863),
.B(n_1393),
.Y(n_8139)
);

INVx1_ASAP7_75t_L g8140 ( 
.A(n_7641),
.Y(n_8140)
);

NAND2xp5_ASAP7_75t_L g8141 ( 
.A(n_7868),
.B(n_1394),
.Y(n_8141)
);

INVx2_ASAP7_75t_L g8142 ( 
.A(n_7644),
.Y(n_8142)
);

INVx1_ASAP7_75t_L g8143 ( 
.A(n_7658),
.Y(n_8143)
);

O2A1O1Ixp33_ASAP7_75t_L g8144 ( 
.A1(n_7792),
.A2(n_299),
.B(n_297),
.C(n_298),
.Y(n_8144)
);

INVx2_ASAP7_75t_L g8145 ( 
.A(n_7668),
.Y(n_8145)
);

INVx1_ASAP7_75t_SL g8146 ( 
.A(n_7690),
.Y(n_8146)
);

AOI22xp5_ASAP7_75t_L g8147 ( 
.A1(n_7850),
.A2(n_299),
.B1(n_297),
.B2(n_298),
.Y(n_8147)
);

A2O1A1Ixp33_ASAP7_75t_L g8148 ( 
.A1(n_7856),
.A2(n_1395),
.B(n_1396),
.C(n_1394),
.Y(n_8148)
);

CKINVDCx9p33_ASAP7_75t_R g8149 ( 
.A(n_7814),
.Y(n_8149)
);

BUFx6f_ASAP7_75t_L g8150 ( 
.A(n_7632),
.Y(n_8150)
);

AOI21xp5_ASAP7_75t_L g8151 ( 
.A1(n_7558),
.A2(n_298),
.B(n_300),
.Y(n_8151)
);

BUFx6f_ASAP7_75t_L g8152 ( 
.A(n_7634),
.Y(n_8152)
);

INVx2_ASAP7_75t_L g8153 ( 
.A(n_7691),
.Y(n_8153)
);

NOR2xp33_ASAP7_75t_L g8154 ( 
.A(n_7912),
.B(n_1396),
.Y(n_8154)
);

AND2x2_ASAP7_75t_L g8155 ( 
.A(n_7888),
.B(n_1397),
.Y(n_8155)
);

A2O1A1Ixp33_ASAP7_75t_L g8156 ( 
.A1(n_7918),
.A2(n_1398),
.B(n_1399),
.C(n_1397),
.Y(n_8156)
);

OAI21xp5_ASAP7_75t_L g8157 ( 
.A1(n_7871),
.A2(n_300),
.B(n_301),
.Y(n_8157)
);

AO31x2_ASAP7_75t_L g8158 ( 
.A1(n_7712),
.A2(n_303),
.A3(n_300),
.B(n_302),
.Y(n_8158)
);

OR2x2_ASAP7_75t_L g8159 ( 
.A(n_7765),
.B(n_1399),
.Y(n_8159)
);

HB1xp67_ASAP7_75t_L g8160 ( 
.A(n_7627),
.Y(n_8160)
);

O2A1O1Ixp33_ASAP7_75t_SL g8161 ( 
.A1(n_7915),
.A2(n_305),
.B(n_303),
.C(n_304),
.Y(n_8161)
);

INVx8_ASAP7_75t_L g8162 ( 
.A(n_7625),
.Y(n_8162)
);

BUFx6f_ASAP7_75t_L g8163 ( 
.A(n_7634),
.Y(n_8163)
);

AOI21xp5_ASAP7_75t_L g8164 ( 
.A1(n_7584),
.A2(n_303),
.B(n_304),
.Y(n_8164)
);

INVx2_ASAP7_75t_SL g8165 ( 
.A(n_7681),
.Y(n_8165)
);

NAND2xp5_ASAP7_75t_L g8166 ( 
.A(n_7635),
.B(n_1400),
.Y(n_8166)
);

INVx1_ASAP7_75t_SL g8167 ( 
.A(n_7725),
.Y(n_8167)
);

AOI22xp5_ASAP7_75t_L g8168 ( 
.A1(n_7904),
.A2(n_306),
.B1(n_304),
.B2(n_305),
.Y(n_8168)
);

BUFx3_ASAP7_75t_L g8169 ( 
.A(n_7542),
.Y(n_8169)
);

AO32x2_ASAP7_75t_L g8170 ( 
.A1(n_7568),
.A2(n_307),
.A3(n_305),
.B1(n_306),
.B2(n_308),
.Y(n_8170)
);

OAI21x1_ASAP7_75t_L g8171 ( 
.A1(n_7697),
.A2(n_306),
.B(n_307),
.Y(n_8171)
);

AOI21xp5_ASAP7_75t_L g8172 ( 
.A1(n_7745),
.A2(n_7754),
.B(n_7919),
.Y(n_8172)
);

O2A1O1Ixp33_ASAP7_75t_L g8173 ( 
.A1(n_7793),
.A2(n_311),
.B(n_309),
.C(n_310),
.Y(n_8173)
);

A2O1A1Ixp33_ASAP7_75t_L g8174 ( 
.A1(n_7781),
.A2(n_1401),
.B(n_1402),
.C(n_1400),
.Y(n_8174)
);

A2O1A1Ixp33_ASAP7_75t_L g8175 ( 
.A1(n_7911),
.A2(n_1403),
.B(n_1404),
.C(n_1401),
.Y(n_8175)
);

INVx1_ASAP7_75t_L g8176 ( 
.A(n_7713),
.Y(n_8176)
);

HB1xp67_ASAP7_75t_L g8177 ( 
.A(n_7740),
.Y(n_8177)
);

AO21x1_ASAP7_75t_L g8178 ( 
.A1(n_7803),
.A2(n_309),
.B(n_310),
.Y(n_8178)
);

AOI22xp33_ASAP7_75t_L g8179 ( 
.A1(n_7904),
.A2(n_312),
.B1(n_309),
.B2(n_311),
.Y(n_8179)
);

BUFx2_ASAP7_75t_L g8180 ( 
.A(n_7842),
.Y(n_8180)
);

BUFx2_ASAP7_75t_L g8181 ( 
.A(n_7842),
.Y(n_8181)
);

INVx2_ASAP7_75t_L g8182 ( 
.A(n_7747),
.Y(n_8182)
);

INVx1_ASAP7_75t_L g8183 ( 
.A(n_7613),
.Y(n_8183)
);

NAND2xp5_ASAP7_75t_L g8184 ( 
.A(n_7891),
.B(n_1404),
.Y(n_8184)
);

A2O1A1Ixp33_ASAP7_75t_L g8185 ( 
.A1(n_7810),
.A2(n_7834),
.B(n_7849),
.C(n_7832),
.Y(n_8185)
);

BUFx12f_ASAP7_75t_L g8186 ( 
.A(n_7653),
.Y(n_8186)
);

AO21x1_ASAP7_75t_L g8187 ( 
.A1(n_7865),
.A2(n_311),
.B(n_312),
.Y(n_8187)
);

INVx1_ASAP7_75t_L g8188 ( 
.A(n_7800),
.Y(n_8188)
);

AOI22xp33_ASAP7_75t_L g8189 ( 
.A1(n_7894),
.A2(n_314),
.B1(n_312),
.B2(n_313),
.Y(n_8189)
);

INVx2_ASAP7_75t_L g8190 ( 
.A(n_7836),
.Y(n_8190)
);

OAI22xp5_ASAP7_75t_L g8191 ( 
.A1(n_7704),
.A2(n_315),
.B1(n_313),
.B2(n_314),
.Y(n_8191)
);

AND2x2_ASAP7_75t_L g8192 ( 
.A(n_7823),
.B(n_1405),
.Y(n_8192)
);

OAI21xp5_ASAP7_75t_SL g8193 ( 
.A1(n_7652),
.A2(n_314),
.B(n_315),
.Y(n_8193)
);

INVxp67_ASAP7_75t_L g8194 ( 
.A(n_7864),
.Y(n_8194)
);

NAND2xp5_ASAP7_75t_L g8195 ( 
.A(n_7875),
.B(n_1405),
.Y(n_8195)
);

OAI21x1_ASAP7_75t_L g8196 ( 
.A1(n_7786),
.A2(n_316),
.B(n_317),
.Y(n_8196)
);

OAI221xp5_ASAP7_75t_L g8197 ( 
.A1(n_7870),
.A2(n_318),
.B1(n_316),
.B2(n_317),
.C(n_319),
.Y(n_8197)
);

NAND3xp33_ASAP7_75t_L g8198 ( 
.A(n_7894),
.B(n_316),
.C(n_317),
.Y(n_8198)
);

AO32x2_ASAP7_75t_L g8199 ( 
.A1(n_7575),
.A2(n_320),
.A3(n_318),
.B1(n_319),
.B2(n_321),
.Y(n_8199)
);

NAND2x1p5_ASAP7_75t_L g8200 ( 
.A(n_7794),
.B(n_1407),
.Y(n_8200)
);

O2A1O1Ixp33_ASAP7_75t_L g8201 ( 
.A1(n_7660),
.A2(n_321),
.B(n_319),
.C(n_320),
.Y(n_8201)
);

AOI21xp5_ASAP7_75t_L g8202 ( 
.A1(n_7895),
.A2(n_320),
.B(n_322),
.Y(n_8202)
);

NAND2xp5_ASAP7_75t_L g8203 ( 
.A(n_7780),
.B(n_1407),
.Y(n_8203)
);

INVxp67_ASAP7_75t_L g8204 ( 
.A(n_7864),
.Y(n_8204)
);

INVx1_ASAP7_75t_L g8205 ( 
.A(n_7848),
.Y(n_8205)
);

INVx1_ASAP7_75t_L g8206 ( 
.A(n_7823),
.Y(n_8206)
);

INVx3_ASAP7_75t_L g8207 ( 
.A(n_7594),
.Y(n_8207)
);

OAI221xp5_ASAP7_75t_SL g8208 ( 
.A1(n_7659),
.A2(n_324),
.B1(n_322),
.B2(n_323),
.C(n_325),
.Y(n_8208)
);

INVx3_ASAP7_75t_L g8209 ( 
.A(n_7594),
.Y(n_8209)
);

HB1xp67_ASAP7_75t_L g8210 ( 
.A(n_7869),
.Y(n_8210)
);

BUFx3_ASAP7_75t_L g8211 ( 
.A(n_7542),
.Y(n_8211)
);

INVx5_ASAP7_75t_L g8212 ( 
.A(n_7645),
.Y(n_8212)
);

NAND2xp5_ASAP7_75t_L g8213 ( 
.A(n_7869),
.B(n_1408),
.Y(n_8213)
);

NAND2xp5_ASAP7_75t_L g8214 ( 
.A(n_7756),
.B(n_1408),
.Y(n_8214)
);

O2A1O1Ixp33_ASAP7_75t_SL g8215 ( 
.A1(n_7687),
.A2(n_324),
.B(n_322),
.C(n_323),
.Y(n_8215)
);

NOR2xp67_ASAP7_75t_SL g8216 ( 
.A(n_7592),
.B(n_323),
.Y(n_8216)
);

AOI21xp5_ASAP7_75t_L g8217 ( 
.A1(n_7603),
.A2(n_325),
.B(n_326),
.Y(n_8217)
);

AO31x2_ASAP7_75t_L g8218 ( 
.A1(n_7719),
.A2(n_327),
.A3(n_325),
.B(n_326),
.Y(n_8218)
);

NOR2xp67_ASAP7_75t_SL g8219 ( 
.A(n_7592),
.B(n_327),
.Y(n_8219)
);

AO32x2_ASAP7_75t_L g8220 ( 
.A1(n_7688),
.A2(n_330),
.A3(n_328),
.B1(n_329),
.B2(n_331),
.Y(n_8220)
);

INVx2_ASAP7_75t_L g8221 ( 
.A(n_7609),
.Y(n_8221)
);

A2O1A1Ixp33_ASAP7_75t_L g8222 ( 
.A1(n_7905),
.A2(n_7787),
.B(n_7816),
.C(n_7646),
.Y(n_8222)
);

O2A1O1Ixp33_ASAP7_75t_SL g8223 ( 
.A1(n_7853),
.A2(n_331),
.B(n_328),
.C(n_329),
.Y(n_8223)
);

OR2x6_ASAP7_75t_L g8224 ( 
.A(n_7623),
.B(n_1409),
.Y(n_8224)
);

NOR2xp33_ASAP7_75t_L g8225 ( 
.A(n_7709),
.B(n_1410),
.Y(n_8225)
);

INVx5_ASAP7_75t_L g8226 ( 
.A(n_7720),
.Y(n_8226)
);

NAND2xp5_ASAP7_75t_SL g8227 ( 
.A(n_7886),
.B(n_1410),
.Y(n_8227)
);

O2A1O1Ixp33_ASAP7_75t_L g8228 ( 
.A1(n_7545),
.A2(n_333),
.B(n_328),
.C(n_332),
.Y(n_8228)
);

INVx1_ASAP7_75t_L g8229 ( 
.A(n_7714),
.Y(n_8229)
);

A2O1A1Ixp33_ASAP7_75t_L g8230 ( 
.A1(n_7772),
.A2(n_1413),
.B(n_1414),
.C(n_1412),
.Y(n_8230)
);

A2O1A1Ixp33_ASAP7_75t_L g8231 ( 
.A1(n_7612),
.A2(n_1414),
.B(n_1415),
.C(n_1413),
.Y(n_8231)
);

INVx2_ASAP7_75t_L g8232 ( 
.A(n_7609),
.Y(n_8232)
);

OAI21xp5_ASAP7_75t_L g8233 ( 
.A1(n_7622),
.A2(n_332),
.B(n_333),
.Y(n_8233)
);

BUFx6f_ASAP7_75t_L g8234 ( 
.A(n_7677),
.Y(n_8234)
);

NOR2xp33_ASAP7_75t_L g8235 ( 
.A(n_7858),
.B(n_1415),
.Y(n_8235)
);

AOI21xp5_ASAP7_75t_L g8236 ( 
.A1(n_7746),
.A2(n_7742),
.B(n_7679),
.Y(n_8236)
);

HB1xp67_ASAP7_75t_L g8237 ( 
.A(n_7968),
.Y(n_8237)
);

INVx1_ASAP7_75t_L g8238 ( 
.A(n_7923),
.Y(n_8238)
);

OAI22xp5_ASAP7_75t_L g8239 ( 
.A1(n_8065),
.A2(n_7788),
.B1(n_7724),
.B2(n_7896),
.Y(n_8239)
);

AND2x4_ASAP7_75t_L g8240 ( 
.A(n_7933),
.B(n_7721),
.Y(n_8240)
);

AOI21xp5_ASAP7_75t_L g8241 ( 
.A1(n_7921),
.A2(n_7695),
.B(n_7743),
.Y(n_8241)
);

INVx2_ASAP7_75t_L g8242 ( 
.A(n_8073),
.Y(n_8242)
);

INVx1_ASAP7_75t_L g8243 ( 
.A(n_7935),
.Y(n_8243)
);

INVx1_ASAP7_75t_L g8244 ( 
.A(n_7941),
.Y(n_8244)
);

INVx1_ASAP7_75t_L g8245 ( 
.A(n_7946),
.Y(n_8245)
);

INVx2_ASAP7_75t_L g8246 ( 
.A(n_8081),
.Y(n_8246)
);

O2A1O1Ixp33_ASAP7_75t_SL g8247 ( 
.A1(n_8227),
.A2(n_7560),
.B(n_7657),
.C(n_7628),
.Y(n_8247)
);

AOI22xp33_ASAP7_75t_SL g8248 ( 
.A1(n_7929),
.A2(n_7955),
.B1(n_7937),
.B2(n_7956),
.Y(n_8248)
);

AOI22xp33_ASAP7_75t_L g8249 ( 
.A1(n_8021),
.A2(n_7729),
.B1(n_7788),
.B2(n_7764),
.Y(n_8249)
);

AND2x2_ASAP7_75t_L g8250 ( 
.A(n_8088),
.B(n_7631),
.Y(n_8250)
);

NAND2x1_ASAP7_75t_L g8251 ( 
.A(n_8082),
.B(n_8084),
.Y(n_8251)
);

AOI22xp33_ASAP7_75t_SL g8252 ( 
.A1(n_7996),
.A2(n_7674),
.B1(n_7736),
.B2(n_7650),
.Y(n_8252)
);

INVx1_ASAP7_75t_L g8253 ( 
.A(n_7947),
.Y(n_8253)
);

HB1xp67_ASAP7_75t_L g8254 ( 
.A(n_8160),
.Y(n_8254)
);

INVx1_ASAP7_75t_SL g8255 ( 
.A(n_8149),
.Y(n_8255)
);

AOI22xp33_ASAP7_75t_L g8256 ( 
.A1(n_8068),
.A2(n_7764),
.B1(n_7731),
.B2(n_7770),
.Y(n_8256)
);

INVx1_ASAP7_75t_L g8257 ( 
.A(n_7952),
.Y(n_8257)
);

BUFx3_ASAP7_75t_L g8258 ( 
.A(n_7982),
.Y(n_8258)
);

AOI22xp33_ASAP7_75t_L g8259 ( 
.A1(n_7922),
.A2(n_7731),
.B1(n_7809),
.B2(n_7777),
.Y(n_8259)
);

OA21x2_ASAP7_75t_L g8260 ( 
.A1(n_8172),
.A2(n_7737),
.B(n_7564),
.Y(n_8260)
);

AND2x2_ASAP7_75t_L g8261 ( 
.A(n_7960),
.B(n_7744),
.Y(n_8261)
);

NAND2xp5_ASAP7_75t_L g8262 ( 
.A(n_7939),
.B(n_7583),
.Y(n_8262)
);

BUFx10_ASAP7_75t_L g8263 ( 
.A(n_8120),
.Y(n_8263)
);

INVx1_ASAP7_75t_L g8264 ( 
.A(n_7959),
.Y(n_8264)
);

INVx1_ASAP7_75t_L g8265 ( 
.A(n_7964),
.Y(n_8265)
);

AOI22xp33_ASAP7_75t_SL g8266 ( 
.A1(n_7958),
.A2(n_7571),
.B1(n_7562),
.B2(n_7591),
.Y(n_8266)
);

AOI22xp33_ASAP7_75t_L g8267 ( 
.A1(n_8197),
.A2(n_7766),
.B1(n_7744),
.B2(n_7715),
.Y(n_8267)
);

OAI21x1_ASAP7_75t_L g8268 ( 
.A1(n_7927),
.A2(n_7708),
.B(n_7559),
.Y(n_8268)
);

INVx1_ASAP7_75t_L g8269 ( 
.A(n_7986),
.Y(n_8269)
);

OAI22xp33_ASAP7_75t_L g8270 ( 
.A1(n_8029),
.A2(n_7766),
.B1(n_7685),
.B2(n_7681),
.Y(n_8270)
);

HB1xp67_ASAP7_75t_L g8271 ( 
.A(n_8177),
.Y(n_8271)
);

INVx2_ASAP7_75t_L g8272 ( 
.A(n_8046),
.Y(n_8272)
);

AND2x4_ASAP7_75t_L g8273 ( 
.A(n_8020),
.B(n_7682),
.Y(n_8273)
);

NAND2xp5_ASAP7_75t_L g8274 ( 
.A(n_8052),
.B(n_7696),
.Y(n_8274)
);

OR2x2_ASAP7_75t_L g8275 ( 
.A(n_7990),
.B(n_7992),
.Y(n_8275)
);

A2O1A1Ixp33_ASAP7_75t_L g8276 ( 
.A1(n_7976),
.A2(n_7710),
.B(n_7572),
.C(n_7579),
.Y(n_8276)
);

AND2x2_ASAP7_75t_L g8277 ( 
.A(n_8180),
.B(n_8181),
.Y(n_8277)
);

HB1xp67_ASAP7_75t_L g8278 ( 
.A(n_7978),
.Y(n_8278)
);

NAND2xp5_ASAP7_75t_L g8279 ( 
.A(n_8188),
.B(n_7548),
.Y(n_8279)
);

NAND2xp5_ASAP7_75t_L g8280 ( 
.A(n_8183),
.B(n_7588),
.Y(n_8280)
);

NAND2xp5_ASAP7_75t_L g8281 ( 
.A(n_8190),
.B(n_7949),
.Y(n_8281)
);

BUFx2_ASAP7_75t_L g8282 ( 
.A(n_8210),
.Y(n_8282)
);

NAND2xp5_ASAP7_75t_L g8283 ( 
.A(n_8085),
.B(n_8086),
.Y(n_8283)
);

INVx2_ASAP7_75t_L g8284 ( 
.A(n_7994),
.Y(n_8284)
);

AOI22xp33_ASAP7_75t_L g8285 ( 
.A1(n_7980),
.A2(n_7752),
.B1(n_7739),
.B2(n_7689),
.Y(n_8285)
);

INVx3_ASAP7_75t_L g8286 ( 
.A(n_8150),
.Y(n_8286)
);

AND2x4_ASAP7_75t_L g8287 ( 
.A(n_8077),
.B(n_8206),
.Y(n_8287)
);

INVx2_ASAP7_75t_L g8288 ( 
.A(n_8004),
.Y(n_8288)
);

OAI22xp5_ASAP7_75t_L g8289 ( 
.A1(n_7995),
.A2(n_7685),
.B1(n_7655),
.B2(n_7649),
.Y(n_8289)
);

INVx2_ASAP7_75t_SL g8290 ( 
.A(n_8162),
.Y(n_8290)
);

INVx1_ASAP7_75t_L g8291 ( 
.A(n_8005),
.Y(n_8291)
);

CKINVDCx12_ASAP7_75t_R g8292 ( 
.A(n_8224),
.Y(n_8292)
);

AOI22xp33_ASAP7_75t_L g8293 ( 
.A1(n_8060),
.A2(n_7567),
.B1(n_7554),
.B2(n_7677),
.Y(n_8293)
);

AOI21xp5_ASAP7_75t_L g8294 ( 
.A1(n_7928),
.A2(n_7930),
.B(n_7934),
.Y(n_8294)
);

AOI222xp33_ASAP7_75t_L g8295 ( 
.A1(n_8091),
.A2(n_7567),
.B1(n_7554),
.B2(n_335),
.C1(n_337),
.C2(n_332),
.Y(n_8295)
);

OAI22xp5_ASAP7_75t_L g8296 ( 
.A1(n_8208),
.A2(n_336),
.B1(n_334),
.B2(n_335),
.Y(n_8296)
);

NOR2xp33_ASAP7_75t_L g8297 ( 
.A(n_7981),
.B(n_1416),
.Y(n_8297)
);

INVx6_ASAP7_75t_L g8298 ( 
.A(n_8043),
.Y(n_8298)
);

AND2x4_ASAP7_75t_L g8299 ( 
.A(n_8044),
.B(n_1417),
.Y(n_8299)
);

AOI22xp33_ASAP7_75t_L g8300 ( 
.A1(n_8049),
.A2(n_1418),
.B1(n_1419),
.B2(n_1417),
.Y(n_8300)
);

OA21x2_ASAP7_75t_L g8301 ( 
.A1(n_7951),
.A2(n_1420),
.B(n_1418),
.Y(n_8301)
);

OAI22xp5_ASAP7_75t_L g8302 ( 
.A1(n_7963),
.A2(n_336),
.B1(n_334),
.B2(n_335),
.Y(n_8302)
);

HB1xp67_ASAP7_75t_L g8303 ( 
.A(n_8011),
.Y(n_8303)
);

INVx1_ASAP7_75t_L g8304 ( 
.A(n_8016),
.Y(n_8304)
);

AOI22xp33_ASAP7_75t_L g8305 ( 
.A1(n_8110),
.A2(n_1422),
.B1(n_1424),
.B2(n_1421),
.Y(n_8305)
);

OAI22xp5_ASAP7_75t_L g8306 ( 
.A1(n_7961),
.A2(n_338),
.B1(n_336),
.B2(n_337),
.Y(n_8306)
);

AND2x2_ASAP7_75t_L g8307 ( 
.A(n_8205),
.B(n_8194),
.Y(n_8307)
);

OAI21xp5_ASAP7_75t_L g8308 ( 
.A1(n_7945),
.A2(n_337),
.B(n_338),
.Y(n_8308)
);

INVx1_ASAP7_75t_L g8309 ( 
.A(n_8019),
.Y(n_8309)
);

INVx1_ASAP7_75t_L g8310 ( 
.A(n_8024),
.Y(n_8310)
);

INVx4_ASAP7_75t_L g8311 ( 
.A(n_8162),
.Y(n_8311)
);

AND2x2_ASAP7_75t_L g8312 ( 
.A(n_8204),
.B(n_1421),
.Y(n_8312)
);

OAI221xp5_ASAP7_75t_L g8313 ( 
.A1(n_8193),
.A2(n_341),
.B1(n_338),
.B2(n_339),
.C(n_342),
.Y(n_8313)
);

AOI22xp33_ASAP7_75t_L g8314 ( 
.A1(n_7974),
.A2(n_1427),
.B1(n_1428),
.B2(n_1422),
.Y(n_8314)
);

INVx3_ASAP7_75t_L g8315 ( 
.A(n_8150),
.Y(n_8315)
);

AOI322xp5_ASAP7_75t_L g8316 ( 
.A1(n_8061),
.A2(n_346),
.A3(n_345),
.B1(n_343),
.B2(n_339),
.C1(n_342),
.C2(n_344),
.Y(n_8316)
);

INVx1_ASAP7_75t_L g8317 ( 
.A(n_8045),
.Y(n_8317)
);

OAI22xp33_ASAP7_75t_L g8318 ( 
.A1(n_7984),
.A2(n_343),
.B1(n_339),
.B2(n_342),
.Y(n_8318)
);

OAI22xp5_ASAP7_75t_L g8319 ( 
.A1(n_7965),
.A2(n_345),
.B1(n_343),
.B2(n_344),
.Y(n_8319)
);

INVx3_ASAP7_75t_L g8320 ( 
.A(n_8152),
.Y(n_8320)
);

AOI22xp33_ASAP7_75t_L g8321 ( 
.A1(n_8076),
.A2(n_1428),
.B1(n_1429),
.B2(n_1427),
.Y(n_8321)
);

INVx2_ASAP7_75t_L g8322 ( 
.A(n_8053),
.Y(n_8322)
);

AOI22xp33_ASAP7_75t_L g8323 ( 
.A1(n_8127),
.A2(n_1430),
.B1(n_1431),
.B2(n_1429),
.Y(n_8323)
);

AOI22xp33_ASAP7_75t_L g8324 ( 
.A1(n_8157),
.A2(n_1432),
.B1(n_1434),
.B2(n_1431),
.Y(n_8324)
);

INVx1_ASAP7_75t_L g8325 ( 
.A(n_8056),
.Y(n_8325)
);

INVx4_ASAP7_75t_SL g8326 ( 
.A(n_8108),
.Y(n_8326)
);

AOI22xp33_ASAP7_75t_L g8327 ( 
.A1(n_8106),
.A2(n_1436),
.B1(n_1437),
.B2(n_1434),
.Y(n_8327)
);

INVx1_ASAP7_75t_L g8328 ( 
.A(n_8058),
.Y(n_8328)
);

AOI22xp33_ASAP7_75t_L g8329 ( 
.A1(n_8003),
.A2(n_1437),
.B1(n_1439),
.B2(n_1436),
.Y(n_8329)
);

OR2x2_ASAP7_75t_L g8330 ( 
.A(n_8062),
.B(n_1439),
.Y(n_8330)
);

O2A1O1Ixp5_ASAP7_75t_L g8331 ( 
.A1(n_8178),
.A2(n_346),
.B(n_344),
.C(n_345),
.Y(n_8331)
);

AND2x2_ASAP7_75t_L g8332 ( 
.A(n_8072),
.B(n_8146),
.Y(n_8332)
);

OAI22xp5_ASAP7_75t_L g8333 ( 
.A1(n_8022),
.A2(n_8137),
.B1(n_8116),
.B2(n_8118),
.Y(n_8333)
);

HB1xp67_ASAP7_75t_L g8334 ( 
.A(n_8090),
.Y(n_8334)
);

INVx4_ASAP7_75t_L g8335 ( 
.A(n_8043),
.Y(n_8335)
);

INVx1_ASAP7_75t_L g8336 ( 
.A(n_8097),
.Y(n_8336)
);

INVx3_ASAP7_75t_L g8337 ( 
.A(n_8152),
.Y(n_8337)
);

AND2x2_ASAP7_75t_L g8338 ( 
.A(n_8229),
.B(n_1440),
.Y(n_8338)
);

OAI22xp33_ASAP7_75t_SL g8339 ( 
.A1(n_8080),
.A2(n_348),
.B1(n_346),
.B2(n_347),
.Y(n_8339)
);

INVx1_ASAP7_75t_L g8340 ( 
.A(n_8126),
.Y(n_8340)
);

INVx1_ASAP7_75t_L g8341 ( 
.A(n_8140),
.Y(n_8341)
);

INVx1_ASAP7_75t_SL g8342 ( 
.A(n_8167),
.Y(n_8342)
);

OAI22xp5_ASAP7_75t_L g8343 ( 
.A1(n_8113),
.A2(n_349),
.B1(n_347),
.B2(n_348),
.Y(n_8343)
);

OAI221xp5_ASAP7_75t_L g8344 ( 
.A1(n_8051),
.A2(n_350),
.B1(n_348),
.B2(n_349),
.C(n_351),
.Y(n_8344)
);

INVx2_ASAP7_75t_L g8345 ( 
.A(n_7975),
.Y(n_8345)
);

AOI22xp33_ASAP7_75t_L g8346 ( 
.A1(n_8047),
.A2(n_7936),
.B1(n_8087),
.B2(n_8025),
.Y(n_8346)
);

INVx6_ASAP7_75t_L g8347 ( 
.A(n_8075),
.Y(n_8347)
);

AND2x4_ASAP7_75t_L g8348 ( 
.A(n_8143),
.B(n_8176),
.Y(n_8348)
);

CKINVDCx5p33_ASAP7_75t_R g8349 ( 
.A(n_8125),
.Y(n_8349)
);

INVx6_ASAP7_75t_L g8350 ( 
.A(n_7987),
.Y(n_8350)
);

BUFx2_ASAP7_75t_L g8351 ( 
.A(n_7972),
.Y(n_8351)
);

AOI22xp33_ASAP7_75t_L g8352 ( 
.A1(n_8031),
.A2(n_1442),
.B1(n_1443),
.B2(n_1441),
.Y(n_8352)
);

INVx2_ASAP7_75t_L g8353 ( 
.A(n_8102),
.Y(n_8353)
);

INVx1_ASAP7_75t_L g8354 ( 
.A(n_8104),
.Y(n_8354)
);

INVx1_ASAP7_75t_L g8355 ( 
.A(n_8109),
.Y(n_8355)
);

OAI22xp5_ASAP7_75t_L g8356 ( 
.A1(n_7931),
.A2(n_352),
.B1(n_350),
.B2(n_351),
.Y(n_8356)
);

OAI22xp5_ASAP7_75t_L g8357 ( 
.A1(n_7931),
.A2(n_353),
.B1(n_351),
.B2(n_352),
.Y(n_8357)
);

INVx1_ASAP7_75t_SL g8358 ( 
.A(n_8121),
.Y(n_8358)
);

INVx6_ASAP7_75t_L g8359 ( 
.A(n_8023),
.Y(n_8359)
);

O2A1O1Ixp33_ASAP7_75t_SL g8360 ( 
.A1(n_8230),
.A2(n_1442),
.B(n_1443),
.C(n_1441),
.Y(n_8360)
);

AOI21xp5_ASAP7_75t_L g8361 ( 
.A1(n_7924),
.A2(n_353),
.B(n_354),
.Y(n_8361)
);

OR2x2_ASAP7_75t_L g8362 ( 
.A(n_7944),
.B(n_1444),
.Y(n_8362)
);

A2O1A1Ixp33_ASAP7_75t_L g8363 ( 
.A1(n_8074),
.A2(n_1446),
.B(n_1447),
.C(n_1445),
.Y(n_8363)
);

INVx2_ASAP7_75t_L g8364 ( 
.A(n_8135),
.Y(n_8364)
);

OAI22xp33_ASAP7_75t_L g8365 ( 
.A1(n_7998),
.A2(n_355),
.B1(n_353),
.B2(n_354),
.Y(n_8365)
);

OAI21x1_ASAP7_75t_L g8366 ( 
.A1(n_7948),
.A2(n_355),
.B(n_356),
.Y(n_8366)
);

HB1xp67_ASAP7_75t_L g8367 ( 
.A(n_8001),
.Y(n_8367)
);

INVx2_ASAP7_75t_L g8368 ( 
.A(n_8138),
.Y(n_8368)
);

INVx2_ASAP7_75t_L g8369 ( 
.A(n_8142),
.Y(n_8369)
);

NAND2xp5_ASAP7_75t_L g8370 ( 
.A(n_8145),
.B(n_1446),
.Y(n_8370)
);

CKINVDCx5p33_ASAP7_75t_R g8371 ( 
.A(n_8038),
.Y(n_8371)
);

OAI22xp5_ASAP7_75t_L g8372 ( 
.A1(n_7997),
.A2(n_357),
.B1(n_355),
.B2(n_356),
.Y(n_8372)
);

OAI22xp33_ASAP7_75t_L g8373 ( 
.A1(n_8080),
.A2(n_8009),
.B1(n_8037),
.B2(n_8147),
.Y(n_8373)
);

INVx5_ASAP7_75t_L g8374 ( 
.A(n_8224),
.Y(n_8374)
);

INVx2_ASAP7_75t_L g8375 ( 
.A(n_8153),
.Y(n_8375)
);

OAI22xp5_ASAP7_75t_L g8376 ( 
.A1(n_8078),
.A2(n_358),
.B1(n_356),
.B2(n_357),
.Y(n_8376)
);

OAI22xp5_ASAP7_75t_L g8377 ( 
.A1(n_7971),
.A2(n_359),
.B1(n_357),
.B2(n_358),
.Y(n_8377)
);

NAND2xp5_ASAP7_75t_L g8378 ( 
.A(n_8182),
.B(n_1449),
.Y(n_8378)
);

AND2x2_ASAP7_75t_L g8379 ( 
.A(n_8192),
.B(n_8010),
.Y(n_8379)
);

AOI22xp33_ASAP7_75t_L g8380 ( 
.A1(n_8187),
.A2(n_1450),
.B1(n_1451),
.B2(n_1449),
.Y(n_8380)
);

AOI22xp33_ASAP7_75t_L g8381 ( 
.A1(n_7979),
.A2(n_1454),
.B1(n_1455),
.B2(n_1453),
.Y(n_8381)
);

INVx1_ASAP7_75t_L g8382 ( 
.A(n_8001),
.Y(n_8382)
);

OAI22xp33_ASAP7_75t_L g8383 ( 
.A1(n_8134),
.A2(n_361),
.B1(n_359),
.B2(n_360),
.Y(n_8383)
);

INVx3_ASAP7_75t_L g8384 ( 
.A(n_8163),
.Y(n_8384)
);

O2A1O1Ixp33_ASAP7_75t_L g8385 ( 
.A1(n_8174),
.A2(n_361),
.B(n_359),
.C(n_360),
.Y(n_8385)
);

BUFx2_ASAP7_75t_L g8386 ( 
.A(n_8226),
.Y(n_8386)
);

CKINVDCx5p33_ASAP7_75t_R g8387 ( 
.A(n_8036),
.Y(n_8387)
);

AND2x4_ASAP7_75t_L g8388 ( 
.A(n_8226),
.B(n_1453),
.Y(n_8388)
);

NAND2xp5_ASAP7_75t_L g8389 ( 
.A(n_8039),
.B(n_1455),
.Y(n_8389)
);

INVx2_ASAP7_75t_L g8390 ( 
.A(n_7985),
.Y(n_8390)
);

INVx2_ASAP7_75t_L g8391 ( 
.A(n_8002),
.Y(n_8391)
);

OAI22xp5_ASAP7_75t_L g8392 ( 
.A1(n_7957),
.A2(n_363),
.B1(n_360),
.B2(n_362),
.Y(n_8392)
);

INVx2_ASAP7_75t_L g8393 ( 
.A(n_7962),
.Y(n_8393)
);

AOI22xp33_ASAP7_75t_L g8394 ( 
.A1(n_8105),
.A2(n_1457),
.B1(n_1458),
.B2(n_1456),
.Y(n_8394)
);

NOR2x1_ASAP7_75t_SL g8395 ( 
.A(n_8212),
.B(n_1457),
.Y(n_8395)
);

AND2x4_ASAP7_75t_L g8396 ( 
.A(n_8221),
.B(n_1458),
.Y(n_8396)
);

NAND2xp5_ASAP7_75t_L g8397 ( 
.A(n_8185),
.B(n_1459),
.Y(n_8397)
);

NAND2xp5_ASAP7_75t_L g8398 ( 
.A(n_8066),
.B(n_8013),
.Y(n_8398)
);

INVx1_ASAP7_75t_L g8399 ( 
.A(n_8030),
.Y(n_8399)
);

CKINVDCx6p67_ASAP7_75t_R g8400 ( 
.A(n_8048),
.Y(n_8400)
);

HB1xp67_ASAP7_75t_L g8401 ( 
.A(n_8070),
.Y(n_8401)
);

AND2x4_ASAP7_75t_L g8402 ( 
.A(n_8232),
.B(n_1459),
.Y(n_8402)
);

INVx3_ASAP7_75t_L g8403 ( 
.A(n_8163),
.Y(n_8403)
);

AOI22xp33_ASAP7_75t_L g8404 ( 
.A1(n_7967),
.A2(n_1463),
.B1(n_1464),
.B2(n_1462),
.Y(n_8404)
);

INVx1_ASAP7_75t_SL g8405 ( 
.A(n_8169),
.Y(n_8405)
);

AOI22xp5_ASAP7_75t_L g8406 ( 
.A1(n_8132),
.A2(n_365),
.B1(n_362),
.B2(n_364),
.Y(n_8406)
);

AOI221xp5_ASAP7_75t_L g8407 ( 
.A1(n_8000),
.A2(n_366),
.B1(n_362),
.B2(n_364),
.C(n_367),
.Y(n_8407)
);

INVx2_ASAP7_75t_L g8408 ( 
.A(n_8071),
.Y(n_8408)
);

OR2x2_ASAP7_75t_L g8409 ( 
.A(n_8026),
.B(n_1462),
.Y(n_8409)
);

OAI22xp5_ASAP7_75t_L g8410 ( 
.A1(n_8148),
.A2(n_368),
.B1(n_364),
.B2(n_367),
.Y(n_8410)
);

INVx1_ASAP7_75t_L g8411 ( 
.A(n_8030),
.Y(n_8411)
);

INVx4_ASAP7_75t_SL g8412 ( 
.A(n_8186),
.Y(n_8412)
);

INVx3_ASAP7_75t_SL g8413 ( 
.A(n_7989),
.Y(n_8413)
);

AO31x2_ASAP7_75t_L g8414 ( 
.A1(n_7991),
.A2(n_370),
.A3(n_368),
.B(n_369),
.Y(n_8414)
);

OAI22xp5_ASAP7_75t_L g8415 ( 
.A1(n_8124),
.A2(n_370),
.B1(n_368),
.B2(n_369),
.Y(n_8415)
);

A2O1A1Ixp33_ASAP7_75t_L g8416 ( 
.A1(n_8201),
.A2(n_1465),
.B(n_1466),
.C(n_1463),
.Y(n_8416)
);

AOI22xp33_ASAP7_75t_L g8417 ( 
.A1(n_7999),
.A2(n_1467),
.B1(n_1468),
.B2(n_1465),
.Y(n_8417)
);

INVx2_ASAP7_75t_SL g8418 ( 
.A(n_8211),
.Y(n_8418)
);

AOI221xp5_ASAP7_75t_L g8419 ( 
.A1(n_8144),
.A2(n_373),
.B1(n_371),
.B2(n_372),
.C(n_374),
.Y(n_8419)
);

INVx2_ASAP7_75t_L g8420 ( 
.A(n_8057),
.Y(n_8420)
);

OAI221xp5_ASAP7_75t_L g8421 ( 
.A1(n_8035),
.A2(n_373),
.B1(n_371),
.B2(n_372),
.C(n_374),
.Y(n_8421)
);

INVx1_ASAP7_75t_L g8422 ( 
.A(n_8114),
.Y(n_8422)
);

HB1xp67_ASAP7_75t_L g8423 ( 
.A(n_7932),
.Y(n_8423)
);

AOI22xp33_ASAP7_75t_L g8424 ( 
.A1(n_8028),
.A2(n_1469),
.B1(n_1470),
.B2(n_1467),
.Y(n_8424)
);

INVx4_ASAP7_75t_L g8425 ( 
.A(n_7943),
.Y(n_8425)
);

NAND2xp5_ASAP7_75t_L g8426 ( 
.A(n_8136),
.B(n_1469),
.Y(n_8426)
);

INVx2_ASAP7_75t_L g8427 ( 
.A(n_8119),
.Y(n_8427)
);

AND2x4_ASAP7_75t_L g8428 ( 
.A(n_8165),
.B(n_1470),
.Y(n_8428)
);

AOI22xp33_ASAP7_75t_L g8429 ( 
.A1(n_8151),
.A2(n_1472),
.B1(n_1473),
.B2(n_1471),
.Y(n_8429)
);

INVx1_ASAP7_75t_L g8430 ( 
.A(n_8114),
.Y(n_8430)
);

BUFx6f_ASAP7_75t_L g8431 ( 
.A(n_8234),
.Y(n_8431)
);

OAI22xp5_ASAP7_75t_L g8432 ( 
.A1(n_8007),
.A2(n_374),
.B1(n_371),
.B2(n_372),
.Y(n_8432)
);

INVx2_ASAP7_75t_L g8433 ( 
.A(n_8213),
.Y(n_8433)
);

INVx2_ASAP7_75t_L g8434 ( 
.A(n_8115),
.Y(n_8434)
);

OAI22xp33_ASAP7_75t_L g8435 ( 
.A1(n_8233),
.A2(n_8198),
.B1(n_8200),
.B2(n_8168),
.Y(n_8435)
);

AND2x2_ASAP7_75t_L g8436 ( 
.A(n_8155),
.B(n_1471),
.Y(n_8436)
);

NAND2xp5_ASAP7_75t_L g8437 ( 
.A(n_8092),
.B(n_8166),
.Y(n_8437)
);

AND2x2_ASAP7_75t_L g8438 ( 
.A(n_8069),
.B(n_1474),
.Y(n_8438)
);

INVx1_ASAP7_75t_L g8439 ( 
.A(n_8115),
.Y(n_8439)
);

INVx1_ASAP7_75t_SL g8440 ( 
.A(n_8234),
.Y(n_8440)
);

INVx4_ASAP7_75t_L g8441 ( 
.A(n_7943),
.Y(n_8441)
);

AOI22xp33_ASAP7_75t_L g8442 ( 
.A1(n_8164),
.A2(n_1475),
.B1(n_1476),
.B2(n_1474),
.Y(n_8442)
);

NOR2xp33_ASAP7_75t_L g8443 ( 
.A(n_8225),
.B(n_8222),
.Y(n_8443)
);

OAI22xp5_ASAP7_75t_L g8444 ( 
.A1(n_8012),
.A2(n_377),
.B1(n_375),
.B2(n_376),
.Y(n_8444)
);

INVx1_ASAP7_75t_L g8445 ( 
.A(n_8158),
.Y(n_8445)
);

AO31x2_ASAP7_75t_L g8446 ( 
.A1(n_8041),
.A2(n_8055),
.A3(n_8156),
.B(n_8175),
.Y(n_8446)
);

INVx3_ASAP7_75t_L g8447 ( 
.A(n_7988),
.Y(n_8447)
);

AOI22xp33_ASAP7_75t_SL g8448 ( 
.A1(n_8111),
.A2(n_377),
.B1(n_375),
.B2(n_376),
.Y(n_8448)
);

INVx1_ASAP7_75t_L g8449 ( 
.A(n_8158),
.Y(n_8449)
);

AOI22xp33_ASAP7_75t_L g8450 ( 
.A1(n_8139),
.A2(n_1477),
.B1(n_1478),
.B2(n_1476),
.Y(n_8450)
);

INVx1_ASAP7_75t_L g8451 ( 
.A(n_7969),
.Y(n_8451)
);

OAI22xp5_ASAP7_75t_L g8452 ( 
.A1(n_8130),
.A2(n_378),
.B1(n_375),
.B2(n_377),
.Y(n_8452)
);

INVx6_ASAP7_75t_L g8453 ( 
.A(n_7993),
.Y(n_8453)
);

AOI22xp33_ASAP7_75t_L g8454 ( 
.A1(n_8040),
.A2(n_1478),
.B1(n_1479),
.B2(n_1477),
.Y(n_8454)
);

CKINVDCx20_ASAP7_75t_R g8455 ( 
.A(n_8033),
.Y(n_8455)
);

INVx1_ASAP7_75t_L g8456 ( 
.A(n_8218),
.Y(n_8456)
);

BUFx3_ASAP7_75t_L g8457 ( 
.A(n_8054),
.Y(n_8457)
);

AOI22xp33_ASAP7_75t_L g8458 ( 
.A1(n_8079),
.A2(n_1480),
.B1(n_1481),
.B2(n_1479),
.Y(n_8458)
);

INVx1_ASAP7_75t_L g8459 ( 
.A(n_8218),
.Y(n_8459)
);

AOI22xp33_ASAP7_75t_L g8460 ( 
.A1(n_7953),
.A2(n_1482),
.B1(n_1483),
.B2(n_1481),
.Y(n_8460)
);

AND2x2_ASAP7_75t_L g8461 ( 
.A(n_8103),
.B(n_1482),
.Y(n_8461)
);

INVx2_ASAP7_75t_L g8462 ( 
.A(n_8018),
.Y(n_8462)
);

AOI22xp33_ASAP7_75t_L g8463 ( 
.A1(n_8064),
.A2(n_1487),
.B1(n_1488),
.B2(n_1485),
.Y(n_8463)
);

INVx3_ASAP7_75t_L g8464 ( 
.A(n_8207),
.Y(n_8464)
);

NAND2xp5_ASAP7_75t_L g8465 ( 
.A(n_8159),
.B(n_1485),
.Y(n_8465)
);

INVx2_ASAP7_75t_L g8466 ( 
.A(n_8209),
.Y(n_8466)
);

INVx1_ASAP7_75t_SL g8467 ( 
.A(n_8203),
.Y(n_8467)
);

INVxp67_ASAP7_75t_L g8468 ( 
.A(n_8089),
.Y(n_8468)
);

NAND2xp5_ASAP7_75t_L g8469 ( 
.A(n_8184),
.B(n_1487),
.Y(n_8469)
);

NAND3xp33_ASAP7_75t_L g8470 ( 
.A(n_8173),
.B(n_378),
.C(n_379),
.Y(n_8470)
);

AOI221xp5_ASAP7_75t_L g8471 ( 
.A1(n_8191),
.A2(n_381),
.B1(n_378),
.B2(n_380),
.C(n_382),
.Y(n_8471)
);

INVx2_ASAP7_75t_L g8472 ( 
.A(n_8059),
.Y(n_8472)
);

INVx3_ASAP7_75t_L g8473 ( 
.A(n_8212),
.Y(n_8473)
);

OAI221xp5_ASAP7_75t_L g8474 ( 
.A1(n_8131),
.A2(n_382),
.B1(n_380),
.B2(n_381),
.C(n_383),
.Y(n_8474)
);

OAI221xp5_ASAP7_75t_L g8475 ( 
.A1(n_8117),
.A2(n_383),
.B1(n_380),
.B2(n_381),
.C(n_384),
.Y(n_8475)
);

A2O1A1Ixp33_ASAP7_75t_L g8476 ( 
.A1(n_7940),
.A2(n_1491),
.B(n_1493),
.C(n_1490),
.Y(n_8476)
);

AOI22xp33_ASAP7_75t_L g8477 ( 
.A1(n_7973),
.A2(n_1491),
.B1(n_1493),
.B2(n_1490),
.Y(n_8477)
);

AOI21xp5_ASAP7_75t_L g8478 ( 
.A1(n_8027),
.A2(n_384),
.B(n_385),
.Y(n_8478)
);

AOI22xp33_ASAP7_75t_L g8479 ( 
.A1(n_8217),
.A2(n_1495),
.B1(n_1496),
.B2(n_1494),
.Y(n_8479)
);

INVx3_ASAP7_75t_L g8480 ( 
.A(n_8099),
.Y(n_8480)
);

AOI22xp33_ASAP7_75t_L g8481 ( 
.A1(n_8034),
.A2(n_8219),
.B1(n_8216),
.B2(n_8050),
.Y(n_8481)
);

OR2x6_ASAP7_75t_L g8482 ( 
.A(n_8236),
.B(n_1496),
.Y(n_8482)
);

BUFx2_ASAP7_75t_L g8483 ( 
.A(n_8032),
.Y(n_8483)
);

AOI211xp5_ASAP7_75t_L g8484 ( 
.A1(n_8223),
.A2(n_386),
.B(n_384),
.C(n_385),
.Y(n_8484)
);

INVx2_ASAP7_75t_L g8485 ( 
.A(n_8067),
.Y(n_8485)
);

AOI21xp5_ASAP7_75t_L g8486 ( 
.A1(n_7938),
.A2(n_385),
.B(n_386),
.Y(n_8486)
);

HB1xp67_ASAP7_75t_L g8487 ( 
.A(n_7926),
.Y(n_8487)
);

INVx1_ASAP7_75t_L g8488 ( 
.A(n_8063),
.Y(n_8488)
);

AOI22xp33_ASAP7_75t_L g8489 ( 
.A1(n_8094),
.A2(n_1499),
.B1(n_1500),
.B2(n_1498),
.Y(n_8489)
);

INVx3_ASAP7_75t_L g8490 ( 
.A(n_7966),
.Y(n_8490)
);

OAI22xp33_ASAP7_75t_SL g8491 ( 
.A1(n_7983),
.A2(n_388),
.B1(n_386),
.B2(n_387),
.Y(n_8491)
);

AOI22xp33_ASAP7_75t_SL g8492 ( 
.A1(n_8202),
.A2(n_389),
.B1(n_387),
.B2(n_388),
.Y(n_8492)
);

OAI22xp33_ASAP7_75t_L g8493 ( 
.A1(n_8095),
.A2(n_391),
.B1(n_388),
.B2(n_390),
.Y(n_8493)
);

O2A1O1Ixp33_ASAP7_75t_L g8494 ( 
.A1(n_8231),
.A2(n_392),
.B(n_390),
.C(n_391),
.Y(n_8494)
);

OAI21xp5_ASAP7_75t_L g8495 ( 
.A1(n_8101),
.A2(n_390),
.B(n_391),
.Y(n_8495)
);

INVx2_ASAP7_75t_L g8496 ( 
.A(n_8096),
.Y(n_8496)
);

AOI22xp33_ASAP7_75t_L g8497 ( 
.A1(n_8098),
.A2(n_1499),
.B1(n_1501),
.B2(n_1498),
.Y(n_8497)
);

AOI22xp33_ASAP7_75t_L g8498 ( 
.A1(n_8123),
.A2(n_8107),
.B1(n_8154),
.B2(n_8129),
.Y(n_8498)
);

AND2x2_ASAP7_75t_L g8499 ( 
.A(n_8235),
.B(n_1502),
.Y(n_8499)
);

AOI21xp33_ASAP7_75t_L g8500 ( 
.A1(n_8133),
.A2(n_392),
.B(n_393),
.Y(n_8500)
);

NAND2xp5_ASAP7_75t_L g8501 ( 
.A(n_8112),
.B(n_1503),
.Y(n_8501)
);

INVx1_ASAP7_75t_L g8502 ( 
.A(n_8100),
.Y(n_8502)
);

OR2x6_ASAP7_75t_L g8503 ( 
.A(n_8228),
.B(n_1503),
.Y(n_8503)
);

AND2x2_ASAP7_75t_L g8504 ( 
.A(n_8195),
.B(n_8017),
.Y(n_8504)
);

BUFx3_ASAP7_75t_L g8505 ( 
.A(n_8214),
.Y(n_8505)
);

OAI22xp5_ASAP7_75t_L g8506 ( 
.A1(n_8083),
.A2(n_394),
.B1(n_392),
.B2(n_393),
.Y(n_8506)
);

AOI22xp33_ASAP7_75t_L g8507 ( 
.A1(n_8179),
.A2(n_1505),
.B1(n_1506),
.B2(n_1504),
.Y(n_8507)
);

OAI211xp5_ASAP7_75t_L g8508 ( 
.A1(n_8093),
.A2(n_395),
.B(n_393),
.C(n_394),
.Y(n_8508)
);

NAND3xp33_ASAP7_75t_L g8509 ( 
.A(n_8042),
.B(n_394),
.C(n_395),
.Y(n_8509)
);

BUFx6f_ASAP7_75t_L g8510 ( 
.A(n_8122),
.Y(n_8510)
);

INVx2_ASAP7_75t_L g8511 ( 
.A(n_8141),
.Y(n_8511)
);

INVx2_ASAP7_75t_L g8512 ( 
.A(n_8196),
.Y(n_8512)
);

NOR2xp33_ASAP7_75t_L g8513 ( 
.A(n_8006),
.B(n_1507),
.Y(n_8513)
);

CKINVDCx5p33_ASAP7_75t_R g8514 ( 
.A(n_8189),
.Y(n_8514)
);

BUFx4f_ASAP7_75t_SL g8515 ( 
.A(n_8161),
.Y(n_8515)
);

OAI22xp33_ASAP7_75t_SL g8516 ( 
.A1(n_8015),
.A2(n_399),
.B1(n_397),
.B2(n_398),
.Y(n_8516)
);

CKINVDCx8_ASAP7_75t_R g8517 ( 
.A(n_8015),
.Y(n_8517)
);

AND2x2_ASAP7_75t_L g8518 ( 
.A(n_8171),
.B(n_1508),
.Y(n_8518)
);

HB1xp67_ASAP7_75t_L g8519 ( 
.A(n_7926),
.Y(n_8519)
);

INVx2_ASAP7_75t_L g8520 ( 
.A(n_7950),
.Y(n_8520)
);

NOR2x1_ASAP7_75t_SL g8521 ( 
.A(n_8220),
.B(n_1509),
.Y(n_8521)
);

INVx1_ASAP7_75t_L g8522 ( 
.A(n_7950),
.Y(n_8522)
);

INVx1_ASAP7_75t_L g8523 ( 
.A(n_8303),
.Y(n_8523)
);

AO21x2_ASAP7_75t_L g8524 ( 
.A1(n_8382),
.A2(n_8215),
.B(n_8014),
.Y(n_8524)
);

AND2x2_ASAP7_75t_L g8525 ( 
.A(n_8282),
.B(n_7925),
.Y(n_8525)
);

INVx1_ASAP7_75t_L g8526 ( 
.A(n_8334),
.Y(n_8526)
);

NOR2x1_ASAP7_75t_SL g8527 ( 
.A(n_8398),
.B(n_8482),
.Y(n_8527)
);

INVx2_ASAP7_75t_SL g8528 ( 
.A(n_8298),
.Y(n_8528)
);

INVx1_ASAP7_75t_L g8529 ( 
.A(n_8238),
.Y(n_8529)
);

INVx2_ASAP7_75t_L g8530 ( 
.A(n_8251),
.Y(n_8530)
);

AND2x2_ASAP7_75t_L g8531 ( 
.A(n_8237),
.B(n_7925),
.Y(n_8531)
);

AOI21xp5_ASAP7_75t_L g8532 ( 
.A1(n_8294),
.A2(n_8308),
.B(n_8248),
.Y(n_8532)
);

AO21x2_ASAP7_75t_L g8533 ( 
.A1(n_8367),
.A2(n_7970),
.B(n_8220),
.Y(n_8533)
);

OAI22xp5_ASAP7_75t_L g8534 ( 
.A1(n_8503),
.A2(n_8346),
.B1(n_8517),
.B2(n_8476),
.Y(n_8534)
);

INVx3_ASAP7_75t_L g8535 ( 
.A(n_8311),
.Y(n_8535)
);

INVx2_ASAP7_75t_SL g8536 ( 
.A(n_8298),
.Y(n_8536)
);

INVx2_ASAP7_75t_L g8537 ( 
.A(n_8275),
.Y(n_8537)
);

BUFx3_ASAP7_75t_L g8538 ( 
.A(n_8258),
.Y(n_8538)
);

INVx2_ASAP7_75t_L g8539 ( 
.A(n_8284),
.Y(n_8539)
);

INVx2_ASAP7_75t_L g8540 ( 
.A(n_8288),
.Y(n_8540)
);

BUFx2_ASAP7_75t_L g8541 ( 
.A(n_8386),
.Y(n_8541)
);

OR2x6_ASAP7_75t_L g8542 ( 
.A(n_8241),
.B(n_8170),
.Y(n_8542)
);

AND2x2_ASAP7_75t_L g8543 ( 
.A(n_8277),
.B(n_8170),
.Y(n_8543)
);

CKINVDCx8_ASAP7_75t_R g8544 ( 
.A(n_8349),
.Y(n_8544)
);

INVx1_ASAP7_75t_L g8545 ( 
.A(n_8243),
.Y(n_8545)
);

AO21x2_ASAP7_75t_L g8546 ( 
.A1(n_8488),
.A2(n_8199),
.B(n_7954),
.Y(n_8546)
);

INVx1_ASAP7_75t_L g8547 ( 
.A(n_8244),
.Y(n_8547)
);

INVx1_ASAP7_75t_L g8548 ( 
.A(n_8245),
.Y(n_8548)
);

NOR2xp33_ASAP7_75t_L g8549 ( 
.A(n_8347),
.B(n_1509),
.Y(n_8549)
);

CKINVDCx5p33_ASAP7_75t_R g8550 ( 
.A(n_8387),
.Y(n_8550)
);

OAI21x1_ASAP7_75t_L g8551 ( 
.A1(n_8520),
.A2(n_8199),
.B(n_7954),
.Y(n_8551)
);

INVx1_ASAP7_75t_L g8552 ( 
.A(n_8253),
.Y(n_8552)
);

BUFx2_ASAP7_75t_L g8553 ( 
.A(n_8271),
.Y(n_8553)
);

INVx1_ASAP7_75t_L g8554 ( 
.A(n_8257),
.Y(n_8554)
);

INVx2_ASAP7_75t_L g8555 ( 
.A(n_8322),
.Y(n_8555)
);

BUFx3_ASAP7_75t_L g8556 ( 
.A(n_8413),
.Y(n_8556)
);

BUFx2_ASAP7_75t_L g8557 ( 
.A(n_8254),
.Y(n_8557)
);

INVx1_ASAP7_75t_L g8558 ( 
.A(n_8264),
.Y(n_8558)
);

INVx1_ASAP7_75t_L g8559 ( 
.A(n_8265),
.Y(n_8559)
);

INVx1_ASAP7_75t_L g8560 ( 
.A(n_8269),
.Y(n_8560)
);

AND2x2_ASAP7_75t_L g8561 ( 
.A(n_8278),
.B(n_7977),
.Y(n_8561)
);

INVx2_ASAP7_75t_L g8562 ( 
.A(n_8291),
.Y(n_8562)
);

NAND2xp5_ASAP7_75t_L g8563 ( 
.A(n_8281),
.B(n_8008),
.Y(n_8563)
);

INVx3_ASAP7_75t_L g8564 ( 
.A(n_8240),
.Y(n_8564)
);

INVx2_ASAP7_75t_L g8565 ( 
.A(n_8304),
.Y(n_8565)
);

INVx1_ASAP7_75t_L g8566 ( 
.A(n_8309),
.Y(n_8566)
);

INVx2_ASAP7_75t_L g8567 ( 
.A(n_8310),
.Y(n_8567)
);

INVx2_ASAP7_75t_L g8568 ( 
.A(n_8317),
.Y(n_8568)
);

INVx1_ASAP7_75t_L g8569 ( 
.A(n_8325),
.Y(n_8569)
);

OAI21xp5_ASAP7_75t_L g8570 ( 
.A1(n_8478),
.A2(n_8128),
.B(n_7977),
.Y(n_8570)
);

AOI22xp33_ASAP7_75t_SL g8571 ( 
.A1(n_8333),
.A2(n_7942),
.B1(n_8128),
.B2(n_8008),
.Y(n_8571)
);

NAND2xp5_ASAP7_75t_L g8572 ( 
.A(n_8332),
.B(n_1510),
.Y(n_8572)
);

AND2x2_ASAP7_75t_L g8573 ( 
.A(n_8250),
.B(n_7942),
.Y(n_8573)
);

INVx1_ASAP7_75t_SL g8574 ( 
.A(n_8255),
.Y(n_8574)
);

INVx3_ASAP7_75t_L g8575 ( 
.A(n_8457),
.Y(n_8575)
);

INVx2_ASAP7_75t_L g8576 ( 
.A(n_8328),
.Y(n_8576)
);

OAI21x1_ASAP7_75t_L g8577 ( 
.A1(n_8268),
.A2(n_398),
.B(n_399),
.Y(n_8577)
);

BUFx3_ASAP7_75t_L g8578 ( 
.A(n_8263),
.Y(n_8578)
);

INVx3_ASAP7_75t_L g8579 ( 
.A(n_8273),
.Y(n_8579)
);

INVx3_ASAP7_75t_L g8580 ( 
.A(n_8287),
.Y(n_8580)
);

INVx2_ASAP7_75t_L g8581 ( 
.A(n_8348),
.Y(n_8581)
);

INVx2_ASAP7_75t_SL g8582 ( 
.A(n_8347),
.Y(n_8582)
);

AOI21xp5_ASAP7_75t_L g8583 ( 
.A1(n_8318),
.A2(n_398),
.B(n_400),
.Y(n_8583)
);

INVx3_ASAP7_75t_L g8584 ( 
.A(n_8335),
.Y(n_8584)
);

BUFx2_ASAP7_75t_L g8585 ( 
.A(n_8473),
.Y(n_8585)
);

NAND2x1p5_ASAP7_75t_L g8586 ( 
.A(n_8260),
.B(n_1510),
.Y(n_8586)
);

BUFx6f_ASAP7_75t_L g8587 ( 
.A(n_8431),
.Y(n_8587)
);

OAI21x1_ASAP7_75t_L g8588 ( 
.A1(n_8434),
.A2(n_400),
.B(n_401),
.Y(n_8588)
);

INVx2_ASAP7_75t_L g8589 ( 
.A(n_8242),
.Y(n_8589)
);

OAI21xp5_ASAP7_75t_L g8590 ( 
.A1(n_8486),
.A2(n_1512),
.B(n_1511),
.Y(n_8590)
);

CKINVDCx20_ASAP7_75t_R g8591 ( 
.A(n_8400),
.Y(n_8591)
);

INVx2_ASAP7_75t_L g8592 ( 
.A(n_8246),
.Y(n_8592)
);

HB1xp67_ASAP7_75t_L g8593 ( 
.A(n_8423),
.Y(n_8593)
);

HB1xp67_ASAP7_75t_L g8594 ( 
.A(n_8390),
.Y(n_8594)
);

NAND2xp5_ASAP7_75t_L g8595 ( 
.A(n_8401),
.B(n_1511),
.Y(n_8595)
);

INVx1_ASAP7_75t_L g8596 ( 
.A(n_8283),
.Y(n_8596)
);

INVx2_ASAP7_75t_L g8597 ( 
.A(n_8272),
.Y(n_8597)
);

AOI22xp33_ASAP7_75t_SL g8598 ( 
.A1(n_8521),
.A2(n_1514),
.B1(n_1515),
.B2(n_1513),
.Y(n_8598)
);

AOI22xp33_ASAP7_75t_L g8599 ( 
.A1(n_8295),
.A2(n_1516),
.B1(n_1517),
.B2(n_1513),
.Y(n_8599)
);

AND2x2_ASAP7_75t_L g8600 ( 
.A(n_8261),
.B(n_400),
.Y(n_8600)
);

INVx1_ASAP7_75t_L g8601 ( 
.A(n_8336),
.Y(n_8601)
);

NOR2xp33_ASAP7_75t_L g8602 ( 
.A(n_8443),
.B(n_1516),
.Y(n_8602)
);

HB1xp67_ASAP7_75t_L g8603 ( 
.A(n_8502),
.Y(n_8603)
);

INVx1_ASAP7_75t_L g8604 ( 
.A(n_8340),
.Y(n_8604)
);

OR2x2_ASAP7_75t_L g8605 ( 
.A(n_8393),
.B(n_401),
.Y(n_8605)
);

INVx2_ASAP7_75t_L g8606 ( 
.A(n_8345),
.Y(n_8606)
);

BUFx2_ASAP7_75t_L g8607 ( 
.A(n_8351),
.Y(n_8607)
);

INVx2_ASAP7_75t_L g8608 ( 
.A(n_8353),
.Y(n_8608)
);

INVx1_ASAP7_75t_L g8609 ( 
.A(n_8341),
.Y(n_8609)
);

AND2x4_ASAP7_75t_L g8610 ( 
.A(n_8307),
.B(n_1517),
.Y(n_8610)
);

INVx2_ASAP7_75t_L g8611 ( 
.A(n_8364),
.Y(n_8611)
);

OAI21xp5_ASAP7_75t_L g8612 ( 
.A1(n_8389),
.A2(n_1519),
.B(n_1518),
.Y(n_8612)
);

NAND2xp5_ASAP7_75t_L g8613 ( 
.A(n_8391),
.B(n_1519),
.Y(n_8613)
);

NOR2xp33_ASAP7_75t_L g8614 ( 
.A(n_8510),
.B(n_1520),
.Y(n_8614)
);

BUFx3_ASAP7_75t_L g8615 ( 
.A(n_8455),
.Y(n_8615)
);

INVx3_ASAP7_75t_L g8616 ( 
.A(n_8453),
.Y(n_8616)
);

INVx2_ASAP7_75t_L g8617 ( 
.A(n_8368),
.Y(n_8617)
);

INVx1_ASAP7_75t_L g8618 ( 
.A(n_8354),
.Y(n_8618)
);

INVx2_ASAP7_75t_L g8619 ( 
.A(n_8369),
.Y(n_8619)
);

INVx2_ASAP7_75t_L g8620 ( 
.A(n_8375),
.Y(n_8620)
);

AOI22xp33_ASAP7_75t_L g8621 ( 
.A1(n_8503),
.A2(n_8470),
.B1(n_8515),
.B2(n_8313),
.Y(n_8621)
);

INVx2_ASAP7_75t_L g8622 ( 
.A(n_8355),
.Y(n_8622)
);

INVx3_ASAP7_75t_L g8623 ( 
.A(n_8453),
.Y(n_8623)
);

INVx2_ASAP7_75t_L g8624 ( 
.A(n_8427),
.Y(n_8624)
);

CKINVDCx6p67_ASAP7_75t_R g8625 ( 
.A(n_8374),
.Y(n_8625)
);

AND2x2_ASAP7_75t_L g8626 ( 
.A(n_8420),
.B(n_401),
.Y(n_8626)
);

BUFx3_ASAP7_75t_L g8627 ( 
.A(n_8371),
.Y(n_8627)
);

AO21x2_ASAP7_75t_L g8628 ( 
.A1(n_8422),
.A2(n_402),
.B(n_403),
.Y(n_8628)
);

AO21x1_ASAP7_75t_L g8629 ( 
.A1(n_8516),
.A2(n_402),
.B(n_403),
.Y(n_8629)
);

INVx2_ASAP7_75t_L g8630 ( 
.A(n_8466),
.Y(n_8630)
);

INVx2_ASAP7_75t_L g8631 ( 
.A(n_8433),
.Y(n_8631)
);

INVx1_ASAP7_75t_L g8632 ( 
.A(n_8399),
.Y(n_8632)
);

AOI22xp33_ASAP7_75t_L g8633 ( 
.A1(n_8407),
.A2(n_1521),
.B1(n_1522),
.B2(n_1520),
.Y(n_8633)
);

INVx1_ASAP7_75t_L g8634 ( 
.A(n_8411),
.Y(n_8634)
);

INVx2_ASAP7_75t_L g8635 ( 
.A(n_8279),
.Y(n_8635)
);

INVx5_ASAP7_75t_L g8636 ( 
.A(n_8482),
.Y(n_8636)
);

INVx1_ASAP7_75t_L g8637 ( 
.A(n_8430),
.Y(n_8637)
);

INVx2_ASAP7_75t_L g8638 ( 
.A(n_8512),
.Y(n_8638)
);

INVx1_ASAP7_75t_L g8639 ( 
.A(n_8439),
.Y(n_8639)
);

INVx1_ASAP7_75t_L g8640 ( 
.A(n_8522),
.Y(n_8640)
);

BUFx6f_ASAP7_75t_L g8641 ( 
.A(n_8431),
.Y(n_8641)
);

AOI21x1_ASAP7_75t_L g8642 ( 
.A1(n_8456),
.A2(n_402),
.B(n_404),
.Y(n_8642)
);

AOI21x1_ASAP7_75t_L g8643 ( 
.A1(n_8459),
.A2(n_405),
.B(n_406),
.Y(n_8643)
);

AND2x2_ASAP7_75t_L g8644 ( 
.A(n_8483),
.B(n_405),
.Y(n_8644)
);

AND2x2_ASAP7_75t_L g8645 ( 
.A(n_8379),
.B(n_406),
.Y(n_8645)
);

INVx1_ASAP7_75t_SL g8646 ( 
.A(n_8342),
.Y(n_8646)
);

INVx1_ASAP7_75t_L g8647 ( 
.A(n_8445),
.Y(n_8647)
);

INVx1_ASAP7_75t_L g8648 ( 
.A(n_8449),
.Y(n_8648)
);

INVx2_ASAP7_75t_L g8649 ( 
.A(n_8408),
.Y(n_8649)
);

INVx1_ASAP7_75t_L g8650 ( 
.A(n_8487),
.Y(n_8650)
);

INVx1_ASAP7_75t_L g8651 ( 
.A(n_8519),
.Y(n_8651)
);

INVx3_ASAP7_75t_L g8652 ( 
.A(n_8447),
.Y(n_8652)
);

OAI21x1_ASAP7_75t_L g8653 ( 
.A1(n_8451),
.A2(n_407),
.B(n_408),
.Y(n_8653)
);

INVx2_ASAP7_75t_L g8654 ( 
.A(n_8472),
.Y(n_8654)
);

INVx1_ASAP7_75t_L g8655 ( 
.A(n_8280),
.Y(n_8655)
);

NAND2xp5_ASAP7_75t_L g8656 ( 
.A(n_8485),
.B(n_1521),
.Y(n_8656)
);

OAI22xp5_ASAP7_75t_L g8657 ( 
.A1(n_8509),
.A2(n_409),
.B1(n_407),
.B2(n_408),
.Y(n_8657)
);

OR2x2_ASAP7_75t_L g8658 ( 
.A(n_8462),
.B(n_407),
.Y(n_8658)
);

INVx2_ASAP7_75t_L g8659 ( 
.A(n_8496),
.Y(n_8659)
);

A2O1A1Ixp33_ASAP7_75t_L g8660 ( 
.A1(n_8361),
.A2(n_1523),
.B(n_1524),
.C(n_1522),
.Y(n_8660)
);

AOI22xp5_ASAP7_75t_L g8661 ( 
.A1(n_8365),
.A2(n_1524),
.B1(n_1525),
.B2(n_1523),
.Y(n_8661)
);

INVx1_ASAP7_75t_L g8662 ( 
.A(n_8330),
.Y(n_8662)
);

INVx3_ASAP7_75t_L g8663 ( 
.A(n_8464),
.Y(n_8663)
);

NAND2xp5_ASAP7_75t_L g8664 ( 
.A(n_8511),
.B(n_1525),
.Y(n_8664)
);

INVx2_ASAP7_75t_L g8665 ( 
.A(n_8510),
.Y(n_8665)
);

INVx2_ASAP7_75t_L g8666 ( 
.A(n_8362),
.Y(n_8666)
);

OAI21x1_ASAP7_75t_L g8667 ( 
.A1(n_8366),
.A2(n_408),
.B(n_409),
.Y(n_8667)
);

OAI21x1_ASAP7_75t_L g8668 ( 
.A1(n_8370),
.A2(n_409),
.B(n_410),
.Y(n_8668)
);

INVx1_ASAP7_75t_L g8669 ( 
.A(n_8378),
.Y(n_8669)
);

OAI21xp5_ASAP7_75t_L g8670 ( 
.A1(n_8397),
.A2(n_1529),
.B(n_1526),
.Y(n_8670)
);

INVx1_ASAP7_75t_L g8671 ( 
.A(n_8301),
.Y(n_8671)
);

INVx1_ASAP7_75t_L g8672 ( 
.A(n_8468),
.Y(n_8672)
);

NAND2xp5_ASAP7_75t_L g8673 ( 
.A(n_8467),
.B(n_1526),
.Y(n_8673)
);

BUFx8_ASAP7_75t_L g8674 ( 
.A(n_8436),
.Y(n_8674)
);

INVx1_ASAP7_75t_L g8675 ( 
.A(n_8262),
.Y(n_8675)
);

INVx2_ASAP7_75t_SL g8676 ( 
.A(n_8350),
.Y(n_8676)
);

OA21x2_ASAP7_75t_L g8677 ( 
.A1(n_8437),
.A2(n_410),
.B(n_411),
.Y(n_8677)
);

HB1xp67_ASAP7_75t_L g8678 ( 
.A(n_8274),
.Y(n_8678)
);

BUFx4f_ASAP7_75t_SL g8679 ( 
.A(n_8425),
.Y(n_8679)
);

CKINVDCx11_ASAP7_75t_R g8680 ( 
.A(n_8326),
.Y(n_8680)
);

OAI21x1_ASAP7_75t_L g8681 ( 
.A1(n_8249),
.A2(n_411),
.B(n_412),
.Y(n_8681)
);

BUFx2_ASAP7_75t_L g8682 ( 
.A(n_8418),
.Y(n_8682)
);

INVx1_ASAP7_75t_L g8683 ( 
.A(n_8409),
.Y(n_8683)
);

AO21x1_ASAP7_75t_SL g8684 ( 
.A1(n_8256),
.A2(n_1530),
.B(n_1529),
.Y(n_8684)
);

INVx2_ASAP7_75t_L g8685 ( 
.A(n_8505),
.Y(n_8685)
);

AOI21x1_ASAP7_75t_L g8686 ( 
.A1(n_8518),
.A2(n_411),
.B(n_412),
.Y(n_8686)
);

INVx2_ASAP7_75t_L g8687 ( 
.A(n_8286),
.Y(n_8687)
);

INVx1_ASAP7_75t_L g8688 ( 
.A(n_8504),
.Y(n_8688)
);

INVx2_ASAP7_75t_L g8689 ( 
.A(n_8315),
.Y(n_8689)
);

NAND2xp5_ASAP7_75t_L g8690 ( 
.A(n_8469),
.B(n_1531),
.Y(n_8690)
);

INVx1_ASAP7_75t_L g8691 ( 
.A(n_8338),
.Y(n_8691)
);

INVx1_ASAP7_75t_L g8692 ( 
.A(n_8465),
.Y(n_8692)
);

AND2x2_ASAP7_75t_L g8693 ( 
.A(n_8405),
.B(n_412),
.Y(n_8693)
);

INVx2_ASAP7_75t_L g8694 ( 
.A(n_8320),
.Y(n_8694)
);

HB1xp67_ASAP7_75t_L g8695 ( 
.A(n_8480),
.Y(n_8695)
);

INVx1_ASAP7_75t_L g8696 ( 
.A(n_8312),
.Y(n_8696)
);

OAI21xp5_ASAP7_75t_L g8697 ( 
.A1(n_8363),
.A2(n_1532),
.B(n_1531),
.Y(n_8697)
);

INVx2_ASAP7_75t_L g8698 ( 
.A(n_8337),
.Y(n_8698)
);

BUFx3_ASAP7_75t_L g8699 ( 
.A(n_8350),
.Y(n_8699)
);

INVx1_ASAP7_75t_L g8700 ( 
.A(n_8414),
.Y(n_8700)
);

INVx1_ASAP7_75t_L g8701 ( 
.A(n_8414),
.Y(n_8701)
);

INVx1_ASAP7_75t_L g8702 ( 
.A(n_8501),
.Y(n_8702)
);

BUFx2_ASAP7_75t_SL g8703 ( 
.A(n_8374),
.Y(n_8703)
);

NOR2xp33_ASAP7_75t_L g8704 ( 
.A(n_8359),
.B(n_1532),
.Y(n_8704)
);

INVx2_ASAP7_75t_L g8705 ( 
.A(n_8384),
.Y(n_8705)
);

INVx1_ASAP7_75t_L g8706 ( 
.A(n_8461),
.Y(n_8706)
);

INVx2_ASAP7_75t_SL g8707 ( 
.A(n_8359),
.Y(n_8707)
);

OR2x2_ASAP7_75t_L g8708 ( 
.A(n_8358),
.B(n_413),
.Y(n_8708)
);

INVx1_ASAP7_75t_L g8709 ( 
.A(n_8403),
.Y(n_8709)
);

INVx1_ASAP7_75t_L g8710 ( 
.A(n_8438),
.Y(n_8710)
);

HB1xp67_ASAP7_75t_L g8711 ( 
.A(n_8440),
.Y(n_8711)
);

INVx1_ASAP7_75t_L g8712 ( 
.A(n_8299),
.Y(n_8712)
);

INVx2_ASAP7_75t_L g8713 ( 
.A(n_8290),
.Y(n_8713)
);

AOI22xp33_ASAP7_75t_L g8714 ( 
.A1(n_8419),
.A2(n_1534),
.B1(n_1535),
.B2(n_1533),
.Y(n_8714)
);

INVx1_ASAP7_75t_L g8715 ( 
.A(n_8446),
.Y(n_8715)
);

INVx2_ASAP7_75t_L g8716 ( 
.A(n_8396),
.Y(n_8716)
);

INVx1_ASAP7_75t_L g8717 ( 
.A(n_8446),
.Y(n_8717)
);

INVx2_ASAP7_75t_L g8718 ( 
.A(n_8402),
.Y(n_8718)
);

INVx1_ASAP7_75t_L g8719 ( 
.A(n_8426),
.Y(n_8719)
);

INVx3_ASAP7_75t_L g8720 ( 
.A(n_8441),
.Y(n_8720)
);

INVx2_ASAP7_75t_L g8721 ( 
.A(n_8490),
.Y(n_8721)
);

INVx1_ASAP7_75t_L g8722 ( 
.A(n_8331),
.Y(n_8722)
);

INVx2_ASAP7_75t_L g8723 ( 
.A(n_8428),
.Y(n_8723)
);

INVx1_ASAP7_75t_L g8724 ( 
.A(n_8297),
.Y(n_8724)
);

AND2x2_ASAP7_75t_L g8725 ( 
.A(n_8412),
.B(n_413),
.Y(n_8725)
);

INVx1_ASAP7_75t_L g8726 ( 
.A(n_8395),
.Y(n_8726)
);

INVx2_ASAP7_75t_L g8727 ( 
.A(n_8388),
.Y(n_8727)
);

INVx1_ASAP7_75t_L g8728 ( 
.A(n_8276),
.Y(n_8728)
);

INVx2_ASAP7_75t_L g8729 ( 
.A(n_8292),
.Y(n_8729)
);

INVx1_ASAP7_75t_L g8730 ( 
.A(n_8247),
.Y(n_8730)
);

AOI21x1_ASAP7_75t_L g8731 ( 
.A1(n_8356),
.A2(n_414),
.B(n_415),
.Y(n_8731)
);

INVx1_ASAP7_75t_L g8732 ( 
.A(n_8513),
.Y(n_8732)
);

AOI22xp33_ASAP7_75t_L g8733 ( 
.A1(n_8373),
.A2(n_1539),
.B1(n_1540),
.B2(n_1538),
.Y(n_8733)
);

INVx1_ASAP7_75t_L g8734 ( 
.A(n_8339),
.Y(n_8734)
);

HB1xp67_ASAP7_75t_L g8735 ( 
.A(n_8289),
.Y(n_8735)
);

INVx2_ASAP7_75t_L g8736 ( 
.A(n_8412),
.Y(n_8736)
);

INVx1_ASAP7_75t_L g8737 ( 
.A(n_8495),
.Y(n_8737)
);

INVx3_ASAP7_75t_L g8738 ( 
.A(n_8499),
.Y(n_8738)
);

INVx3_ASAP7_75t_L g8739 ( 
.A(n_8326),
.Y(n_8739)
);

INVx1_ASAP7_75t_L g8740 ( 
.A(n_8491),
.Y(n_8740)
);

OR2x6_ASAP7_75t_L g8741 ( 
.A(n_8385),
.B(n_1540),
.Y(n_8741)
);

INVx4_ASAP7_75t_L g8742 ( 
.A(n_8514),
.Y(n_8742)
);

INVx1_ASAP7_75t_L g8743 ( 
.A(n_8293),
.Y(n_8743)
);

NAND2xp5_ASAP7_75t_L g8744 ( 
.A(n_8498),
.B(n_1541),
.Y(n_8744)
);

INVx3_ASAP7_75t_L g8745 ( 
.A(n_8259),
.Y(n_8745)
);

INVx1_ASAP7_75t_L g8746 ( 
.A(n_8270),
.Y(n_8746)
);

OAI21x1_ASAP7_75t_L g8747 ( 
.A1(n_8494),
.A2(n_414),
.B(n_415),
.Y(n_8747)
);

AND2x2_ASAP7_75t_L g8748 ( 
.A(n_8285),
.B(n_416),
.Y(n_8748)
);

INVx1_ASAP7_75t_L g8749 ( 
.A(n_8493),
.Y(n_8749)
);

INVx2_ASAP7_75t_L g8750 ( 
.A(n_8406),
.Y(n_8750)
);

NAND2xp5_ASAP7_75t_L g8751 ( 
.A(n_8266),
.B(n_1541),
.Y(n_8751)
);

AND2x2_ASAP7_75t_L g8752 ( 
.A(n_8481),
.B(n_416),
.Y(n_8752)
);

HB1xp67_ASAP7_75t_L g8753 ( 
.A(n_8357),
.Y(n_8753)
);

OAI21x1_ASAP7_75t_L g8754 ( 
.A1(n_8377),
.A2(n_8306),
.B(n_8267),
.Y(n_8754)
);

AND2x2_ASAP7_75t_L g8755 ( 
.A(n_8252),
.B(n_417),
.Y(n_8755)
);

INVx3_ASAP7_75t_L g8756 ( 
.A(n_8435),
.Y(n_8756)
);

INVx2_ASAP7_75t_L g8757 ( 
.A(n_8239),
.Y(n_8757)
);

AND2x2_ASAP7_75t_L g8758 ( 
.A(n_8492),
.B(n_417),
.Y(n_8758)
);

INVx1_ASAP7_75t_L g8759 ( 
.A(n_8360),
.Y(n_8759)
);

INVx2_ASAP7_75t_L g8760 ( 
.A(n_8432),
.Y(n_8760)
);

NAND2x1_ASAP7_75t_L g8761 ( 
.A(n_8380),
.B(n_417),
.Y(n_8761)
);

BUFx6f_ASAP7_75t_L g8762 ( 
.A(n_8484),
.Y(n_8762)
);

AOI22xp33_ASAP7_75t_L g8763 ( 
.A1(n_8344),
.A2(n_1544),
.B1(n_1545),
.B2(n_1543),
.Y(n_8763)
);

INVx1_ASAP7_75t_L g8764 ( 
.A(n_8416),
.Y(n_8764)
);

INVx1_ASAP7_75t_L g8765 ( 
.A(n_8508),
.Y(n_8765)
);

INVx1_ASAP7_75t_L g8766 ( 
.A(n_8383),
.Y(n_8766)
);

AOI221xp5_ASAP7_75t_L g8767 ( 
.A1(n_8532),
.A2(n_8296),
.B1(n_8500),
.B2(n_8421),
.C(n_8474),
.Y(n_8767)
);

INVx1_ASAP7_75t_L g8768 ( 
.A(n_8647),
.Y(n_8768)
);

INVx1_ASAP7_75t_SL g8769 ( 
.A(n_8680),
.Y(n_8769)
);

BUFx2_ASAP7_75t_L g8770 ( 
.A(n_8541),
.Y(n_8770)
);

INVx2_ASAP7_75t_L g8771 ( 
.A(n_8530),
.Y(n_8771)
);

AND2x2_ASAP7_75t_L g8772 ( 
.A(n_8585),
.B(n_8424),
.Y(n_8772)
);

INVx3_ASAP7_75t_L g8773 ( 
.A(n_8739),
.Y(n_8773)
);

AOI22xp33_ASAP7_75t_L g8774 ( 
.A1(n_8756),
.A2(n_8300),
.B1(n_8372),
.B2(n_8343),
.Y(n_8774)
);

OAI22xp5_ASAP7_75t_L g8775 ( 
.A1(n_8571),
.A2(n_8305),
.B1(n_8314),
.B2(n_8324),
.Y(n_8775)
);

AOI22xp33_ASAP7_75t_L g8776 ( 
.A1(n_8732),
.A2(n_8376),
.B1(n_8452),
.B2(n_8415),
.Y(n_8776)
);

OAI222xp33_ASAP7_75t_L g8777 ( 
.A1(n_8534),
.A2(n_8448),
.B1(n_8475),
.B2(n_8444),
.C1(n_8450),
.C2(n_8497),
.Y(n_8777)
);

NAND3xp33_ASAP7_75t_L g8778 ( 
.A(n_8715),
.B(n_8471),
.C(n_8316),
.Y(n_8778)
);

NAND2xp5_ASAP7_75t_L g8779 ( 
.A(n_8561),
.B(n_8429),
.Y(n_8779)
);

OAI22xp33_ASAP7_75t_L g8780 ( 
.A1(n_8542),
.A2(n_8410),
.B1(n_8302),
.B2(n_8319),
.Y(n_8780)
);

AOI22xp33_ASAP7_75t_L g8781 ( 
.A1(n_8762),
.A2(n_8327),
.B1(n_8323),
.B2(n_8321),
.Y(n_8781)
);

AOI222xp33_ASAP7_75t_L g8782 ( 
.A1(n_8762),
.A2(n_8417),
.B1(n_8442),
.B2(n_8404),
.C1(n_8392),
.C2(n_8506),
.Y(n_8782)
);

INVx1_ASAP7_75t_L g8783 ( 
.A(n_8648),
.Y(n_8783)
);

AND2x2_ASAP7_75t_L g8784 ( 
.A(n_8564),
.B(n_8479),
.Y(n_8784)
);

AOI22xp33_ASAP7_75t_L g8785 ( 
.A1(n_8766),
.A2(n_8394),
.B1(n_8352),
.B2(n_8329),
.Y(n_8785)
);

AOI21xp5_ASAP7_75t_L g8786 ( 
.A1(n_8590),
.A2(n_8489),
.B(n_8460),
.Y(n_8786)
);

AOI22xp33_ASAP7_75t_SL g8787 ( 
.A1(n_8527),
.A2(n_8636),
.B1(n_8570),
.B2(n_8737),
.Y(n_8787)
);

AND2x4_ASAP7_75t_L g8788 ( 
.A(n_8584),
.B(n_8463),
.Y(n_8788)
);

AOI22xp33_ASAP7_75t_L g8789 ( 
.A1(n_8741),
.A2(n_8381),
.B1(n_8458),
.B2(n_8454),
.Y(n_8789)
);

AOI22xp33_ASAP7_75t_SL g8790 ( 
.A1(n_8636),
.A2(n_8477),
.B1(n_8507),
.B2(n_1544),
.Y(n_8790)
);

AOI22xp33_ASAP7_75t_L g8791 ( 
.A1(n_8741),
.A2(n_1546),
.B1(n_1547),
.B2(n_1543),
.Y(n_8791)
);

AOI22xp5_ASAP7_75t_L g8792 ( 
.A1(n_8764),
.A2(n_420),
.B1(n_418),
.B2(n_419),
.Y(n_8792)
);

INVx4_ASAP7_75t_L g8793 ( 
.A(n_8556),
.Y(n_8793)
);

NOR2xp33_ASAP7_75t_L g8794 ( 
.A(n_8544),
.B(n_1547),
.Y(n_8794)
);

BUFx3_ASAP7_75t_L g8795 ( 
.A(n_8627),
.Y(n_8795)
);

AND2x2_ASAP7_75t_L g8796 ( 
.A(n_8580),
.B(n_418),
.Y(n_8796)
);

OAI22xp5_ASAP7_75t_L g8797 ( 
.A1(n_8621),
.A2(n_421),
.B1(n_419),
.B2(n_420),
.Y(n_8797)
);

NOR2xp33_ASAP7_75t_L g8798 ( 
.A(n_8742),
.B(n_1548),
.Y(n_8798)
);

AOI22xp33_ASAP7_75t_L g8799 ( 
.A1(n_8733),
.A2(n_1549),
.B1(n_1550),
.B2(n_1548),
.Y(n_8799)
);

BUFx4f_ASAP7_75t_SL g8800 ( 
.A(n_8591),
.Y(n_8800)
);

INVx2_ASAP7_75t_L g8801 ( 
.A(n_8593),
.Y(n_8801)
);

AND2x2_ASAP7_75t_L g8802 ( 
.A(n_8579),
.B(n_419),
.Y(n_8802)
);

OAI21x1_ASAP7_75t_L g8803 ( 
.A1(n_8717),
.A2(n_420),
.B(n_421),
.Y(n_8803)
);

OAI221xp5_ASAP7_75t_L g8804 ( 
.A1(n_8612),
.A2(n_423),
.B1(n_421),
.B2(n_422),
.C(n_424),
.Y(n_8804)
);

AOI21xp5_ASAP7_75t_L g8805 ( 
.A1(n_8697),
.A2(n_1552),
.B(n_1551),
.Y(n_8805)
);

AOI22xp33_ASAP7_75t_L g8806 ( 
.A1(n_8765),
.A2(n_1554),
.B1(n_1555),
.B2(n_1553),
.Y(n_8806)
);

OAI332xp33_ASAP7_75t_L g8807 ( 
.A1(n_8734),
.A2(n_427),
.A3(n_426),
.B1(n_424),
.B2(n_428),
.B3(n_422),
.C1(n_423),
.C2(n_425),
.Y(n_8807)
);

AOI21xp5_ASAP7_75t_L g8808 ( 
.A1(n_8583),
.A2(n_1554),
.B(n_1553),
.Y(n_8808)
);

OAI21x1_ASAP7_75t_L g8809 ( 
.A1(n_8671),
.A2(n_422),
.B(n_424),
.Y(n_8809)
);

CKINVDCx8_ASAP7_75t_R g8810 ( 
.A(n_8703),
.Y(n_8810)
);

AOI21xp5_ASAP7_75t_L g8811 ( 
.A1(n_8660),
.A2(n_1557),
.B(n_1556),
.Y(n_8811)
);

A2O1A1Ixp33_ASAP7_75t_L g8812 ( 
.A1(n_8602),
.A2(n_428),
.B(n_425),
.C(n_427),
.Y(n_8812)
);

NAND2xp5_ASAP7_75t_L g8813 ( 
.A(n_8655),
.B(n_1556),
.Y(n_8813)
);

AND2x2_ASAP7_75t_L g8814 ( 
.A(n_8666),
.B(n_425),
.Y(n_8814)
);

INVx1_ASAP7_75t_L g8815 ( 
.A(n_8640),
.Y(n_8815)
);

AOI22xp33_ASAP7_75t_L g8816 ( 
.A1(n_8722),
.A2(n_1558),
.B1(n_1559),
.B2(n_1557),
.Y(n_8816)
);

AO21x2_ASAP7_75t_L g8817 ( 
.A1(n_8650),
.A2(n_428),
.B(n_429),
.Y(n_8817)
);

INVx1_ASAP7_75t_L g8818 ( 
.A(n_8632),
.Y(n_8818)
);

INVx2_ASAP7_75t_L g8819 ( 
.A(n_8638),
.Y(n_8819)
);

AND2x2_ASAP7_75t_L g8820 ( 
.A(n_8678),
.B(n_429),
.Y(n_8820)
);

INVx1_ASAP7_75t_L g8821 ( 
.A(n_8634),
.Y(n_8821)
);

INVx1_ASAP7_75t_L g8822 ( 
.A(n_8637),
.Y(n_8822)
);

AOI22xp33_ASAP7_75t_SL g8823 ( 
.A1(n_8735),
.A2(n_1560),
.B1(n_1561),
.B2(n_1558),
.Y(n_8823)
);

AOI221xp5_ASAP7_75t_L g8824 ( 
.A1(n_8657),
.A2(n_431),
.B1(n_429),
.B2(n_430),
.C(n_432),
.Y(n_8824)
);

AOI22xp33_ASAP7_75t_L g8825 ( 
.A1(n_8760),
.A2(n_1562),
.B1(n_1563),
.B2(n_1561),
.Y(n_8825)
);

INVx1_ASAP7_75t_L g8826 ( 
.A(n_8639),
.Y(n_8826)
);

AOI22xp33_ASAP7_75t_L g8827 ( 
.A1(n_8745),
.A2(n_1563),
.B1(n_1564),
.B2(n_1562),
.Y(n_8827)
);

INVx1_ASAP7_75t_L g8828 ( 
.A(n_8529),
.Y(n_8828)
);

AOI222xp33_ASAP7_75t_L g8829 ( 
.A1(n_8670),
.A2(n_432),
.B1(n_434),
.B2(n_430),
.C1(n_431),
.C2(n_433),
.Y(n_8829)
);

AOI22xp33_ASAP7_75t_L g8830 ( 
.A1(n_8757),
.A2(n_1565),
.B1(n_1566),
.B2(n_1564),
.Y(n_8830)
);

OA21x2_ASAP7_75t_L g8831 ( 
.A1(n_8651),
.A2(n_433),
.B(n_434),
.Y(n_8831)
);

AOI22xp33_ASAP7_75t_L g8832 ( 
.A1(n_8749),
.A2(n_8599),
.B1(n_8542),
.B2(n_8750),
.Y(n_8832)
);

OAI22xp5_ASAP7_75t_L g8833 ( 
.A1(n_8661),
.A2(n_436),
.B1(n_433),
.B2(n_435),
.Y(n_8833)
);

INVx3_ASAP7_75t_L g8834 ( 
.A(n_8736),
.Y(n_8834)
);

INVx2_ASAP7_75t_L g8835 ( 
.A(n_8562),
.Y(n_8835)
);

AND2x2_ASAP7_75t_L g8836 ( 
.A(n_8553),
.B(n_437),
.Y(n_8836)
);

INVx1_ASAP7_75t_L g8837 ( 
.A(n_8545),
.Y(n_8837)
);

OAI22xp33_ASAP7_75t_L g8838 ( 
.A1(n_8625),
.A2(n_8586),
.B1(n_8728),
.B2(n_8746),
.Y(n_8838)
);

INVx1_ASAP7_75t_L g8839 ( 
.A(n_8547),
.Y(n_8839)
);

INVx1_ASAP7_75t_L g8840 ( 
.A(n_8548),
.Y(n_8840)
);

AOI22xp33_ASAP7_75t_L g8841 ( 
.A1(n_8753),
.A2(n_1566),
.B1(n_1567),
.B2(n_1565),
.Y(n_8841)
);

OAI21x1_ASAP7_75t_L g8842 ( 
.A1(n_8551),
.A2(n_438),
.B(n_439),
.Y(n_8842)
);

AO21x1_ASAP7_75t_L g8843 ( 
.A1(n_8726),
.A2(n_438),
.B(n_439),
.Y(n_8843)
);

AOI22xp33_ASAP7_75t_L g8844 ( 
.A1(n_8629),
.A2(n_1568),
.B1(n_1569),
.B2(n_1567),
.Y(n_8844)
);

OAI21xp33_ASAP7_75t_L g8845 ( 
.A1(n_8598),
.A2(n_8763),
.B(n_8714),
.Y(n_8845)
);

OAI21x1_ASAP7_75t_SL g8846 ( 
.A1(n_8528),
.A2(n_439),
.B(n_440),
.Y(n_8846)
);

AOI33xp33_ASAP7_75t_L g8847 ( 
.A1(n_8740),
.A2(n_442),
.A3(n_444),
.B1(n_440),
.B2(n_441),
.B3(n_443),
.Y(n_8847)
);

OAI22xp5_ASAP7_75t_L g8848 ( 
.A1(n_8633),
.A2(n_8759),
.B1(n_8730),
.B2(n_8743),
.Y(n_8848)
);

OAI221xp5_ASAP7_75t_L g8849 ( 
.A1(n_8751),
.A2(n_442),
.B1(n_440),
.B2(n_441),
.C(n_443),
.Y(n_8849)
);

BUFx3_ASAP7_75t_L g8850 ( 
.A(n_8615),
.Y(n_8850)
);

OAI33xp33_ASAP7_75t_L g8851 ( 
.A1(n_8744),
.A2(n_443),
.A3(n_445),
.B1(n_441),
.B2(n_442),
.B3(n_444),
.Y(n_8851)
);

OAI211xp5_ASAP7_75t_SL g8852 ( 
.A1(n_8669),
.A2(n_446),
.B(n_444),
.C(n_445),
.Y(n_8852)
);

AOI22xp33_ASAP7_75t_L g8853 ( 
.A1(n_8754),
.A2(n_8752),
.B1(n_8675),
.B2(n_8761),
.Y(n_8853)
);

AND2x2_ASAP7_75t_L g8854 ( 
.A(n_8557),
.B(n_446),
.Y(n_8854)
);

OAI21x1_ASAP7_75t_L g8855 ( 
.A1(n_8525),
.A2(n_446),
.B(n_447),
.Y(n_8855)
);

NAND2xp5_ASAP7_75t_L g8856 ( 
.A(n_8635),
.B(n_1568),
.Y(n_8856)
);

INVx1_ASAP7_75t_L g8857 ( 
.A(n_8552),
.Y(n_8857)
);

AOI22xp33_ASAP7_75t_L g8858 ( 
.A1(n_8719),
.A2(n_8755),
.B1(n_8683),
.B2(n_8533),
.Y(n_8858)
);

INVx3_ASAP7_75t_L g8859 ( 
.A(n_8699),
.Y(n_8859)
);

HB1xp67_ASAP7_75t_L g8860 ( 
.A(n_8531),
.Y(n_8860)
);

AOI22xp5_ASAP7_75t_L g8861 ( 
.A1(n_8573),
.A2(n_449),
.B1(n_447),
.B2(n_448),
.Y(n_8861)
);

OAI22xp5_ASAP7_75t_SL g8862 ( 
.A1(n_8679),
.A2(n_8677),
.B1(n_8574),
.B2(n_8729),
.Y(n_8862)
);

AOI221xp5_ASAP7_75t_L g8863 ( 
.A1(n_8700),
.A2(n_450),
.B1(n_448),
.B2(n_449),
.C(n_451),
.Y(n_8863)
);

AOI221xp5_ASAP7_75t_L g8864 ( 
.A1(n_8701),
.A2(n_451),
.B1(n_448),
.B2(n_449),
.C(n_452),
.Y(n_8864)
);

AOI221xp5_ASAP7_75t_L g8865 ( 
.A1(n_8758),
.A2(n_453),
.B1(n_451),
.B2(n_452),
.C(n_454),
.Y(n_8865)
);

INVx1_ASAP7_75t_SL g8866 ( 
.A(n_8607),
.Y(n_8866)
);

AOI22xp33_ASAP7_75t_L g8867 ( 
.A1(n_8748),
.A2(n_1570),
.B1(n_1571),
.B2(n_1569),
.Y(n_8867)
);

OR2x6_ASAP7_75t_L g8868 ( 
.A(n_8582),
.B(n_1571),
.Y(n_8868)
);

AOI22xp33_ASAP7_75t_L g8869 ( 
.A1(n_8702),
.A2(n_8692),
.B1(n_8724),
.B2(n_8688),
.Y(n_8869)
);

AND2x2_ASAP7_75t_L g8870 ( 
.A(n_8682),
.B(n_452),
.Y(n_8870)
);

AOI22xp33_ASAP7_75t_L g8871 ( 
.A1(n_8546),
.A2(n_1573),
.B1(n_1574),
.B2(n_1572),
.Y(n_8871)
);

OAI221xp5_ASAP7_75t_SL g8872 ( 
.A1(n_8595),
.A2(n_8690),
.B1(n_8673),
.B2(n_8725),
.C(n_8614),
.Y(n_8872)
);

INVx1_ASAP7_75t_L g8873 ( 
.A(n_8554),
.Y(n_8873)
);

AOI22xp33_ASAP7_75t_L g8874 ( 
.A1(n_8524),
.A2(n_1574),
.B1(n_1575),
.B2(n_1572),
.Y(n_8874)
);

OAI22xp5_ASAP7_75t_L g8875 ( 
.A1(n_8536),
.A2(n_455),
.B1(n_453),
.B2(n_454),
.Y(n_8875)
);

OAI22xp33_ASAP7_75t_L g8876 ( 
.A1(n_8563),
.A2(n_456),
.B1(n_453),
.B2(n_455),
.Y(n_8876)
);

OAI22xp33_ASAP7_75t_L g8877 ( 
.A1(n_8646),
.A2(n_459),
.B1(n_456),
.B2(n_457),
.Y(n_8877)
);

AOI22xp33_ASAP7_75t_L g8878 ( 
.A1(n_8684),
.A2(n_1577),
.B1(n_1578),
.B2(n_1575),
.Y(n_8878)
);

NAND3xp33_ASAP7_75t_L g8879 ( 
.A(n_8603),
.B(n_457),
.C(n_459),
.Y(n_8879)
);

AND2x2_ASAP7_75t_L g8880 ( 
.A(n_8581),
.B(n_457),
.Y(n_8880)
);

AOI22xp33_ASAP7_75t_L g8881 ( 
.A1(n_8747),
.A2(n_1579),
.B1(n_1580),
.B2(n_1578),
.Y(n_8881)
);

AND2x2_ASAP7_75t_L g8882 ( 
.A(n_8652),
.B(n_459),
.Y(n_8882)
);

OAI22xp5_ASAP7_75t_L g8883 ( 
.A1(n_8695),
.A2(n_462),
.B1(n_460),
.B2(n_461),
.Y(n_8883)
);

AOI22xp33_ASAP7_75t_L g8884 ( 
.A1(n_8672),
.A2(n_1580),
.B1(n_1581),
.B2(n_1579),
.Y(n_8884)
);

AOI22xp33_ASAP7_75t_L g8885 ( 
.A1(n_8685),
.A2(n_1583),
.B1(n_1584),
.B2(n_1582),
.Y(n_8885)
);

OAI22xp5_ASAP7_75t_L g8886 ( 
.A1(n_8721),
.A2(n_462),
.B1(n_460),
.B2(n_461),
.Y(n_8886)
);

CKINVDCx20_ASAP7_75t_R g8887 ( 
.A(n_8550),
.Y(n_8887)
);

AOI22xp33_ASAP7_75t_L g8888 ( 
.A1(n_8738),
.A2(n_1584),
.B1(n_1585),
.B2(n_1582),
.Y(n_8888)
);

INVx1_ASAP7_75t_L g8889 ( 
.A(n_8558),
.Y(n_8889)
);

INVx1_ASAP7_75t_L g8890 ( 
.A(n_8559),
.Y(n_8890)
);

AOI221xp5_ASAP7_75t_L g8891 ( 
.A1(n_8662),
.A2(n_464),
.B1(n_460),
.B2(n_463),
.C(n_465),
.Y(n_8891)
);

OAI221xp5_ASAP7_75t_L g8892 ( 
.A1(n_8549),
.A2(n_465),
.B1(n_463),
.B2(n_464),
.C(n_466),
.Y(n_8892)
);

INVx2_ASAP7_75t_L g8893 ( 
.A(n_8565),
.Y(n_8893)
);

OAI22xp5_ASAP7_75t_L g8894 ( 
.A1(n_8676),
.A2(n_465),
.B1(n_463),
.B2(n_464),
.Y(n_8894)
);

AND2x2_ASAP7_75t_L g8895 ( 
.A(n_8663),
.B(n_466),
.Y(n_8895)
);

AND2x2_ASAP7_75t_L g8896 ( 
.A(n_8665),
.B(n_466),
.Y(n_8896)
);

INVx1_ASAP7_75t_L g8897 ( 
.A(n_8560),
.Y(n_8897)
);

OAI22xp33_ASAP7_75t_L g8898 ( 
.A1(n_8727),
.A2(n_469),
.B1(n_467),
.B2(n_468),
.Y(n_8898)
);

OAI21x1_ASAP7_75t_L g8899 ( 
.A1(n_8577),
.A2(n_467),
.B(n_468),
.Y(n_8899)
);

AOI221xp5_ASAP7_75t_L g8900 ( 
.A1(n_8613),
.A2(n_469),
.B1(n_467),
.B2(n_468),
.C(n_470),
.Y(n_8900)
);

AOI22xp33_ASAP7_75t_L g8901 ( 
.A1(n_8696),
.A2(n_1586),
.B1(n_1587),
.B2(n_1585),
.Y(n_8901)
);

OAI22xp5_ASAP7_75t_L g8902 ( 
.A1(n_8707),
.A2(n_471),
.B1(n_469),
.B2(n_470),
.Y(n_8902)
);

AND2x4_ASAP7_75t_L g8903 ( 
.A(n_8687),
.B(n_1586),
.Y(n_8903)
);

OAI22xp5_ASAP7_75t_L g8904 ( 
.A1(n_8713),
.A2(n_8623),
.B1(n_8616),
.B2(n_8712),
.Y(n_8904)
);

AND2x2_ASAP7_75t_L g8905 ( 
.A(n_8711),
.B(n_470),
.Y(n_8905)
);

AOI22xp5_ASAP7_75t_L g8906 ( 
.A1(n_8704),
.A2(n_473),
.B1(n_471),
.B2(n_472),
.Y(n_8906)
);

OAI21xp5_ASAP7_75t_L g8907 ( 
.A1(n_8668),
.A2(n_471),
.B(n_472),
.Y(n_8907)
);

OR2x2_ASAP7_75t_L g8908 ( 
.A(n_8594),
.B(n_8537),
.Y(n_8908)
);

INVx3_ASAP7_75t_L g8909 ( 
.A(n_8538),
.Y(n_8909)
);

AND2x2_ASAP7_75t_L g8910 ( 
.A(n_8575),
.B(n_472),
.Y(n_8910)
);

INVx1_ASAP7_75t_L g8911 ( 
.A(n_8566),
.Y(n_8911)
);

AOI22xp33_ASAP7_75t_L g8912 ( 
.A1(n_8706),
.A2(n_1588),
.B1(n_1589),
.B2(n_1587),
.Y(n_8912)
);

AOI22xp33_ASAP7_75t_SL g8913 ( 
.A1(n_8628),
.A2(n_1589),
.B1(n_1590),
.B2(n_1588),
.Y(n_8913)
);

OAI22xp33_ASAP7_75t_L g8914 ( 
.A1(n_8658),
.A2(n_8572),
.B1(n_8694),
.B2(n_8689),
.Y(n_8914)
);

AOI21xp5_ASAP7_75t_L g8915 ( 
.A1(n_8656),
.A2(n_1593),
.B(n_1590),
.Y(n_8915)
);

AOI22xp33_ASAP7_75t_L g8916 ( 
.A1(n_8716),
.A2(n_1594),
.B1(n_1595),
.B2(n_1593),
.Y(n_8916)
);

INVx1_ASAP7_75t_L g8917 ( 
.A(n_8569),
.Y(n_8917)
);

BUFx3_ASAP7_75t_R g8918 ( 
.A(n_8674),
.Y(n_8918)
);

INVx1_ASAP7_75t_L g8919 ( 
.A(n_8567),
.Y(n_8919)
);

INVx1_ASAP7_75t_L g8920 ( 
.A(n_8568),
.Y(n_8920)
);

OAI21xp33_ASAP7_75t_L g8921 ( 
.A1(n_8731),
.A2(n_473),
.B(n_474),
.Y(n_8921)
);

BUFx12f_ASAP7_75t_L g8922 ( 
.A(n_8708),
.Y(n_8922)
);

INVx2_ASAP7_75t_SL g8923 ( 
.A(n_8578),
.Y(n_8923)
);

AOI22xp33_ASAP7_75t_L g8924 ( 
.A1(n_8718),
.A2(n_8710),
.B1(n_8691),
.B2(n_8681),
.Y(n_8924)
);

OAI22xp5_ASAP7_75t_L g8925 ( 
.A1(n_8723),
.A2(n_475),
.B1(n_473),
.B2(n_474),
.Y(n_8925)
);

INVx1_ASAP7_75t_SL g8926 ( 
.A(n_8644),
.Y(n_8926)
);

NOR2x1_ASAP7_75t_R g8927 ( 
.A(n_8610),
.B(n_474),
.Y(n_8927)
);

OAI221xp5_ASAP7_75t_SL g8928 ( 
.A1(n_8605),
.A2(n_477),
.B1(n_475),
.B2(n_476),
.C(n_478),
.Y(n_8928)
);

INVx2_ASAP7_75t_L g8929 ( 
.A(n_8576),
.Y(n_8929)
);

INVx2_ASAP7_75t_L g8930 ( 
.A(n_8622),
.Y(n_8930)
);

AOI22xp5_ASAP7_75t_L g8931 ( 
.A1(n_8543),
.A2(n_479),
.B1(n_476),
.B2(n_477),
.Y(n_8931)
);

OR2x2_ASAP7_75t_L g8932 ( 
.A(n_8523),
.B(n_476),
.Y(n_8932)
);

INVx1_ASAP7_75t_L g8933 ( 
.A(n_8601),
.Y(n_8933)
);

AOI221xp5_ASAP7_75t_L g8934 ( 
.A1(n_8664),
.A2(n_8596),
.B1(n_8526),
.B2(n_8659),
.C(n_8649),
.Y(n_8934)
);

NAND2xp5_ASAP7_75t_L g8935 ( 
.A(n_8654),
.B(n_1596),
.Y(n_8935)
);

AND2x2_ASAP7_75t_L g8936 ( 
.A(n_8698),
.B(n_479),
.Y(n_8936)
);

AND2x4_ASAP7_75t_L g8937 ( 
.A(n_8705),
.B(n_1598),
.Y(n_8937)
);

INVx4_ASAP7_75t_L g8938 ( 
.A(n_8587),
.Y(n_8938)
);

OAI22xp33_ASAP7_75t_L g8939 ( 
.A1(n_8709),
.A2(n_481),
.B1(n_479),
.B2(n_480),
.Y(n_8939)
);

AND2x2_ASAP7_75t_L g8940 ( 
.A(n_8624),
.B(n_480),
.Y(n_8940)
);

OAI21xp5_ASAP7_75t_L g8941 ( 
.A1(n_8667),
.A2(n_480),
.B(n_481),
.Y(n_8941)
);

OAI221xp5_ASAP7_75t_L g8942 ( 
.A1(n_8686),
.A2(n_483),
.B1(n_481),
.B2(n_482),
.C(n_484),
.Y(n_8942)
);

OAI21x1_ASAP7_75t_L g8943 ( 
.A1(n_8642),
.A2(n_482),
.B(n_483),
.Y(n_8943)
);

AOI22xp33_ASAP7_75t_L g8944 ( 
.A1(n_8535),
.A2(n_1600),
.B1(n_1601),
.B2(n_1599),
.Y(n_8944)
);

AOI221xp5_ASAP7_75t_L g8945 ( 
.A1(n_8626),
.A2(n_484),
.B1(n_482),
.B2(n_483),
.C(n_485),
.Y(n_8945)
);

AOI222xp33_ASAP7_75t_L g8946 ( 
.A1(n_8645),
.A2(n_486),
.B1(n_489),
.B2(n_484),
.C1(n_485),
.C2(n_488),
.Y(n_8946)
);

OAI21x1_ASAP7_75t_L g8947 ( 
.A1(n_8643),
.A2(n_485),
.B(n_486),
.Y(n_8947)
);

INVx1_ASAP7_75t_L g8948 ( 
.A(n_8604),
.Y(n_8948)
);

CKINVDCx5p33_ASAP7_75t_R g8949 ( 
.A(n_8587),
.Y(n_8949)
);

AOI22xp33_ASAP7_75t_L g8950 ( 
.A1(n_8631),
.A2(n_1600),
.B1(n_1601),
.B2(n_1599),
.Y(n_8950)
);

INVx1_ASAP7_75t_L g8951 ( 
.A(n_8609),
.Y(n_8951)
);

AOI22xp33_ASAP7_75t_L g8952 ( 
.A1(n_8600),
.A2(n_1603),
.B1(n_1605),
.B2(n_1602),
.Y(n_8952)
);

OAI22xp33_ASAP7_75t_L g8953 ( 
.A1(n_8630),
.A2(n_489),
.B1(n_486),
.B2(n_488),
.Y(n_8953)
);

OA21x2_ASAP7_75t_L g8954 ( 
.A1(n_8618),
.A2(n_490),
.B(n_489),
.Y(n_8954)
);

INVxp67_ASAP7_75t_L g8955 ( 
.A(n_8693),
.Y(n_8955)
);

AND2x2_ASAP7_75t_L g8956 ( 
.A(n_8589),
.B(n_488),
.Y(n_8956)
);

OAI22xp5_ASAP7_75t_L g8957 ( 
.A1(n_8641),
.A2(n_492),
.B1(n_490),
.B2(n_491),
.Y(n_8957)
);

NAND2xp33_ASAP7_75t_R g8958 ( 
.A(n_8720),
.B(n_8597),
.Y(n_8958)
);

AOI22xp33_ASAP7_75t_SL g8959 ( 
.A1(n_8653),
.A2(n_1605),
.B1(n_1607),
.B2(n_1603),
.Y(n_8959)
);

OAI22xp5_ASAP7_75t_L g8960 ( 
.A1(n_8641),
.A2(n_493),
.B1(n_491),
.B2(n_492),
.Y(n_8960)
);

AOI21xp5_ASAP7_75t_L g8961 ( 
.A1(n_8539),
.A2(n_1609),
.B(n_1607),
.Y(n_8961)
);

AOI22xp33_ASAP7_75t_L g8962 ( 
.A1(n_8606),
.A2(n_1610),
.B1(n_1611),
.B2(n_1609),
.Y(n_8962)
);

OAI22xp33_ASAP7_75t_SL g8963 ( 
.A1(n_8608),
.A2(n_493),
.B1(n_491),
.B2(n_492),
.Y(n_8963)
);

OAI22xp5_ASAP7_75t_L g8964 ( 
.A1(n_8540),
.A2(n_495),
.B1(n_493),
.B2(n_494),
.Y(n_8964)
);

AOI22xp33_ASAP7_75t_L g8965 ( 
.A1(n_8620),
.A2(n_1611),
.B1(n_1612),
.B2(n_1610),
.Y(n_8965)
);

BUFx6f_ASAP7_75t_L g8966 ( 
.A(n_8588),
.Y(n_8966)
);

NAND3xp33_ASAP7_75t_L g8967 ( 
.A(n_8611),
.B(n_494),
.C(n_496),
.Y(n_8967)
);

INVx1_ASAP7_75t_L g8968 ( 
.A(n_8555),
.Y(n_8968)
);

AOI22xp5_ASAP7_75t_L g8969 ( 
.A1(n_8617),
.A2(n_497),
.B1(n_494),
.B2(n_496),
.Y(n_8969)
);

INVx1_ASAP7_75t_L g8970 ( 
.A(n_8592),
.Y(n_8970)
);

AOI22xp33_ASAP7_75t_L g8971 ( 
.A1(n_8619),
.A2(n_1613),
.B1(n_1614),
.B2(n_1612),
.Y(n_8971)
);

OAI22xp33_ASAP7_75t_L g8972 ( 
.A1(n_8532),
.A2(n_499),
.B1(n_497),
.B2(n_498),
.Y(n_8972)
);

AND2x2_ASAP7_75t_L g8973 ( 
.A(n_8541),
.B(n_497),
.Y(n_8973)
);

AOI22xp33_ASAP7_75t_L g8974 ( 
.A1(n_8532),
.A2(n_1614),
.B1(n_1615),
.B2(n_1613),
.Y(n_8974)
);

BUFx2_ASAP7_75t_L g8975 ( 
.A(n_8541),
.Y(n_8975)
);

INVx1_ASAP7_75t_L g8976 ( 
.A(n_8647),
.Y(n_8976)
);

OAI221xp5_ASAP7_75t_L g8977 ( 
.A1(n_8532),
.A2(n_500),
.B1(n_498),
.B2(n_499),
.C(n_501),
.Y(n_8977)
);

HB1xp67_ASAP7_75t_L g8978 ( 
.A(n_8531),
.Y(n_8978)
);

INVx1_ASAP7_75t_L g8979 ( 
.A(n_8647),
.Y(n_8979)
);

AOI22xp33_ASAP7_75t_L g8980 ( 
.A1(n_8532),
.A2(n_1616),
.B1(n_1617),
.B2(n_1615),
.Y(n_8980)
);

AOI22xp33_ASAP7_75t_L g8981 ( 
.A1(n_8532),
.A2(n_1618),
.B1(n_1619),
.B2(n_1616),
.Y(n_8981)
);

AOI22xp33_ASAP7_75t_L g8982 ( 
.A1(n_8532),
.A2(n_1620),
.B1(n_1621),
.B2(n_1618),
.Y(n_8982)
);

AND2x2_ASAP7_75t_L g8983 ( 
.A(n_8541),
.B(n_501),
.Y(n_8983)
);

AND2x2_ASAP7_75t_L g8984 ( 
.A(n_8541),
.B(n_501),
.Y(n_8984)
);

INVx1_ASAP7_75t_L g8985 ( 
.A(n_8647),
.Y(n_8985)
);

OAI22xp5_ASAP7_75t_L g8986 ( 
.A1(n_8571),
.A2(n_504),
.B1(n_502),
.B2(n_503),
.Y(n_8986)
);

NAND3xp33_ASAP7_75t_L g8987 ( 
.A(n_8532),
.B(n_502),
.C(n_505),
.Y(n_8987)
);

HB1xp67_ASAP7_75t_L g8988 ( 
.A(n_8531),
.Y(n_8988)
);

INVx1_ASAP7_75t_L g8989 ( 
.A(n_8647),
.Y(n_8989)
);

OAI211xp5_ASAP7_75t_L g8990 ( 
.A1(n_8532),
.A2(n_506),
.B(n_502),
.C(n_505),
.Y(n_8990)
);

OAI222xp33_ASAP7_75t_L g8991 ( 
.A1(n_8532),
.A2(n_507),
.B1(n_509),
.B2(n_505),
.C1(n_506),
.C2(n_508),
.Y(n_8991)
);

AOI33xp33_ASAP7_75t_L g8992 ( 
.A1(n_8571),
.A2(n_509),
.A3(n_511),
.B1(n_506),
.B2(n_507),
.B3(n_510),
.Y(n_8992)
);

OAI22xp5_ASAP7_75t_L g8993 ( 
.A1(n_8571),
.A2(n_510),
.B1(n_507),
.B2(n_509),
.Y(n_8993)
);

AOI22xp33_ASAP7_75t_SL g8994 ( 
.A1(n_8532),
.A2(n_1621),
.B1(n_1622),
.B2(n_1620),
.Y(n_8994)
);

AOI22xp33_ASAP7_75t_L g8995 ( 
.A1(n_8532),
.A2(n_1624),
.B1(n_1625),
.B2(n_1623),
.Y(n_8995)
);

OAI211xp5_ASAP7_75t_SL g8996 ( 
.A1(n_8532),
.A2(n_512),
.B(n_510),
.C(n_511),
.Y(n_8996)
);

CKINVDCx6p67_ASAP7_75t_R g8997 ( 
.A(n_8680),
.Y(n_8997)
);

OAI22xp5_ASAP7_75t_L g8998 ( 
.A1(n_8571),
.A2(n_513),
.B1(n_511),
.B2(n_512),
.Y(n_8998)
);

BUFx3_ASAP7_75t_L g8999 ( 
.A(n_8556),
.Y(n_8999)
);

AOI22xp33_ASAP7_75t_L g9000 ( 
.A1(n_8532),
.A2(n_1625),
.B1(n_1626),
.B2(n_1624),
.Y(n_9000)
);

NAND2xp5_ASAP7_75t_L g9001 ( 
.A(n_8561),
.B(n_1627),
.Y(n_9001)
);

AOI22xp33_ASAP7_75t_SL g9002 ( 
.A1(n_8532),
.A2(n_1628),
.B1(n_1630),
.B2(n_1627),
.Y(n_9002)
);

OAI22xp33_ASAP7_75t_L g9003 ( 
.A1(n_8532),
.A2(n_515),
.B1(n_512),
.B2(n_513),
.Y(n_9003)
);

OR2x2_ASAP7_75t_L g9004 ( 
.A(n_8594),
.B(n_515),
.Y(n_9004)
);

OAI22xp33_ASAP7_75t_L g9005 ( 
.A1(n_8532),
.A2(n_517),
.B1(n_515),
.B2(n_516),
.Y(n_9005)
);

INVx1_ASAP7_75t_L g9006 ( 
.A(n_8647),
.Y(n_9006)
);

AOI221xp5_ASAP7_75t_L g9007 ( 
.A1(n_8532),
.A2(n_518),
.B1(n_516),
.B2(n_517),
.C(n_519),
.Y(n_9007)
);

NOR2xp33_ASAP7_75t_L g9008 ( 
.A(n_8739),
.B(n_2252),
.Y(n_9008)
);

INVx1_ASAP7_75t_L g9009 ( 
.A(n_8647),
.Y(n_9009)
);

AOI221xp5_ASAP7_75t_L g9010 ( 
.A1(n_8532),
.A2(n_518),
.B1(n_516),
.B2(n_517),
.C(n_519),
.Y(n_9010)
);

OAI22xp5_ASAP7_75t_L g9011 ( 
.A1(n_8571),
.A2(n_520),
.B1(n_518),
.B2(n_519),
.Y(n_9011)
);

AOI22xp33_ASAP7_75t_L g9012 ( 
.A1(n_8532),
.A2(n_1630),
.B1(n_1631),
.B2(n_1628),
.Y(n_9012)
);

AOI22xp33_ASAP7_75t_L g9013 ( 
.A1(n_8532),
.A2(n_1632),
.B1(n_1633),
.B2(n_1631),
.Y(n_9013)
);

AOI22xp5_ASAP7_75t_L g9014 ( 
.A1(n_8534),
.A2(n_522),
.B1(n_520),
.B2(n_521),
.Y(n_9014)
);

HB1xp67_ASAP7_75t_L g9015 ( 
.A(n_8531),
.Y(n_9015)
);

INVx3_ASAP7_75t_L g9016 ( 
.A(n_8739),
.Y(n_9016)
);

AO21x2_ASAP7_75t_L g9017 ( 
.A1(n_8671),
.A2(n_521),
.B(n_522),
.Y(n_9017)
);

AND2x2_ASAP7_75t_L g9018 ( 
.A(n_8541),
.B(n_521),
.Y(n_9018)
);

INVx1_ASAP7_75t_L g9019 ( 
.A(n_8647),
.Y(n_9019)
);

NAND3xp33_ASAP7_75t_L g9020 ( 
.A(n_8532),
.B(n_523),
.C(n_524),
.Y(n_9020)
);

AOI22xp33_ASAP7_75t_SL g9021 ( 
.A1(n_8532),
.A2(n_1635),
.B1(n_1636),
.B2(n_1634),
.Y(n_9021)
);

BUFx4f_ASAP7_75t_SL g9022 ( 
.A(n_8591),
.Y(n_9022)
);

AOI22xp5_ASAP7_75t_L g9023 ( 
.A1(n_8534),
.A2(n_525),
.B1(n_523),
.B2(n_524),
.Y(n_9023)
);

AND2x4_ASAP7_75t_L g9024 ( 
.A(n_8541),
.B(n_1634),
.Y(n_9024)
);

INVx1_ASAP7_75t_SL g9025 ( 
.A(n_8680),
.Y(n_9025)
);

OAI221xp5_ASAP7_75t_L g9026 ( 
.A1(n_8532),
.A2(n_525),
.B1(n_523),
.B2(n_524),
.C(n_526),
.Y(n_9026)
);

BUFx12f_ASAP7_75t_L g9027 ( 
.A(n_8680),
.Y(n_9027)
);

OAI22xp33_ASAP7_75t_L g9028 ( 
.A1(n_8532),
.A2(n_527),
.B1(n_525),
.B2(n_526),
.Y(n_9028)
);

BUFx12f_ASAP7_75t_L g9029 ( 
.A(n_8680),
.Y(n_9029)
);

OAI22xp33_ASAP7_75t_L g9030 ( 
.A1(n_8532),
.A2(n_529),
.B1(n_527),
.B2(n_528),
.Y(n_9030)
);

OR2x2_ASAP7_75t_L g9031 ( 
.A(n_8594),
.B(n_528),
.Y(n_9031)
);

HB1xp67_ASAP7_75t_L g9032 ( 
.A(n_8831),
.Y(n_9032)
);

AOI22xp33_ASAP7_75t_SL g9033 ( 
.A1(n_8862),
.A2(n_536),
.B1(n_544),
.B2(n_528),
.Y(n_9033)
);

HB1xp67_ASAP7_75t_L g9034 ( 
.A(n_8831),
.Y(n_9034)
);

INVx1_ASAP7_75t_L g9035 ( 
.A(n_8768),
.Y(n_9035)
);

AO21x2_ASAP7_75t_L g9036 ( 
.A1(n_9001),
.A2(n_529),
.B(n_530),
.Y(n_9036)
);

BUFx3_ASAP7_75t_L g9037 ( 
.A(n_9027),
.Y(n_9037)
);

INVx1_ASAP7_75t_L g9038 ( 
.A(n_8783),
.Y(n_9038)
);

INVx3_ASAP7_75t_L g9039 ( 
.A(n_8810),
.Y(n_9039)
);

BUFx2_ASAP7_75t_L g9040 ( 
.A(n_8770),
.Y(n_9040)
);

AND2x2_ASAP7_75t_L g9041 ( 
.A(n_8975),
.B(n_530),
.Y(n_9041)
);

INVx1_ASAP7_75t_L g9042 ( 
.A(n_8815),
.Y(n_9042)
);

AND2x2_ASAP7_75t_SL g9043 ( 
.A(n_8992),
.B(n_530),
.Y(n_9043)
);

INVx3_ASAP7_75t_L g9044 ( 
.A(n_9029),
.Y(n_9044)
);

AND2x4_ASAP7_75t_L g9045 ( 
.A(n_8773),
.B(n_531),
.Y(n_9045)
);

AND2x4_ASAP7_75t_L g9046 ( 
.A(n_9016),
.B(n_532),
.Y(n_9046)
);

HB1xp67_ASAP7_75t_L g9047 ( 
.A(n_8954),
.Y(n_9047)
);

INVx2_ASAP7_75t_L g9048 ( 
.A(n_8834),
.Y(n_9048)
);

OAI221xp5_ASAP7_75t_L g9049 ( 
.A1(n_8787),
.A2(n_534),
.B1(n_532),
.B2(n_533),
.C(n_535),
.Y(n_9049)
);

AND2x2_ASAP7_75t_L g9050 ( 
.A(n_8866),
.B(n_533),
.Y(n_9050)
);

AND2x2_ASAP7_75t_L g9051 ( 
.A(n_8772),
.B(n_8801),
.Y(n_9051)
);

INVx2_ASAP7_75t_L g9052 ( 
.A(n_8771),
.Y(n_9052)
);

INVx1_ASAP7_75t_L g9053 ( 
.A(n_8818),
.Y(n_9053)
);

NAND2xp5_ASAP7_75t_L g9054 ( 
.A(n_8934),
.B(n_1635),
.Y(n_9054)
);

OR2x2_ASAP7_75t_L g9055 ( 
.A(n_8908),
.B(n_534),
.Y(n_9055)
);

NAND2xp5_ASAP7_75t_L g9056 ( 
.A(n_8858),
.B(n_1636),
.Y(n_9056)
);

NOR2xp33_ASAP7_75t_L g9057 ( 
.A(n_8997),
.B(n_1637),
.Y(n_9057)
);

INVx1_ASAP7_75t_L g9058 ( 
.A(n_8821),
.Y(n_9058)
);

INVx2_ASAP7_75t_L g9059 ( 
.A(n_8835),
.Y(n_9059)
);

INVx2_ASAP7_75t_L g9060 ( 
.A(n_8893),
.Y(n_9060)
);

INVx2_ASAP7_75t_L g9061 ( 
.A(n_8929),
.Y(n_9061)
);

INVx1_ASAP7_75t_L g9062 ( 
.A(n_8822),
.Y(n_9062)
);

BUFx2_ASAP7_75t_L g9063 ( 
.A(n_8793),
.Y(n_9063)
);

INVx1_ASAP7_75t_L g9064 ( 
.A(n_8826),
.Y(n_9064)
);

AND2x2_ASAP7_75t_L g9065 ( 
.A(n_8784),
.B(n_534),
.Y(n_9065)
);

AND2x2_ASAP7_75t_L g9066 ( 
.A(n_8926),
.B(n_8859),
.Y(n_9066)
);

INVx1_ASAP7_75t_L g9067 ( 
.A(n_8976),
.Y(n_9067)
);

INVx1_ASAP7_75t_L g9068 ( 
.A(n_8979),
.Y(n_9068)
);

AND2x2_ASAP7_75t_L g9069 ( 
.A(n_8860),
.B(n_535),
.Y(n_9069)
);

INVx1_ASAP7_75t_L g9070 ( 
.A(n_8985),
.Y(n_9070)
);

AND2x2_ASAP7_75t_L g9071 ( 
.A(n_8978),
.B(n_535),
.Y(n_9071)
);

INVx2_ASAP7_75t_L g9072 ( 
.A(n_8930),
.Y(n_9072)
);

INVx2_ASAP7_75t_L g9073 ( 
.A(n_8819),
.Y(n_9073)
);

AND2x2_ASAP7_75t_L g9074 ( 
.A(n_8988),
.B(n_536),
.Y(n_9074)
);

INVx2_ASAP7_75t_L g9075 ( 
.A(n_8966),
.Y(n_9075)
);

AOI22xp33_ASAP7_75t_L g9076 ( 
.A1(n_8845),
.A2(n_1639),
.B1(n_1640),
.B2(n_1637),
.Y(n_9076)
);

INVx1_ASAP7_75t_L g9077 ( 
.A(n_8989),
.Y(n_9077)
);

INVx1_ASAP7_75t_L g9078 ( 
.A(n_9006),
.Y(n_9078)
);

BUFx3_ASAP7_75t_L g9079 ( 
.A(n_8887),
.Y(n_9079)
);

OR2x2_ASAP7_75t_L g9080 ( 
.A(n_8869),
.B(n_536),
.Y(n_9080)
);

AND2x2_ASAP7_75t_L g9081 ( 
.A(n_9015),
.B(n_537),
.Y(n_9081)
);

HB1xp67_ASAP7_75t_L g9082 ( 
.A(n_8954),
.Y(n_9082)
);

NAND2xp5_ASAP7_75t_L g9083 ( 
.A(n_8914),
.B(n_1640),
.Y(n_9083)
);

INVx3_ASAP7_75t_L g9084 ( 
.A(n_8999),
.Y(n_9084)
);

INVx3_ASAP7_75t_L g9085 ( 
.A(n_8938),
.Y(n_9085)
);

NOR2xp33_ASAP7_75t_L g9086 ( 
.A(n_8769),
.B(n_1641),
.Y(n_9086)
);

INVx1_ASAP7_75t_L g9087 ( 
.A(n_9009),
.Y(n_9087)
);

INVx2_ASAP7_75t_L g9088 ( 
.A(n_8966),
.Y(n_9088)
);

AND2x2_ASAP7_75t_L g9089 ( 
.A(n_8955),
.B(n_537),
.Y(n_9089)
);

INVx1_ASAP7_75t_L g9090 ( 
.A(n_9019),
.Y(n_9090)
);

INVx3_ASAP7_75t_L g9091 ( 
.A(n_8909),
.Y(n_9091)
);

AO21x2_ASAP7_75t_L g9092 ( 
.A1(n_8876),
.A2(n_537),
.B(n_538),
.Y(n_9092)
);

INVx2_ASAP7_75t_L g9093 ( 
.A(n_8970),
.Y(n_9093)
);

AND2x2_ASAP7_75t_L g9094 ( 
.A(n_8923),
.B(n_539),
.Y(n_9094)
);

OR2x2_ASAP7_75t_SL g9095 ( 
.A(n_8987),
.B(n_539),
.Y(n_9095)
);

INVx1_ASAP7_75t_L g9096 ( 
.A(n_8828),
.Y(n_9096)
);

AND2x2_ASAP7_75t_L g9097 ( 
.A(n_8924),
.B(n_539),
.Y(n_9097)
);

INVx1_ASAP7_75t_L g9098 ( 
.A(n_8837),
.Y(n_9098)
);

HB1xp67_ASAP7_75t_L g9099 ( 
.A(n_8842),
.Y(n_9099)
);

AND2x2_ASAP7_75t_L g9100 ( 
.A(n_8904),
.B(n_540),
.Y(n_9100)
);

AND2x2_ASAP7_75t_L g9101 ( 
.A(n_8968),
.B(n_540),
.Y(n_9101)
);

INVx2_ASAP7_75t_L g9102 ( 
.A(n_8919),
.Y(n_9102)
);

INVx2_ASAP7_75t_L g9103 ( 
.A(n_8920),
.Y(n_9103)
);

INVx1_ASAP7_75t_L g9104 ( 
.A(n_8839),
.Y(n_9104)
);

BUFx2_ASAP7_75t_L g9105 ( 
.A(n_8922),
.Y(n_9105)
);

OR2x2_ASAP7_75t_L g9106 ( 
.A(n_8779),
.B(n_540),
.Y(n_9106)
);

INVx1_ASAP7_75t_L g9107 ( 
.A(n_8840),
.Y(n_9107)
);

INVx2_ASAP7_75t_SL g9108 ( 
.A(n_9025),
.Y(n_9108)
);

AND2x2_ASAP7_75t_L g9109 ( 
.A(n_8820),
.B(n_8853),
.Y(n_9109)
);

NAND2x1_ASAP7_75t_L g9110 ( 
.A(n_8857),
.B(n_541),
.Y(n_9110)
);

INVx2_ASAP7_75t_L g9111 ( 
.A(n_8873),
.Y(n_9111)
);

OR2x2_ASAP7_75t_L g9112 ( 
.A(n_8932),
.B(n_542),
.Y(n_9112)
);

INVx1_ASAP7_75t_L g9113 ( 
.A(n_8889),
.Y(n_9113)
);

AND2x2_ASAP7_75t_L g9114 ( 
.A(n_8836),
.B(n_542),
.Y(n_9114)
);

INVx2_ASAP7_75t_L g9115 ( 
.A(n_8890),
.Y(n_9115)
);

AND2x4_ASAP7_75t_L g9116 ( 
.A(n_8850),
.B(n_542),
.Y(n_9116)
);

NAND2xp5_ASAP7_75t_L g9117 ( 
.A(n_8813),
.B(n_1641),
.Y(n_9117)
);

AND2x2_ASAP7_75t_L g9118 ( 
.A(n_8854),
.B(n_543),
.Y(n_9118)
);

NAND2xp5_ASAP7_75t_L g9119 ( 
.A(n_8856),
.B(n_1643),
.Y(n_9119)
);

OA21x2_ASAP7_75t_L g9120 ( 
.A1(n_8855),
.A2(n_543),
.B(n_544),
.Y(n_9120)
);

OR2x2_ASAP7_75t_L g9121 ( 
.A(n_9004),
.B(n_9031),
.Y(n_9121)
);

AND2x2_ASAP7_75t_L g9122 ( 
.A(n_8788),
.B(n_544),
.Y(n_9122)
);

INVx1_ASAP7_75t_L g9123 ( 
.A(n_8897),
.Y(n_9123)
);

AOI22xp33_ASAP7_75t_L g9124 ( 
.A1(n_8767),
.A2(n_1644),
.B1(n_1645),
.B2(n_1643),
.Y(n_9124)
);

AND2x4_ASAP7_75t_L g9125 ( 
.A(n_8795),
.B(n_8882),
.Y(n_9125)
);

INVx1_ASAP7_75t_L g9126 ( 
.A(n_8911),
.Y(n_9126)
);

BUFx3_ASAP7_75t_L g9127 ( 
.A(n_8800),
.Y(n_9127)
);

NAND2xp5_ASAP7_75t_L g9128 ( 
.A(n_8917),
.B(n_1644),
.Y(n_9128)
);

INVx3_ASAP7_75t_L g9129 ( 
.A(n_9022),
.Y(n_9129)
);

NOR2x1_ASAP7_75t_SL g9130 ( 
.A(n_8868),
.B(n_545),
.Y(n_9130)
);

OR2x2_ASAP7_75t_L g9131 ( 
.A(n_8933),
.B(n_545),
.Y(n_9131)
);

INVx2_ASAP7_75t_L g9132 ( 
.A(n_8948),
.Y(n_9132)
);

AND2x2_ASAP7_75t_L g9133 ( 
.A(n_8951),
.B(n_545),
.Y(n_9133)
);

BUFx2_ASAP7_75t_L g9134 ( 
.A(n_9024),
.Y(n_9134)
);

AND2x2_ASAP7_75t_L g9135 ( 
.A(n_8973),
.B(n_546),
.Y(n_9135)
);

NAND2xp5_ASAP7_75t_L g9136 ( 
.A(n_8940),
.B(n_1646),
.Y(n_9136)
);

INVx2_ASAP7_75t_L g9137 ( 
.A(n_8956),
.Y(n_9137)
);

INVx4_ASAP7_75t_L g9138 ( 
.A(n_8949),
.Y(n_9138)
);

HB1xp67_ASAP7_75t_L g9139 ( 
.A(n_8958),
.Y(n_9139)
);

AOI22xp33_ASAP7_75t_L g9140 ( 
.A1(n_8775),
.A2(n_1647),
.B1(n_1648),
.B2(n_1646),
.Y(n_9140)
);

BUFx3_ASAP7_75t_L g9141 ( 
.A(n_8910),
.Y(n_9141)
);

BUFx3_ASAP7_75t_L g9142 ( 
.A(n_8870),
.Y(n_9142)
);

BUFx2_ASAP7_75t_L g9143 ( 
.A(n_8983),
.Y(n_9143)
);

INVxp67_ASAP7_75t_L g9144 ( 
.A(n_8927),
.Y(n_9144)
);

INVx1_ASAP7_75t_L g9145 ( 
.A(n_8935),
.Y(n_9145)
);

INVx2_ASAP7_75t_L g9146 ( 
.A(n_8895),
.Y(n_9146)
);

AND2x2_ASAP7_75t_L g9147 ( 
.A(n_8984),
.B(n_9018),
.Y(n_9147)
);

INVx1_ASAP7_75t_L g9148 ( 
.A(n_8817),
.Y(n_9148)
);

INVx2_ASAP7_75t_L g9149 ( 
.A(n_8809),
.Y(n_9149)
);

INVx1_ASAP7_75t_L g9150 ( 
.A(n_9017),
.Y(n_9150)
);

INVx1_ASAP7_75t_L g9151 ( 
.A(n_8814),
.Y(n_9151)
);

NAND2xp5_ASAP7_75t_L g9152 ( 
.A(n_8832),
.B(n_1648),
.Y(n_9152)
);

INVx3_ASAP7_75t_L g9153 ( 
.A(n_8903),
.Y(n_9153)
);

INVx2_ASAP7_75t_L g9154 ( 
.A(n_8936),
.Y(n_9154)
);

INVx2_ASAP7_75t_L g9155 ( 
.A(n_8802),
.Y(n_9155)
);

BUFx2_ASAP7_75t_L g9156 ( 
.A(n_8868),
.Y(n_9156)
);

INVx1_ASAP7_75t_L g9157 ( 
.A(n_8880),
.Y(n_9157)
);

INVx1_ASAP7_75t_L g9158 ( 
.A(n_8803),
.Y(n_9158)
);

INVx3_ASAP7_75t_L g9159 ( 
.A(n_8937),
.Y(n_9159)
);

AND2x2_ASAP7_75t_L g9160 ( 
.A(n_8796),
.B(n_547),
.Y(n_9160)
);

AND2x2_ASAP7_75t_L g9161 ( 
.A(n_8905),
.B(n_548),
.Y(n_9161)
);

AND2x2_ASAP7_75t_L g9162 ( 
.A(n_8896),
.B(n_548),
.Y(n_9162)
);

AND2x2_ASAP7_75t_L g9163 ( 
.A(n_9008),
.B(n_549),
.Y(n_9163)
);

NOR2xp33_ASAP7_75t_L g9164 ( 
.A(n_8872),
.B(n_1649),
.Y(n_9164)
);

INVx2_ASAP7_75t_L g9165 ( 
.A(n_8899),
.Y(n_9165)
);

INVx1_ASAP7_75t_L g9166 ( 
.A(n_8943),
.Y(n_9166)
);

INVx2_ASAP7_75t_L g9167 ( 
.A(n_8947),
.Y(n_9167)
);

INVx2_ASAP7_75t_L g9168 ( 
.A(n_8846),
.Y(n_9168)
);

INVx2_ASAP7_75t_L g9169 ( 
.A(n_8848),
.Y(n_9169)
);

AND2x4_ASAP7_75t_L g9170 ( 
.A(n_8907),
.B(n_549),
.Y(n_9170)
);

INVx1_ASAP7_75t_L g9171 ( 
.A(n_8843),
.Y(n_9171)
);

INVx2_ASAP7_75t_L g9172 ( 
.A(n_8879),
.Y(n_9172)
);

OR2x2_ASAP7_75t_L g9173 ( 
.A(n_8778),
.B(n_549),
.Y(n_9173)
);

INVx2_ASAP7_75t_L g9174 ( 
.A(n_8967),
.Y(n_9174)
);

INVx1_ASAP7_75t_L g9175 ( 
.A(n_8963),
.Y(n_9175)
);

AND2x4_ASAP7_75t_L g9176 ( 
.A(n_8941),
.B(n_550),
.Y(n_9176)
);

AND2x2_ASAP7_75t_L g9177 ( 
.A(n_8798),
.B(n_550),
.Y(n_9177)
);

INVxp67_ASAP7_75t_SL g9178 ( 
.A(n_8838),
.Y(n_9178)
);

INVx2_ASAP7_75t_L g9179 ( 
.A(n_8861),
.Y(n_9179)
);

INVx2_ASAP7_75t_L g9180 ( 
.A(n_9014),
.Y(n_9180)
);

AND2x2_ASAP7_75t_L g9181 ( 
.A(n_9023),
.B(n_551),
.Y(n_9181)
);

BUFx2_ASAP7_75t_L g9182 ( 
.A(n_8918),
.Y(n_9182)
);

INVx1_ASAP7_75t_L g9183 ( 
.A(n_8931),
.Y(n_9183)
);

AND2x2_ASAP7_75t_L g9184 ( 
.A(n_8794),
.B(n_551),
.Y(n_9184)
);

AND2x2_ASAP7_75t_L g9185 ( 
.A(n_8915),
.B(n_551),
.Y(n_9185)
);

NAND2xp5_ASAP7_75t_L g9186 ( 
.A(n_9020),
.B(n_1650),
.Y(n_9186)
);

INVx2_ASAP7_75t_L g9187 ( 
.A(n_8942),
.Y(n_9187)
);

OR2x2_ASAP7_75t_L g9188 ( 
.A(n_8780),
.B(n_552),
.Y(n_9188)
);

INVx1_ASAP7_75t_L g9189 ( 
.A(n_8921),
.Y(n_9189)
);

BUFx2_ASAP7_75t_L g9190 ( 
.A(n_8883),
.Y(n_9190)
);

INVx2_ASAP7_75t_L g9191 ( 
.A(n_8969),
.Y(n_9191)
);

INVx2_ASAP7_75t_L g9192 ( 
.A(n_8849),
.Y(n_9192)
);

AND2x4_ASAP7_75t_SL g9193 ( 
.A(n_8791),
.B(n_552),
.Y(n_9193)
);

INVx2_ASAP7_75t_L g9194 ( 
.A(n_8977),
.Y(n_9194)
);

INVx1_ASAP7_75t_L g9195 ( 
.A(n_8986),
.Y(n_9195)
);

INVx1_ASAP7_75t_L g9196 ( 
.A(n_8993),
.Y(n_9196)
);

INVx2_ASAP7_75t_L g9197 ( 
.A(n_9026),
.Y(n_9197)
);

INVx1_ASAP7_75t_L g9198 ( 
.A(n_8998),
.Y(n_9198)
);

INVx5_ASAP7_75t_SL g9199 ( 
.A(n_8991),
.Y(n_9199)
);

BUFx3_ASAP7_75t_L g9200 ( 
.A(n_8906),
.Y(n_9200)
);

NOR2x1_ASAP7_75t_SL g9201 ( 
.A(n_8990),
.B(n_552),
.Y(n_9201)
);

INVx2_ASAP7_75t_L g9202 ( 
.A(n_9011),
.Y(n_9202)
);

INVx2_ASAP7_75t_L g9203 ( 
.A(n_8792),
.Y(n_9203)
);

INVx2_ASAP7_75t_L g9204 ( 
.A(n_8964),
.Y(n_9204)
);

AND2x2_ASAP7_75t_L g9205 ( 
.A(n_8776),
.B(n_553),
.Y(n_9205)
);

INVx1_ASAP7_75t_L g9206 ( 
.A(n_8939),
.Y(n_9206)
);

INVx2_ASAP7_75t_L g9207 ( 
.A(n_8886),
.Y(n_9207)
);

INVx2_ASAP7_75t_L g9208 ( 
.A(n_8892),
.Y(n_9208)
);

INVx1_ASAP7_75t_L g9209 ( 
.A(n_8847),
.Y(n_9209)
);

HB1xp67_ASAP7_75t_L g9210 ( 
.A(n_8961),
.Y(n_9210)
);

CKINVDCx5p33_ASAP7_75t_R g9211 ( 
.A(n_8875),
.Y(n_9211)
);

OR2x2_ASAP7_75t_L g9212 ( 
.A(n_8928),
.B(n_8925),
.Y(n_9212)
);

OR2x6_ASAP7_75t_L g9213 ( 
.A(n_8805),
.B(n_1650),
.Y(n_9213)
);

AND2x2_ASAP7_75t_L g9214 ( 
.A(n_8774),
.B(n_553),
.Y(n_9214)
);

INVx1_ASAP7_75t_L g9215 ( 
.A(n_8953),
.Y(n_9215)
);

AND2x2_ASAP7_75t_L g9216 ( 
.A(n_8785),
.B(n_553),
.Y(n_9216)
);

AND2x2_ASAP7_75t_L g9217 ( 
.A(n_8871),
.B(n_554),
.Y(n_9217)
);

AND2x2_ASAP7_75t_L g9218 ( 
.A(n_8959),
.B(n_555),
.Y(n_9218)
);

INVx2_ASAP7_75t_SL g9219 ( 
.A(n_8894),
.Y(n_9219)
);

INVx2_ASAP7_75t_L g9220 ( 
.A(n_8804),
.Y(n_9220)
);

INVx1_ASAP7_75t_L g9221 ( 
.A(n_8898),
.Y(n_9221)
);

NAND2xp5_ASAP7_75t_L g9222 ( 
.A(n_8972),
.B(n_1652),
.Y(n_9222)
);

AND2x2_ASAP7_75t_L g9223 ( 
.A(n_8789),
.B(n_8786),
.Y(n_9223)
);

OAI31xp33_ASAP7_75t_SL g9224 ( 
.A1(n_9003),
.A2(n_557),
.A3(n_555),
.B(n_556),
.Y(n_9224)
);

AND2x2_ASAP7_75t_L g9225 ( 
.A(n_8874),
.B(n_555),
.Y(n_9225)
);

AND2x2_ASAP7_75t_L g9226 ( 
.A(n_8881),
.B(n_556),
.Y(n_9226)
);

AND2x2_ASAP7_75t_L g9227 ( 
.A(n_8913),
.B(n_557),
.Y(n_9227)
);

AND2x4_ASAP7_75t_L g9228 ( 
.A(n_8808),
.B(n_8812),
.Y(n_9228)
);

BUFx2_ASAP7_75t_SL g9229 ( 
.A(n_8902),
.Y(n_9229)
);

INVx1_ASAP7_75t_L g9230 ( 
.A(n_9005),
.Y(n_9230)
);

INVx2_ASAP7_75t_L g9231 ( 
.A(n_8797),
.Y(n_9231)
);

INVx3_ASAP7_75t_L g9232 ( 
.A(n_8877),
.Y(n_9232)
);

INVx2_ASAP7_75t_L g9233 ( 
.A(n_8957),
.Y(n_9233)
);

INVx2_ASAP7_75t_SL g9234 ( 
.A(n_8960),
.Y(n_9234)
);

AND2x2_ASAP7_75t_L g9235 ( 
.A(n_8952),
.B(n_557),
.Y(n_9235)
);

AND2x2_ASAP7_75t_L g9236 ( 
.A(n_8946),
.B(n_8844),
.Y(n_9236)
);

INVx1_ASAP7_75t_L g9237 ( 
.A(n_9028),
.Y(n_9237)
);

NAND2xp5_ASAP7_75t_L g9238 ( 
.A(n_9030),
.B(n_1652),
.Y(n_9238)
);

INVx2_ASAP7_75t_L g9239 ( 
.A(n_8833),
.Y(n_9239)
);

INVx2_ASAP7_75t_L g9240 ( 
.A(n_8851),
.Y(n_9240)
);

INVx2_ASAP7_75t_L g9241 ( 
.A(n_8852),
.Y(n_9241)
);

INVx4_ASAP7_75t_R g9242 ( 
.A(n_8807),
.Y(n_9242)
);

AND2x2_ASAP7_75t_L g9243 ( 
.A(n_8867),
.B(n_558),
.Y(n_9243)
);

INVx2_ASAP7_75t_SL g9244 ( 
.A(n_8823),
.Y(n_9244)
);

OR2x2_ASAP7_75t_L g9245 ( 
.A(n_8841),
.B(n_558),
.Y(n_9245)
);

INVx4_ASAP7_75t_L g9246 ( 
.A(n_8994),
.Y(n_9246)
);

INVx1_ASAP7_75t_L g9247 ( 
.A(n_8996),
.Y(n_9247)
);

AND2x2_ASAP7_75t_L g9248 ( 
.A(n_8878),
.B(n_558),
.Y(n_9248)
);

INVx4_ASAP7_75t_R g9249 ( 
.A(n_9002),
.Y(n_9249)
);

INVx2_ASAP7_75t_L g9250 ( 
.A(n_9021),
.Y(n_9250)
);

INVx2_ASAP7_75t_L g9251 ( 
.A(n_8829),
.Y(n_9251)
);

INVx2_ASAP7_75t_L g9252 ( 
.A(n_8863),
.Y(n_9252)
);

INVx2_ASAP7_75t_L g9253 ( 
.A(n_8864),
.Y(n_9253)
);

INVx1_ASAP7_75t_L g9254 ( 
.A(n_8900),
.Y(n_9254)
);

BUFx6f_ASAP7_75t_L g9255 ( 
.A(n_8945),
.Y(n_9255)
);

NAND2xp5_ASAP7_75t_L g9256 ( 
.A(n_9007),
.B(n_1653),
.Y(n_9256)
);

BUFx2_ASAP7_75t_L g9257 ( 
.A(n_8865),
.Y(n_9257)
);

NOR2x1_ASAP7_75t_L g9258 ( 
.A(n_8777),
.B(n_559),
.Y(n_9258)
);

NAND4xp25_ASAP7_75t_L g9259 ( 
.A(n_9010),
.B(n_561),
.C(n_559),
.D(n_560),
.Y(n_9259)
);

AND2x2_ASAP7_75t_L g9260 ( 
.A(n_8888),
.B(n_559),
.Y(n_9260)
);

BUFx2_ASAP7_75t_L g9261 ( 
.A(n_8891),
.Y(n_9261)
);

INVx1_ASAP7_75t_L g9262 ( 
.A(n_8811),
.Y(n_9262)
);

OR2x2_ASAP7_75t_L g9263 ( 
.A(n_8912),
.B(n_560),
.Y(n_9263)
);

OR2x2_ASAP7_75t_L g9264 ( 
.A(n_8901),
.B(n_8916),
.Y(n_9264)
);

AND2x2_ASAP7_75t_L g9265 ( 
.A(n_8790),
.B(n_560),
.Y(n_9265)
);

INVx1_ASAP7_75t_L g9266 ( 
.A(n_8950),
.Y(n_9266)
);

INVx2_ASAP7_75t_L g9267 ( 
.A(n_8974),
.Y(n_9267)
);

NAND2xp5_ASAP7_75t_L g9268 ( 
.A(n_8980),
.B(n_8981),
.Y(n_9268)
);

NOR2x1_ASAP7_75t_SL g9269 ( 
.A(n_8982),
.B(n_561),
.Y(n_9269)
);

INVx1_ASAP7_75t_L g9270 ( 
.A(n_8884),
.Y(n_9270)
);

AND2x2_ASAP7_75t_L g9271 ( 
.A(n_8781),
.B(n_8782),
.Y(n_9271)
);

OR2x6_ASAP7_75t_L g9272 ( 
.A(n_8995),
.B(n_1653),
.Y(n_9272)
);

BUFx6f_ASAP7_75t_L g9273 ( 
.A(n_8944),
.Y(n_9273)
);

AND2x2_ASAP7_75t_L g9274 ( 
.A(n_9000),
.B(n_561),
.Y(n_9274)
);

INVx1_ASAP7_75t_L g9275 ( 
.A(n_8962),
.Y(n_9275)
);

BUFx2_ASAP7_75t_L g9276 ( 
.A(n_8824),
.Y(n_9276)
);

INVx2_ASAP7_75t_L g9277 ( 
.A(n_9012),
.Y(n_9277)
);

INVx1_ASAP7_75t_L g9278 ( 
.A(n_8965),
.Y(n_9278)
);

AND2x2_ASAP7_75t_L g9279 ( 
.A(n_9013),
.B(n_562),
.Y(n_9279)
);

BUFx2_ASAP7_75t_L g9280 ( 
.A(n_8971),
.Y(n_9280)
);

INVx2_ASAP7_75t_L g9281 ( 
.A(n_8816),
.Y(n_9281)
);

INVx1_ASAP7_75t_L g9282 ( 
.A(n_8825),
.Y(n_9282)
);

INVx2_ASAP7_75t_SL g9283 ( 
.A(n_8827),
.Y(n_9283)
);

INVx1_ASAP7_75t_L g9284 ( 
.A(n_8806),
.Y(n_9284)
);

INVx1_ASAP7_75t_L g9285 ( 
.A(n_8830),
.Y(n_9285)
);

AND2x2_ASAP7_75t_L g9286 ( 
.A(n_8885),
.B(n_562),
.Y(n_9286)
);

HB1xp67_ASAP7_75t_L g9287 ( 
.A(n_8799),
.Y(n_9287)
);

INVx2_ASAP7_75t_L g9288 ( 
.A(n_8770),
.Y(n_9288)
);

INVx1_ASAP7_75t_L g9289 ( 
.A(n_8768),
.Y(n_9289)
);

INVx1_ASAP7_75t_L g9290 ( 
.A(n_8768),
.Y(n_9290)
);

AND2x2_ASAP7_75t_L g9291 ( 
.A(n_8770),
.B(n_562),
.Y(n_9291)
);

AND2x2_ASAP7_75t_L g9292 ( 
.A(n_8770),
.B(n_563),
.Y(n_9292)
);

INVx1_ASAP7_75t_L g9293 ( 
.A(n_8768),
.Y(n_9293)
);

BUFx2_ASAP7_75t_L g9294 ( 
.A(n_8770),
.Y(n_9294)
);

INVx2_ASAP7_75t_L g9295 ( 
.A(n_8770),
.Y(n_9295)
);

INVx2_ASAP7_75t_L g9296 ( 
.A(n_8770),
.Y(n_9296)
);

AND2x2_ASAP7_75t_L g9297 ( 
.A(n_8770),
.B(n_563),
.Y(n_9297)
);

BUFx2_ASAP7_75t_L g9298 ( 
.A(n_8770),
.Y(n_9298)
);

HB1xp67_ASAP7_75t_L g9299 ( 
.A(n_8831),
.Y(n_9299)
);

NAND2xp5_ASAP7_75t_L g9300 ( 
.A(n_8934),
.B(n_1654),
.Y(n_9300)
);

INVx5_ASAP7_75t_L g9301 ( 
.A(n_9027),
.Y(n_9301)
);

NAND2xp5_ASAP7_75t_L g9302 ( 
.A(n_8934),
.B(n_1654),
.Y(n_9302)
);

INVx2_ASAP7_75t_L g9303 ( 
.A(n_8770),
.Y(n_9303)
);

NOR2xp33_ASAP7_75t_L g9304 ( 
.A(n_8997),
.B(n_1655),
.Y(n_9304)
);

INVx1_ASAP7_75t_L g9305 ( 
.A(n_8768),
.Y(n_9305)
);

INVx2_ASAP7_75t_L g9306 ( 
.A(n_8770),
.Y(n_9306)
);

INVx1_ASAP7_75t_L g9307 ( 
.A(n_8768),
.Y(n_9307)
);

INVx2_ASAP7_75t_L g9308 ( 
.A(n_8770),
.Y(n_9308)
);

AND2x2_ASAP7_75t_L g9309 ( 
.A(n_8770),
.B(n_564),
.Y(n_9309)
);

INVx1_ASAP7_75t_L g9310 ( 
.A(n_8768),
.Y(n_9310)
);

AND2x2_ASAP7_75t_L g9311 ( 
.A(n_8770),
.B(n_564),
.Y(n_9311)
);

HB1xp67_ASAP7_75t_L g9312 ( 
.A(n_8831),
.Y(n_9312)
);

INVx1_ASAP7_75t_L g9313 ( 
.A(n_8768),
.Y(n_9313)
);

AND2x4_ASAP7_75t_L g9314 ( 
.A(n_8773),
.B(n_565),
.Y(n_9314)
);

INVxp67_ASAP7_75t_SL g9315 ( 
.A(n_8770),
.Y(n_9315)
);

NOR2xp33_ASAP7_75t_L g9316 ( 
.A(n_8997),
.B(n_1655),
.Y(n_9316)
);

INVx3_ASAP7_75t_L g9317 ( 
.A(n_8810),
.Y(n_9317)
);

AND2x2_ASAP7_75t_L g9318 ( 
.A(n_8770),
.B(n_565),
.Y(n_9318)
);

AND2x2_ASAP7_75t_L g9319 ( 
.A(n_8770),
.B(n_565),
.Y(n_9319)
);

NAND2xp5_ASAP7_75t_L g9320 ( 
.A(n_8934),
.B(n_1656),
.Y(n_9320)
);

INVx1_ASAP7_75t_L g9321 ( 
.A(n_8768),
.Y(n_9321)
);

AND2x2_ASAP7_75t_L g9322 ( 
.A(n_8770),
.B(n_566),
.Y(n_9322)
);

OR2x2_ASAP7_75t_L g9323 ( 
.A(n_8908),
.B(n_566),
.Y(n_9323)
);

AND2x4_ASAP7_75t_L g9324 ( 
.A(n_8773),
.B(n_567),
.Y(n_9324)
);

INVx2_ASAP7_75t_L g9325 ( 
.A(n_8770),
.Y(n_9325)
);

AND2x4_ASAP7_75t_L g9326 ( 
.A(n_8773),
.B(n_567),
.Y(n_9326)
);

INVx2_ASAP7_75t_SL g9327 ( 
.A(n_9027),
.Y(n_9327)
);

AND2x2_ASAP7_75t_L g9328 ( 
.A(n_8770),
.B(n_567),
.Y(n_9328)
);

INVx2_ASAP7_75t_L g9329 ( 
.A(n_8770),
.Y(n_9329)
);

AND2x2_ASAP7_75t_L g9330 ( 
.A(n_8770),
.B(n_568),
.Y(n_9330)
);

INVx2_ASAP7_75t_L g9331 ( 
.A(n_8770),
.Y(n_9331)
);

INVx1_ASAP7_75t_L g9332 ( 
.A(n_8768),
.Y(n_9332)
);

AND2x2_ASAP7_75t_L g9333 ( 
.A(n_8770),
.B(n_568),
.Y(n_9333)
);

OAI33xp33_ASAP7_75t_L g9334 ( 
.A1(n_9171),
.A2(n_571),
.A3(n_574),
.B1(n_569),
.B2(n_570),
.B3(n_572),
.Y(n_9334)
);

OAI31xp33_ASAP7_75t_L g9335 ( 
.A1(n_9049),
.A2(n_571),
.A3(n_572),
.B(n_570),
.Y(n_9335)
);

OR2x2_ASAP7_75t_L g9336 ( 
.A(n_9288),
.B(n_569),
.Y(n_9336)
);

AOI211xp5_ASAP7_75t_SL g9337 ( 
.A1(n_9139),
.A2(n_571),
.B(n_569),
.C(n_570),
.Y(n_9337)
);

OAI22xp5_ASAP7_75t_L g9338 ( 
.A1(n_9199),
.A2(n_575),
.B1(n_572),
.B2(n_574),
.Y(n_9338)
);

NAND2xp5_ASAP7_75t_L g9339 ( 
.A(n_9223),
.B(n_575),
.Y(n_9339)
);

OAI22xp33_ASAP7_75t_L g9340 ( 
.A1(n_9246),
.A2(n_9258),
.B1(n_9178),
.B2(n_9034),
.Y(n_9340)
);

AO31x2_ASAP7_75t_L g9341 ( 
.A1(n_9148),
.A2(n_577),
.A3(n_575),
.B(n_576),
.Y(n_9341)
);

INVx2_ASAP7_75t_L g9342 ( 
.A(n_9063),
.Y(n_9342)
);

BUFx3_ASAP7_75t_L g9343 ( 
.A(n_9301),
.Y(n_9343)
);

INVx1_ASAP7_75t_L g9344 ( 
.A(n_9035),
.Y(n_9344)
);

OAI22xp5_ASAP7_75t_L g9345 ( 
.A1(n_9199),
.A2(n_578),
.B1(n_576),
.B2(n_577),
.Y(n_9345)
);

INVx2_ASAP7_75t_L g9346 ( 
.A(n_9105),
.Y(n_9346)
);

AOI22xp33_ASAP7_75t_SL g9347 ( 
.A1(n_9229),
.A2(n_578),
.B1(n_576),
.B2(n_577),
.Y(n_9347)
);

INVx2_ASAP7_75t_L g9348 ( 
.A(n_9108),
.Y(n_9348)
);

OAI22xp5_ASAP7_75t_L g9349 ( 
.A1(n_9033),
.A2(n_581),
.B1(n_579),
.B2(n_580),
.Y(n_9349)
);

INVx2_ASAP7_75t_L g9350 ( 
.A(n_9040),
.Y(n_9350)
);

OAI221xp5_ASAP7_75t_L g9351 ( 
.A1(n_9276),
.A2(n_581),
.B1(n_579),
.B2(n_580),
.C(n_582),
.Y(n_9351)
);

OA21x2_ASAP7_75t_L g9352 ( 
.A1(n_9182),
.A2(n_579),
.B(n_582),
.Y(n_9352)
);

HB1xp67_ASAP7_75t_L g9353 ( 
.A(n_9294),
.Y(n_9353)
);

INVx1_ASAP7_75t_L g9354 ( 
.A(n_9038),
.Y(n_9354)
);

OAI33xp33_ASAP7_75t_L g9355 ( 
.A1(n_9150),
.A2(n_584),
.A3(n_586),
.B1(n_582),
.B2(n_583),
.B3(n_585),
.Y(n_9355)
);

BUFx3_ASAP7_75t_L g9356 ( 
.A(n_9301),
.Y(n_9356)
);

AOI22xp33_ASAP7_75t_L g9357 ( 
.A1(n_9251),
.A2(n_585),
.B1(n_583),
.B2(n_584),
.Y(n_9357)
);

AND2x2_ASAP7_75t_L g9358 ( 
.A(n_9298),
.B(n_584),
.Y(n_9358)
);

AND2x2_ASAP7_75t_L g9359 ( 
.A(n_9051),
.B(n_587),
.Y(n_9359)
);

NAND2xp5_ASAP7_75t_L g9360 ( 
.A(n_9262),
.B(n_587),
.Y(n_9360)
);

OAI22xp33_ASAP7_75t_L g9361 ( 
.A1(n_9032),
.A2(n_9312),
.B1(n_9299),
.B2(n_9169),
.Y(n_9361)
);

AND2x2_ASAP7_75t_L g9362 ( 
.A(n_9066),
.B(n_587),
.Y(n_9362)
);

OAI31xp33_ASAP7_75t_L g9363 ( 
.A1(n_9261),
.A2(n_590),
.A3(n_591),
.B(n_589),
.Y(n_9363)
);

INVx2_ASAP7_75t_L g9364 ( 
.A(n_9091),
.Y(n_9364)
);

OAI211xp5_ASAP7_75t_L g9365 ( 
.A1(n_9224),
.A2(n_597),
.B(n_605),
.C(n_588),
.Y(n_9365)
);

OAI22xp5_ASAP7_75t_L g9366 ( 
.A1(n_9190),
.A2(n_590),
.B1(n_588),
.B2(n_589),
.Y(n_9366)
);

OAI22xp5_ASAP7_75t_L g9367 ( 
.A1(n_9257),
.A2(n_594),
.B1(n_592),
.B2(n_593),
.Y(n_9367)
);

NAND2xp5_ASAP7_75t_L g9368 ( 
.A(n_9210),
.B(n_592),
.Y(n_9368)
);

AND2x2_ASAP7_75t_L g9369 ( 
.A(n_9315),
.B(n_592),
.Y(n_9369)
);

INVx2_ASAP7_75t_L g9370 ( 
.A(n_9085),
.Y(n_9370)
);

INVx1_ASAP7_75t_L g9371 ( 
.A(n_9042),
.Y(n_9371)
);

AOI21xp5_ASAP7_75t_L g9372 ( 
.A1(n_9056),
.A2(n_593),
.B(n_594),
.Y(n_9372)
);

NAND3xp33_ASAP7_75t_L g9373 ( 
.A(n_9047),
.B(n_593),
.C(n_595),
.Y(n_9373)
);

AOI22xp33_ASAP7_75t_L g9374 ( 
.A1(n_9255),
.A2(n_597),
.B1(n_595),
.B2(n_596),
.Y(n_9374)
);

OA21x2_ASAP7_75t_L g9375 ( 
.A1(n_9175),
.A2(n_595),
.B(n_596),
.Y(n_9375)
);

AOI22xp33_ASAP7_75t_L g9376 ( 
.A1(n_9255),
.A2(n_599),
.B1(n_596),
.B2(n_598),
.Y(n_9376)
);

AND2x2_ASAP7_75t_L g9377 ( 
.A(n_9295),
.B(n_598),
.Y(n_9377)
);

AND2x2_ASAP7_75t_L g9378 ( 
.A(n_9296),
.B(n_599),
.Y(n_9378)
);

NOR2xp33_ASAP7_75t_L g9379 ( 
.A(n_9044),
.B(n_600),
.Y(n_9379)
);

AND2x2_ASAP7_75t_L g9380 ( 
.A(n_9303),
.B(n_600),
.Y(n_9380)
);

AOI22xp33_ASAP7_75t_L g9381 ( 
.A1(n_9271),
.A2(n_603),
.B1(n_601),
.B2(n_602),
.Y(n_9381)
);

AOI221xp5_ASAP7_75t_L g9382 ( 
.A1(n_9164),
.A2(n_603),
.B1(n_601),
.B2(n_602),
.C(n_604),
.Y(n_9382)
);

AND2x4_ASAP7_75t_L g9383 ( 
.A(n_9039),
.B(n_601),
.Y(n_9383)
);

AOI22xp5_ASAP7_75t_L g9384 ( 
.A1(n_9228),
.A2(n_605),
.B1(n_602),
.B2(n_604),
.Y(n_9384)
);

OAI211xp5_ASAP7_75t_L g9385 ( 
.A1(n_9140),
.A2(n_614),
.B(n_623),
.C(n_606),
.Y(n_9385)
);

OR2x2_ASAP7_75t_L g9386 ( 
.A(n_9306),
.B(n_606),
.Y(n_9386)
);

INVx2_ASAP7_75t_L g9387 ( 
.A(n_9317),
.Y(n_9387)
);

OAI22xp33_ASAP7_75t_L g9388 ( 
.A1(n_9213),
.A2(n_609),
.B1(n_607),
.B2(n_608),
.Y(n_9388)
);

NAND3xp33_ASAP7_75t_L g9389 ( 
.A(n_9082),
.B(n_9124),
.C(n_9259),
.Y(n_9389)
);

INVx1_ASAP7_75t_L g9390 ( 
.A(n_9053),
.Y(n_9390)
);

NAND2xp5_ASAP7_75t_L g9391 ( 
.A(n_9174),
.B(n_9149),
.Y(n_9391)
);

INVx1_ASAP7_75t_L g9392 ( 
.A(n_9058),
.Y(n_9392)
);

BUFx2_ASAP7_75t_L g9393 ( 
.A(n_9156),
.Y(n_9393)
);

OAI221xp5_ASAP7_75t_L g9394 ( 
.A1(n_9220),
.A2(n_9173),
.B1(n_9083),
.B2(n_9192),
.C(n_9254),
.Y(n_9394)
);

AND2x4_ASAP7_75t_L g9395 ( 
.A(n_9327),
.B(n_607),
.Y(n_9395)
);

AOI221xp5_ASAP7_75t_L g9396 ( 
.A1(n_9054),
.A2(n_609),
.B1(n_607),
.B2(n_608),
.C(n_610),
.Y(n_9396)
);

AOI22xp33_ASAP7_75t_L g9397 ( 
.A1(n_9200),
.A2(n_612),
.B1(n_610),
.B2(n_611),
.Y(n_9397)
);

AO21x2_ASAP7_75t_L g9398 ( 
.A1(n_9300),
.A2(n_610),
.B(n_611),
.Y(n_9398)
);

OAI211xp5_ASAP7_75t_SL g9399 ( 
.A1(n_9194),
.A2(n_9197),
.B(n_9208),
.C(n_9187),
.Y(n_9399)
);

OAI21xp5_ASAP7_75t_L g9400 ( 
.A1(n_9302),
.A2(n_612),
.B(n_613),
.Y(n_9400)
);

NAND2xp5_ASAP7_75t_L g9401 ( 
.A(n_9158),
.B(n_612),
.Y(n_9401)
);

AND2x4_ASAP7_75t_SL g9402 ( 
.A(n_9138),
.B(n_613),
.Y(n_9402)
);

AOI22xp33_ASAP7_75t_L g9403 ( 
.A1(n_9280),
.A2(n_615),
.B1(n_613),
.B2(n_614),
.Y(n_9403)
);

INVxp67_ASAP7_75t_SL g9404 ( 
.A(n_9130),
.Y(n_9404)
);

OAI22xp33_ASAP7_75t_L g9405 ( 
.A1(n_9213),
.A2(n_9253),
.B1(n_9252),
.B2(n_9320),
.Y(n_9405)
);

INVxp67_ASAP7_75t_SL g9406 ( 
.A(n_9110),
.Y(n_9406)
);

OAI21xp33_ASAP7_75t_L g9407 ( 
.A1(n_9043),
.A2(n_615),
.B(n_616),
.Y(n_9407)
);

OAI31xp33_ASAP7_75t_L g9408 ( 
.A1(n_9236),
.A2(n_617),
.A3(n_619),
.B(n_616),
.Y(n_9408)
);

OA21x2_ASAP7_75t_L g9409 ( 
.A1(n_9075),
.A2(n_615),
.B(n_619),
.Y(n_9409)
);

OAI22xp33_ASAP7_75t_L g9410 ( 
.A1(n_9188),
.A2(n_621),
.B1(n_619),
.B2(n_620),
.Y(n_9410)
);

AOI22xp33_ASAP7_75t_L g9411 ( 
.A1(n_9287),
.A2(n_622),
.B1(n_620),
.B2(n_621),
.Y(n_9411)
);

INVx2_ASAP7_75t_L g9412 ( 
.A(n_9084),
.Y(n_9412)
);

INVx2_ASAP7_75t_L g9413 ( 
.A(n_9308),
.Y(n_9413)
);

NAND4xp25_ASAP7_75t_L g9414 ( 
.A(n_9076),
.B(n_624),
.C(n_622),
.D(n_623),
.Y(n_9414)
);

AOI22xp33_ASAP7_75t_L g9415 ( 
.A1(n_9273),
.A2(n_625),
.B1(n_623),
.B2(n_624),
.Y(n_9415)
);

OAI22xp5_ASAP7_75t_L g9416 ( 
.A1(n_9232),
.A2(n_626),
.B1(n_624),
.B2(n_625),
.Y(n_9416)
);

AOI33xp33_ASAP7_75t_L g9417 ( 
.A1(n_9242),
.A2(n_628),
.A3(n_630),
.B1(n_626),
.B2(n_627),
.B3(n_629),
.Y(n_9417)
);

OAI21xp5_ASAP7_75t_L g9418 ( 
.A1(n_9256),
.A2(n_628),
.B(n_629),
.Y(n_9418)
);

OA332x1_ASAP7_75t_L g9419 ( 
.A1(n_9249),
.A2(n_9095),
.A3(n_9212),
.B1(n_9244),
.B2(n_9209),
.B3(n_9201),
.C1(n_9195),
.C2(n_9198),
.Y(n_9419)
);

INVx2_ASAP7_75t_L g9420 ( 
.A(n_9325),
.Y(n_9420)
);

AOI221xp5_ASAP7_75t_L g9421 ( 
.A1(n_9196),
.A2(n_631),
.B1(n_628),
.B2(n_630),
.C(n_632),
.Y(n_9421)
);

INVx2_ASAP7_75t_L g9422 ( 
.A(n_9329),
.Y(n_9422)
);

NOR2xp33_ASAP7_75t_L g9423 ( 
.A(n_9037),
.B(n_631),
.Y(n_9423)
);

HB1xp67_ASAP7_75t_L g9424 ( 
.A(n_9143),
.Y(n_9424)
);

INVx1_ASAP7_75t_L g9425 ( 
.A(n_9062),
.Y(n_9425)
);

OAI33xp33_ASAP7_75t_L g9426 ( 
.A1(n_9230),
.A2(n_633),
.A3(n_635),
.B1(n_631),
.B2(n_632),
.B3(n_634),
.Y(n_9426)
);

BUFx6f_ASAP7_75t_L g9427 ( 
.A(n_9127),
.Y(n_9427)
);

INVx2_ASAP7_75t_L g9428 ( 
.A(n_9331),
.Y(n_9428)
);

INVx1_ASAP7_75t_L g9429 ( 
.A(n_9064),
.Y(n_9429)
);

BUFx3_ASAP7_75t_L g9430 ( 
.A(n_9129),
.Y(n_9430)
);

AOI33xp33_ASAP7_75t_L g9431 ( 
.A1(n_9247),
.A2(n_634),
.A3(n_636),
.B1(n_632),
.B2(n_633),
.B3(n_635),
.Y(n_9431)
);

OA222x2_ASAP7_75t_L g9432 ( 
.A1(n_9080),
.A2(n_635),
.B1(n_637),
.B2(n_633),
.C1(n_634),
.C2(n_636),
.Y(n_9432)
);

AOI21xp5_ASAP7_75t_L g9433 ( 
.A1(n_9268),
.A2(n_636),
.B(n_637),
.Y(n_9433)
);

AND2x2_ASAP7_75t_L g9434 ( 
.A(n_9048),
.B(n_638),
.Y(n_9434)
);

INVx1_ASAP7_75t_L g9435 ( 
.A(n_9067),
.Y(n_9435)
);

AOI22xp33_ASAP7_75t_L g9436 ( 
.A1(n_9273),
.A2(n_640),
.B1(n_638),
.B2(n_639),
.Y(n_9436)
);

INVx1_ASAP7_75t_L g9437 ( 
.A(n_9068),
.Y(n_9437)
);

BUFx2_ASAP7_75t_L g9438 ( 
.A(n_9134),
.Y(n_9438)
);

AOI221xp5_ASAP7_75t_L g9439 ( 
.A1(n_9240),
.A2(n_9172),
.B1(n_9189),
.B2(n_9237),
.C(n_9250),
.Y(n_9439)
);

INVx1_ASAP7_75t_L g9440 ( 
.A(n_9070),
.Y(n_9440)
);

AND2x4_ASAP7_75t_L g9441 ( 
.A(n_9141),
.B(n_638),
.Y(n_9441)
);

AOI211xp5_ASAP7_75t_SL g9442 ( 
.A1(n_9222),
.A2(n_641),
.B(n_639),
.C(n_640),
.Y(n_9442)
);

OR2x2_ASAP7_75t_L g9443 ( 
.A(n_9055),
.B(n_639),
.Y(n_9443)
);

OAI21xp5_ASAP7_75t_SL g9444 ( 
.A1(n_9176),
.A2(n_644),
.B(n_643),
.Y(n_9444)
);

AND2x4_ASAP7_75t_L g9445 ( 
.A(n_9125),
.B(n_642),
.Y(n_9445)
);

AOI22xp5_ASAP7_75t_L g9446 ( 
.A1(n_9092),
.A2(n_644),
.B1(n_642),
.B2(n_643),
.Y(n_9446)
);

OAI31xp33_ASAP7_75t_L g9447 ( 
.A1(n_9097),
.A2(n_645),
.A3(n_646),
.B(n_643),
.Y(n_9447)
);

AND2x2_ASAP7_75t_L g9448 ( 
.A(n_9146),
.B(n_642),
.Y(n_9448)
);

AND2x4_ASAP7_75t_L g9449 ( 
.A(n_9155),
.B(n_645),
.Y(n_9449)
);

AOI21xp5_ASAP7_75t_L g9450 ( 
.A1(n_9186),
.A2(n_645),
.B(n_646),
.Y(n_9450)
);

AOI21xp5_ASAP7_75t_L g9451 ( 
.A1(n_9152),
.A2(n_646),
.B(n_647),
.Y(n_9451)
);

INVx1_ASAP7_75t_L g9452 ( 
.A(n_9077),
.Y(n_9452)
);

NAND3xp33_ASAP7_75t_L g9453 ( 
.A(n_9241),
.B(n_647),
.C(n_648),
.Y(n_9453)
);

AOI22xp33_ASAP7_75t_L g9454 ( 
.A1(n_9202),
.A2(n_650),
.B1(n_648),
.B2(n_649),
.Y(n_9454)
);

AOI22xp33_ASAP7_75t_L g9455 ( 
.A1(n_9267),
.A2(n_650),
.B1(n_648),
.B2(n_649),
.Y(n_9455)
);

INVx1_ASAP7_75t_L g9456 ( 
.A(n_9078),
.Y(n_9456)
);

INVx1_ASAP7_75t_L g9457 ( 
.A(n_9087),
.Y(n_9457)
);

BUFx2_ASAP7_75t_L g9458 ( 
.A(n_9142),
.Y(n_9458)
);

OAI211xp5_ASAP7_75t_SL g9459 ( 
.A1(n_9284),
.A2(n_651),
.B(n_649),
.C(n_650),
.Y(n_9459)
);

INVx1_ASAP7_75t_L g9460 ( 
.A(n_9090),
.Y(n_9460)
);

AOI221xp5_ASAP7_75t_L g9461 ( 
.A1(n_9183),
.A2(n_654),
.B1(n_651),
.B2(n_652),
.C(n_655),
.Y(n_9461)
);

INVx1_ASAP7_75t_L g9462 ( 
.A(n_9096),
.Y(n_9462)
);

OAI21xp33_ASAP7_75t_L g9463 ( 
.A1(n_9238),
.A2(n_654),
.B(n_656),
.Y(n_9463)
);

AND2x2_ASAP7_75t_L g9464 ( 
.A(n_9088),
.B(n_9137),
.Y(n_9464)
);

AND2x4_ASAP7_75t_L g9465 ( 
.A(n_9154),
.B(n_654),
.Y(n_9465)
);

NAND2xp5_ASAP7_75t_L g9466 ( 
.A(n_9036),
.B(n_656),
.Y(n_9466)
);

AND2x2_ASAP7_75t_L g9467 ( 
.A(n_9109),
.B(n_656),
.Y(n_9467)
);

INVx2_ASAP7_75t_SL g9468 ( 
.A(n_9045),
.Y(n_9468)
);

AND2x2_ASAP7_75t_L g9469 ( 
.A(n_9145),
.B(n_657),
.Y(n_9469)
);

HB1xp67_ASAP7_75t_L g9470 ( 
.A(n_9099),
.Y(n_9470)
);

BUFx2_ASAP7_75t_L g9471 ( 
.A(n_9168),
.Y(n_9471)
);

OR2x2_ASAP7_75t_L g9472 ( 
.A(n_9323),
.B(n_657),
.Y(n_9472)
);

OAI221xp5_ASAP7_75t_L g9473 ( 
.A1(n_9283),
.A2(n_9231),
.B1(n_9144),
.B2(n_9277),
.C(n_9270),
.Y(n_9473)
);

INVx2_ASAP7_75t_L g9474 ( 
.A(n_9052),
.Y(n_9474)
);

INVx1_ASAP7_75t_L g9475 ( 
.A(n_9098),
.Y(n_9475)
);

INVx2_ASAP7_75t_L g9476 ( 
.A(n_9153),
.Y(n_9476)
);

AOI22xp33_ASAP7_75t_L g9477 ( 
.A1(n_9281),
.A2(n_659),
.B1(n_657),
.B2(n_658),
.Y(n_9477)
);

NAND2x1_ASAP7_75t_L g9478 ( 
.A(n_9165),
.B(n_658),
.Y(n_9478)
);

AND2x2_ASAP7_75t_L g9479 ( 
.A(n_9147),
.B(n_658),
.Y(n_9479)
);

AOI221xp5_ASAP7_75t_L g9480 ( 
.A1(n_9206),
.A2(n_661),
.B1(n_659),
.B2(n_660),
.C(n_662),
.Y(n_9480)
);

AND2x4_ASAP7_75t_L g9481 ( 
.A(n_9159),
.B(n_659),
.Y(n_9481)
);

OR2x6_ASAP7_75t_L g9482 ( 
.A(n_9046),
.B(n_9314),
.Y(n_9482)
);

AOI222xp33_ASAP7_75t_L g9483 ( 
.A1(n_9265),
.A2(n_662),
.B1(n_664),
.B2(n_660),
.C1(n_661),
.C2(n_663),
.Y(n_9483)
);

NAND4xp25_ASAP7_75t_L g9484 ( 
.A(n_9216),
.B(n_664),
.C(n_661),
.D(n_663),
.Y(n_9484)
);

AOI22xp33_ASAP7_75t_SL g9485 ( 
.A1(n_9170),
.A2(n_665),
.B1(n_663),
.B2(n_664),
.Y(n_9485)
);

AOI221xp5_ASAP7_75t_L g9486 ( 
.A1(n_9282),
.A2(n_667),
.B1(n_665),
.B2(n_666),
.C(n_668),
.Y(n_9486)
);

INVx1_ASAP7_75t_L g9487 ( 
.A(n_9104),
.Y(n_9487)
);

AND2x2_ASAP7_75t_L g9488 ( 
.A(n_9151),
.B(n_665),
.Y(n_9488)
);

INVx2_ASAP7_75t_L g9489 ( 
.A(n_9073),
.Y(n_9489)
);

OAI221xp5_ASAP7_75t_L g9490 ( 
.A1(n_9285),
.A2(n_668),
.B1(n_666),
.B2(n_667),
.C(n_669),
.Y(n_9490)
);

AOI22xp33_ASAP7_75t_L g9491 ( 
.A1(n_9180),
.A2(n_670),
.B1(n_666),
.B2(n_669),
.Y(n_9491)
);

OA21x2_ASAP7_75t_L g9492 ( 
.A1(n_9167),
.A2(n_672),
.B(n_671),
.Y(n_9492)
);

INVx1_ASAP7_75t_L g9493 ( 
.A(n_9107),
.Y(n_9493)
);

AND2x4_ASAP7_75t_L g9494 ( 
.A(n_9157),
.B(n_670),
.Y(n_9494)
);

INVx1_ASAP7_75t_L g9495 ( 
.A(n_9113),
.Y(n_9495)
);

NAND2xp5_ASAP7_75t_L g9496 ( 
.A(n_9239),
.B(n_671),
.Y(n_9496)
);

NAND4xp25_ASAP7_75t_L g9497 ( 
.A(n_9214),
.B(n_673),
.C(n_671),
.D(n_672),
.Y(n_9497)
);

AOI22xp33_ASAP7_75t_L g9498 ( 
.A1(n_9191),
.A2(n_674),
.B1(n_672),
.B2(n_673),
.Y(n_9498)
);

OAI221xp5_ASAP7_75t_L g9499 ( 
.A1(n_9266),
.A2(n_675),
.B1(n_673),
.B2(n_674),
.C(n_676),
.Y(n_9499)
);

OAI22xp5_ASAP7_75t_L g9500 ( 
.A1(n_9215),
.A2(n_677),
.B1(n_675),
.B2(n_676),
.Y(n_9500)
);

INVx2_ASAP7_75t_SL g9501 ( 
.A(n_9324),
.Y(n_9501)
);

OR2x2_ASAP7_75t_L g9502 ( 
.A(n_9121),
.B(n_675),
.Y(n_9502)
);

NAND2xp5_ASAP7_75t_SL g9503 ( 
.A(n_9079),
.B(n_677),
.Y(n_9503)
);

AND2x2_ASAP7_75t_L g9504 ( 
.A(n_9204),
.B(n_678),
.Y(n_9504)
);

INVxp67_ASAP7_75t_L g9505 ( 
.A(n_9106),
.Y(n_9505)
);

AOI22xp33_ASAP7_75t_L g9506 ( 
.A1(n_9275),
.A2(n_680),
.B1(n_678),
.B2(n_679),
.Y(n_9506)
);

NAND2xp5_ASAP7_75t_L g9507 ( 
.A(n_9166),
.B(n_678),
.Y(n_9507)
);

INVx1_ASAP7_75t_L g9508 ( 
.A(n_9123),
.Y(n_9508)
);

OAI33xp33_ASAP7_75t_L g9509 ( 
.A1(n_9221),
.A2(n_682),
.A3(n_684),
.B1(n_680),
.B2(n_681),
.B3(n_683),
.Y(n_9509)
);

OA21x2_ASAP7_75t_L g9510 ( 
.A1(n_9179),
.A2(n_683),
.B(n_681),
.Y(n_9510)
);

OAI221xp5_ASAP7_75t_L g9511 ( 
.A1(n_9278),
.A2(n_683),
.B1(n_680),
.B2(n_681),
.C(n_684),
.Y(n_9511)
);

INVx3_ASAP7_75t_L g9512 ( 
.A(n_9326),
.Y(n_9512)
);

NAND3xp33_ASAP7_75t_L g9513 ( 
.A(n_9264),
.B(n_9203),
.C(n_9185),
.Y(n_9513)
);

A2O1A1Ixp33_ASAP7_75t_L g9514 ( 
.A1(n_9227),
.A2(n_686),
.B(n_687),
.C(n_685),
.Y(n_9514)
);

OAI22xp5_ASAP7_75t_L g9515 ( 
.A1(n_9211),
.A2(n_686),
.B1(n_684),
.B2(n_685),
.Y(n_9515)
);

OR2x2_ASAP7_75t_L g9516 ( 
.A(n_9059),
.B(n_685),
.Y(n_9516)
);

OAI33xp33_ASAP7_75t_L g9517 ( 
.A1(n_9126),
.A2(n_688),
.A3(n_690),
.B1(n_686),
.B2(n_687),
.B3(n_689),
.Y(n_9517)
);

AOI33xp33_ASAP7_75t_L g9518 ( 
.A1(n_9181),
.A2(n_689),
.A3(n_691),
.B1(n_687),
.B2(n_688),
.B3(n_690),
.Y(n_9518)
);

NAND3xp33_ASAP7_75t_L g9519 ( 
.A(n_9272),
.B(n_689),
.C(n_690),
.Y(n_9519)
);

INVx1_ASAP7_75t_L g9520 ( 
.A(n_9289),
.Y(n_9520)
);

NAND2xp5_ASAP7_75t_L g9521 ( 
.A(n_9207),
.B(n_9100),
.Y(n_9521)
);

OAI211xp5_ASAP7_75t_L g9522 ( 
.A1(n_9218),
.A2(n_699),
.B(n_707),
.C(n_691),
.Y(n_9522)
);

INVx2_ASAP7_75t_L g9523 ( 
.A(n_9060),
.Y(n_9523)
);

INVx1_ASAP7_75t_L g9524 ( 
.A(n_9290),
.Y(n_9524)
);

OAI22xp5_ASAP7_75t_L g9525 ( 
.A1(n_9219),
.A2(n_693),
.B1(n_691),
.B2(n_692),
.Y(n_9525)
);

AOI22xp5_ASAP7_75t_L g9526 ( 
.A1(n_9272),
.A2(n_694),
.B1(n_692),
.B2(n_693),
.Y(n_9526)
);

AOI22xp33_ASAP7_75t_SL g9527 ( 
.A1(n_9269),
.A2(n_695),
.B1(n_693),
.B2(n_694),
.Y(n_9527)
);

INVx2_ASAP7_75t_L g9528 ( 
.A(n_9061),
.Y(n_9528)
);

AOI221xp5_ASAP7_75t_L g9529 ( 
.A1(n_9205),
.A2(n_696),
.B1(n_694),
.B2(n_695),
.C(n_697),
.Y(n_9529)
);

OAI22xp33_ASAP7_75t_L g9530 ( 
.A1(n_9245),
.A2(n_697),
.B1(n_695),
.B2(n_696),
.Y(n_9530)
);

INVx2_ASAP7_75t_L g9531 ( 
.A(n_9072),
.Y(n_9531)
);

AND2x2_ASAP7_75t_L g9532 ( 
.A(n_9069),
.B(n_696),
.Y(n_9532)
);

AO21x2_ASAP7_75t_L g9533 ( 
.A1(n_9071),
.A2(n_698),
.B(n_699),
.Y(n_9533)
);

INVx2_ASAP7_75t_L g9534 ( 
.A(n_9111),
.Y(n_9534)
);

AOI22xp33_ASAP7_75t_L g9535 ( 
.A1(n_9233),
.A2(n_700),
.B1(n_698),
.B2(n_699),
.Y(n_9535)
);

AOI22xp5_ASAP7_75t_L g9536 ( 
.A1(n_9234),
.A2(n_702),
.B1(n_698),
.B2(n_701),
.Y(n_9536)
);

AND2x2_ASAP7_75t_L g9537 ( 
.A(n_9074),
.B(n_701),
.Y(n_9537)
);

OAI22xp5_ASAP7_75t_L g9538 ( 
.A1(n_9120),
.A2(n_703),
.B1(n_701),
.B2(n_702),
.Y(n_9538)
);

AOI22xp33_ASAP7_75t_L g9539 ( 
.A1(n_9217),
.A2(n_704),
.B1(n_702),
.B2(n_703),
.Y(n_9539)
);

OAI33xp33_ASAP7_75t_L g9540 ( 
.A1(n_9293),
.A2(n_9313),
.A3(n_9305),
.B1(n_9310),
.B2(n_9307),
.B3(n_9321),
.Y(n_9540)
);

AND2x2_ASAP7_75t_L g9541 ( 
.A(n_9081),
.B(n_704),
.Y(n_9541)
);

AND2x4_ASAP7_75t_L g9542 ( 
.A(n_9041),
.B(n_704),
.Y(n_9542)
);

OAI22xp33_ASAP7_75t_L g9543 ( 
.A1(n_9263),
.A2(n_707),
.B1(n_705),
.B2(n_706),
.Y(n_9543)
);

OAI211xp5_ASAP7_75t_L g9544 ( 
.A1(n_9225),
.A2(n_714),
.B(n_722),
.C(n_705),
.Y(n_9544)
);

AOI22xp33_ASAP7_75t_L g9545 ( 
.A1(n_9274),
.A2(n_709),
.B1(n_706),
.B2(n_708),
.Y(n_9545)
);

AOI22xp33_ASAP7_75t_L g9546 ( 
.A1(n_9279),
.A2(n_710),
.B1(n_708),
.B2(n_709),
.Y(n_9546)
);

OAI21x1_ASAP7_75t_L g9547 ( 
.A1(n_9115),
.A2(n_708),
.B(n_709),
.Y(n_9547)
);

OAI22xp33_ASAP7_75t_L g9548 ( 
.A1(n_9128),
.A2(n_712),
.B1(n_710),
.B2(n_711),
.Y(n_9548)
);

OAI22xp5_ASAP7_75t_L g9549 ( 
.A1(n_9131),
.A2(n_713),
.B1(n_711),
.B2(n_712),
.Y(n_9549)
);

INVx2_ASAP7_75t_L g9550 ( 
.A(n_9132),
.Y(n_9550)
);

NAND2x1p5_ASAP7_75t_L g9551 ( 
.A(n_9291),
.B(n_713),
.Y(n_9551)
);

NOR2x1_ASAP7_75t_L g9552 ( 
.A(n_9292),
.B(n_9297),
.Y(n_9552)
);

AOI22xp33_ASAP7_75t_L g9553 ( 
.A1(n_9226),
.A2(n_715),
.B1(n_712),
.B2(n_714),
.Y(n_9553)
);

INVx2_ASAP7_75t_L g9554 ( 
.A(n_9093),
.Y(n_9554)
);

OAI22xp33_ASAP7_75t_L g9555 ( 
.A1(n_9112),
.A2(n_9332),
.B1(n_9103),
.B2(n_9102),
.Y(n_9555)
);

INVx1_ASAP7_75t_L g9556 ( 
.A(n_9101),
.Y(n_9556)
);

INVx1_ASAP7_75t_SL g9557 ( 
.A(n_9309),
.Y(n_9557)
);

NOR2xp33_ASAP7_75t_L g9558 ( 
.A(n_9057),
.B(n_715),
.Y(n_9558)
);

OAI21xp33_ASAP7_75t_L g9559 ( 
.A1(n_9286),
.A2(n_716),
.B(n_717),
.Y(n_9559)
);

OAI22xp33_ASAP7_75t_L g9560 ( 
.A1(n_9119),
.A2(n_718),
.B1(n_716),
.B2(n_717),
.Y(n_9560)
);

INVx2_ASAP7_75t_SL g9561 ( 
.A(n_9311),
.Y(n_9561)
);

INVx1_ASAP7_75t_L g9562 ( 
.A(n_9133),
.Y(n_9562)
);

INVx1_ASAP7_75t_L g9563 ( 
.A(n_9089),
.Y(n_9563)
);

INVx1_ASAP7_75t_L g9564 ( 
.A(n_9318),
.Y(n_9564)
);

OAI221xp5_ASAP7_75t_SL g9565 ( 
.A1(n_9243),
.A2(n_719),
.B1(n_721),
.B2(n_718),
.C(n_720),
.Y(n_9565)
);

NOR2xp33_ASAP7_75t_L g9566 ( 
.A(n_9304),
.B(n_717),
.Y(n_9566)
);

INVx1_ASAP7_75t_L g9567 ( 
.A(n_9319),
.Y(n_9567)
);

OAI221xp5_ASAP7_75t_L g9568 ( 
.A1(n_9316),
.A2(n_721),
.B1(n_719),
.B2(n_720),
.C(n_722),
.Y(n_9568)
);

AOI22xp33_ASAP7_75t_L g9569 ( 
.A1(n_9260),
.A2(n_721),
.B1(n_719),
.B2(n_720),
.Y(n_9569)
);

BUFx3_ASAP7_75t_L g9570 ( 
.A(n_9116),
.Y(n_9570)
);

NOR2xp33_ASAP7_75t_L g9571 ( 
.A(n_9065),
.B(n_723),
.Y(n_9571)
);

AOI21xp33_ASAP7_75t_L g9572 ( 
.A1(n_9235),
.A2(n_723),
.B(n_724),
.Y(n_9572)
);

INVx2_ASAP7_75t_L g9573 ( 
.A(n_9094),
.Y(n_9573)
);

NAND3xp33_ASAP7_75t_L g9574 ( 
.A(n_9248),
.B(n_723),
.C(n_724),
.Y(n_9574)
);

AOI22xp33_ASAP7_75t_SL g9575 ( 
.A1(n_9193),
.A2(n_726),
.B1(n_724),
.B2(n_725),
.Y(n_9575)
);

OAI221xp5_ASAP7_75t_L g9576 ( 
.A1(n_9086),
.A2(n_727),
.B1(n_725),
.B2(n_726),
.C(n_728),
.Y(n_9576)
);

NAND2xp5_ASAP7_75t_L g9577 ( 
.A(n_9322),
.B(n_725),
.Y(n_9577)
);

INVx2_ASAP7_75t_L g9578 ( 
.A(n_9122),
.Y(n_9578)
);

INVx1_ASAP7_75t_L g9579 ( 
.A(n_9328),
.Y(n_9579)
);

OR2x6_ASAP7_75t_L g9580 ( 
.A(n_9330),
.B(n_727),
.Y(n_9580)
);

AO22x1_ASAP7_75t_L g9581 ( 
.A1(n_9333),
.A2(n_729),
.B1(n_727),
.B2(n_728),
.Y(n_9581)
);

INVx1_ASAP7_75t_L g9582 ( 
.A(n_9050),
.Y(n_9582)
);

AOI221xp5_ASAP7_75t_L g9583 ( 
.A1(n_9117),
.A2(n_730),
.B1(n_728),
.B2(n_729),
.C(n_731),
.Y(n_9583)
);

INVx1_ASAP7_75t_SL g9584 ( 
.A(n_9135),
.Y(n_9584)
);

OAI21x1_ASAP7_75t_L g9585 ( 
.A1(n_9136),
.A2(n_729),
.B(n_730),
.Y(n_9585)
);

AND2x2_ASAP7_75t_L g9586 ( 
.A(n_9161),
.B(n_731),
.Y(n_9586)
);

AND2x2_ASAP7_75t_L g9587 ( 
.A(n_9114),
.B(n_731),
.Y(n_9587)
);

OAI211xp5_ASAP7_75t_L g9588 ( 
.A1(n_9177),
.A2(n_740),
.B(n_748),
.C(n_732),
.Y(n_9588)
);

AOI222xp33_ASAP7_75t_L g9589 ( 
.A1(n_9184),
.A2(n_734),
.B1(n_736),
.B2(n_732),
.C1(n_733),
.C2(n_735),
.Y(n_9589)
);

OAI221xp5_ASAP7_75t_SL g9590 ( 
.A1(n_9163),
.A2(n_735),
.B1(n_737),
.B2(n_734),
.C(n_736),
.Y(n_9590)
);

AND2x2_ASAP7_75t_L g9591 ( 
.A(n_9118),
.B(n_733),
.Y(n_9591)
);

OAI22xp5_ASAP7_75t_L g9592 ( 
.A1(n_9160),
.A2(n_735),
.B1(n_733),
.B2(n_734),
.Y(n_9592)
);

OA21x2_ASAP7_75t_L g9593 ( 
.A1(n_9162),
.A2(n_736),
.B(n_738),
.Y(n_9593)
);

OAI211xp5_ASAP7_75t_SL g9594 ( 
.A1(n_9258),
.A2(n_741),
.B(n_739),
.C(n_740),
.Y(n_9594)
);

AOI22xp33_ASAP7_75t_SL g9595 ( 
.A1(n_9199),
.A2(n_741),
.B1(n_739),
.B2(n_740),
.Y(n_9595)
);

OAI22xp5_ASAP7_75t_L g9596 ( 
.A1(n_9199),
.A2(n_742),
.B1(n_739),
.B2(n_741),
.Y(n_9596)
);

OR2x2_ASAP7_75t_L g9597 ( 
.A(n_9288),
.B(n_742),
.Y(n_9597)
);

AND2x2_ASAP7_75t_L g9598 ( 
.A(n_9139),
.B(n_742),
.Y(n_9598)
);

NAND2xp5_ASAP7_75t_L g9599 ( 
.A(n_9223),
.B(n_743),
.Y(n_9599)
);

AOI22xp33_ASAP7_75t_L g9600 ( 
.A1(n_9246),
.A2(n_745),
.B1(n_743),
.B2(n_744),
.Y(n_9600)
);

INVx1_ASAP7_75t_L g9601 ( 
.A(n_9035),
.Y(n_9601)
);

AOI322xp5_ASAP7_75t_L g9602 ( 
.A1(n_9258),
.A2(n_749),
.A3(n_748),
.B1(n_746),
.B2(n_744),
.C1(n_745),
.C2(n_747),
.Y(n_9602)
);

OAI211xp5_ASAP7_75t_SL g9603 ( 
.A1(n_9258),
.A2(n_748),
.B(n_744),
.C(n_746),
.Y(n_9603)
);

AOI22xp33_ASAP7_75t_SL g9604 ( 
.A1(n_9199),
.A2(n_751),
.B1(n_749),
.B2(n_750),
.Y(n_9604)
);

AND2x2_ASAP7_75t_L g9605 ( 
.A(n_9139),
.B(n_750),
.Y(n_9605)
);

INVx3_ASAP7_75t_L g9606 ( 
.A(n_9037),
.Y(n_9606)
);

AOI22xp33_ASAP7_75t_L g9607 ( 
.A1(n_9246),
.A2(n_753),
.B1(n_750),
.B2(n_752),
.Y(n_9607)
);

OAI33xp33_ASAP7_75t_L g9608 ( 
.A1(n_9171),
.A2(n_755),
.A3(n_757),
.B1(n_752),
.B2(n_753),
.B3(n_756),
.Y(n_9608)
);

OAI22xp5_ASAP7_75t_L g9609 ( 
.A1(n_9199),
.A2(n_756),
.B1(n_753),
.B2(n_755),
.Y(n_9609)
);

AOI221xp5_ASAP7_75t_L g9610 ( 
.A1(n_9246),
.A2(n_757),
.B1(n_755),
.B2(n_756),
.C(n_758),
.Y(n_9610)
);

OAI22xp33_ASAP7_75t_L g9611 ( 
.A1(n_9139),
.A2(n_759),
.B1(n_757),
.B2(n_758),
.Y(n_9611)
);

AND2x2_ASAP7_75t_L g9612 ( 
.A(n_9139),
.B(n_759),
.Y(n_9612)
);

NAND2xp5_ASAP7_75t_L g9613 ( 
.A(n_9223),
.B(n_760),
.Y(n_9613)
);

BUFx6f_ASAP7_75t_L g9614 ( 
.A(n_9037),
.Y(n_9614)
);

INVx2_ASAP7_75t_L g9615 ( 
.A(n_9063),
.Y(n_9615)
);

AND2x2_ASAP7_75t_L g9616 ( 
.A(n_9139),
.B(n_760),
.Y(n_9616)
);

AOI22xp33_ASAP7_75t_L g9617 ( 
.A1(n_9246),
.A2(n_763),
.B1(n_761),
.B2(n_762),
.Y(n_9617)
);

OAI31xp33_ASAP7_75t_L g9618 ( 
.A1(n_9049),
.A2(n_764),
.A3(n_765),
.B(n_763),
.Y(n_9618)
);

INVx1_ASAP7_75t_L g9619 ( 
.A(n_9035),
.Y(n_9619)
);

NAND2xp5_ASAP7_75t_L g9620 ( 
.A(n_9223),
.B(n_761),
.Y(n_9620)
);

OAI211xp5_ASAP7_75t_L g9621 ( 
.A1(n_9258),
.A2(n_772),
.B(n_780),
.C(n_764),
.Y(n_9621)
);

OAI31xp33_ASAP7_75t_L g9622 ( 
.A1(n_9049),
.A2(n_766),
.A3(n_767),
.B(n_765),
.Y(n_9622)
);

BUFx3_ASAP7_75t_L g9623 ( 
.A(n_9301),
.Y(n_9623)
);

OA21x2_ASAP7_75t_L g9624 ( 
.A1(n_9171),
.A2(n_764),
.B(n_765),
.Y(n_9624)
);

NAND2xp5_ASAP7_75t_L g9625 ( 
.A(n_9223),
.B(n_766),
.Y(n_9625)
);

HB1xp67_ASAP7_75t_L g9626 ( 
.A(n_9040),
.Y(n_9626)
);

OR2x2_ASAP7_75t_L g9627 ( 
.A(n_9288),
.B(n_766),
.Y(n_9627)
);

OAI211xp5_ASAP7_75t_L g9628 ( 
.A1(n_9258),
.A2(n_775),
.B(n_783),
.C(n_767),
.Y(n_9628)
);

BUFx2_ASAP7_75t_L g9629 ( 
.A(n_9182),
.Y(n_9629)
);

NAND2xp5_ASAP7_75t_L g9630 ( 
.A(n_9223),
.B(n_767),
.Y(n_9630)
);

OAI31xp33_ASAP7_75t_L g9631 ( 
.A1(n_9049),
.A2(n_770),
.A3(n_771),
.B(n_769),
.Y(n_9631)
);

AOI31xp33_ASAP7_75t_L g9632 ( 
.A1(n_9258),
.A2(n_770),
.A3(n_768),
.B(n_769),
.Y(n_9632)
);

AOI21x1_ASAP7_75t_L g9633 ( 
.A1(n_9182),
.A2(n_768),
.B(n_769),
.Y(n_9633)
);

OAI33xp33_ASAP7_75t_L g9634 ( 
.A1(n_9171),
.A2(n_772),
.A3(n_774),
.B1(n_768),
.B2(n_771),
.B3(n_773),
.Y(n_9634)
);

INVx2_ASAP7_75t_L g9635 ( 
.A(n_9063),
.Y(n_9635)
);

AOI21xp5_ASAP7_75t_L g9636 ( 
.A1(n_9258),
.A2(n_771),
.B(n_772),
.Y(n_9636)
);

INVx2_ASAP7_75t_L g9637 ( 
.A(n_9063),
.Y(n_9637)
);

AOI221xp5_ASAP7_75t_L g9638 ( 
.A1(n_9246),
.A2(n_776),
.B1(n_773),
.B2(n_775),
.C(n_777),
.Y(n_9638)
);

OAI31xp33_ASAP7_75t_L g9639 ( 
.A1(n_9049),
.A2(n_777),
.A3(n_778),
.B(n_776),
.Y(n_9639)
);

A2O1A1Ixp33_ASAP7_75t_L g9640 ( 
.A1(n_9258),
.A2(n_777),
.B(n_778),
.C(n_776),
.Y(n_9640)
);

AOI22xp5_ASAP7_75t_L g9641 ( 
.A1(n_9258),
.A2(n_779),
.B1(n_773),
.B2(n_778),
.Y(n_9641)
);

AND2x2_ASAP7_75t_L g9642 ( 
.A(n_9139),
.B(n_779),
.Y(n_9642)
);

NAND4xp25_ASAP7_75t_SL g9643 ( 
.A(n_9258),
.B(n_782),
.C(n_780),
.D(n_781),
.Y(n_9643)
);

INVx1_ASAP7_75t_L g9644 ( 
.A(n_9035),
.Y(n_9644)
);

OAI22xp5_ASAP7_75t_L g9645 ( 
.A1(n_9199),
.A2(n_782),
.B1(n_780),
.B2(n_781),
.Y(n_9645)
);

INVx2_ASAP7_75t_L g9646 ( 
.A(n_9063),
.Y(n_9646)
);

OAI31xp33_ASAP7_75t_L g9647 ( 
.A1(n_9049),
.A2(n_783),
.A3(n_784),
.B(n_782),
.Y(n_9647)
);

OR2x6_ASAP7_75t_L g9648 ( 
.A(n_9182),
.B(n_781),
.Y(n_9648)
);

AOI33xp33_ASAP7_75t_L g9649 ( 
.A1(n_9033),
.A2(n_785),
.A3(n_788),
.B1(n_783),
.B2(n_784),
.B3(n_786),
.Y(n_9649)
);

OAI21xp5_ASAP7_75t_SL g9650 ( 
.A1(n_9258),
.A2(n_788),
.B(n_786),
.Y(n_9650)
);

INVx1_ASAP7_75t_L g9651 ( 
.A(n_9035),
.Y(n_9651)
);

AOI22xp33_ASAP7_75t_L g9652 ( 
.A1(n_9246),
.A2(n_789),
.B1(n_784),
.B2(n_788),
.Y(n_9652)
);

AND2x4_ASAP7_75t_L g9653 ( 
.A(n_9063),
.B(n_789),
.Y(n_9653)
);

AO21x2_ASAP7_75t_L g9654 ( 
.A1(n_9032),
.A2(n_790),
.B(n_791),
.Y(n_9654)
);

NOR2xp33_ASAP7_75t_SL g9655 ( 
.A(n_9643),
.B(n_790),
.Y(n_9655)
);

INVx1_ASAP7_75t_L g9656 ( 
.A(n_9424),
.Y(n_9656)
);

INVx1_ASAP7_75t_L g9657 ( 
.A(n_9438),
.Y(n_9657)
);

AND2x2_ASAP7_75t_L g9658 ( 
.A(n_9629),
.B(n_790),
.Y(n_9658)
);

HB1xp67_ASAP7_75t_L g9659 ( 
.A(n_9353),
.Y(n_9659)
);

INVx1_ASAP7_75t_L g9660 ( 
.A(n_9516),
.Y(n_9660)
);

INVx2_ASAP7_75t_L g9661 ( 
.A(n_9430),
.Y(n_9661)
);

OR2x2_ASAP7_75t_L g9662 ( 
.A(n_9393),
.B(n_791),
.Y(n_9662)
);

INVx1_ASAP7_75t_L g9663 ( 
.A(n_9626),
.Y(n_9663)
);

INVx1_ASAP7_75t_L g9664 ( 
.A(n_9562),
.Y(n_9664)
);

INVx1_ASAP7_75t_L g9665 ( 
.A(n_9556),
.Y(n_9665)
);

INVx1_ASAP7_75t_L g9666 ( 
.A(n_9344),
.Y(n_9666)
);

OR2x2_ASAP7_75t_L g9667 ( 
.A(n_9557),
.B(n_792),
.Y(n_9667)
);

HB1xp67_ASAP7_75t_L g9668 ( 
.A(n_9458),
.Y(n_9668)
);

INVx2_ASAP7_75t_L g9669 ( 
.A(n_9343),
.Y(n_9669)
);

NAND2xp5_ASAP7_75t_L g9670 ( 
.A(n_9340),
.B(n_9404),
.Y(n_9670)
);

HB1xp67_ASAP7_75t_L g9671 ( 
.A(n_9552),
.Y(n_9671)
);

AND2x2_ASAP7_75t_L g9672 ( 
.A(n_9346),
.B(n_792),
.Y(n_9672)
);

INVx1_ASAP7_75t_L g9673 ( 
.A(n_9354),
.Y(n_9673)
);

AND2x2_ASAP7_75t_L g9674 ( 
.A(n_9387),
.B(n_792),
.Y(n_9674)
);

INVx1_ASAP7_75t_L g9675 ( 
.A(n_9371),
.Y(n_9675)
);

HB1xp67_ASAP7_75t_L g9676 ( 
.A(n_9561),
.Y(n_9676)
);

NOR2x1_ASAP7_75t_L g9677 ( 
.A(n_9654),
.B(n_793),
.Y(n_9677)
);

INVx1_ASAP7_75t_L g9678 ( 
.A(n_9390),
.Y(n_9678)
);

INVx1_ASAP7_75t_L g9679 ( 
.A(n_9392),
.Y(n_9679)
);

AND2x2_ASAP7_75t_L g9680 ( 
.A(n_9606),
.B(n_793),
.Y(n_9680)
);

AND2x2_ASAP7_75t_L g9681 ( 
.A(n_9348),
.B(n_793),
.Y(n_9681)
);

INVx1_ASAP7_75t_L g9682 ( 
.A(n_9425),
.Y(n_9682)
);

INVx1_ASAP7_75t_L g9683 ( 
.A(n_9429),
.Y(n_9683)
);

AND2x2_ASAP7_75t_SL g9684 ( 
.A(n_9417),
.B(n_794),
.Y(n_9684)
);

AOI22xp33_ASAP7_75t_L g9685 ( 
.A1(n_9389),
.A2(n_796),
.B1(n_794),
.B2(n_795),
.Y(n_9685)
);

INVx2_ASAP7_75t_L g9686 ( 
.A(n_9356),
.Y(n_9686)
);

OR2x2_ASAP7_75t_L g9687 ( 
.A(n_9584),
.B(n_794),
.Y(n_9687)
);

OR2x2_ASAP7_75t_L g9688 ( 
.A(n_9521),
.B(n_9391),
.Y(n_9688)
);

AND2x2_ASAP7_75t_L g9689 ( 
.A(n_9342),
.B(n_9615),
.Y(n_9689)
);

INVx2_ASAP7_75t_L g9690 ( 
.A(n_9623),
.Y(n_9690)
);

AND2x2_ASAP7_75t_L g9691 ( 
.A(n_9635),
.B(n_795),
.Y(n_9691)
);

AND2x2_ASAP7_75t_L g9692 ( 
.A(n_9637),
.B(n_795),
.Y(n_9692)
);

INVx1_ASAP7_75t_L g9693 ( 
.A(n_9435),
.Y(n_9693)
);

INVxp67_ASAP7_75t_SL g9694 ( 
.A(n_9478),
.Y(n_9694)
);

HB1xp67_ASAP7_75t_L g9695 ( 
.A(n_9470),
.Y(n_9695)
);

INVxp67_ASAP7_75t_SL g9696 ( 
.A(n_9406),
.Y(n_9696)
);

AND2x4_ASAP7_75t_L g9697 ( 
.A(n_9646),
.B(n_796),
.Y(n_9697)
);

INVx2_ASAP7_75t_L g9698 ( 
.A(n_9614),
.Y(n_9698)
);

OR2x2_ASAP7_75t_L g9699 ( 
.A(n_9350),
.B(n_797),
.Y(n_9699)
);

AND2x2_ASAP7_75t_L g9700 ( 
.A(n_9412),
.B(n_9370),
.Y(n_9700)
);

INVx1_ASAP7_75t_L g9701 ( 
.A(n_9437),
.Y(n_9701)
);

INVx2_ASAP7_75t_L g9702 ( 
.A(n_9614),
.Y(n_9702)
);

AND2x2_ASAP7_75t_L g9703 ( 
.A(n_9578),
.B(n_797),
.Y(n_9703)
);

BUFx2_ASAP7_75t_L g9704 ( 
.A(n_9648),
.Y(n_9704)
);

INVx1_ASAP7_75t_L g9705 ( 
.A(n_9440),
.Y(n_9705)
);

INVx1_ASAP7_75t_L g9706 ( 
.A(n_9452),
.Y(n_9706)
);

BUFx3_ASAP7_75t_L g9707 ( 
.A(n_9427),
.Y(n_9707)
);

OR2x2_ASAP7_75t_L g9708 ( 
.A(n_9582),
.B(n_798),
.Y(n_9708)
);

INVx1_ASAP7_75t_L g9709 ( 
.A(n_9456),
.Y(n_9709)
);

AND2x2_ASAP7_75t_L g9710 ( 
.A(n_9364),
.B(n_799),
.Y(n_9710)
);

INVx2_ASAP7_75t_L g9711 ( 
.A(n_9427),
.Y(n_9711)
);

AND2x4_ASAP7_75t_L g9712 ( 
.A(n_9570),
.B(n_799),
.Y(n_9712)
);

OR2x2_ASAP7_75t_L g9713 ( 
.A(n_9564),
.B(n_800),
.Y(n_9713)
);

OR2x2_ASAP7_75t_L g9714 ( 
.A(n_9567),
.B(n_800),
.Y(n_9714)
);

AND2x2_ASAP7_75t_L g9715 ( 
.A(n_9573),
.B(n_9476),
.Y(n_9715)
);

INVx1_ASAP7_75t_L g9716 ( 
.A(n_9457),
.Y(n_9716)
);

INVx2_ASAP7_75t_L g9717 ( 
.A(n_9512),
.Y(n_9717)
);

OR2x2_ASAP7_75t_L g9718 ( 
.A(n_9579),
.B(n_801),
.Y(n_9718)
);

NAND2xp5_ASAP7_75t_L g9719 ( 
.A(n_9598),
.B(n_801),
.Y(n_9719)
);

AND2x2_ASAP7_75t_L g9720 ( 
.A(n_9464),
.B(n_9563),
.Y(n_9720)
);

NAND2xp5_ASAP7_75t_L g9721 ( 
.A(n_9605),
.B(n_9612),
.Y(n_9721)
);

NAND2xp5_ASAP7_75t_L g9722 ( 
.A(n_9616),
.B(n_801),
.Y(n_9722)
);

AND2x4_ASAP7_75t_L g9723 ( 
.A(n_9468),
.B(n_802),
.Y(n_9723)
);

HB1xp67_ASAP7_75t_L g9724 ( 
.A(n_9492),
.Y(n_9724)
);

INVx2_ASAP7_75t_L g9725 ( 
.A(n_9501),
.Y(n_9725)
);

INVxp67_ASAP7_75t_SL g9726 ( 
.A(n_9338),
.Y(n_9726)
);

INVx2_ASAP7_75t_L g9727 ( 
.A(n_9471),
.Y(n_9727)
);

INVx1_ASAP7_75t_L g9728 ( 
.A(n_9460),
.Y(n_9728)
);

INVx1_ASAP7_75t_L g9729 ( 
.A(n_9462),
.Y(n_9729)
);

AND2x4_ASAP7_75t_L g9730 ( 
.A(n_9482),
.B(n_802),
.Y(n_9730)
);

NOR2x1_ASAP7_75t_SL g9731 ( 
.A(n_9633),
.B(n_9482),
.Y(n_9731)
);

INVx1_ASAP7_75t_L g9732 ( 
.A(n_9475),
.Y(n_9732)
);

INVx1_ASAP7_75t_L g9733 ( 
.A(n_9487),
.Y(n_9733)
);

INVx1_ASAP7_75t_L g9734 ( 
.A(n_9493),
.Y(n_9734)
);

AND2x2_ASAP7_75t_L g9735 ( 
.A(n_9642),
.B(n_804),
.Y(n_9735)
);

AND2x2_ASAP7_75t_L g9736 ( 
.A(n_9505),
.B(n_804),
.Y(n_9736)
);

OR2x2_ASAP7_75t_L g9737 ( 
.A(n_9513),
.B(n_805),
.Y(n_9737)
);

AND2x4_ASAP7_75t_L g9738 ( 
.A(n_9413),
.B(n_9420),
.Y(n_9738)
);

HB1xp67_ASAP7_75t_L g9739 ( 
.A(n_9492),
.Y(n_9739)
);

INVx2_ASAP7_75t_L g9740 ( 
.A(n_9648),
.Y(n_9740)
);

INVx2_ASAP7_75t_L g9741 ( 
.A(n_9336),
.Y(n_9741)
);

OR2x2_ASAP7_75t_L g9742 ( 
.A(n_9422),
.B(n_805),
.Y(n_9742)
);

HB1xp67_ASAP7_75t_L g9743 ( 
.A(n_9352),
.Y(n_9743)
);

INVx2_ASAP7_75t_L g9744 ( 
.A(n_9386),
.Y(n_9744)
);

INVx1_ASAP7_75t_L g9745 ( 
.A(n_9495),
.Y(n_9745)
);

AND2x2_ASAP7_75t_L g9746 ( 
.A(n_9428),
.B(n_806),
.Y(n_9746)
);

NOR2xp67_ASAP7_75t_L g9747 ( 
.A(n_9636),
.B(n_806),
.Y(n_9747)
);

INVx1_ASAP7_75t_L g9748 ( 
.A(n_9508),
.Y(n_9748)
);

INVx2_ASAP7_75t_L g9749 ( 
.A(n_9597),
.Y(n_9749)
);

INVx1_ASAP7_75t_L g9750 ( 
.A(n_9520),
.Y(n_9750)
);

INVx1_ASAP7_75t_SL g9751 ( 
.A(n_9402),
.Y(n_9751)
);

NAND2xp5_ASAP7_75t_L g9752 ( 
.A(n_9398),
.B(n_806),
.Y(n_9752)
);

INVx1_ASAP7_75t_L g9753 ( 
.A(n_9524),
.Y(n_9753)
);

INVx3_ASAP7_75t_L g9754 ( 
.A(n_9653),
.Y(n_9754)
);

AND2x4_ASAP7_75t_L g9755 ( 
.A(n_9481),
.B(n_807),
.Y(n_9755)
);

HB1xp67_ASAP7_75t_L g9756 ( 
.A(n_9375),
.Y(n_9756)
);

BUFx2_ASAP7_75t_L g9757 ( 
.A(n_9409),
.Y(n_9757)
);

HB1xp67_ASAP7_75t_L g9758 ( 
.A(n_9624),
.Y(n_9758)
);

AND2x2_ASAP7_75t_L g9759 ( 
.A(n_9362),
.B(n_807),
.Y(n_9759)
);

AND2x4_ASAP7_75t_L g9760 ( 
.A(n_9445),
.B(n_807),
.Y(n_9760)
);

AND2x2_ASAP7_75t_L g9761 ( 
.A(n_9359),
.B(n_808),
.Y(n_9761)
);

NAND3xp33_ASAP7_75t_L g9762 ( 
.A(n_9595),
.B(n_808),
.C(n_809),
.Y(n_9762)
);

INVx3_ASAP7_75t_L g9763 ( 
.A(n_9383),
.Y(n_9763)
);

INVx2_ASAP7_75t_L g9764 ( 
.A(n_9627),
.Y(n_9764)
);

AND2x2_ASAP7_75t_L g9765 ( 
.A(n_9467),
.B(n_808),
.Y(n_9765)
);

AND2x2_ASAP7_75t_L g9766 ( 
.A(n_9504),
.B(n_809),
.Y(n_9766)
);

AND2x2_ASAP7_75t_L g9767 ( 
.A(n_9479),
.B(n_810),
.Y(n_9767)
);

INVx1_ASAP7_75t_L g9768 ( 
.A(n_9601),
.Y(n_9768)
);

OR2x2_ASAP7_75t_L g9769 ( 
.A(n_9473),
.B(n_810),
.Y(n_9769)
);

INVx1_ASAP7_75t_L g9770 ( 
.A(n_9619),
.Y(n_9770)
);

NAND2x1p5_ASAP7_75t_L g9771 ( 
.A(n_9593),
.B(n_810),
.Y(n_9771)
);

INVx1_ASAP7_75t_SL g9772 ( 
.A(n_9395),
.Y(n_9772)
);

AND2x2_ASAP7_75t_L g9773 ( 
.A(n_9358),
.B(n_811),
.Y(n_9773)
);

INVx2_ASAP7_75t_L g9774 ( 
.A(n_9377),
.Y(n_9774)
);

BUFx2_ASAP7_75t_L g9775 ( 
.A(n_9580),
.Y(n_9775)
);

AND2x2_ASAP7_75t_L g9776 ( 
.A(n_9369),
.B(n_811),
.Y(n_9776)
);

AND2x2_ASAP7_75t_L g9777 ( 
.A(n_9488),
.B(n_811),
.Y(n_9777)
);

HB1xp67_ASAP7_75t_L g9778 ( 
.A(n_9510),
.Y(n_9778)
);

AND2x2_ASAP7_75t_L g9779 ( 
.A(n_9502),
.B(n_812),
.Y(n_9779)
);

AND2x2_ASAP7_75t_L g9780 ( 
.A(n_9378),
.B(n_812),
.Y(n_9780)
);

BUFx2_ASAP7_75t_L g9781 ( 
.A(n_9580),
.Y(n_9781)
);

NAND2xp5_ASAP7_75t_L g9782 ( 
.A(n_9337),
.B(n_812),
.Y(n_9782)
);

INVxp67_ASAP7_75t_L g9783 ( 
.A(n_9533),
.Y(n_9783)
);

INVx1_ASAP7_75t_L g9784 ( 
.A(n_9644),
.Y(n_9784)
);

NAND2xp5_ASAP7_75t_L g9785 ( 
.A(n_9439),
.B(n_9604),
.Y(n_9785)
);

NAND2xp5_ASAP7_75t_L g9786 ( 
.A(n_9347),
.B(n_813),
.Y(n_9786)
);

NAND2xp5_ASAP7_75t_L g9787 ( 
.A(n_9372),
.B(n_813),
.Y(n_9787)
);

INVx1_ASAP7_75t_L g9788 ( 
.A(n_9651),
.Y(n_9788)
);

AND2x2_ASAP7_75t_L g9789 ( 
.A(n_9380),
.B(n_813),
.Y(n_9789)
);

INVx2_ASAP7_75t_L g9790 ( 
.A(n_9474),
.Y(n_9790)
);

OR2x2_ASAP7_75t_L g9791 ( 
.A(n_9401),
.B(n_814),
.Y(n_9791)
);

INVx2_ASAP7_75t_L g9792 ( 
.A(n_9489),
.Y(n_9792)
);

INVx4_ASAP7_75t_L g9793 ( 
.A(n_9441),
.Y(n_9793)
);

INVx2_ASAP7_75t_L g9794 ( 
.A(n_9523),
.Y(n_9794)
);

AND2x2_ASAP7_75t_L g9795 ( 
.A(n_9469),
.B(n_814),
.Y(n_9795)
);

INVx1_ASAP7_75t_L g9796 ( 
.A(n_9534),
.Y(n_9796)
);

AND2x4_ASAP7_75t_L g9797 ( 
.A(n_9434),
.B(n_814),
.Y(n_9797)
);

INVx1_ASAP7_75t_L g9798 ( 
.A(n_9550),
.Y(n_9798)
);

INVx2_ASAP7_75t_L g9799 ( 
.A(n_9528),
.Y(n_9799)
);

HB1xp67_ASAP7_75t_L g9800 ( 
.A(n_9510),
.Y(n_9800)
);

NAND2xp33_ASAP7_75t_R g9801 ( 
.A(n_9433),
.B(n_815),
.Y(n_9801)
);

AND2x2_ASAP7_75t_L g9802 ( 
.A(n_9531),
.B(n_816),
.Y(n_9802)
);

INVx3_ASAP7_75t_L g9803 ( 
.A(n_9494),
.Y(n_9803)
);

INVx1_ASAP7_75t_L g9804 ( 
.A(n_9554),
.Y(n_9804)
);

INVx1_ASAP7_75t_L g9805 ( 
.A(n_9448),
.Y(n_9805)
);

AND2x2_ASAP7_75t_L g9806 ( 
.A(n_9551),
.B(n_9532),
.Y(n_9806)
);

AND2x4_ASAP7_75t_L g9807 ( 
.A(n_9465),
.B(n_816),
.Y(n_9807)
);

INVx2_ASAP7_75t_L g9808 ( 
.A(n_9449),
.Y(n_9808)
);

AND2x2_ASAP7_75t_L g9809 ( 
.A(n_9537),
.B(n_816),
.Y(n_9809)
);

AND2x2_ASAP7_75t_L g9810 ( 
.A(n_9541),
.B(n_817),
.Y(n_9810)
);

INVx1_ASAP7_75t_L g9811 ( 
.A(n_9341),
.Y(n_9811)
);

INVx2_ASAP7_75t_SL g9812 ( 
.A(n_9542),
.Y(n_9812)
);

AND2x2_ASAP7_75t_L g9813 ( 
.A(n_9496),
.B(n_817),
.Y(n_9813)
);

INVx2_ASAP7_75t_L g9814 ( 
.A(n_9341),
.Y(n_9814)
);

BUFx3_ASAP7_75t_L g9815 ( 
.A(n_9587),
.Y(n_9815)
);

NAND2xp5_ASAP7_75t_L g9816 ( 
.A(n_9650),
.B(n_817),
.Y(n_9816)
);

INVx1_ASAP7_75t_L g9817 ( 
.A(n_9368),
.Y(n_9817)
);

AND2x2_ASAP7_75t_L g9818 ( 
.A(n_9586),
.B(n_818),
.Y(n_9818)
);

AND2x2_ASAP7_75t_L g9819 ( 
.A(n_9591),
.B(n_818),
.Y(n_9819)
);

AND2x2_ASAP7_75t_L g9820 ( 
.A(n_9585),
.B(n_818),
.Y(n_9820)
);

INVx1_ASAP7_75t_L g9821 ( 
.A(n_9507),
.Y(n_9821)
);

NAND2x1_ASAP7_75t_L g9822 ( 
.A(n_9632),
.B(n_819),
.Y(n_9822)
);

AND2x2_ASAP7_75t_L g9823 ( 
.A(n_9360),
.B(n_819),
.Y(n_9823)
);

INVx2_ASAP7_75t_L g9824 ( 
.A(n_9547),
.Y(n_9824)
);

INVx1_ASAP7_75t_L g9825 ( 
.A(n_9443),
.Y(n_9825)
);

NAND2xp5_ASAP7_75t_L g9826 ( 
.A(n_9405),
.B(n_819),
.Y(n_9826)
);

AND2x2_ASAP7_75t_L g9827 ( 
.A(n_9571),
.B(n_820),
.Y(n_9827)
);

INVx1_ASAP7_75t_SL g9828 ( 
.A(n_9472),
.Y(n_9828)
);

AND2x2_ASAP7_75t_L g9829 ( 
.A(n_9379),
.B(n_820),
.Y(n_9829)
);

NAND2xp5_ASAP7_75t_L g9830 ( 
.A(n_9581),
.B(n_821),
.Y(n_9830)
);

INVx1_ASAP7_75t_L g9831 ( 
.A(n_9466),
.Y(n_9831)
);

AND4x1_ASAP7_75t_L g9832 ( 
.A(n_9408),
.B(n_823),
.C(n_821),
.D(n_822),
.Y(n_9832)
);

INVx2_ASAP7_75t_L g9833 ( 
.A(n_9339),
.Y(n_9833)
);

AND2x2_ASAP7_75t_L g9834 ( 
.A(n_9432),
.B(n_9599),
.Y(n_9834)
);

AND2x2_ASAP7_75t_L g9835 ( 
.A(n_9613),
.B(n_822),
.Y(n_9835)
);

AND2x2_ASAP7_75t_L g9836 ( 
.A(n_9620),
.B(n_823),
.Y(n_9836)
);

NAND2xp5_ASAP7_75t_L g9837 ( 
.A(n_9451),
.B(n_9555),
.Y(n_9837)
);

INVx1_ASAP7_75t_L g9838 ( 
.A(n_9625),
.Y(n_9838)
);

HB1xp67_ASAP7_75t_L g9839 ( 
.A(n_9345),
.Y(n_9839)
);

INVx2_ASAP7_75t_L g9840 ( 
.A(n_9630),
.Y(n_9840)
);

INVx1_ASAP7_75t_L g9841 ( 
.A(n_9373),
.Y(n_9841)
);

INVx1_ASAP7_75t_L g9842 ( 
.A(n_9538),
.Y(n_9842)
);

AND2x2_ASAP7_75t_L g9843 ( 
.A(n_9400),
.B(n_824),
.Y(n_9843)
);

INVx1_ASAP7_75t_L g9844 ( 
.A(n_9577),
.Y(n_9844)
);

NAND2xp5_ASAP7_75t_L g9845 ( 
.A(n_9596),
.B(n_824),
.Y(n_9845)
);

INVx2_ASAP7_75t_SL g9846 ( 
.A(n_9503),
.Y(n_9846)
);

NAND2xp5_ASAP7_75t_L g9847 ( 
.A(n_9609),
.B(n_824),
.Y(n_9847)
);

INVx2_ASAP7_75t_L g9848 ( 
.A(n_9423),
.Y(n_9848)
);

AND2x2_ASAP7_75t_L g9849 ( 
.A(n_9418),
.B(n_825),
.Y(n_9849)
);

OR2x2_ASAP7_75t_L g9850 ( 
.A(n_9361),
.B(n_825),
.Y(n_9850)
);

NAND2xp5_ASAP7_75t_L g9851 ( 
.A(n_9645),
.B(n_825),
.Y(n_9851)
);

AND2x2_ASAP7_75t_L g9852 ( 
.A(n_9641),
.B(n_826),
.Y(n_9852)
);

INVx2_ASAP7_75t_L g9853 ( 
.A(n_9453),
.Y(n_9853)
);

INVx2_ASAP7_75t_L g9854 ( 
.A(n_9394),
.Y(n_9854)
);

HB1xp67_ASAP7_75t_L g9855 ( 
.A(n_9416),
.Y(n_9855)
);

INVx1_ASAP7_75t_L g9856 ( 
.A(n_9446),
.Y(n_9856)
);

NAND4xp25_ASAP7_75t_L g9857 ( 
.A(n_9610),
.B(n_828),
.C(n_826),
.D(n_827),
.Y(n_9857)
);

NAND2xp5_ASAP7_75t_L g9858 ( 
.A(n_9611),
.B(n_826),
.Y(n_9858)
);

NAND2xp5_ASAP7_75t_L g9859 ( 
.A(n_9450),
.B(n_827),
.Y(n_9859)
);

NAND2xp5_ASAP7_75t_L g9860 ( 
.A(n_9444),
.B(n_827),
.Y(n_9860)
);

OR2x2_ASAP7_75t_L g9861 ( 
.A(n_9500),
.B(n_828),
.Y(n_9861)
);

AOI21xp33_ASAP7_75t_L g9862 ( 
.A1(n_9621),
.A2(n_828),
.B(n_829),
.Y(n_9862)
);

INVx2_ASAP7_75t_L g9863 ( 
.A(n_9574),
.Y(n_9863)
);

NAND2xp5_ASAP7_75t_L g9864 ( 
.A(n_9410),
.B(n_829),
.Y(n_9864)
);

NAND2xp5_ASAP7_75t_L g9865 ( 
.A(n_9548),
.B(n_829),
.Y(n_9865)
);

INVx4_ASAP7_75t_L g9866 ( 
.A(n_9419),
.Y(n_9866)
);

BUFx2_ASAP7_75t_L g9867 ( 
.A(n_9640),
.Y(n_9867)
);

INVx1_ASAP7_75t_L g9868 ( 
.A(n_9549),
.Y(n_9868)
);

HB1xp67_ASAP7_75t_L g9869 ( 
.A(n_9366),
.Y(n_9869)
);

INVx1_ASAP7_75t_L g9870 ( 
.A(n_9525),
.Y(n_9870)
);

NAND2xp5_ASAP7_75t_L g9871 ( 
.A(n_9442),
.B(n_830),
.Y(n_9871)
);

OR2x2_ASAP7_75t_L g9872 ( 
.A(n_9497),
.B(n_830),
.Y(n_9872)
);

INVx2_ASAP7_75t_L g9873 ( 
.A(n_9519),
.Y(n_9873)
);

INVx1_ASAP7_75t_L g9874 ( 
.A(n_9592),
.Y(n_9874)
);

OAI22xp5_ASAP7_75t_L g9875 ( 
.A1(n_9365),
.A2(n_832),
.B1(n_830),
.B2(n_831),
.Y(n_9875)
);

INVx1_ASAP7_75t_L g9876 ( 
.A(n_9536),
.Y(n_9876)
);

NAND2xp5_ASAP7_75t_L g9877 ( 
.A(n_9463),
.B(n_831),
.Y(n_9877)
);

INVx1_ASAP7_75t_L g9878 ( 
.A(n_9518),
.Y(n_9878)
);

INVx1_ASAP7_75t_L g9879 ( 
.A(n_9560),
.Y(n_9879)
);

AND2x2_ASAP7_75t_SL g9880 ( 
.A(n_9649),
.B(n_831),
.Y(n_9880)
);

AND2x2_ASAP7_75t_L g9881 ( 
.A(n_9558),
.B(n_832),
.Y(n_9881)
);

BUFx2_ASAP7_75t_L g9882 ( 
.A(n_9514),
.Y(n_9882)
);

OR2x2_ASAP7_75t_L g9883 ( 
.A(n_9484),
.B(n_9590),
.Y(n_9883)
);

NOR2xp33_ASAP7_75t_L g9884 ( 
.A(n_9399),
.B(n_832),
.Y(n_9884)
);

INVx1_ASAP7_75t_L g9885 ( 
.A(n_9588),
.Y(n_9885)
);

INVx1_ASAP7_75t_L g9886 ( 
.A(n_9384),
.Y(n_9886)
);

NAND2x1p5_ASAP7_75t_SL g9887 ( 
.A(n_9335),
.B(n_833),
.Y(n_9887)
);

INVx2_ASAP7_75t_L g9888 ( 
.A(n_9566),
.Y(n_9888)
);

BUFx2_ASAP7_75t_L g9889 ( 
.A(n_9388),
.Y(n_9889)
);

INVxp67_ASAP7_75t_L g9890 ( 
.A(n_9628),
.Y(n_9890)
);

INVx1_ASAP7_75t_L g9891 ( 
.A(n_9559),
.Y(n_9891)
);

INVx2_ASAP7_75t_L g9892 ( 
.A(n_9490),
.Y(n_9892)
);

OR2x2_ASAP7_75t_L g9893 ( 
.A(n_9515),
.B(n_833),
.Y(n_9893)
);

NAND2xp5_ASAP7_75t_L g9894 ( 
.A(n_9602),
.B(n_834),
.Y(n_9894)
);

AND2x2_ASAP7_75t_L g9895 ( 
.A(n_9485),
.B(n_834),
.Y(n_9895)
);

NAND2xp5_ASAP7_75t_L g9896 ( 
.A(n_9447),
.B(n_835),
.Y(n_9896)
);

AND2x2_ASAP7_75t_L g9897 ( 
.A(n_9572),
.B(n_835),
.Y(n_9897)
);

NAND2xp5_ASAP7_75t_L g9898 ( 
.A(n_9704),
.B(n_9407),
.Y(n_9898)
);

NAND4xp25_ASAP7_75t_SL g9899 ( 
.A(n_9834),
.B(n_9670),
.C(n_9785),
.D(n_9638),
.Y(n_9899)
);

NAND2xp5_ASAP7_75t_SL g9900 ( 
.A(n_9661),
.B(n_9527),
.Y(n_9900)
);

INVx2_ASAP7_75t_L g9901 ( 
.A(n_9707),
.Y(n_9901)
);

OAI33xp33_ASAP7_75t_L g9902 ( 
.A1(n_9783),
.A2(n_9349),
.A3(n_9530),
.B1(n_9543),
.B2(n_9367),
.B3(n_9594),
.Y(n_9902)
);

HB1xp67_ASAP7_75t_L g9903 ( 
.A(n_9775),
.Y(n_9903)
);

AND2x2_ASAP7_75t_L g9904 ( 
.A(n_9781),
.B(n_9600),
.Y(n_9904)
);

AOI22xp33_ASAP7_75t_L g9905 ( 
.A1(n_9866),
.A2(n_9603),
.B1(n_9382),
.B2(n_9618),
.Y(n_9905)
);

INVx1_ASAP7_75t_L g9906 ( 
.A(n_9659),
.Y(n_9906)
);

AOI22xp5_ASAP7_75t_L g9907 ( 
.A1(n_9867),
.A2(n_9608),
.B1(n_9634),
.B2(n_9334),
.Y(n_9907)
);

OAI21xp5_ASAP7_75t_L g9908 ( 
.A1(n_9677),
.A2(n_9756),
.B(n_9743),
.Y(n_9908)
);

BUFx2_ASAP7_75t_L g9909 ( 
.A(n_9696),
.Y(n_9909)
);

AND2x2_ASAP7_75t_L g9910 ( 
.A(n_9740),
.B(n_9806),
.Y(n_9910)
);

OAI221xp5_ASAP7_75t_L g9911 ( 
.A1(n_9882),
.A2(n_9607),
.B1(n_9652),
.B2(n_9617),
.C(n_9631),
.Y(n_9911)
);

OR2x2_ASAP7_75t_L g9912 ( 
.A(n_9721),
.B(n_9565),
.Y(n_9912)
);

AND2x2_ASAP7_75t_L g9913 ( 
.A(n_9772),
.B(n_9357),
.Y(n_9913)
);

AND2x2_ASAP7_75t_L g9914 ( 
.A(n_9669),
.B(n_9575),
.Y(n_9914)
);

OAI22xp5_ASAP7_75t_L g9915 ( 
.A1(n_9889),
.A2(n_9526),
.B1(n_9480),
.B2(n_9403),
.Y(n_9915)
);

AOI33xp33_ASAP7_75t_L g9916 ( 
.A1(n_9685),
.A2(n_9381),
.A3(n_9411),
.B1(n_9397),
.B2(n_9539),
.B3(n_9553),
.Y(n_9916)
);

AND4x1_ASAP7_75t_L g9917 ( 
.A(n_9655),
.B(n_9363),
.C(n_9639),
.D(n_9622),
.Y(n_9917)
);

HB1xp67_ASAP7_75t_L g9918 ( 
.A(n_9668),
.Y(n_9918)
);

OAI22xp5_ASAP7_75t_L g9919 ( 
.A1(n_9879),
.A2(n_9499),
.B1(n_9511),
.B2(n_9351),
.Y(n_9919)
);

AND2x2_ASAP7_75t_L g9920 ( 
.A(n_9686),
.B(n_9589),
.Y(n_9920)
);

NOR2xp33_ASAP7_75t_L g9921 ( 
.A(n_9793),
.B(n_9751),
.Y(n_9921)
);

AND2x2_ASAP7_75t_L g9922 ( 
.A(n_9690),
.B(n_9415),
.Y(n_9922)
);

OR2x2_ASAP7_75t_L g9923 ( 
.A(n_9828),
.B(n_9522),
.Y(n_9923)
);

INVx2_ASAP7_75t_L g9924 ( 
.A(n_9763),
.Y(n_9924)
);

INVx1_ASAP7_75t_L g9925 ( 
.A(n_9695),
.Y(n_9925)
);

NAND4xp25_ASAP7_75t_L g9926 ( 
.A(n_9837),
.B(n_9647),
.C(n_9396),
.D(n_9421),
.Y(n_9926)
);

HB1xp67_ASAP7_75t_L g9927 ( 
.A(n_9671),
.Y(n_9927)
);

AOI22xp33_ASAP7_75t_L g9928 ( 
.A1(n_9854),
.A2(n_9414),
.B1(n_9540),
.B2(n_9426),
.Y(n_9928)
);

AOI221xp5_ASAP7_75t_L g9929 ( 
.A1(n_9758),
.A2(n_9887),
.B1(n_9726),
.B2(n_9757),
.C(n_9862),
.Y(n_9929)
);

OAI22xp5_ASAP7_75t_L g9930 ( 
.A1(n_9842),
.A2(n_9454),
.B1(n_9455),
.B2(n_9568),
.Y(n_9930)
);

OAI321xp33_ASAP7_75t_L g9931 ( 
.A1(n_9857),
.A2(n_9459),
.A3(n_9486),
.B1(n_9385),
.B2(n_9461),
.C(n_9544),
.Y(n_9931)
);

OR2x2_ASAP7_75t_L g9932 ( 
.A(n_9657),
.B(n_9576),
.Y(n_9932)
);

INVx1_ASAP7_75t_L g9933 ( 
.A(n_9724),
.Y(n_9933)
);

NAND4xp25_ASAP7_75t_L g9934 ( 
.A(n_9689),
.B(n_9483),
.C(n_9529),
.D(n_9431),
.Y(n_9934)
);

AND2x2_ASAP7_75t_L g9935 ( 
.A(n_9698),
.B(n_9436),
.Y(n_9935)
);

AO21x2_ASAP7_75t_L g9936 ( 
.A1(n_9731),
.A2(n_9355),
.B(n_9509),
.Y(n_9936)
);

HB1xp67_ASAP7_75t_L g9937 ( 
.A(n_9739),
.Y(n_9937)
);

AOI22xp33_ASAP7_75t_L g9938 ( 
.A1(n_9839),
.A2(n_9517),
.B1(n_9583),
.B2(n_9477),
.Y(n_9938)
);

BUFx2_ASAP7_75t_L g9939 ( 
.A(n_9694),
.Y(n_9939)
);

INVx1_ASAP7_75t_L g9940 ( 
.A(n_9778),
.Y(n_9940)
);

INVx1_ASAP7_75t_L g9941 ( 
.A(n_9800),
.Y(n_9941)
);

OAI33xp33_ASAP7_75t_L g9942 ( 
.A1(n_9811),
.A2(n_9875),
.A3(n_9656),
.B1(n_9663),
.B2(n_9850),
.B3(n_9856),
.Y(n_9942)
);

AND2x2_ASAP7_75t_L g9943 ( 
.A(n_9702),
.B(n_9535),
.Y(n_9943)
);

INVx2_ASAP7_75t_L g9944 ( 
.A(n_9754),
.Y(n_9944)
);

OAI22xp5_ASAP7_75t_L g9945 ( 
.A1(n_9869),
.A2(n_9506),
.B1(n_9498),
.B2(n_9545),
.Y(n_9945)
);

INVx2_ASAP7_75t_L g9946 ( 
.A(n_9815),
.Y(n_9946)
);

OAI22xp5_ASAP7_75t_L g9947 ( 
.A1(n_9855),
.A2(n_9546),
.B1(n_9569),
.B2(n_9491),
.Y(n_9947)
);

INVx2_ASAP7_75t_L g9948 ( 
.A(n_9730),
.Y(n_9948)
);

AND2x2_ASAP7_75t_L g9949 ( 
.A(n_9711),
.B(n_9374),
.Y(n_9949)
);

INVx2_ASAP7_75t_L g9950 ( 
.A(n_9803),
.Y(n_9950)
);

INVx1_ASAP7_75t_L g9951 ( 
.A(n_9691),
.Y(n_9951)
);

OAI22xp33_ASAP7_75t_L g9952 ( 
.A1(n_9822),
.A2(n_9376),
.B1(n_837),
.B2(n_838),
.Y(n_9952)
);

OR2x2_ASAP7_75t_L g9953 ( 
.A(n_9774),
.B(n_835),
.Y(n_9953)
);

NAND4xp25_ASAP7_75t_SL g9954 ( 
.A(n_9762),
.B(n_9894),
.C(n_9883),
.D(n_9885),
.Y(n_9954)
);

AND2x2_ASAP7_75t_L g9955 ( 
.A(n_9812),
.B(n_9725),
.Y(n_9955)
);

INVx1_ASAP7_75t_L g9956 ( 
.A(n_9692),
.Y(n_9956)
);

INVx1_ASAP7_75t_L g9957 ( 
.A(n_9742),
.Y(n_9957)
);

INVx1_ASAP7_75t_L g9958 ( 
.A(n_9662),
.Y(n_9958)
);

OR2x2_ASAP7_75t_L g9959 ( 
.A(n_9870),
.B(n_836),
.Y(n_9959)
);

OR2x2_ASAP7_75t_L g9960 ( 
.A(n_9805),
.B(n_836),
.Y(n_9960)
);

BUFx2_ASAP7_75t_L g9961 ( 
.A(n_9676),
.Y(n_9961)
);

INVx2_ASAP7_75t_L g9962 ( 
.A(n_9717),
.Y(n_9962)
);

OR2x2_ASAP7_75t_L g9963 ( 
.A(n_9688),
.B(n_837),
.Y(n_9963)
);

INVx3_ASAP7_75t_L g9964 ( 
.A(n_9712),
.Y(n_9964)
);

INVx1_ASAP7_75t_L g9965 ( 
.A(n_9746),
.Y(n_9965)
);

AND2x2_ASAP7_75t_L g9966 ( 
.A(n_9700),
.B(n_838),
.Y(n_9966)
);

INVx1_ASAP7_75t_L g9967 ( 
.A(n_9672),
.Y(n_9967)
);

AOI221x1_ASAP7_75t_L g9968 ( 
.A1(n_9826),
.A2(n_840),
.B1(n_838),
.B2(n_839),
.C(n_841),
.Y(n_9968)
);

AND2x2_ASAP7_75t_SL g9969 ( 
.A(n_9684),
.B(n_840),
.Y(n_9969)
);

INVx2_ASAP7_75t_L g9970 ( 
.A(n_9808),
.Y(n_9970)
);

OAI221xp5_ASAP7_75t_L g9971 ( 
.A1(n_9890),
.A2(n_841),
.B1(n_839),
.B2(n_840),
.C(n_842),
.Y(n_9971)
);

INVx1_ASAP7_75t_L g9972 ( 
.A(n_9658),
.Y(n_9972)
);

AOI22xp5_ASAP7_75t_L g9973 ( 
.A1(n_9801),
.A2(n_842),
.B1(n_839),
.B2(n_841),
.Y(n_9973)
);

OR2x2_ASAP7_75t_L g9974 ( 
.A(n_9825),
.B(n_843),
.Y(n_9974)
);

OR2x2_ASAP7_75t_L g9975 ( 
.A(n_9741),
.B(n_843),
.Y(n_9975)
);

AND2x2_ASAP7_75t_L g9976 ( 
.A(n_9720),
.B(n_844),
.Y(n_9976)
);

INVx2_ASAP7_75t_L g9977 ( 
.A(n_9727),
.Y(n_9977)
);

OR2x2_ASAP7_75t_L g9978 ( 
.A(n_9744),
.B(n_844),
.Y(n_9978)
);

INVx5_ASAP7_75t_L g9979 ( 
.A(n_9680),
.Y(n_9979)
);

NAND2xp5_ASAP7_75t_L g9980 ( 
.A(n_9846),
.B(n_9747),
.Y(n_9980)
);

BUFx3_ASAP7_75t_L g9981 ( 
.A(n_9723),
.Y(n_9981)
);

NAND2xp5_ASAP7_75t_L g9982 ( 
.A(n_9891),
.B(n_845),
.Y(n_9982)
);

INVx1_ASAP7_75t_SL g9983 ( 
.A(n_9735),
.Y(n_9983)
);

INVx1_ASAP7_75t_L g9984 ( 
.A(n_9802),
.Y(n_9984)
);

INVx1_ASAP7_75t_L g9985 ( 
.A(n_9699),
.Y(n_9985)
);

HB1xp67_ASAP7_75t_L g9986 ( 
.A(n_9771),
.Y(n_9986)
);

OR2x2_ASAP7_75t_L g9987 ( 
.A(n_9749),
.B(n_845),
.Y(n_9987)
);

OAI211xp5_ASAP7_75t_L g9988 ( 
.A1(n_9782),
.A2(n_9871),
.B(n_9841),
.C(n_9878),
.Y(n_9988)
);

INVx1_ASAP7_75t_L g9989 ( 
.A(n_9764),
.Y(n_9989)
);

BUFx2_ASAP7_75t_L g9990 ( 
.A(n_9738),
.Y(n_9990)
);

NOR3xp33_ASAP7_75t_L g9991 ( 
.A(n_9831),
.B(n_854),
.C(n_846),
.Y(n_9991)
);

AND2x2_ASAP7_75t_L g9992 ( 
.A(n_9848),
.B(n_846),
.Y(n_9992)
);

NAND2xp5_ASAP7_75t_L g9993 ( 
.A(n_9863),
.B(n_846),
.Y(n_9993)
);

NAND2xp5_ASAP7_75t_L g9994 ( 
.A(n_9873),
.B(n_847),
.Y(n_9994)
);

INVx2_ASAP7_75t_L g9995 ( 
.A(n_9697),
.Y(n_9995)
);

OR2x2_ASAP7_75t_L g9996 ( 
.A(n_9868),
.B(n_847),
.Y(n_9996)
);

OR2x2_ASAP7_75t_L g9997 ( 
.A(n_9874),
.B(n_847),
.Y(n_9997)
);

INVx1_ASAP7_75t_L g9998 ( 
.A(n_9660),
.Y(n_9998)
);

OAI211xp5_ASAP7_75t_L g9999 ( 
.A1(n_9896),
.A2(n_850),
.B(n_848),
.C(n_849),
.Y(n_9999)
);

NOR2xp33_ASAP7_75t_L g10000 ( 
.A(n_9853),
.B(n_848),
.Y(n_10000)
);

NAND2xp5_ASAP7_75t_L g10001 ( 
.A(n_9892),
.B(n_848),
.Y(n_10001)
);

AND2x2_ASAP7_75t_L g10002 ( 
.A(n_9715),
.B(n_849),
.Y(n_10002)
);

OR2x2_ASAP7_75t_L g10003 ( 
.A(n_9769),
.B(n_849),
.Y(n_10003)
);

OAI22xp5_ASAP7_75t_L g10004 ( 
.A1(n_9876),
.A2(n_852),
.B1(n_850),
.B2(n_851),
.Y(n_10004)
);

INVx1_ASAP7_75t_L g10005 ( 
.A(n_9687),
.Y(n_10005)
);

INVx1_ASAP7_75t_L g10006 ( 
.A(n_9703),
.Y(n_10006)
);

INVx1_ASAP7_75t_L g10007 ( 
.A(n_9667),
.Y(n_10007)
);

NAND2xp5_ASAP7_75t_L g10008 ( 
.A(n_9833),
.B(n_851),
.Y(n_10008)
);

AOI22xp33_ASAP7_75t_L g10009 ( 
.A1(n_9886),
.A2(n_854),
.B1(n_852),
.B2(n_853),
.Y(n_10009)
);

INVx4_ASAP7_75t_L g10010 ( 
.A(n_9755),
.Y(n_10010)
);

INVx1_ASAP7_75t_L g10011 ( 
.A(n_9681),
.Y(n_10011)
);

HB1xp67_ASAP7_75t_L g10012 ( 
.A(n_9814),
.Y(n_10012)
);

INVx1_ASAP7_75t_L g10013 ( 
.A(n_9708),
.Y(n_10013)
);

INVx1_ASAP7_75t_L g10014 ( 
.A(n_9713),
.Y(n_10014)
);

AND2x2_ASAP7_75t_L g10015 ( 
.A(n_9840),
.B(n_852),
.Y(n_10015)
);

AND2x2_ASAP7_75t_L g10016 ( 
.A(n_9844),
.B(n_853),
.Y(n_10016)
);

AO21x2_ASAP7_75t_L g10017 ( 
.A1(n_9752),
.A2(n_854),
.B(n_855),
.Y(n_10017)
);

NAND2xp5_ASAP7_75t_L g10018 ( 
.A(n_9838),
.B(n_855),
.Y(n_10018)
);

INVx2_ASAP7_75t_L g10019 ( 
.A(n_9710),
.Y(n_10019)
);

NAND3xp33_ASAP7_75t_L g10020 ( 
.A(n_9832),
.B(n_855),
.C(n_856),
.Y(n_10020)
);

INVx1_ASAP7_75t_L g10021 ( 
.A(n_9714),
.Y(n_10021)
);

AND2x2_ASAP7_75t_L g10022 ( 
.A(n_9817),
.B(n_856),
.Y(n_10022)
);

AO21x2_ASAP7_75t_L g10023 ( 
.A1(n_9830),
.A2(n_856),
.B(n_857),
.Y(n_10023)
);

AOI22xp33_ASAP7_75t_L g10024 ( 
.A1(n_9888),
.A2(n_859),
.B1(n_857),
.B2(n_858),
.Y(n_10024)
);

NAND2xp5_ASAP7_75t_L g10025 ( 
.A(n_9824),
.B(n_857),
.Y(n_10025)
);

AOI21xp5_ASAP7_75t_L g10026 ( 
.A1(n_9859),
.A2(n_858),
.B(n_859),
.Y(n_10026)
);

AO21x2_ASAP7_75t_L g10027 ( 
.A1(n_9737),
.A2(n_858),
.B(n_860),
.Y(n_10027)
);

AND2x2_ASAP7_75t_L g10028 ( 
.A(n_9821),
.B(n_860),
.Y(n_10028)
);

INVx1_ASAP7_75t_L g10029 ( 
.A(n_9718),
.Y(n_10029)
);

NAND2xp5_ASAP7_75t_L g10030 ( 
.A(n_9884),
.B(n_9835),
.Y(n_10030)
);

OR2x2_ASAP7_75t_L g10031 ( 
.A(n_9664),
.B(n_861),
.Y(n_10031)
);

INVx1_ASAP7_75t_L g10032 ( 
.A(n_9674),
.Y(n_10032)
);

AND2x2_ASAP7_75t_L g10033 ( 
.A(n_9836),
.B(n_861),
.Y(n_10033)
);

OAI33xp33_ASAP7_75t_L g10034 ( 
.A1(n_9665),
.A2(n_864),
.A3(n_866),
.B1(n_862),
.B2(n_863),
.B3(n_865),
.Y(n_10034)
);

AND2x2_ASAP7_75t_L g10035 ( 
.A(n_9765),
.B(n_862),
.Y(n_10035)
);

BUFx3_ASAP7_75t_L g10036 ( 
.A(n_9760),
.Y(n_10036)
);

AOI21xp33_ASAP7_75t_L g10037 ( 
.A1(n_9796),
.A2(n_9804),
.B(n_9798),
.Y(n_10037)
);

OAI31xp33_ASAP7_75t_L g10038 ( 
.A1(n_9865),
.A2(n_864),
.A3(n_862),
.B(n_863),
.Y(n_10038)
);

INVx2_ASAP7_75t_L g10039 ( 
.A(n_9797),
.Y(n_10039)
);

INVx2_ASAP7_75t_L g10040 ( 
.A(n_9790),
.Y(n_10040)
);

OAI22xp5_ASAP7_75t_L g10041 ( 
.A1(n_9893),
.A2(n_867),
.B1(n_865),
.B2(n_866),
.Y(n_10041)
);

OAI221xp5_ASAP7_75t_L g10042 ( 
.A1(n_9816),
.A2(n_867),
.B1(n_865),
.B2(n_866),
.C(n_868),
.Y(n_10042)
);

AND2x4_ASAP7_75t_L g10043 ( 
.A(n_9736),
.B(n_867),
.Y(n_10043)
);

AND2x2_ASAP7_75t_L g10044 ( 
.A(n_9813),
.B(n_868),
.Y(n_10044)
);

AND2x2_ASAP7_75t_L g10045 ( 
.A(n_9766),
.B(n_868),
.Y(n_10045)
);

INVx3_ASAP7_75t_L g10046 ( 
.A(n_9807),
.Y(n_10046)
);

AND2x2_ASAP7_75t_L g10047 ( 
.A(n_9776),
.B(n_869),
.Y(n_10047)
);

AOI22xp5_ASAP7_75t_L g10048 ( 
.A1(n_9880),
.A2(n_871),
.B1(n_869),
.B2(n_870),
.Y(n_10048)
);

AO221x2_ASAP7_75t_L g10049 ( 
.A1(n_9860),
.A2(n_886),
.B1(n_894),
.B2(n_878),
.C(n_869),
.Y(n_10049)
);

INVx2_ASAP7_75t_SL g10050 ( 
.A(n_9818),
.Y(n_10050)
);

INVx2_ASAP7_75t_L g10051 ( 
.A(n_9792),
.Y(n_10051)
);

AOI33xp33_ASAP7_75t_L g10052 ( 
.A1(n_9895),
.A2(n_872),
.A3(n_875),
.B1(n_870),
.B2(n_871),
.B3(n_873),
.Y(n_10052)
);

AOI22xp5_ASAP7_75t_L g10053 ( 
.A1(n_9852),
.A2(n_872),
.B1(n_870),
.B2(n_871),
.Y(n_10053)
);

AO21x2_ASAP7_75t_L g10054 ( 
.A1(n_9858),
.A2(n_872),
.B(n_873),
.Y(n_10054)
);

AND2x2_ASAP7_75t_L g10055 ( 
.A(n_9823),
.B(n_875),
.Y(n_10055)
);

OAI21x1_ASAP7_75t_L g10056 ( 
.A1(n_9794),
.A2(n_876),
.B(n_877),
.Y(n_10056)
);

OR2x2_ASAP7_75t_L g10057 ( 
.A(n_9799),
.B(n_876),
.Y(n_10057)
);

NOR3xp33_ASAP7_75t_L g10058 ( 
.A(n_9787),
.B(n_884),
.C(n_876),
.Y(n_10058)
);

INVx3_ASAP7_75t_L g10059 ( 
.A(n_9780),
.Y(n_10059)
);

AND2x4_ASAP7_75t_SL g10060 ( 
.A(n_9759),
.B(n_877),
.Y(n_10060)
);

INVx1_ASAP7_75t_L g10061 ( 
.A(n_9666),
.Y(n_10061)
);

INVx3_ASAP7_75t_L g10062 ( 
.A(n_9789),
.Y(n_10062)
);

INVx1_ASAP7_75t_L g10063 ( 
.A(n_9673),
.Y(n_10063)
);

AND2x2_ASAP7_75t_L g10064 ( 
.A(n_9761),
.B(n_877),
.Y(n_10064)
);

INVx1_ASAP7_75t_L g10065 ( 
.A(n_9675),
.Y(n_10065)
);

INVx1_ASAP7_75t_L g10066 ( 
.A(n_9678),
.Y(n_10066)
);

INVx2_ASAP7_75t_L g10067 ( 
.A(n_9779),
.Y(n_10067)
);

NOR2x1_ASAP7_75t_L g10068 ( 
.A(n_9845),
.B(n_878),
.Y(n_10068)
);

AND2x2_ASAP7_75t_L g10069 ( 
.A(n_9773),
.B(n_879),
.Y(n_10069)
);

INVx1_ASAP7_75t_L g10070 ( 
.A(n_9679),
.Y(n_10070)
);

OR2x2_ASAP7_75t_L g10071 ( 
.A(n_9791),
.B(n_879),
.Y(n_10071)
);

NAND2xp5_ASAP7_75t_L g10072 ( 
.A(n_9820),
.B(n_879),
.Y(n_10072)
);

INVx1_ASAP7_75t_L g10073 ( 
.A(n_9682),
.Y(n_10073)
);

NAND2xp5_ASAP7_75t_L g10074 ( 
.A(n_9795),
.B(n_880),
.Y(n_10074)
);

NAND2xp5_ASAP7_75t_L g10075 ( 
.A(n_9827),
.B(n_880),
.Y(n_10075)
);

NOR2xp33_ASAP7_75t_L g10076 ( 
.A(n_9872),
.B(n_880),
.Y(n_10076)
);

OR2x2_ASAP7_75t_L g10077 ( 
.A(n_9861),
.B(n_881),
.Y(n_10077)
);

INVx2_ASAP7_75t_L g10078 ( 
.A(n_9683),
.Y(n_10078)
);

INVx1_ASAP7_75t_L g10079 ( 
.A(n_9693),
.Y(n_10079)
);

OAI31xp33_ASAP7_75t_L g10080 ( 
.A1(n_9864),
.A2(n_883),
.A3(n_881),
.B(n_882),
.Y(n_10080)
);

AOI33xp33_ASAP7_75t_L g10081 ( 
.A1(n_9701),
.A2(n_883),
.A3(n_885),
.B1(n_881),
.B2(n_882),
.B3(n_884),
.Y(n_10081)
);

INVx1_ASAP7_75t_L g10082 ( 
.A(n_9705),
.Y(n_10082)
);

INVx1_ASAP7_75t_L g10083 ( 
.A(n_9706),
.Y(n_10083)
);

INVx3_ASAP7_75t_L g10084 ( 
.A(n_9809),
.Y(n_10084)
);

INVx3_ASAP7_75t_L g10085 ( 
.A(n_9810),
.Y(n_10085)
);

NAND2xp5_ASAP7_75t_L g10086 ( 
.A(n_9881),
.B(n_882),
.Y(n_10086)
);

OR2x2_ASAP7_75t_L g10087 ( 
.A(n_9898),
.B(n_9719),
.Y(n_10087)
);

INVx2_ASAP7_75t_L g10088 ( 
.A(n_9981),
.Y(n_10088)
);

INVx1_ASAP7_75t_L g10089 ( 
.A(n_9918),
.Y(n_10089)
);

INVx2_ASAP7_75t_L g10090 ( 
.A(n_9961),
.Y(n_10090)
);

INVx2_ASAP7_75t_L g10091 ( 
.A(n_9979),
.Y(n_10091)
);

INVx2_ASAP7_75t_L g10092 ( 
.A(n_9979),
.Y(n_10092)
);

AND2x4_ASAP7_75t_L g10093 ( 
.A(n_9979),
.B(n_9819),
.Y(n_10093)
);

OR2x2_ASAP7_75t_L g10094 ( 
.A(n_9903),
.B(n_9722),
.Y(n_10094)
);

INVx1_ASAP7_75t_L g10095 ( 
.A(n_9909),
.Y(n_10095)
);

NAND2xp5_ASAP7_75t_L g10096 ( 
.A(n_9969),
.B(n_9777),
.Y(n_10096)
);

AND2x2_ASAP7_75t_L g10097 ( 
.A(n_9910),
.B(n_9767),
.Y(n_10097)
);

INVx1_ASAP7_75t_L g10098 ( 
.A(n_9937),
.Y(n_10098)
);

OR2x2_ASAP7_75t_L g10099 ( 
.A(n_9923),
.B(n_9847),
.Y(n_10099)
);

NAND2x1p5_ASAP7_75t_L g10100 ( 
.A(n_10010),
.B(n_9829),
.Y(n_10100)
);

NAND2xp5_ASAP7_75t_L g10101 ( 
.A(n_9939),
.B(n_9843),
.Y(n_10101)
);

AND2x2_ASAP7_75t_L g10102 ( 
.A(n_9955),
.B(n_9897),
.Y(n_10102)
);

INVx1_ASAP7_75t_L g10103 ( 
.A(n_10012),
.Y(n_10103)
);

OR2x2_ASAP7_75t_L g10104 ( 
.A(n_9983),
.B(n_9851),
.Y(n_10104)
);

INVx1_ASAP7_75t_L g10105 ( 
.A(n_10002),
.Y(n_10105)
);

AND2x2_ASAP7_75t_L g10106 ( 
.A(n_9964),
.B(n_9921),
.Y(n_10106)
);

INVx1_ASAP7_75t_L g10107 ( 
.A(n_9966),
.Y(n_10107)
);

NAND2xp5_ASAP7_75t_L g10108 ( 
.A(n_9936),
.B(n_9849),
.Y(n_10108)
);

NAND2xp5_ASAP7_75t_L g10109 ( 
.A(n_9929),
.B(n_10046),
.Y(n_10109)
);

AND2x4_ASAP7_75t_L g10110 ( 
.A(n_10036),
.B(n_9709),
.Y(n_10110)
);

NAND2xp5_ASAP7_75t_L g10111 ( 
.A(n_9907),
.B(n_9716),
.Y(n_10111)
);

INVxp67_ASAP7_75t_SL g10112 ( 
.A(n_9927),
.Y(n_10112)
);

INVx1_ASAP7_75t_L g10113 ( 
.A(n_9906),
.Y(n_10113)
);

AND2x2_ASAP7_75t_L g10114 ( 
.A(n_9948),
.B(n_9914),
.Y(n_10114)
);

NAND2xp5_ASAP7_75t_L g10115 ( 
.A(n_9986),
.B(n_9904),
.Y(n_10115)
);

NAND2xp5_ASAP7_75t_L g10116 ( 
.A(n_9920),
.B(n_9728),
.Y(n_10116)
);

OR2x2_ASAP7_75t_L g10117 ( 
.A(n_9980),
.B(n_9729),
.Y(n_10117)
);

INVx1_ASAP7_75t_L g10118 ( 
.A(n_9933),
.Y(n_10118)
);

NOR2xp67_ASAP7_75t_L g10119 ( 
.A(n_10059),
.B(n_9732),
.Y(n_10119)
);

INVx2_ASAP7_75t_L g10120 ( 
.A(n_9990),
.Y(n_10120)
);

OR2x2_ASAP7_75t_L g10121 ( 
.A(n_9995),
.B(n_9733),
.Y(n_10121)
);

INVx1_ASAP7_75t_L g10122 ( 
.A(n_9940),
.Y(n_10122)
);

NAND2x1_ASAP7_75t_L g10123 ( 
.A(n_10084),
.B(n_9734),
.Y(n_10123)
);

AND2x2_ASAP7_75t_L g10124 ( 
.A(n_9944),
.B(n_9745),
.Y(n_10124)
);

INVx1_ASAP7_75t_L g10125 ( 
.A(n_9941),
.Y(n_10125)
);

OR2x2_ASAP7_75t_L g10126 ( 
.A(n_10050),
.B(n_9748),
.Y(n_10126)
);

NAND2xp5_ASAP7_75t_L g10127 ( 
.A(n_10085),
.B(n_9750),
.Y(n_10127)
);

AOI22xp5_ASAP7_75t_L g10128 ( 
.A1(n_9899),
.A2(n_9786),
.B1(n_9877),
.B2(n_9768),
.Y(n_10128)
);

INVx1_ASAP7_75t_L g10129 ( 
.A(n_9976),
.Y(n_10129)
);

INVx1_ASAP7_75t_L g10130 ( 
.A(n_9925),
.Y(n_10130)
);

INVx2_ASAP7_75t_L g10131 ( 
.A(n_10062),
.Y(n_10131)
);

OR2x2_ASAP7_75t_L g10132 ( 
.A(n_9972),
.B(n_9753),
.Y(n_10132)
);

INVx1_ASAP7_75t_L g10133 ( 
.A(n_10057),
.Y(n_10133)
);

NOR2x1_ASAP7_75t_L g10134 ( 
.A(n_9908),
.B(n_9770),
.Y(n_10134)
);

AND2x2_ASAP7_75t_L g10135 ( 
.A(n_9901),
.B(n_9784),
.Y(n_10135)
);

OR2x2_ASAP7_75t_L g10136 ( 
.A(n_10039),
.B(n_9788),
.Y(n_10136)
);

AND2x4_ASAP7_75t_L g10137 ( 
.A(n_9950),
.B(n_883),
.Y(n_10137)
);

AND2x2_ASAP7_75t_L g10138 ( 
.A(n_9924),
.B(n_885),
.Y(n_10138)
);

INVx2_ASAP7_75t_L g10139 ( 
.A(n_9946),
.Y(n_10139)
);

OAI22xp5_ASAP7_75t_L g10140 ( 
.A1(n_9905),
.A2(n_888),
.B1(n_886),
.B2(n_887),
.Y(n_10140)
);

AND2x2_ASAP7_75t_L g10141 ( 
.A(n_9922),
.B(n_887),
.Y(n_10141)
);

INVx2_ASAP7_75t_L g10142 ( 
.A(n_10043),
.Y(n_10142)
);

INVx1_ASAP7_75t_L g10143 ( 
.A(n_9953),
.Y(n_10143)
);

HB1xp67_ASAP7_75t_L g10144 ( 
.A(n_10027),
.Y(n_10144)
);

AND2x2_ASAP7_75t_L g10145 ( 
.A(n_9949),
.B(n_887),
.Y(n_10145)
);

AND2x2_ASAP7_75t_L g10146 ( 
.A(n_9943),
.B(n_888),
.Y(n_10146)
);

OR2x2_ASAP7_75t_L g10147 ( 
.A(n_9932),
.B(n_888),
.Y(n_10147)
);

OR2x2_ASAP7_75t_L g10148 ( 
.A(n_10030),
.B(n_9997),
.Y(n_10148)
);

OR2x2_ASAP7_75t_L g10149 ( 
.A(n_9996),
.B(n_889),
.Y(n_10149)
);

INVx1_ASAP7_75t_L g10150 ( 
.A(n_9975),
.Y(n_10150)
);

OAI21xp33_ASAP7_75t_SL g10151 ( 
.A1(n_9928),
.A2(n_889),
.B(n_890),
.Y(n_10151)
);

NAND2xp5_ASAP7_75t_L g10152 ( 
.A(n_9913),
.B(n_889),
.Y(n_10152)
);

AND2x2_ASAP7_75t_L g10153 ( 
.A(n_9935),
.B(n_890),
.Y(n_10153)
);

AND2x2_ASAP7_75t_L g10154 ( 
.A(n_10067),
.B(n_891),
.Y(n_10154)
);

AND2x2_ASAP7_75t_L g10155 ( 
.A(n_10019),
.B(n_891),
.Y(n_10155)
);

INVx1_ASAP7_75t_L g10156 ( 
.A(n_9978),
.Y(n_10156)
);

AND2x4_ASAP7_75t_L g10157 ( 
.A(n_9970),
.B(n_9977),
.Y(n_10157)
);

INVx1_ASAP7_75t_L g10158 ( 
.A(n_9987),
.Y(n_10158)
);

INVx1_ASAP7_75t_L g10159 ( 
.A(n_9992),
.Y(n_10159)
);

INVx1_ASAP7_75t_L g10160 ( 
.A(n_9951),
.Y(n_10160)
);

NAND3xp33_ASAP7_75t_SL g10161 ( 
.A(n_9917),
.B(n_891),
.C(n_892),
.Y(n_10161)
);

OAI21xp5_ASAP7_75t_L g10162 ( 
.A1(n_9915),
.A2(n_892),
.B(n_893),
.Y(n_10162)
);

AND2x2_ASAP7_75t_L g10163 ( 
.A(n_9956),
.B(n_9967),
.Y(n_10163)
);

AOI221xp5_ASAP7_75t_L g10164 ( 
.A1(n_9942),
.A2(n_895),
.B1(n_897),
.B2(n_894),
.C(n_896),
.Y(n_10164)
);

NAND2xp5_ASAP7_75t_L g10165 ( 
.A(n_9973),
.B(n_892),
.Y(n_10165)
);

INVx2_ASAP7_75t_L g10166 ( 
.A(n_10060),
.Y(n_10166)
);

HB1xp67_ASAP7_75t_L g10167 ( 
.A(n_9958),
.Y(n_10167)
);

AND2x2_ASAP7_75t_L g10168 ( 
.A(n_10032),
.B(n_894),
.Y(n_10168)
);

INVx1_ASAP7_75t_L g10169 ( 
.A(n_10015),
.Y(n_10169)
);

NAND2x1p5_ASAP7_75t_L g10170 ( 
.A(n_10068),
.B(n_895),
.Y(n_10170)
);

NAND2xp5_ASAP7_75t_L g10171 ( 
.A(n_10023),
.B(n_895),
.Y(n_10171)
);

INVx1_ASAP7_75t_L g10172 ( 
.A(n_10011),
.Y(n_10172)
);

OR2x2_ASAP7_75t_SL g10173 ( 
.A(n_10020),
.B(n_896),
.Y(n_10173)
);

AND2x2_ASAP7_75t_L g10174 ( 
.A(n_10006),
.B(n_896),
.Y(n_10174)
);

NAND2xp5_ASAP7_75t_L g10175 ( 
.A(n_9968),
.B(n_897),
.Y(n_10175)
);

OR2x2_ASAP7_75t_L g10176 ( 
.A(n_9959),
.B(n_897),
.Y(n_10176)
);

NAND2xp5_ASAP7_75t_L g10177 ( 
.A(n_9938),
.B(n_898),
.Y(n_10177)
);

AND2x2_ASAP7_75t_L g10178 ( 
.A(n_10005),
.B(n_898),
.Y(n_10178)
);

AND2x2_ASAP7_75t_L g10179 ( 
.A(n_10007),
.B(n_898),
.Y(n_10179)
);

INVx1_ASAP7_75t_L g10180 ( 
.A(n_9965),
.Y(n_10180)
);

INVx2_ASAP7_75t_L g10181 ( 
.A(n_9962),
.Y(n_10181)
);

AND2x2_ASAP7_75t_L g10182 ( 
.A(n_9984),
.B(n_899),
.Y(n_10182)
);

INVx1_ASAP7_75t_L g10183 ( 
.A(n_9985),
.Y(n_10183)
);

OR2x2_ASAP7_75t_L g10184 ( 
.A(n_9912),
.B(n_900),
.Y(n_10184)
);

INVx1_ASAP7_75t_L g10185 ( 
.A(n_9960),
.Y(n_10185)
);

OR2x2_ASAP7_75t_L g10186 ( 
.A(n_10003),
.B(n_900),
.Y(n_10186)
);

INVx1_ASAP7_75t_L g10187 ( 
.A(n_10071),
.Y(n_10187)
);

INVx1_ASAP7_75t_L g10188 ( 
.A(n_10013),
.Y(n_10188)
);

AND2x2_ASAP7_75t_L g10189 ( 
.A(n_10014),
.B(n_10021),
.Y(n_10189)
);

NAND2xp5_ASAP7_75t_L g10190 ( 
.A(n_10026),
.B(n_900),
.Y(n_10190)
);

HB1xp67_ASAP7_75t_L g10191 ( 
.A(n_10017),
.Y(n_10191)
);

OR2x2_ASAP7_75t_L g10192 ( 
.A(n_9900),
.B(n_901),
.Y(n_10192)
);

AND2x4_ASAP7_75t_L g10193 ( 
.A(n_9989),
.B(n_901),
.Y(n_10193)
);

AND2x2_ASAP7_75t_L g10194 ( 
.A(n_10029),
.B(n_901),
.Y(n_10194)
);

INVx2_ASAP7_75t_L g10195 ( 
.A(n_10045),
.Y(n_10195)
);

INVx1_ASAP7_75t_L g10196 ( 
.A(n_9974),
.Y(n_10196)
);

AND2x2_ASAP7_75t_L g10197 ( 
.A(n_9957),
.B(n_902),
.Y(n_10197)
);

OR2x2_ASAP7_75t_L g10198 ( 
.A(n_9954),
.B(n_10054),
.Y(n_10198)
);

AND2x2_ASAP7_75t_L g10199 ( 
.A(n_10033),
.B(n_10055),
.Y(n_10199)
);

INVx2_ASAP7_75t_L g10200 ( 
.A(n_10047),
.Y(n_10200)
);

INVx2_ASAP7_75t_L g10201 ( 
.A(n_10035),
.Y(n_10201)
);

INVx1_ASAP7_75t_L g10202 ( 
.A(n_10031),
.Y(n_10202)
);

AND2x4_ASAP7_75t_L g10203 ( 
.A(n_9998),
.B(n_10064),
.Y(n_10203)
);

AND2x2_ASAP7_75t_L g10204 ( 
.A(n_10044),
.B(n_902),
.Y(n_10204)
);

AND2x4_ASAP7_75t_L g10205 ( 
.A(n_10069),
.B(n_10040),
.Y(n_10205)
);

INVx1_ASAP7_75t_L g10206 ( 
.A(n_10028),
.Y(n_10206)
);

OR2x2_ASAP7_75t_L g10207 ( 
.A(n_9963),
.B(n_902),
.Y(n_10207)
);

INVx1_ASAP7_75t_L g10208 ( 
.A(n_10016),
.Y(n_10208)
);

INVx1_ASAP7_75t_L g10209 ( 
.A(n_10022),
.Y(n_10209)
);

AND2x2_ASAP7_75t_L g10210 ( 
.A(n_10076),
.B(n_903),
.Y(n_10210)
);

INVx2_ASAP7_75t_L g10211 ( 
.A(n_10056),
.Y(n_10211)
);

OR2x2_ASAP7_75t_L g10212 ( 
.A(n_9988),
.B(n_904),
.Y(n_10212)
);

INVx1_ASAP7_75t_L g10213 ( 
.A(n_10074),
.Y(n_10213)
);

NOR3xp33_ASAP7_75t_L g10214 ( 
.A(n_9926),
.B(n_904),
.C(n_905),
.Y(n_10214)
);

AND2x2_ASAP7_75t_L g10215 ( 
.A(n_9982),
.B(n_905),
.Y(n_10215)
);

NAND2xp5_ASAP7_75t_L g10216 ( 
.A(n_10058),
.B(n_905),
.Y(n_10216)
);

AOI22xp5_ASAP7_75t_L g10217 ( 
.A1(n_9902),
.A2(n_9945),
.B1(n_9947),
.B2(n_9919),
.Y(n_10217)
);

OR2x2_ASAP7_75t_L g10218 ( 
.A(n_10077),
.B(n_906),
.Y(n_10218)
);

AND2x2_ASAP7_75t_L g10219 ( 
.A(n_10051),
.B(n_906),
.Y(n_10219)
);

OR2x2_ASAP7_75t_L g10220 ( 
.A(n_9934),
.B(n_907),
.Y(n_10220)
);

AND2x2_ASAP7_75t_L g10221 ( 
.A(n_10000),
.B(n_908),
.Y(n_10221)
);

INVx1_ASAP7_75t_L g10222 ( 
.A(n_10086),
.Y(n_10222)
);

OR2x2_ASAP7_75t_L g10223 ( 
.A(n_10001),
.B(n_908),
.Y(n_10223)
);

AND2x2_ASAP7_75t_L g10224 ( 
.A(n_10048),
.B(n_908),
.Y(n_10224)
);

AND2x2_ASAP7_75t_L g10225 ( 
.A(n_9994),
.B(n_909),
.Y(n_10225)
);

INVx1_ASAP7_75t_L g10226 ( 
.A(n_10075),
.Y(n_10226)
);

NAND2xp5_ASAP7_75t_L g10227 ( 
.A(n_10080),
.B(n_909),
.Y(n_10227)
);

OR2x2_ASAP7_75t_L g10228 ( 
.A(n_10025),
.B(n_909),
.Y(n_10228)
);

INVx1_ASAP7_75t_L g10229 ( 
.A(n_10008),
.Y(n_10229)
);

OR2x2_ASAP7_75t_L g10230 ( 
.A(n_10018),
.B(n_910),
.Y(n_10230)
);

OR2x2_ASAP7_75t_L g10231 ( 
.A(n_9993),
.B(n_910),
.Y(n_10231)
);

INVx1_ASAP7_75t_L g10232 ( 
.A(n_10072),
.Y(n_10232)
);

NAND2xp5_ASAP7_75t_L g10233 ( 
.A(n_10038),
.B(n_911),
.Y(n_10233)
);

INVxp67_ASAP7_75t_L g10234 ( 
.A(n_9971),
.Y(n_10234)
);

AND2x2_ASAP7_75t_L g10235 ( 
.A(n_10106),
.B(n_10078),
.Y(n_10235)
);

AND2x2_ASAP7_75t_L g10236 ( 
.A(n_10097),
.B(n_10049),
.Y(n_10236)
);

AND2x2_ASAP7_75t_L g10237 ( 
.A(n_10114),
.B(n_10049),
.Y(n_10237)
);

NAND2xp5_ASAP7_75t_L g10238 ( 
.A(n_10093),
.B(n_9952),
.Y(n_10238)
);

AND2x2_ASAP7_75t_L g10239 ( 
.A(n_10166),
.B(n_10061),
.Y(n_10239)
);

NOR3xp33_ASAP7_75t_L g10240 ( 
.A(n_10108),
.B(n_9999),
.C(n_10042),
.Y(n_10240)
);

OR2x2_ASAP7_75t_L g10241 ( 
.A(n_10096),
.B(n_9930),
.Y(n_10241)
);

OAI21xp5_ASAP7_75t_L g10242 ( 
.A1(n_10134),
.A2(n_9931),
.B(n_9911),
.Y(n_10242)
);

OR2x2_ASAP7_75t_L g10243 ( 
.A(n_10120),
.B(n_10090),
.Y(n_10243)
);

INVxp67_ASAP7_75t_L g10244 ( 
.A(n_10144),
.Y(n_10244)
);

INVx1_ASAP7_75t_L g10245 ( 
.A(n_10170),
.Y(n_10245)
);

INVxp67_ASAP7_75t_SL g10246 ( 
.A(n_10100),
.Y(n_10246)
);

INVx2_ASAP7_75t_L g10247 ( 
.A(n_10091),
.Y(n_10247)
);

INVx1_ASAP7_75t_L g10248 ( 
.A(n_10199),
.Y(n_10248)
);

HB1xp67_ASAP7_75t_L g10249 ( 
.A(n_10092),
.Y(n_10249)
);

AOI22xp33_ASAP7_75t_L g10250 ( 
.A1(n_10164),
.A2(n_9991),
.B1(n_10037),
.B2(n_10063),
.Y(n_10250)
);

OR2x2_ASAP7_75t_L g10251 ( 
.A(n_10101),
.B(n_10065),
.Y(n_10251)
);

AND2x2_ASAP7_75t_L g10252 ( 
.A(n_10102),
.B(n_10066),
.Y(n_10252)
);

INVx2_ASAP7_75t_L g10253 ( 
.A(n_10123),
.Y(n_10253)
);

AND2x2_ASAP7_75t_L g10254 ( 
.A(n_10088),
.B(n_10070),
.Y(n_10254)
);

AND2x2_ASAP7_75t_L g10255 ( 
.A(n_10146),
.B(n_10073),
.Y(n_10255)
);

INVx1_ASAP7_75t_L g10256 ( 
.A(n_10167),
.Y(n_10256)
);

AND2x2_ASAP7_75t_L g10257 ( 
.A(n_10142),
.B(n_10079),
.Y(n_10257)
);

AND2x2_ASAP7_75t_L g10258 ( 
.A(n_10145),
.B(n_10082),
.Y(n_10258)
);

INVx1_ASAP7_75t_L g10259 ( 
.A(n_10112),
.Y(n_10259)
);

BUFx2_ASAP7_75t_L g10260 ( 
.A(n_10095),
.Y(n_10260)
);

NOR2xp33_ASAP7_75t_L g10261 ( 
.A(n_10151),
.B(n_10053),
.Y(n_10261)
);

NAND3xp33_ASAP7_75t_L g10262 ( 
.A(n_10217),
.B(n_10009),
.C(n_10024),
.Y(n_10262)
);

AND2x2_ASAP7_75t_L g10263 ( 
.A(n_10153),
.B(n_10083),
.Y(n_10263)
);

INVx1_ASAP7_75t_L g10264 ( 
.A(n_10204),
.Y(n_10264)
);

BUFx2_ASAP7_75t_L g10265 ( 
.A(n_10191),
.Y(n_10265)
);

INVx2_ASAP7_75t_SL g10266 ( 
.A(n_10110),
.Y(n_10266)
);

INVx1_ASAP7_75t_L g10267 ( 
.A(n_10089),
.Y(n_10267)
);

AND2x2_ASAP7_75t_L g10268 ( 
.A(n_10141),
.B(n_10041),
.Y(n_10268)
);

INVx1_ASAP7_75t_SL g10269 ( 
.A(n_10147),
.Y(n_10269)
);

NAND2xp5_ASAP7_75t_L g10270 ( 
.A(n_10214),
.B(n_10052),
.Y(n_10270)
);

INVx1_ASAP7_75t_L g10271 ( 
.A(n_10189),
.Y(n_10271)
);

INVx1_ASAP7_75t_L g10272 ( 
.A(n_10138),
.Y(n_10272)
);

NAND2xp5_ASAP7_75t_L g10273 ( 
.A(n_10119),
.B(n_10081),
.Y(n_10273)
);

INVx2_ASAP7_75t_L g10274 ( 
.A(n_10137),
.Y(n_10274)
);

INVx1_ASAP7_75t_L g10275 ( 
.A(n_10194),
.Y(n_10275)
);

OAI222xp33_ASAP7_75t_L g10276 ( 
.A1(n_10128),
.A2(n_10111),
.B1(n_10198),
.B2(n_10109),
.C1(n_10099),
.C2(n_10116),
.Y(n_10276)
);

NAND4xp25_ASAP7_75t_L g10277 ( 
.A(n_10115),
.B(n_9916),
.C(n_10004),
.D(n_10034),
.Y(n_10277)
);

NAND2xp5_ASAP7_75t_L g10278 ( 
.A(n_10205),
.B(n_911),
.Y(n_10278)
);

OR2x2_ASAP7_75t_L g10279 ( 
.A(n_10173),
.B(n_911),
.Y(n_10279)
);

INVx2_ASAP7_75t_L g10280 ( 
.A(n_10195),
.Y(n_10280)
);

BUFx3_ASAP7_75t_L g10281 ( 
.A(n_10203),
.Y(n_10281)
);

OR2x2_ASAP7_75t_L g10282 ( 
.A(n_10212),
.B(n_912),
.Y(n_10282)
);

INVx1_ASAP7_75t_L g10283 ( 
.A(n_10178),
.Y(n_10283)
);

AND2x2_ASAP7_75t_L g10284 ( 
.A(n_10200),
.B(n_912),
.Y(n_10284)
);

AND2x2_ASAP7_75t_L g10285 ( 
.A(n_10201),
.B(n_10131),
.Y(n_10285)
);

INVx1_ASAP7_75t_L g10286 ( 
.A(n_10179),
.Y(n_10286)
);

AND2x2_ASAP7_75t_L g10287 ( 
.A(n_10163),
.B(n_912),
.Y(n_10287)
);

INVx1_ASAP7_75t_L g10288 ( 
.A(n_10197),
.Y(n_10288)
);

AND2x2_ASAP7_75t_L g10289 ( 
.A(n_10129),
.B(n_913),
.Y(n_10289)
);

OR2x2_ASAP7_75t_L g10290 ( 
.A(n_10184),
.B(n_913),
.Y(n_10290)
);

AND2x2_ASAP7_75t_L g10291 ( 
.A(n_10105),
.B(n_913),
.Y(n_10291)
);

INVx2_ASAP7_75t_L g10292 ( 
.A(n_10157),
.Y(n_10292)
);

AND2x2_ASAP7_75t_L g10293 ( 
.A(n_10107),
.B(n_914),
.Y(n_10293)
);

OAI211xp5_ASAP7_75t_SL g10294 ( 
.A1(n_10177),
.A2(n_922),
.B(n_930),
.C(n_914),
.Y(n_10294)
);

AND2x2_ASAP7_75t_SL g10295 ( 
.A(n_10148),
.B(n_914),
.Y(n_10295)
);

NAND2xp5_ASAP7_75t_L g10296 ( 
.A(n_10206),
.B(n_915),
.Y(n_10296)
);

NAND2xp5_ASAP7_75t_L g10297 ( 
.A(n_10208),
.B(n_915),
.Y(n_10297)
);

INVx2_ASAP7_75t_L g10298 ( 
.A(n_10218),
.Y(n_10298)
);

OR2x2_ASAP7_75t_L g10299 ( 
.A(n_10220),
.B(n_916),
.Y(n_10299)
);

INVx1_ASAP7_75t_L g10300 ( 
.A(n_10098),
.Y(n_10300)
);

AND4x1_ASAP7_75t_L g10301 ( 
.A(n_10162),
.B(n_10152),
.C(n_10187),
.D(n_10159),
.Y(n_10301)
);

INVx1_ASAP7_75t_L g10302 ( 
.A(n_10168),
.Y(n_10302)
);

NAND2xp5_ASAP7_75t_L g10303 ( 
.A(n_10209),
.B(n_916),
.Y(n_10303)
);

NOR3xp33_ASAP7_75t_L g10304 ( 
.A(n_10161),
.B(n_917),
.C(n_918),
.Y(n_10304)
);

AND2x2_ASAP7_75t_L g10305 ( 
.A(n_10139),
.B(n_917),
.Y(n_10305)
);

AND2x2_ASAP7_75t_L g10306 ( 
.A(n_10169),
.B(n_917),
.Y(n_10306)
);

INVx1_ASAP7_75t_L g10307 ( 
.A(n_10174),
.Y(n_10307)
);

INVx1_ASAP7_75t_L g10308 ( 
.A(n_10182),
.Y(n_10308)
);

AND2x2_ASAP7_75t_L g10309 ( 
.A(n_10135),
.B(n_918),
.Y(n_10309)
);

OR2x2_ASAP7_75t_L g10310 ( 
.A(n_10094),
.B(n_918),
.Y(n_10310)
);

NAND3xp33_ASAP7_75t_L g10311 ( 
.A(n_10234),
.B(n_919),
.C(n_920),
.Y(n_10311)
);

INVx2_ASAP7_75t_L g10312 ( 
.A(n_10154),
.Y(n_10312)
);

AOI22xp5_ASAP7_75t_L g10313 ( 
.A1(n_10140),
.A2(n_921),
.B1(n_919),
.B2(n_920),
.Y(n_10313)
);

OR2x2_ASAP7_75t_L g10314 ( 
.A(n_10104),
.B(n_919),
.Y(n_10314)
);

INVxp67_ASAP7_75t_SL g10315 ( 
.A(n_10171),
.Y(n_10315)
);

INVx1_ASAP7_75t_L g10316 ( 
.A(n_10103),
.Y(n_10316)
);

OR2x2_ASAP7_75t_L g10317 ( 
.A(n_10192),
.B(n_920),
.Y(n_10317)
);

INVxp67_ASAP7_75t_L g10318 ( 
.A(n_10175),
.Y(n_10318)
);

AND2x2_ASAP7_75t_L g10319 ( 
.A(n_10211),
.B(n_921),
.Y(n_10319)
);

INVx1_ASAP7_75t_L g10320 ( 
.A(n_10186),
.Y(n_10320)
);

INVx1_ASAP7_75t_SL g10321 ( 
.A(n_10149),
.Y(n_10321)
);

INVx1_ASAP7_75t_L g10322 ( 
.A(n_10155),
.Y(n_10322)
);

INVx1_ASAP7_75t_L g10323 ( 
.A(n_10207),
.Y(n_10323)
);

NAND2xp5_ASAP7_75t_L g10324 ( 
.A(n_10193),
.B(n_921),
.Y(n_10324)
);

INVx1_ASAP7_75t_L g10325 ( 
.A(n_10126),
.Y(n_10325)
);

OR2x2_ASAP7_75t_L g10326 ( 
.A(n_10136),
.B(n_922),
.Y(n_10326)
);

NAND2xp5_ASAP7_75t_L g10327 ( 
.A(n_10215),
.B(n_923),
.Y(n_10327)
);

INVx1_ASAP7_75t_L g10328 ( 
.A(n_10176),
.Y(n_10328)
);

INVx1_ASAP7_75t_L g10329 ( 
.A(n_10121),
.Y(n_10329)
);

AOI22xp5_ASAP7_75t_L g10330 ( 
.A1(n_10227),
.A2(n_925),
.B1(n_923),
.B2(n_924),
.Y(n_10330)
);

INVx1_ASAP7_75t_SL g10331 ( 
.A(n_10221),
.Y(n_10331)
);

NAND4xp25_ASAP7_75t_SL g10332 ( 
.A(n_10233),
.B(n_925),
.C(n_923),
.D(n_924),
.Y(n_10332)
);

INVxp67_ASAP7_75t_SL g10333 ( 
.A(n_10190),
.Y(n_10333)
);

AND2x2_ASAP7_75t_L g10334 ( 
.A(n_10196),
.B(n_10124),
.Y(n_10334)
);

AND2x2_ASAP7_75t_L g10335 ( 
.A(n_10185),
.B(n_926),
.Y(n_10335)
);

BUFx2_ASAP7_75t_L g10336 ( 
.A(n_10202),
.Y(n_10336)
);

AND2x2_ASAP7_75t_L g10337 ( 
.A(n_10150),
.B(n_926),
.Y(n_10337)
);

AND2x2_ASAP7_75t_L g10338 ( 
.A(n_10156),
.B(n_10158),
.Y(n_10338)
);

NOR3xp33_ASAP7_75t_SL g10339 ( 
.A(n_10127),
.B(n_926),
.C(n_927),
.Y(n_10339)
);

NAND3xp33_ASAP7_75t_L g10340 ( 
.A(n_10113),
.B(n_927),
.C(n_928),
.Y(n_10340)
);

OR2x2_ASAP7_75t_L g10341 ( 
.A(n_10087),
.B(n_928),
.Y(n_10341)
);

AND2x2_ASAP7_75t_L g10342 ( 
.A(n_10143),
.B(n_10133),
.Y(n_10342)
);

HB1xp67_ASAP7_75t_L g10343 ( 
.A(n_10219),
.Y(n_10343)
);

HB1xp67_ASAP7_75t_L g10344 ( 
.A(n_10188),
.Y(n_10344)
);

INVx1_ASAP7_75t_L g10345 ( 
.A(n_10132),
.Y(n_10345)
);

INVx1_ASAP7_75t_L g10346 ( 
.A(n_10117),
.Y(n_10346)
);

NOR3xp33_ASAP7_75t_L g10347 ( 
.A(n_10222),
.B(n_928),
.C(n_929),
.Y(n_10347)
);

NAND3xp33_ASAP7_75t_L g10348 ( 
.A(n_10130),
.B(n_929),
.C(n_930),
.Y(n_10348)
);

AOI211xp5_ASAP7_75t_L g10349 ( 
.A1(n_10183),
.A2(n_932),
.B(n_930),
.C(n_931),
.Y(n_10349)
);

OR2x2_ASAP7_75t_L g10350 ( 
.A(n_10160),
.B(n_932),
.Y(n_10350)
);

OAI31xp33_ASAP7_75t_L g10351 ( 
.A1(n_10216),
.A2(n_10224),
.A3(n_10165),
.B(n_10122),
.Y(n_10351)
);

INVx2_ASAP7_75t_L g10352 ( 
.A(n_10118),
.Y(n_10352)
);

NAND2xp5_ASAP7_75t_L g10353 ( 
.A(n_10225),
.B(n_10210),
.Y(n_10353)
);

AND2x2_ASAP7_75t_L g10354 ( 
.A(n_10226),
.B(n_932),
.Y(n_10354)
);

INVx2_ASAP7_75t_L g10355 ( 
.A(n_10125),
.Y(n_10355)
);

CKINVDCx16_ASAP7_75t_R g10356 ( 
.A(n_10223),
.Y(n_10356)
);

AND2x4_ASAP7_75t_L g10357 ( 
.A(n_10181),
.B(n_933),
.Y(n_10357)
);

NAND2xp5_ASAP7_75t_L g10358 ( 
.A(n_10232),
.B(n_933),
.Y(n_10358)
);

AO22x1_ASAP7_75t_L g10359 ( 
.A1(n_10172),
.A2(n_935),
.B1(n_933),
.B2(n_934),
.Y(n_10359)
);

OR2x2_ASAP7_75t_L g10360 ( 
.A(n_10180),
.B(n_934),
.Y(n_10360)
);

OR2x2_ASAP7_75t_L g10361 ( 
.A(n_10213),
.B(n_934),
.Y(n_10361)
);

AND2x2_ASAP7_75t_L g10362 ( 
.A(n_10236),
.B(n_10229),
.Y(n_10362)
);

NAND2x1p5_ASAP7_75t_L g10363 ( 
.A(n_10245),
.B(n_10231),
.Y(n_10363)
);

INVx3_ASAP7_75t_L g10364 ( 
.A(n_10281),
.Y(n_10364)
);

NAND2x1p5_ASAP7_75t_L g10365 ( 
.A(n_10266),
.B(n_10228),
.Y(n_10365)
);

NOR2xp33_ASAP7_75t_L g10366 ( 
.A(n_10318),
.B(n_10356),
.Y(n_10366)
);

OAI22xp33_ASAP7_75t_L g10367 ( 
.A1(n_10242),
.A2(n_10230),
.B1(n_937),
.B2(n_935),
.Y(n_10367)
);

OR2x2_ASAP7_75t_L g10368 ( 
.A(n_10273),
.B(n_935),
.Y(n_10368)
);

AND2x2_ASAP7_75t_L g10369 ( 
.A(n_10237),
.B(n_936),
.Y(n_10369)
);

AND2x4_ASAP7_75t_L g10370 ( 
.A(n_10246),
.B(n_936),
.Y(n_10370)
);

INVx1_ASAP7_75t_L g10371 ( 
.A(n_10249),
.Y(n_10371)
);

INVx1_ASAP7_75t_L g10372 ( 
.A(n_10260),
.Y(n_10372)
);

OR2x2_ASAP7_75t_L g10373 ( 
.A(n_10243),
.B(n_10241),
.Y(n_10373)
);

NAND2xp5_ASAP7_75t_L g10374 ( 
.A(n_10295),
.B(n_936),
.Y(n_10374)
);

NAND3xp33_ASAP7_75t_L g10375 ( 
.A(n_10240),
.B(n_937),
.C(n_938),
.Y(n_10375)
);

NAND2xp5_ASAP7_75t_L g10376 ( 
.A(n_10359),
.B(n_938),
.Y(n_10376)
);

OR2x2_ASAP7_75t_L g10377 ( 
.A(n_10248),
.B(n_938),
.Y(n_10377)
);

AND2x2_ASAP7_75t_SL g10378 ( 
.A(n_10304),
.B(n_10336),
.Y(n_10378)
);

INVx1_ASAP7_75t_L g10379 ( 
.A(n_10265),
.Y(n_10379)
);

OR2x2_ASAP7_75t_L g10380 ( 
.A(n_10331),
.B(n_939),
.Y(n_10380)
);

AND2x2_ASAP7_75t_L g10381 ( 
.A(n_10235),
.B(n_939),
.Y(n_10381)
);

AOI21xp33_ASAP7_75t_L g10382 ( 
.A1(n_10238),
.A2(n_939),
.B(n_940),
.Y(n_10382)
);

INVx1_ASAP7_75t_L g10383 ( 
.A(n_10343),
.Y(n_10383)
);

NAND2xp5_ASAP7_75t_L g10384 ( 
.A(n_10261),
.B(n_940),
.Y(n_10384)
);

AND2x4_ASAP7_75t_L g10385 ( 
.A(n_10274),
.B(n_941),
.Y(n_10385)
);

INVx1_ASAP7_75t_L g10386 ( 
.A(n_10287),
.Y(n_10386)
);

NOR2xp33_ASAP7_75t_L g10387 ( 
.A(n_10276),
.B(n_941),
.Y(n_10387)
);

OAI321xp33_ASAP7_75t_L g10388 ( 
.A1(n_10277),
.A2(n_943),
.A3(n_945),
.B1(n_941),
.B2(n_942),
.C(n_944),
.Y(n_10388)
);

AND2x4_ASAP7_75t_SL g10389 ( 
.A(n_10292),
.B(n_942),
.Y(n_10389)
);

AND2x2_ASAP7_75t_L g10390 ( 
.A(n_10334),
.B(n_943),
.Y(n_10390)
);

INVx1_ASAP7_75t_L g10391 ( 
.A(n_10259),
.Y(n_10391)
);

OR2x2_ASAP7_75t_L g10392 ( 
.A(n_10269),
.B(n_943),
.Y(n_10392)
);

INVx2_ASAP7_75t_SL g10393 ( 
.A(n_10253),
.Y(n_10393)
);

OR2x2_ASAP7_75t_L g10394 ( 
.A(n_10353),
.B(n_944),
.Y(n_10394)
);

NAND2xp5_ASAP7_75t_L g10395 ( 
.A(n_10268),
.B(n_10319),
.Y(n_10395)
);

OAI21xp5_ASAP7_75t_L g10396 ( 
.A1(n_10262),
.A2(n_952),
.B(n_944),
.Y(n_10396)
);

AND2x2_ASAP7_75t_L g10397 ( 
.A(n_10239),
.B(n_945),
.Y(n_10397)
);

NOR2xp33_ASAP7_75t_L g10398 ( 
.A(n_10332),
.B(n_945),
.Y(n_10398)
);

INVx1_ASAP7_75t_L g10399 ( 
.A(n_10309),
.Y(n_10399)
);

AND2x2_ASAP7_75t_L g10400 ( 
.A(n_10285),
.B(n_946),
.Y(n_10400)
);

INVx2_ASAP7_75t_L g10401 ( 
.A(n_10357),
.Y(n_10401)
);

A2O1A1Ixp33_ASAP7_75t_L g10402 ( 
.A1(n_10339),
.A2(n_948),
.B(n_946),
.C(n_947),
.Y(n_10402)
);

INVx2_ASAP7_75t_L g10403 ( 
.A(n_10357),
.Y(n_10403)
);

NOR2xp33_ASAP7_75t_L g10404 ( 
.A(n_10279),
.B(n_948),
.Y(n_10404)
);

AND2x4_ASAP7_75t_L g10405 ( 
.A(n_10271),
.B(n_948),
.Y(n_10405)
);

INVx1_ASAP7_75t_SL g10406 ( 
.A(n_10290),
.Y(n_10406)
);

AOI211x1_ASAP7_75t_L g10407 ( 
.A1(n_10301),
.A2(n_951),
.B(n_949),
.C(n_950),
.Y(n_10407)
);

INVx1_ASAP7_75t_L g10408 ( 
.A(n_10252),
.Y(n_10408)
);

INVx1_ASAP7_75t_L g10409 ( 
.A(n_10289),
.Y(n_10409)
);

INVx1_ASAP7_75t_L g10410 ( 
.A(n_10291),
.Y(n_10410)
);

NAND2xp5_ASAP7_75t_L g10411 ( 
.A(n_10247),
.B(n_949),
.Y(n_10411)
);

INVx2_ASAP7_75t_L g10412 ( 
.A(n_10326),
.Y(n_10412)
);

INVx1_ASAP7_75t_L g10413 ( 
.A(n_10293),
.Y(n_10413)
);

INVx1_ASAP7_75t_L g10414 ( 
.A(n_10335),
.Y(n_10414)
);

AND2x2_ASAP7_75t_L g10415 ( 
.A(n_10255),
.B(n_950),
.Y(n_10415)
);

NAND2xp5_ASAP7_75t_L g10416 ( 
.A(n_10256),
.B(n_950),
.Y(n_10416)
);

NAND2xp5_ASAP7_75t_L g10417 ( 
.A(n_10264),
.B(n_951),
.Y(n_10417)
);

NOR2xp67_ASAP7_75t_L g10418 ( 
.A(n_10244),
.B(n_951),
.Y(n_10418)
);

AND2x4_ASAP7_75t_L g10419 ( 
.A(n_10338),
.B(n_952),
.Y(n_10419)
);

OR2x2_ASAP7_75t_L g10420 ( 
.A(n_10299),
.B(n_953),
.Y(n_10420)
);

INVx1_ASAP7_75t_L g10421 ( 
.A(n_10258),
.Y(n_10421)
);

INVx1_ASAP7_75t_L g10422 ( 
.A(n_10263),
.Y(n_10422)
);

INVx1_ASAP7_75t_L g10423 ( 
.A(n_10337),
.Y(n_10423)
);

AND2x4_ASAP7_75t_SL g10424 ( 
.A(n_10312),
.B(n_953),
.Y(n_10424)
);

INVx2_ASAP7_75t_L g10425 ( 
.A(n_10306),
.Y(n_10425)
);

AND2x2_ASAP7_75t_L g10426 ( 
.A(n_10342),
.B(n_954),
.Y(n_10426)
);

INVxp67_ASAP7_75t_L g10427 ( 
.A(n_10282),
.Y(n_10427)
);

INVx1_ASAP7_75t_L g10428 ( 
.A(n_10284),
.Y(n_10428)
);

INVx1_ASAP7_75t_L g10429 ( 
.A(n_10278),
.Y(n_10429)
);

AND2x2_ASAP7_75t_L g10430 ( 
.A(n_10275),
.B(n_954),
.Y(n_10430)
);

NAND2xp5_ASAP7_75t_L g10431 ( 
.A(n_10321),
.B(n_954),
.Y(n_10431)
);

INVx2_ASAP7_75t_L g10432 ( 
.A(n_10350),
.Y(n_10432)
);

INVx1_ASAP7_75t_L g10433 ( 
.A(n_10310),
.Y(n_10433)
);

INVx1_ASAP7_75t_L g10434 ( 
.A(n_10344),
.Y(n_10434)
);

INVx1_ASAP7_75t_L g10435 ( 
.A(n_10305),
.Y(n_10435)
);

AND2x2_ASAP7_75t_SL g10436 ( 
.A(n_10325),
.B(n_955),
.Y(n_10436)
);

AND2x2_ASAP7_75t_L g10437 ( 
.A(n_10283),
.B(n_955),
.Y(n_10437)
);

OR2x2_ASAP7_75t_L g10438 ( 
.A(n_10314),
.B(n_956),
.Y(n_10438)
);

AND2x2_ASAP7_75t_L g10439 ( 
.A(n_10286),
.B(n_956),
.Y(n_10439)
);

AND2x2_ASAP7_75t_L g10440 ( 
.A(n_10288),
.B(n_956),
.Y(n_10440)
);

BUFx2_ASAP7_75t_L g10441 ( 
.A(n_10345),
.Y(n_10441)
);

INVx1_ASAP7_75t_SL g10442 ( 
.A(n_10317),
.Y(n_10442)
);

INVx1_ASAP7_75t_SL g10443 ( 
.A(n_10341),
.Y(n_10443)
);

AND2x2_ASAP7_75t_L g10444 ( 
.A(n_10302),
.B(n_957),
.Y(n_10444)
);

NAND2xp5_ASAP7_75t_L g10445 ( 
.A(n_10250),
.B(n_957),
.Y(n_10445)
);

AND2x2_ASAP7_75t_L g10446 ( 
.A(n_10307),
.B(n_957),
.Y(n_10446)
);

NAND2xp5_ASAP7_75t_L g10447 ( 
.A(n_10308),
.B(n_958),
.Y(n_10447)
);

NAND2xp5_ASAP7_75t_L g10448 ( 
.A(n_10272),
.B(n_10315),
.Y(n_10448)
);

INVx1_ASAP7_75t_L g10449 ( 
.A(n_10257),
.Y(n_10449)
);

AND2x2_ASAP7_75t_L g10450 ( 
.A(n_10322),
.B(n_958),
.Y(n_10450)
);

INVx1_ASAP7_75t_SL g10451 ( 
.A(n_10354),
.Y(n_10451)
);

OAI22xp33_ASAP7_75t_L g10452 ( 
.A1(n_10270),
.A2(n_961),
.B1(n_959),
.B2(n_960),
.Y(n_10452)
);

INVx1_ASAP7_75t_L g10453 ( 
.A(n_10360),
.Y(n_10453)
);

NAND2xp5_ASAP7_75t_L g10454 ( 
.A(n_10349),
.B(n_959),
.Y(n_10454)
);

INVx2_ASAP7_75t_SL g10455 ( 
.A(n_10254),
.Y(n_10455)
);

OR2x2_ASAP7_75t_L g10456 ( 
.A(n_10280),
.B(n_10298),
.Y(n_10456)
);

OR2x2_ASAP7_75t_L g10457 ( 
.A(n_10329),
.B(n_959),
.Y(n_10457)
);

OAI22xp5_ASAP7_75t_L g10458 ( 
.A1(n_10330),
.A2(n_962),
.B1(n_960),
.B2(n_961),
.Y(n_10458)
);

OR2x6_ASAP7_75t_L g10459 ( 
.A(n_10328),
.B(n_961),
.Y(n_10459)
);

AND2x2_ASAP7_75t_L g10460 ( 
.A(n_10333),
.B(n_10320),
.Y(n_10460)
);

INVx1_ASAP7_75t_L g10461 ( 
.A(n_10324),
.Y(n_10461)
);

NAND2xp5_ASAP7_75t_L g10462 ( 
.A(n_10323),
.B(n_960),
.Y(n_10462)
);

NOR2xp33_ASAP7_75t_L g10463 ( 
.A(n_10294),
.B(n_962),
.Y(n_10463)
);

OR2x6_ASAP7_75t_L g10464 ( 
.A(n_10346),
.B(n_10327),
.Y(n_10464)
);

NAND2xp5_ASAP7_75t_L g10465 ( 
.A(n_10347),
.B(n_10313),
.Y(n_10465)
);

AND2x2_ASAP7_75t_L g10466 ( 
.A(n_10267),
.B(n_962),
.Y(n_10466)
);

INVx3_ASAP7_75t_L g10467 ( 
.A(n_10352),
.Y(n_10467)
);

INVx2_ASAP7_75t_L g10468 ( 
.A(n_10361),
.Y(n_10468)
);

INVx2_ASAP7_75t_L g10469 ( 
.A(n_10251),
.Y(n_10469)
);

NAND2xp5_ASAP7_75t_L g10470 ( 
.A(n_10364),
.B(n_10300),
.Y(n_10470)
);

NAND2xp5_ASAP7_75t_SL g10471 ( 
.A(n_10378),
.B(n_10351),
.Y(n_10471)
);

NAND2xp5_ASAP7_75t_L g10472 ( 
.A(n_10369),
.B(n_10316),
.Y(n_10472)
);

INVx1_ASAP7_75t_L g10473 ( 
.A(n_10365),
.Y(n_10473)
);

OR2x2_ASAP7_75t_L g10474 ( 
.A(n_10395),
.B(n_10296),
.Y(n_10474)
);

NAND2xp5_ASAP7_75t_L g10475 ( 
.A(n_10436),
.B(n_10355),
.Y(n_10475)
);

AND2x2_ASAP7_75t_L g10476 ( 
.A(n_10362),
.B(n_10297),
.Y(n_10476)
);

NAND2xp5_ASAP7_75t_L g10477 ( 
.A(n_10407),
.B(n_10418),
.Y(n_10477)
);

AND2x2_ASAP7_75t_L g10478 ( 
.A(n_10408),
.B(n_10303),
.Y(n_10478)
);

AND2x2_ASAP7_75t_L g10479 ( 
.A(n_10363),
.B(n_10358),
.Y(n_10479)
);

AND2x2_ASAP7_75t_L g10480 ( 
.A(n_10421),
.B(n_10311),
.Y(n_10480)
);

OAI211xp5_ASAP7_75t_L g10481 ( 
.A1(n_10387),
.A2(n_10348),
.B(n_10340),
.C(n_965),
.Y(n_10481)
);

INVx1_ASAP7_75t_L g10482 ( 
.A(n_10389),
.Y(n_10482)
);

INVx1_ASAP7_75t_L g10483 ( 
.A(n_10390),
.Y(n_10483)
);

AND2x2_ASAP7_75t_L g10484 ( 
.A(n_10422),
.B(n_963),
.Y(n_10484)
);

NAND2xp5_ASAP7_75t_L g10485 ( 
.A(n_10401),
.B(n_963),
.Y(n_10485)
);

AND2x2_ASAP7_75t_L g10486 ( 
.A(n_10455),
.B(n_963),
.Y(n_10486)
);

AND2x2_ASAP7_75t_L g10487 ( 
.A(n_10460),
.B(n_964),
.Y(n_10487)
);

OAI21x1_ASAP7_75t_SL g10488 ( 
.A1(n_10376),
.A2(n_972),
.B(n_964),
.Y(n_10488)
);

INVxp67_ASAP7_75t_L g10489 ( 
.A(n_10366),
.Y(n_10489)
);

INVx1_ASAP7_75t_L g10490 ( 
.A(n_10424),
.Y(n_10490)
);

INVx2_ASAP7_75t_SL g10491 ( 
.A(n_10403),
.Y(n_10491)
);

OA21x2_ASAP7_75t_SL g10492 ( 
.A1(n_10451),
.A2(n_964),
.B(n_965),
.Y(n_10492)
);

INVx1_ASAP7_75t_L g10493 ( 
.A(n_10426),
.Y(n_10493)
);

HB1xp67_ASAP7_75t_L g10494 ( 
.A(n_10459),
.Y(n_10494)
);

AND2x2_ASAP7_75t_L g10495 ( 
.A(n_10425),
.B(n_966),
.Y(n_10495)
);

NAND2xp33_ASAP7_75t_L g10496 ( 
.A(n_10402),
.B(n_966),
.Y(n_10496)
);

OAI21xp5_ASAP7_75t_SL g10497 ( 
.A1(n_10372),
.A2(n_967),
.B(n_968),
.Y(n_10497)
);

NAND2xp5_ASAP7_75t_L g10498 ( 
.A(n_10370),
.B(n_967),
.Y(n_10498)
);

NAND2xp5_ASAP7_75t_L g10499 ( 
.A(n_10393),
.B(n_10371),
.Y(n_10499)
);

NOR2xp33_ASAP7_75t_L g10500 ( 
.A(n_10373),
.B(n_10427),
.Y(n_10500)
);

AND2x2_ASAP7_75t_L g10501 ( 
.A(n_10386),
.B(n_967),
.Y(n_10501)
);

NOR2x1_ASAP7_75t_L g10502 ( 
.A(n_10375),
.B(n_968),
.Y(n_10502)
);

NAND2xp5_ASAP7_75t_L g10503 ( 
.A(n_10385),
.B(n_969),
.Y(n_10503)
);

AND2x4_ASAP7_75t_L g10504 ( 
.A(n_10441),
.B(n_969),
.Y(n_10504)
);

NAND2xp5_ASAP7_75t_L g10505 ( 
.A(n_10415),
.B(n_969),
.Y(n_10505)
);

INVx1_ASAP7_75t_L g10506 ( 
.A(n_10381),
.Y(n_10506)
);

NAND2xp5_ASAP7_75t_L g10507 ( 
.A(n_10419),
.B(n_970),
.Y(n_10507)
);

OR2x2_ASAP7_75t_L g10508 ( 
.A(n_10384),
.B(n_970),
.Y(n_10508)
);

OR2x2_ASAP7_75t_L g10509 ( 
.A(n_10380),
.B(n_971),
.Y(n_10509)
);

INVx1_ASAP7_75t_L g10510 ( 
.A(n_10397),
.Y(n_10510)
);

AND2x2_ASAP7_75t_L g10511 ( 
.A(n_10399),
.B(n_971),
.Y(n_10511)
);

INVx2_ASAP7_75t_L g10512 ( 
.A(n_10459),
.Y(n_10512)
);

INVx2_ASAP7_75t_L g10513 ( 
.A(n_10392),
.Y(n_10513)
);

INVx1_ASAP7_75t_L g10514 ( 
.A(n_10400),
.Y(n_10514)
);

OAI21x1_ASAP7_75t_L g10515 ( 
.A1(n_10374),
.A2(n_971),
.B(n_972),
.Y(n_10515)
);

AND2x4_ASAP7_75t_L g10516 ( 
.A(n_10383),
.B(n_973),
.Y(n_10516)
);

NAND2xp5_ASAP7_75t_L g10517 ( 
.A(n_10398),
.B(n_973),
.Y(n_10517)
);

OAI21xp33_ASAP7_75t_L g10518 ( 
.A1(n_10465),
.A2(n_973),
.B(n_974),
.Y(n_10518)
);

NAND2xp5_ASAP7_75t_SL g10519 ( 
.A(n_10388),
.B(n_974),
.Y(n_10519)
);

INVx1_ASAP7_75t_SL g10520 ( 
.A(n_10443),
.Y(n_10520)
);

BUFx2_ASAP7_75t_L g10521 ( 
.A(n_10464),
.Y(n_10521)
);

BUFx3_ASAP7_75t_L g10522 ( 
.A(n_10449),
.Y(n_10522)
);

NAND2xp5_ASAP7_75t_SL g10523 ( 
.A(n_10442),
.B(n_975),
.Y(n_10523)
);

INVx1_ASAP7_75t_L g10524 ( 
.A(n_10377),
.Y(n_10524)
);

AND2x2_ASAP7_75t_L g10525 ( 
.A(n_10414),
.B(n_975),
.Y(n_10525)
);

INVx1_ASAP7_75t_L g10526 ( 
.A(n_10430),
.Y(n_10526)
);

INVx1_ASAP7_75t_SL g10527 ( 
.A(n_10406),
.Y(n_10527)
);

INVx1_ASAP7_75t_L g10528 ( 
.A(n_10437),
.Y(n_10528)
);

INVx3_ASAP7_75t_SL g10529 ( 
.A(n_10405),
.Y(n_10529)
);

HB1xp67_ASAP7_75t_L g10530 ( 
.A(n_10464),
.Y(n_10530)
);

INVx1_ASAP7_75t_L g10531 ( 
.A(n_10439),
.Y(n_10531)
);

INVx1_ASAP7_75t_L g10532 ( 
.A(n_10440),
.Y(n_10532)
);

INVx1_ASAP7_75t_L g10533 ( 
.A(n_10444),
.Y(n_10533)
);

INVx1_ASAP7_75t_L g10534 ( 
.A(n_10446),
.Y(n_10534)
);

AOI222xp33_ASAP7_75t_L g10535 ( 
.A1(n_10396),
.A2(n_977),
.B1(n_979),
.B2(n_975),
.C1(n_976),
.C2(n_978),
.Y(n_10535)
);

INVx1_ASAP7_75t_SL g10536 ( 
.A(n_10456),
.Y(n_10536)
);

INVx2_ASAP7_75t_L g10537 ( 
.A(n_10420),
.Y(n_10537)
);

NAND2xp5_ASAP7_75t_L g10538 ( 
.A(n_10463),
.B(n_976),
.Y(n_10538)
);

NAND2xp5_ASAP7_75t_L g10539 ( 
.A(n_10379),
.B(n_976),
.Y(n_10539)
);

HB1xp67_ASAP7_75t_L g10540 ( 
.A(n_10438),
.Y(n_10540)
);

INVx1_ASAP7_75t_L g10541 ( 
.A(n_10450),
.Y(n_10541)
);

INVx2_ASAP7_75t_L g10542 ( 
.A(n_10457),
.Y(n_10542)
);

NOR2xp33_ASAP7_75t_L g10543 ( 
.A(n_10423),
.B(n_977),
.Y(n_10543)
);

INVx2_ASAP7_75t_SL g10544 ( 
.A(n_10434),
.Y(n_10544)
);

NAND2x1p5_ASAP7_75t_L g10545 ( 
.A(n_10467),
.B(n_10433),
.Y(n_10545)
);

AND2x2_ASAP7_75t_L g10546 ( 
.A(n_10409),
.B(n_978),
.Y(n_10546)
);

INVx1_ASAP7_75t_L g10547 ( 
.A(n_10431),
.Y(n_10547)
);

NAND2xp5_ASAP7_75t_L g10548 ( 
.A(n_10410),
.B(n_978),
.Y(n_10548)
);

AND4x1_ASAP7_75t_L g10549 ( 
.A(n_10404),
.B(n_981),
.C(n_979),
.D(n_980),
.Y(n_10549)
);

NAND2xp5_ASAP7_75t_L g10550 ( 
.A(n_10413),
.B(n_979),
.Y(n_10550)
);

OR2x2_ASAP7_75t_L g10551 ( 
.A(n_10394),
.B(n_980),
.Y(n_10551)
);

INVx1_ASAP7_75t_L g10552 ( 
.A(n_10466),
.Y(n_10552)
);

OR2x6_ASAP7_75t_L g10553 ( 
.A(n_10469),
.B(n_980),
.Y(n_10553)
);

INVx1_ASAP7_75t_L g10554 ( 
.A(n_10411),
.Y(n_10554)
);

AOI221xp5_ASAP7_75t_L g10555 ( 
.A1(n_10367),
.A2(n_984),
.B1(n_981),
.B2(n_983),
.C(n_985),
.Y(n_10555)
);

NAND2xp5_ASAP7_75t_L g10556 ( 
.A(n_10428),
.B(n_981),
.Y(n_10556)
);

AOI221xp5_ASAP7_75t_L g10557 ( 
.A1(n_10382),
.A2(n_986),
.B1(n_983),
.B2(n_985),
.C(n_987),
.Y(n_10557)
);

INVx2_ASAP7_75t_SL g10558 ( 
.A(n_10412),
.Y(n_10558)
);

AOI22xp33_ASAP7_75t_L g10559 ( 
.A1(n_10445),
.A2(n_987),
.B1(n_985),
.B2(n_986),
.Y(n_10559)
);

NAND2xp5_ASAP7_75t_L g10560 ( 
.A(n_10435),
.B(n_987),
.Y(n_10560)
);

INVx1_ASAP7_75t_L g10561 ( 
.A(n_10417),
.Y(n_10561)
);

INVx2_ASAP7_75t_L g10562 ( 
.A(n_10468),
.Y(n_10562)
);

INVx1_ASAP7_75t_L g10563 ( 
.A(n_10462),
.Y(n_10563)
);

INVx2_ASAP7_75t_SL g10564 ( 
.A(n_10432),
.Y(n_10564)
);

AND2x4_ASAP7_75t_SL g10565 ( 
.A(n_10453),
.B(n_989),
.Y(n_10565)
);

XOR2xp5_ASAP7_75t_L g10566 ( 
.A(n_10368),
.B(n_989),
.Y(n_10566)
);

NAND2xp5_ASAP7_75t_L g10567 ( 
.A(n_10391),
.B(n_989),
.Y(n_10567)
);

AND2x2_ASAP7_75t_L g10568 ( 
.A(n_10429),
.B(n_990),
.Y(n_10568)
);

NAND2xp5_ASAP7_75t_L g10569 ( 
.A(n_10452),
.B(n_990),
.Y(n_10569)
);

INVx2_ASAP7_75t_L g10570 ( 
.A(n_10461),
.Y(n_10570)
);

AND2x2_ASAP7_75t_L g10571 ( 
.A(n_10448),
.B(n_990),
.Y(n_10571)
);

AND2x2_ASAP7_75t_L g10572 ( 
.A(n_10454),
.B(n_991),
.Y(n_10572)
);

INVx1_ASAP7_75t_L g10573 ( 
.A(n_10447),
.Y(n_10573)
);

NAND2xp5_ASAP7_75t_L g10574 ( 
.A(n_10458),
.B(n_991),
.Y(n_10574)
);

OAI21xp5_ASAP7_75t_SL g10575 ( 
.A1(n_10416),
.A2(n_992),
.B(n_993),
.Y(n_10575)
);

NAND2x2_ASAP7_75t_L g10576 ( 
.A(n_10455),
.B(n_992),
.Y(n_10576)
);

AND3x2_ASAP7_75t_L g10577 ( 
.A(n_10441),
.B(n_992),
.C(n_993),
.Y(n_10577)
);

NAND4xp25_ASAP7_75t_L g10578 ( 
.A(n_10366),
.B(n_995),
.C(n_993),
.D(n_994),
.Y(n_10578)
);

OR2x2_ASAP7_75t_L g10579 ( 
.A(n_10365),
.B(n_994),
.Y(n_10579)
);

INVx1_ASAP7_75t_SL g10580 ( 
.A(n_10389),
.Y(n_10580)
);

NAND2xp5_ASAP7_75t_L g10581 ( 
.A(n_10577),
.B(n_995),
.Y(n_10581)
);

AND2x2_ASAP7_75t_L g10582 ( 
.A(n_10529),
.B(n_995),
.Y(n_10582)
);

OAI21xp5_ASAP7_75t_L g10583 ( 
.A1(n_10471),
.A2(n_996),
.B(n_997),
.Y(n_10583)
);

AOI21xp33_ASAP7_75t_SL g10584 ( 
.A1(n_10545),
.A2(n_996),
.B(n_997),
.Y(n_10584)
);

OAI22xp5_ASAP7_75t_L g10585 ( 
.A1(n_10576),
.A2(n_999),
.B1(n_997),
.B2(n_998),
.Y(n_10585)
);

OAI21xp5_ASAP7_75t_SL g10586 ( 
.A1(n_10536),
.A2(n_999),
.B(n_1000),
.Y(n_10586)
);

INVx1_ASAP7_75t_L g10587 ( 
.A(n_10494),
.Y(n_10587)
);

INVx1_ASAP7_75t_L g10588 ( 
.A(n_10579),
.Y(n_10588)
);

INVx1_ASAP7_75t_L g10589 ( 
.A(n_10530),
.Y(n_10589)
);

NAND2xp5_ASAP7_75t_L g10590 ( 
.A(n_10580),
.B(n_999),
.Y(n_10590)
);

A2O1A1Ixp33_ASAP7_75t_L g10591 ( 
.A1(n_10500),
.A2(n_1003),
.B(n_1001),
.C(n_1002),
.Y(n_10591)
);

OAI221xp5_ASAP7_75t_L g10592 ( 
.A1(n_10489),
.A2(n_10527),
.B1(n_10520),
.B2(n_10491),
.C(n_10473),
.Y(n_10592)
);

A2O1A1Ixp33_ASAP7_75t_L g10593 ( 
.A1(n_10497),
.A2(n_1003),
.B(n_1001),
.C(n_1002),
.Y(n_10593)
);

NOR2xp33_ASAP7_75t_L g10594 ( 
.A(n_10549),
.B(n_1002),
.Y(n_10594)
);

HB1xp67_ASAP7_75t_L g10595 ( 
.A(n_10553),
.Y(n_10595)
);

OAI21xp5_ASAP7_75t_L g10596 ( 
.A1(n_10477),
.A2(n_1003),
.B(n_1004),
.Y(n_10596)
);

AO221x1_ASAP7_75t_L g10597 ( 
.A1(n_10488),
.A2(n_1006),
.B1(n_1004),
.B2(n_1005),
.C(n_1007),
.Y(n_10597)
);

AOI22xp5_ASAP7_75t_L g10598 ( 
.A1(n_10482),
.A2(n_1008),
.B1(n_1005),
.B2(n_1006),
.Y(n_10598)
);

NOR2xp33_ASAP7_75t_SL g10599 ( 
.A(n_10521),
.B(n_1005),
.Y(n_10599)
);

NOR2xp33_ASAP7_75t_L g10600 ( 
.A(n_10578),
.B(n_1006),
.Y(n_10600)
);

NAND2xp5_ASAP7_75t_L g10601 ( 
.A(n_10504),
.B(n_1008),
.Y(n_10601)
);

AOI22xp5_ASAP7_75t_L g10602 ( 
.A1(n_10558),
.A2(n_1010),
.B1(n_1008),
.B2(n_1009),
.Y(n_10602)
);

NAND2xp5_ASAP7_75t_L g10603 ( 
.A(n_10512),
.B(n_1009),
.Y(n_10603)
);

INVx1_ASAP7_75t_L g10604 ( 
.A(n_10565),
.Y(n_10604)
);

AOI221xp5_ASAP7_75t_L g10605 ( 
.A1(n_10481),
.A2(n_1011),
.B1(n_1009),
.B2(n_1010),
.C(n_1012),
.Y(n_10605)
);

INVx1_ASAP7_75t_L g10606 ( 
.A(n_10487),
.Y(n_10606)
);

AND2x2_ASAP7_75t_L g10607 ( 
.A(n_10490),
.B(n_1011),
.Y(n_10607)
);

AOI21xp5_ASAP7_75t_L g10608 ( 
.A1(n_10519),
.A2(n_1013),
.B(n_1014),
.Y(n_10608)
);

BUFx2_ASAP7_75t_L g10609 ( 
.A(n_10553),
.Y(n_10609)
);

OAI21xp33_ASAP7_75t_L g10610 ( 
.A1(n_10499),
.A2(n_1013),
.B(n_1014),
.Y(n_10610)
);

INVxp67_ASAP7_75t_SL g10611 ( 
.A(n_10475),
.Y(n_10611)
);

INVx1_ASAP7_75t_L g10612 ( 
.A(n_10566),
.Y(n_10612)
);

INVx2_ASAP7_75t_L g10613 ( 
.A(n_10516),
.Y(n_10613)
);

INVx1_ASAP7_75t_L g10614 ( 
.A(n_10486),
.Y(n_10614)
);

AOI22xp33_ASAP7_75t_SL g10615 ( 
.A1(n_10522),
.A2(n_1022),
.B1(n_1030),
.B2(n_1014),
.Y(n_10615)
);

NOR2xp33_ASAP7_75t_L g10616 ( 
.A(n_10483),
.B(n_1015),
.Y(n_10616)
);

INVx1_ASAP7_75t_L g10617 ( 
.A(n_10540),
.Y(n_10617)
);

AOI21xp5_ASAP7_75t_SL g10618 ( 
.A1(n_10523),
.A2(n_1015),
.B(n_1016),
.Y(n_10618)
);

AND2x2_ASAP7_75t_L g10619 ( 
.A(n_10479),
.B(n_1015),
.Y(n_10619)
);

AOI211xp5_ASAP7_75t_SL g10620 ( 
.A1(n_10496),
.A2(n_1024),
.B(n_1032),
.C(n_1016),
.Y(n_10620)
);

INVx2_ASAP7_75t_SL g10621 ( 
.A(n_10516),
.Y(n_10621)
);

OR2x2_ASAP7_75t_L g10622 ( 
.A(n_10472),
.B(n_1016),
.Y(n_10622)
);

AOI22xp5_ASAP7_75t_L g10623 ( 
.A1(n_10564),
.A2(n_1019),
.B1(n_1017),
.B2(n_1018),
.Y(n_10623)
);

AOI21xp33_ASAP7_75t_L g10624 ( 
.A1(n_10470),
.A2(n_1017),
.B(n_1018),
.Y(n_10624)
);

AOI22xp5_ASAP7_75t_L g10625 ( 
.A1(n_10480),
.A2(n_1021),
.B1(n_1019),
.B2(n_1020),
.Y(n_10625)
);

AND2x2_ASAP7_75t_L g10626 ( 
.A(n_10476),
.B(n_1019),
.Y(n_10626)
);

NOR2xp33_ASAP7_75t_L g10627 ( 
.A(n_10506),
.B(n_1020),
.Y(n_10627)
);

AND2x2_ASAP7_75t_L g10628 ( 
.A(n_10514),
.B(n_1020),
.Y(n_10628)
);

AOI211xp5_ASAP7_75t_SL g10629 ( 
.A1(n_10493),
.A2(n_1029),
.B(n_1037),
.C(n_1021),
.Y(n_10629)
);

OR2x2_ASAP7_75t_L g10630 ( 
.A(n_10485),
.B(n_1021),
.Y(n_10630)
);

OR2x2_ASAP7_75t_L g10631 ( 
.A(n_10510),
.B(n_1022),
.Y(n_10631)
);

NAND2xp33_ASAP7_75t_L g10632 ( 
.A(n_10502),
.B(n_1022),
.Y(n_10632)
);

INVx1_ASAP7_75t_L g10633 ( 
.A(n_10501),
.Y(n_10633)
);

AND2x4_ASAP7_75t_L g10634 ( 
.A(n_10513),
.B(n_10495),
.Y(n_10634)
);

AOI22xp5_ASAP7_75t_L g10635 ( 
.A1(n_10544),
.A2(n_1025),
.B1(n_1023),
.B2(n_1024),
.Y(n_10635)
);

INVx1_ASAP7_75t_L g10636 ( 
.A(n_10511),
.Y(n_10636)
);

INVx1_ASAP7_75t_L g10637 ( 
.A(n_10484),
.Y(n_10637)
);

INVx1_ASAP7_75t_L g10638 ( 
.A(n_10509),
.Y(n_10638)
);

INVx2_ASAP7_75t_L g10639 ( 
.A(n_10551),
.Y(n_10639)
);

NAND2xp5_ASAP7_75t_L g10640 ( 
.A(n_10525),
.B(n_1023),
.Y(n_10640)
);

INVx1_ASAP7_75t_L g10641 ( 
.A(n_10546),
.Y(n_10641)
);

NOR2xp33_ASAP7_75t_L g10642 ( 
.A(n_10518),
.B(n_1023),
.Y(n_10642)
);

INVx1_ASAP7_75t_L g10643 ( 
.A(n_10498),
.Y(n_10643)
);

INVx1_ASAP7_75t_L g10644 ( 
.A(n_10503),
.Y(n_10644)
);

NAND2xp5_ASAP7_75t_L g10645 ( 
.A(n_10526),
.B(n_10528),
.Y(n_10645)
);

OAI21xp33_ASAP7_75t_SL g10646 ( 
.A1(n_10524),
.A2(n_1025),
.B(n_1026),
.Y(n_10646)
);

NOR2xp33_ASAP7_75t_L g10647 ( 
.A(n_10531),
.B(n_10532),
.Y(n_10647)
);

AOI221xp5_ASAP7_75t_L g10648 ( 
.A1(n_10533),
.A2(n_1027),
.B1(n_1025),
.B2(n_1026),
.C(n_1028),
.Y(n_10648)
);

INVx1_ASAP7_75t_L g10649 ( 
.A(n_10505),
.Y(n_10649)
);

INVx1_ASAP7_75t_L g10650 ( 
.A(n_10507),
.Y(n_10650)
);

OAI32xp33_ASAP7_75t_L g10651 ( 
.A1(n_10539),
.A2(n_1028),
.A3(n_1026),
.B1(n_1027),
.B2(n_1029),
.Y(n_10651)
);

INVxp67_ASAP7_75t_L g10652 ( 
.A(n_10543),
.Y(n_10652)
);

AOI221xp5_ASAP7_75t_L g10653 ( 
.A1(n_10534),
.A2(n_10541),
.B1(n_10562),
.B2(n_10552),
.C(n_10555),
.Y(n_10653)
);

NAND2xp5_ASAP7_75t_SL g10654 ( 
.A(n_10535),
.B(n_1027),
.Y(n_10654)
);

XNOR2xp5_ASAP7_75t_L g10655 ( 
.A(n_10478),
.B(n_1030),
.Y(n_10655)
);

NAND2xp5_ASAP7_75t_L g10656 ( 
.A(n_10571),
.B(n_1031),
.Y(n_10656)
);

INVx1_ASAP7_75t_L g10657 ( 
.A(n_10508),
.Y(n_10657)
);

AOI22xp5_ASAP7_75t_L g10658 ( 
.A1(n_10572),
.A2(n_1033),
.B1(n_1031),
.B2(n_1032),
.Y(n_10658)
);

NAND2xp5_ASAP7_75t_L g10659 ( 
.A(n_10568),
.B(n_10537),
.Y(n_10659)
);

INVx1_ASAP7_75t_L g10660 ( 
.A(n_10515),
.Y(n_10660)
);

OR2x2_ASAP7_75t_L g10661 ( 
.A(n_10517),
.B(n_1031),
.Y(n_10661)
);

XNOR2x2_ASAP7_75t_L g10662 ( 
.A(n_10569),
.B(n_1032),
.Y(n_10662)
);

OAI22xp33_ASAP7_75t_L g10663 ( 
.A1(n_10538),
.A2(n_1035),
.B1(n_1033),
.B2(n_1034),
.Y(n_10663)
);

INVx1_ASAP7_75t_L g10664 ( 
.A(n_10548),
.Y(n_10664)
);

AOI21xp5_ASAP7_75t_L g10665 ( 
.A1(n_10575),
.A2(n_1034),
.B(n_1035),
.Y(n_10665)
);

OR2x2_ASAP7_75t_L g10666 ( 
.A(n_10550),
.B(n_1034),
.Y(n_10666)
);

INVx1_ASAP7_75t_L g10667 ( 
.A(n_10556),
.Y(n_10667)
);

INVx1_ASAP7_75t_L g10668 ( 
.A(n_10560),
.Y(n_10668)
);

AOI22xp33_ASAP7_75t_L g10669 ( 
.A1(n_10547),
.A2(n_1037),
.B1(n_1035),
.B2(n_1036),
.Y(n_10669)
);

AOI322xp5_ASAP7_75t_L g10670 ( 
.A1(n_10557),
.A2(n_1041),
.A3(n_1040),
.B1(n_1038),
.B2(n_1036),
.C1(n_1037),
.C2(n_1039),
.Y(n_10670)
);

AOI21xp33_ASAP7_75t_SL g10671 ( 
.A1(n_10542),
.A2(n_10474),
.B(n_10574),
.Y(n_10671)
);

OAI211xp5_ASAP7_75t_SL g10672 ( 
.A1(n_10563),
.A2(n_1041),
.B(n_1039),
.C(n_1040),
.Y(n_10672)
);

OAI21xp33_ASAP7_75t_L g10673 ( 
.A1(n_10561),
.A2(n_10573),
.B(n_10554),
.Y(n_10673)
);

NOR2xp33_ASAP7_75t_L g10674 ( 
.A(n_10570),
.B(n_1039),
.Y(n_10674)
);

OAI21xp33_ASAP7_75t_L g10675 ( 
.A1(n_10567),
.A2(n_10559),
.B(n_10492),
.Y(n_10675)
);

OAI32xp33_ASAP7_75t_L g10676 ( 
.A1(n_10576),
.A2(n_1042),
.A3(n_1040),
.B1(n_1041),
.B2(n_1043),
.Y(n_10676)
);

INVx1_ASAP7_75t_L g10677 ( 
.A(n_10494),
.Y(n_10677)
);

AOI221xp5_ASAP7_75t_L g10678 ( 
.A1(n_10471),
.A2(n_1044),
.B1(n_1042),
.B2(n_1043),
.C(n_1045),
.Y(n_10678)
);

INVx1_ASAP7_75t_L g10679 ( 
.A(n_10494),
.Y(n_10679)
);

INVx1_ASAP7_75t_L g10680 ( 
.A(n_10494),
.Y(n_10680)
);

NAND2xp5_ASAP7_75t_L g10681 ( 
.A(n_10577),
.B(n_1042),
.Y(n_10681)
);

INVx2_ASAP7_75t_SL g10682 ( 
.A(n_10565),
.Y(n_10682)
);

INVx1_ASAP7_75t_L g10683 ( 
.A(n_10494),
.Y(n_10683)
);

OAI21xp5_ASAP7_75t_L g10684 ( 
.A1(n_10471),
.A2(n_1043),
.B(n_1044),
.Y(n_10684)
);

AOI21xp5_ASAP7_75t_L g10685 ( 
.A1(n_10471),
.A2(n_1044),
.B(n_1045),
.Y(n_10685)
);

INVx1_ASAP7_75t_L g10686 ( 
.A(n_10494),
.Y(n_10686)
);

AOI21xp33_ASAP7_75t_L g10687 ( 
.A1(n_10473),
.A2(n_1046),
.B(n_1657),
.Y(n_10687)
);

AOI211xp5_ASAP7_75t_L g10688 ( 
.A1(n_10471),
.A2(n_1046),
.B(n_1659),
.C(n_1657),
.Y(n_10688)
);

OAI21xp33_ASAP7_75t_SL g10689 ( 
.A1(n_10471),
.A2(n_1660),
.B(n_1661),
.Y(n_10689)
);

INVx1_ASAP7_75t_L g10690 ( 
.A(n_10494),
.Y(n_10690)
);

NAND2xp5_ASAP7_75t_L g10691 ( 
.A(n_10577),
.B(n_1661),
.Y(n_10691)
);

NAND2xp5_ASAP7_75t_L g10692 ( 
.A(n_10577),
.B(n_1662),
.Y(n_10692)
);

AOI21xp33_ASAP7_75t_L g10693 ( 
.A1(n_10473),
.A2(n_1665),
.B(n_1664),
.Y(n_10693)
);

AOI22xp5_ASAP7_75t_L g10694 ( 
.A1(n_10520),
.A2(n_1665),
.B1(n_1663),
.B2(n_1664),
.Y(n_10694)
);

INVx1_ASAP7_75t_L g10695 ( 
.A(n_10494),
.Y(n_10695)
);

OAI221xp5_ASAP7_75t_L g10696 ( 
.A1(n_10471),
.A2(n_1667),
.B1(n_1663),
.B2(n_1666),
.C(n_1668),
.Y(n_10696)
);

INVx2_ASAP7_75t_L g10697 ( 
.A(n_10545),
.Y(n_10697)
);

INVx2_ASAP7_75t_L g10698 ( 
.A(n_10545),
.Y(n_10698)
);

OR2x2_ASAP7_75t_L g10699 ( 
.A(n_10477),
.B(n_1667),
.Y(n_10699)
);

INVx1_ASAP7_75t_L g10700 ( 
.A(n_10494),
.Y(n_10700)
);

INVx1_ASAP7_75t_SL g10701 ( 
.A(n_10529),
.Y(n_10701)
);

OR2x2_ASAP7_75t_L g10702 ( 
.A(n_10477),
.B(n_1668),
.Y(n_10702)
);

INVx1_ASAP7_75t_L g10703 ( 
.A(n_10494),
.Y(n_10703)
);

OAI22xp33_ASAP7_75t_L g10704 ( 
.A1(n_10576),
.A2(n_1672),
.B1(n_1669),
.B2(n_1671),
.Y(n_10704)
);

INVx1_ASAP7_75t_L g10705 ( 
.A(n_10494),
.Y(n_10705)
);

INVx1_ASAP7_75t_L g10706 ( 
.A(n_10494),
.Y(n_10706)
);

AND2x2_ASAP7_75t_L g10707 ( 
.A(n_10529),
.B(n_1669),
.Y(n_10707)
);

NAND2xp5_ASAP7_75t_L g10708 ( 
.A(n_10577),
.B(n_1671),
.Y(n_10708)
);

OAI22xp5_ASAP7_75t_L g10709 ( 
.A1(n_10576),
.A2(n_1674),
.B1(n_1672),
.B2(n_1673),
.Y(n_10709)
);

NAND3xp33_ASAP7_75t_L g10710 ( 
.A(n_10473),
.B(n_2254),
.C(n_2253),
.Y(n_10710)
);

INVxp67_ASAP7_75t_L g10711 ( 
.A(n_10494),
.Y(n_10711)
);

AND2x2_ASAP7_75t_L g10712 ( 
.A(n_10529),
.B(n_1673),
.Y(n_10712)
);

AOI22xp33_ASAP7_75t_L g10713 ( 
.A1(n_10471),
.A2(n_1676),
.B1(n_1674),
.B2(n_1675),
.Y(n_10713)
);

AOI221xp5_ASAP7_75t_L g10714 ( 
.A1(n_10592),
.A2(n_1677),
.B1(n_1675),
.B2(n_1676),
.C(n_1678),
.Y(n_10714)
);

NAND2xp5_ASAP7_75t_L g10715 ( 
.A(n_10701),
.B(n_10621),
.Y(n_10715)
);

NAND2xp5_ASAP7_75t_L g10716 ( 
.A(n_10582),
.B(n_1679),
.Y(n_10716)
);

NAND2xp5_ASAP7_75t_L g10717 ( 
.A(n_10707),
.B(n_1681),
.Y(n_10717)
);

NOR2x1_ASAP7_75t_L g10718 ( 
.A(n_10586),
.B(n_1681),
.Y(n_10718)
);

AOI21xp33_ASAP7_75t_SL g10719 ( 
.A1(n_10704),
.A2(n_1682),
.B(n_1683),
.Y(n_10719)
);

HB1xp67_ASAP7_75t_L g10720 ( 
.A(n_10595),
.Y(n_10720)
);

OAI22xp33_ASAP7_75t_L g10721 ( 
.A1(n_10599),
.A2(n_1685),
.B1(n_1686),
.B2(n_1684),
.Y(n_10721)
);

NAND2xp5_ASAP7_75t_L g10722 ( 
.A(n_10712),
.B(n_1683),
.Y(n_10722)
);

INVx1_ASAP7_75t_L g10723 ( 
.A(n_10609),
.Y(n_10723)
);

INVx1_ASAP7_75t_L g10724 ( 
.A(n_10607),
.Y(n_10724)
);

INVxp67_ASAP7_75t_L g10725 ( 
.A(n_10594),
.Y(n_10725)
);

INVx2_ASAP7_75t_L g10726 ( 
.A(n_10613),
.Y(n_10726)
);

AOI21xp5_ASAP7_75t_L g10727 ( 
.A1(n_10632),
.A2(n_1685),
.B(n_1686),
.Y(n_10727)
);

NAND2xp5_ASAP7_75t_L g10728 ( 
.A(n_10629),
.B(n_1687),
.Y(n_10728)
);

NAND3xp33_ASAP7_75t_SL g10729 ( 
.A(n_10688),
.B(n_1687),
.C(n_1688),
.Y(n_10729)
);

INVx1_ASAP7_75t_L g10730 ( 
.A(n_10655),
.Y(n_10730)
);

OR2x2_ASAP7_75t_L g10731 ( 
.A(n_10682),
.B(n_1688),
.Y(n_10731)
);

OAI221xp5_ASAP7_75t_SL g10732 ( 
.A1(n_10711),
.A2(n_1691),
.B1(n_1689),
.B2(n_1690),
.C(n_1692),
.Y(n_10732)
);

INVx1_ASAP7_75t_L g10733 ( 
.A(n_10581),
.Y(n_10733)
);

OAI211xp5_ASAP7_75t_L g10734 ( 
.A1(n_10689),
.A2(n_1699),
.B(n_1707),
.C(n_1689),
.Y(n_10734)
);

NOR3xp33_ASAP7_75t_L g10735 ( 
.A(n_10587),
.B(n_1692),
.C(n_1693),
.Y(n_10735)
);

INVx1_ASAP7_75t_L g10736 ( 
.A(n_10681),
.Y(n_10736)
);

NAND2xp5_ASAP7_75t_L g10737 ( 
.A(n_10597),
.B(n_1693),
.Y(n_10737)
);

INVxp67_ASAP7_75t_L g10738 ( 
.A(n_10691),
.Y(n_10738)
);

NOR2x1_ASAP7_75t_SL g10739 ( 
.A(n_10697),
.B(n_1694),
.Y(n_10739)
);

NAND5xp2_ASAP7_75t_L g10740 ( 
.A(n_10653),
.B(n_1710),
.C(n_1718),
.D(n_1702),
.E(n_1694),
.Y(n_10740)
);

AND2x2_ASAP7_75t_L g10741 ( 
.A(n_10604),
.B(n_1695),
.Y(n_10741)
);

AND2x2_ASAP7_75t_L g10742 ( 
.A(n_10677),
.B(n_10679),
.Y(n_10742)
);

OR2x2_ASAP7_75t_L g10743 ( 
.A(n_10590),
.B(n_10585),
.Y(n_10743)
);

NAND2xp5_ASAP7_75t_L g10744 ( 
.A(n_10619),
.B(n_1695),
.Y(n_10744)
);

NAND4xp25_ASAP7_75t_L g10745 ( 
.A(n_10589),
.B(n_1698),
.C(n_1696),
.D(n_1697),
.Y(n_10745)
);

INVx1_ASAP7_75t_SL g10746 ( 
.A(n_10692),
.Y(n_10746)
);

NAND2xp5_ASAP7_75t_L g10747 ( 
.A(n_10584),
.B(n_10615),
.Y(n_10747)
);

INVx1_ASAP7_75t_L g10748 ( 
.A(n_10708),
.Y(n_10748)
);

NAND2xp5_ASAP7_75t_L g10749 ( 
.A(n_10680),
.B(n_1696),
.Y(n_10749)
);

AOI222xp33_ASAP7_75t_L g10750 ( 
.A1(n_10583),
.A2(n_1700),
.B1(n_1702),
.B2(n_1698),
.C1(n_1699),
.C2(n_1701),
.Y(n_10750)
);

AOI22xp33_ASAP7_75t_SL g10751 ( 
.A1(n_10698),
.A2(n_1704),
.B1(n_1700),
.B2(n_1703),
.Y(n_10751)
);

AND2x2_ASAP7_75t_L g10752 ( 
.A(n_10683),
.B(n_1703),
.Y(n_10752)
);

INVx1_ASAP7_75t_L g10753 ( 
.A(n_10628),
.Y(n_10753)
);

AND2x2_ASAP7_75t_L g10754 ( 
.A(n_10686),
.B(n_1704),
.Y(n_10754)
);

AND2x2_ASAP7_75t_L g10755 ( 
.A(n_10690),
.B(n_1705),
.Y(n_10755)
);

INVx1_ASAP7_75t_L g10756 ( 
.A(n_10631),
.Y(n_10756)
);

AOI211x1_ASAP7_75t_L g10757 ( 
.A1(n_10684),
.A2(n_1707),
.B(n_1705),
.C(n_1706),
.Y(n_10757)
);

INVx1_ASAP7_75t_L g10758 ( 
.A(n_10626),
.Y(n_10758)
);

AND2x2_ASAP7_75t_L g10759 ( 
.A(n_10695),
.B(n_1708),
.Y(n_10759)
);

AND2x2_ASAP7_75t_L g10760 ( 
.A(n_10700),
.B(n_1708),
.Y(n_10760)
);

NAND2xp5_ASAP7_75t_L g10761 ( 
.A(n_10703),
.B(n_1709),
.Y(n_10761)
);

BUFx12f_ASAP7_75t_L g10762 ( 
.A(n_10634),
.Y(n_10762)
);

INVx1_ASAP7_75t_L g10763 ( 
.A(n_10699),
.Y(n_10763)
);

INVx1_ASAP7_75t_L g10764 ( 
.A(n_10702),
.Y(n_10764)
);

INVx1_ASAP7_75t_L g10765 ( 
.A(n_10705),
.Y(n_10765)
);

AND2x2_ASAP7_75t_L g10766 ( 
.A(n_10706),
.B(n_1709),
.Y(n_10766)
);

NAND2xp5_ASAP7_75t_L g10767 ( 
.A(n_10620),
.B(n_1710),
.Y(n_10767)
);

INVx1_ASAP7_75t_L g10768 ( 
.A(n_10601),
.Y(n_10768)
);

AOI21xp5_ASAP7_75t_SL g10769 ( 
.A1(n_10593),
.A2(n_1711),
.B(n_1712),
.Y(n_10769)
);

NOR2xp67_ASAP7_75t_L g10770 ( 
.A(n_10646),
.B(n_2260),
.Y(n_10770)
);

INVx1_ASAP7_75t_L g10771 ( 
.A(n_10640),
.Y(n_10771)
);

AND2x2_ASAP7_75t_L g10772 ( 
.A(n_10606),
.B(n_10634),
.Y(n_10772)
);

NAND2xp33_ASAP7_75t_R g10773 ( 
.A(n_10660),
.B(n_1711),
.Y(n_10773)
);

INVx1_ASAP7_75t_L g10774 ( 
.A(n_10617),
.Y(n_10774)
);

XOR2x2_ASAP7_75t_L g10775 ( 
.A(n_10662),
.B(n_10709),
.Y(n_10775)
);

NAND2xp5_ASAP7_75t_L g10776 ( 
.A(n_10614),
.B(n_1712),
.Y(n_10776)
);

INVx1_ASAP7_75t_SL g10777 ( 
.A(n_10622),
.Y(n_10777)
);

NAND3xp33_ASAP7_75t_SL g10778 ( 
.A(n_10678),
.B(n_1713),
.C(n_1714),
.Y(n_10778)
);

NOR2xp33_ASAP7_75t_L g10779 ( 
.A(n_10676),
.B(n_1713),
.Y(n_10779)
);

OAI21xp5_ASAP7_75t_SL g10780 ( 
.A1(n_10713),
.A2(n_2263),
.B(n_1714),
.Y(n_10780)
);

AND2x2_ASAP7_75t_L g10781 ( 
.A(n_10633),
.B(n_1715),
.Y(n_10781)
);

INVx1_ASAP7_75t_L g10782 ( 
.A(n_10603),
.Y(n_10782)
);

NOR4xp25_ASAP7_75t_L g10783 ( 
.A(n_10675),
.B(n_10673),
.C(n_10654),
.D(n_10696),
.Y(n_10783)
);

NAND2xp5_ASAP7_75t_L g10784 ( 
.A(n_10670),
.B(n_1715),
.Y(n_10784)
);

INVx1_ASAP7_75t_L g10785 ( 
.A(n_10656),
.Y(n_10785)
);

OAI22xp33_ASAP7_75t_L g10786 ( 
.A1(n_10625),
.A2(n_1719),
.B1(n_1720),
.B2(n_1717),
.Y(n_10786)
);

HB1xp67_ASAP7_75t_L g10787 ( 
.A(n_10588),
.Y(n_10787)
);

INVx2_ASAP7_75t_L g10788 ( 
.A(n_10661),
.Y(n_10788)
);

INVx1_ASAP7_75t_L g10789 ( 
.A(n_10659),
.Y(n_10789)
);

INVx1_ASAP7_75t_L g10790 ( 
.A(n_10611),
.Y(n_10790)
);

INVx1_ASAP7_75t_L g10791 ( 
.A(n_10636),
.Y(n_10791)
);

NAND2xp5_ASAP7_75t_L g10792 ( 
.A(n_10637),
.B(n_10641),
.Y(n_10792)
);

NOR2xp33_ASAP7_75t_L g10793 ( 
.A(n_10672),
.B(n_1716),
.Y(n_10793)
);

AND2x2_ASAP7_75t_L g10794 ( 
.A(n_10639),
.B(n_1717),
.Y(n_10794)
);

OR2x6_ASAP7_75t_L g10795 ( 
.A(n_10618),
.B(n_1719),
.Y(n_10795)
);

INVx1_ASAP7_75t_L g10796 ( 
.A(n_10616),
.Y(n_10796)
);

XNOR2x2_ASAP7_75t_L g10797 ( 
.A(n_10605),
.B(n_1720),
.Y(n_10797)
);

NAND2xp5_ASAP7_75t_L g10798 ( 
.A(n_10627),
.B(n_1721),
.Y(n_10798)
);

OA211x2_ASAP7_75t_L g10799 ( 
.A1(n_10610),
.A2(n_1723),
.B(n_1721),
.C(n_1722),
.Y(n_10799)
);

INVxp67_ASAP7_75t_L g10800 ( 
.A(n_10600),
.Y(n_10800)
);

INVx2_ASAP7_75t_L g10801 ( 
.A(n_10630),
.Y(n_10801)
);

NAND2xp5_ASAP7_75t_L g10802 ( 
.A(n_10669),
.B(n_1722),
.Y(n_10802)
);

AND2x2_ASAP7_75t_L g10803 ( 
.A(n_10638),
.B(n_1723),
.Y(n_10803)
);

NAND2xp5_ASAP7_75t_SL g10804 ( 
.A(n_10663),
.B(n_1724),
.Y(n_10804)
);

NAND2xp5_ASAP7_75t_L g10805 ( 
.A(n_10665),
.B(n_1725),
.Y(n_10805)
);

INVx1_ASAP7_75t_L g10806 ( 
.A(n_10645),
.Y(n_10806)
);

INVx1_ASAP7_75t_L g10807 ( 
.A(n_10666),
.Y(n_10807)
);

NAND2x1p5_ASAP7_75t_L g10808 ( 
.A(n_10657),
.B(n_1727),
.Y(n_10808)
);

NAND2xp5_ASAP7_75t_L g10809 ( 
.A(n_10598),
.B(n_1726),
.Y(n_10809)
);

OAI21xp5_ASAP7_75t_SL g10810 ( 
.A1(n_10608),
.A2(n_2258),
.B(n_2257),
.Y(n_10810)
);

INVx2_ASAP7_75t_L g10811 ( 
.A(n_10612),
.Y(n_10811)
);

INVx1_ASAP7_75t_L g10812 ( 
.A(n_10602),
.Y(n_10812)
);

NAND4xp25_ASAP7_75t_L g10813 ( 
.A(n_10647),
.B(n_10685),
.C(n_10671),
.D(n_10652),
.Y(n_10813)
);

INVx1_ASAP7_75t_L g10814 ( 
.A(n_10623),
.Y(n_10814)
);

INVx1_ASAP7_75t_L g10815 ( 
.A(n_10635),
.Y(n_10815)
);

NAND2xp5_ASAP7_75t_L g10816 ( 
.A(n_10694),
.B(n_1726),
.Y(n_10816)
);

NAND2xp5_ASAP7_75t_SL g10817 ( 
.A(n_10596),
.B(n_1727),
.Y(n_10817)
);

INVx1_ASAP7_75t_L g10818 ( 
.A(n_10658),
.Y(n_10818)
);

OAI21xp33_ASAP7_75t_SL g10819 ( 
.A1(n_10643),
.A2(n_1728),
.B(n_1729),
.Y(n_10819)
);

INVx2_ASAP7_75t_L g10820 ( 
.A(n_10649),
.Y(n_10820)
);

NAND2xp5_ASAP7_75t_L g10821 ( 
.A(n_10642),
.B(n_1730),
.Y(n_10821)
);

INVx1_ASAP7_75t_L g10822 ( 
.A(n_10710),
.Y(n_10822)
);

INVx1_ASAP7_75t_L g10823 ( 
.A(n_10674),
.Y(n_10823)
);

INVx1_ASAP7_75t_L g10824 ( 
.A(n_10651),
.Y(n_10824)
);

HB1xp67_ASAP7_75t_L g10825 ( 
.A(n_10591),
.Y(n_10825)
);

AND3x1_ASAP7_75t_L g10826 ( 
.A(n_10648),
.B(n_1740),
.C(n_1730),
.Y(n_10826)
);

NAND2xp5_ASAP7_75t_L g10827 ( 
.A(n_10650),
.B(n_1731),
.Y(n_10827)
);

XNOR2xp5_ASAP7_75t_L g10828 ( 
.A(n_10644),
.B(n_1731),
.Y(n_10828)
);

INVx1_ASAP7_75t_L g10829 ( 
.A(n_10664),
.Y(n_10829)
);

NAND3xp33_ASAP7_75t_L g10830 ( 
.A(n_10687),
.B(n_1732),
.C(n_1735),
.Y(n_10830)
);

NAND2xp5_ASAP7_75t_L g10831 ( 
.A(n_10667),
.B(n_10668),
.Y(n_10831)
);

NAND2xp5_ASAP7_75t_L g10832 ( 
.A(n_10624),
.B(n_1736),
.Y(n_10832)
);

INVxp67_ASAP7_75t_L g10833 ( 
.A(n_10693),
.Y(n_10833)
);

INVx1_ASAP7_75t_L g10834 ( 
.A(n_10582),
.Y(n_10834)
);

XOR2xp5_ASAP7_75t_L g10835 ( 
.A(n_10775),
.B(n_1736),
.Y(n_10835)
);

NAND2xp5_ASAP7_75t_L g10836 ( 
.A(n_10770),
.B(n_1737),
.Y(n_10836)
);

XNOR2xp5_ASAP7_75t_L g10837 ( 
.A(n_10826),
.B(n_1738),
.Y(n_10837)
);

AND2x2_ASAP7_75t_L g10838 ( 
.A(n_10772),
.B(n_1738),
.Y(n_10838)
);

INVx1_ASAP7_75t_L g10839 ( 
.A(n_10720),
.Y(n_10839)
);

INVx2_ASAP7_75t_L g10840 ( 
.A(n_10739),
.Y(n_10840)
);

OAI22xp33_ASAP7_75t_L g10841 ( 
.A1(n_10795),
.A2(n_1741),
.B1(n_1739),
.B2(n_1740),
.Y(n_10841)
);

OAI21xp5_ASAP7_75t_L g10842 ( 
.A1(n_10715),
.A2(n_1743),
.B(n_1742),
.Y(n_10842)
);

NOR2xp33_ASAP7_75t_L g10843 ( 
.A(n_10762),
.B(n_1739),
.Y(n_10843)
);

AND2x2_ASAP7_75t_L g10844 ( 
.A(n_10726),
.B(n_1744),
.Y(n_10844)
);

NAND2xp5_ASAP7_75t_L g10845 ( 
.A(n_10834),
.B(n_1744),
.Y(n_10845)
);

NAND2xp5_ASAP7_75t_SL g10846 ( 
.A(n_10819),
.B(n_1745),
.Y(n_10846)
);

OAI21xp5_ASAP7_75t_SL g10847 ( 
.A1(n_10723),
.A2(n_1745),
.B(n_1746),
.Y(n_10847)
);

INVx1_ASAP7_75t_L g10848 ( 
.A(n_10731),
.Y(n_10848)
);

AOI21xp5_ASAP7_75t_L g10849 ( 
.A1(n_10727),
.A2(n_1746),
.B(n_1747),
.Y(n_10849)
);

AND2x2_ASAP7_75t_L g10850 ( 
.A(n_10741),
.B(n_1747),
.Y(n_10850)
);

OR2x2_ASAP7_75t_L g10851 ( 
.A(n_10795),
.B(n_1748),
.Y(n_10851)
);

INVx1_ASAP7_75t_L g10852 ( 
.A(n_10742),
.Y(n_10852)
);

AOI322xp5_ASAP7_75t_L g10853 ( 
.A1(n_10824),
.A2(n_1754),
.A3(n_1753),
.B1(n_1750),
.B2(n_1748),
.C1(n_1749),
.C2(n_1752),
.Y(n_10853)
);

INVx1_ASAP7_75t_L g10854 ( 
.A(n_10787),
.Y(n_10854)
);

INVx1_ASAP7_75t_L g10855 ( 
.A(n_10808),
.Y(n_10855)
);

INVx2_ASAP7_75t_L g10856 ( 
.A(n_10752),
.Y(n_10856)
);

OAI22xp33_ASAP7_75t_L g10857 ( 
.A1(n_10728),
.A2(n_1755),
.B1(n_1752),
.B2(n_1753),
.Y(n_10857)
);

NOR2xp33_ASAP7_75t_L g10858 ( 
.A(n_10740),
.B(n_1755),
.Y(n_10858)
);

AOI22xp33_ASAP7_75t_L g10859 ( 
.A1(n_10765),
.A2(n_10774),
.B1(n_10790),
.B2(n_10811),
.Y(n_10859)
);

XNOR2xp5_ASAP7_75t_L g10860 ( 
.A(n_10828),
.B(n_1756),
.Y(n_10860)
);

OAI31xp33_ASAP7_75t_L g10861 ( 
.A1(n_10734),
.A2(n_1759),
.A3(n_1757),
.B(n_1758),
.Y(n_10861)
);

INVx1_ASAP7_75t_L g10862 ( 
.A(n_10754),
.Y(n_10862)
);

AND2x2_ASAP7_75t_L g10863 ( 
.A(n_10724),
.B(n_1757),
.Y(n_10863)
);

INVx1_ASAP7_75t_L g10864 ( 
.A(n_10755),
.Y(n_10864)
);

NAND2xp5_ASAP7_75t_L g10865 ( 
.A(n_10759),
.B(n_1759),
.Y(n_10865)
);

OAI22xp5_ASAP7_75t_L g10866 ( 
.A1(n_10725),
.A2(n_1762),
.B1(n_1760),
.B2(n_1761),
.Y(n_10866)
);

INVx2_ASAP7_75t_L g10867 ( 
.A(n_10760),
.Y(n_10867)
);

AOI21xp33_ASAP7_75t_SL g10868 ( 
.A1(n_10773),
.A2(n_1761),
.B(n_1763),
.Y(n_10868)
);

INVx2_ASAP7_75t_L g10869 ( 
.A(n_10766),
.Y(n_10869)
);

AOI21xp33_ASAP7_75t_SL g10870 ( 
.A1(n_10737),
.A2(n_1763),
.B(n_1764),
.Y(n_10870)
);

INVx1_ASAP7_75t_L g10871 ( 
.A(n_10716),
.Y(n_10871)
);

INVx1_ASAP7_75t_L g10872 ( 
.A(n_10717),
.Y(n_10872)
);

INVx1_ASAP7_75t_L g10873 ( 
.A(n_10722),
.Y(n_10873)
);

NAND2xp5_ASAP7_75t_L g10874 ( 
.A(n_10751),
.B(n_1765),
.Y(n_10874)
);

INVxp67_ASAP7_75t_L g10875 ( 
.A(n_10779),
.Y(n_10875)
);

OAI222xp33_ASAP7_75t_L g10876 ( 
.A1(n_10718),
.A2(n_1767),
.B1(n_1769),
.B2(n_1765),
.C1(n_1766),
.C2(n_1768),
.Y(n_10876)
);

INVx1_ASAP7_75t_L g10877 ( 
.A(n_10803),
.Y(n_10877)
);

NAND2xp5_ASAP7_75t_L g10878 ( 
.A(n_10758),
.B(n_1766),
.Y(n_10878)
);

AOI21xp33_ASAP7_75t_L g10879 ( 
.A1(n_10743),
.A2(n_1768),
.B(n_1770),
.Y(n_10879)
);

AOI221x1_ASAP7_75t_L g10880 ( 
.A1(n_10813),
.A2(n_2260),
.B1(n_2251),
.B2(n_1772),
.C(n_1770),
.Y(n_10880)
);

INVx1_ASAP7_75t_L g10881 ( 
.A(n_10767),
.Y(n_10881)
);

NAND2xp5_ASAP7_75t_L g10882 ( 
.A(n_10781),
.B(n_1771),
.Y(n_10882)
);

OAI22x1_ASAP7_75t_L g10883 ( 
.A1(n_10753),
.A2(n_1776),
.B1(n_1773),
.B2(n_1775),
.Y(n_10883)
);

INVx2_ASAP7_75t_L g10884 ( 
.A(n_10794),
.Y(n_10884)
);

INVx3_ASAP7_75t_SL g10885 ( 
.A(n_10777),
.Y(n_10885)
);

HB1xp67_ASAP7_75t_L g10886 ( 
.A(n_10799),
.Y(n_10886)
);

INVx1_ASAP7_75t_L g10887 ( 
.A(n_10744),
.Y(n_10887)
);

INVx1_ASAP7_75t_L g10888 ( 
.A(n_10747),
.Y(n_10888)
);

NOR2xp33_ASAP7_75t_L g10889 ( 
.A(n_10745),
.B(n_1775),
.Y(n_10889)
);

NAND2xp5_ASAP7_75t_SL g10890 ( 
.A(n_10719),
.B(n_1776),
.Y(n_10890)
);

OR2x2_ASAP7_75t_L g10891 ( 
.A(n_10784),
.B(n_1777),
.Y(n_10891)
);

INVx1_ASAP7_75t_L g10892 ( 
.A(n_10749),
.Y(n_10892)
);

INVx2_ASAP7_75t_L g10893 ( 
.A(n_10733),
.Y(n_10893)
);

INVx2_ASAP7_75t_L g10894 ( 
.A(n_10736),
.Y(n_10894)
);

AOI221xp5_ASAP7_75t_L g10895 ( 
.A1(n_10783),
.A2(n_1780),
.B1(n_1777),
.B2(n_1778),
.C(n_1781),
.Y(n_10895)
);

AND2x2_ASAP7_75t_L g10896 ( 
.A(n_10746),
.B(n_1778),
.Y(n_10896)
);

AND2x2_ASAP7_75t_L g10897 ( 
.A(n_10748),
.B(n_1780),
.Y(n_10897)
);

OAI22xp5_ASAP7_75t_SL g10898 ( 
.A1(n_10757),
.A2(n_1783),
.B1(n_1781),
.B2(n_1782),
.Y(n_10898)
);

INVxp67_ASAP7_75t_L g10899 ( 
.A(n_10793),
.Y(n_10899)
);

A2O1A1Ixp33_ASAP7_75t_L g10900 ( 
.A1(n_10714),
.A2(n_1785),
.B(n_1782),
.C(n_1784),
.Y(n_10900)
);

OAI21xp5_ASAP7_75t_L g10901 ( 
.A1(n_10830),
.A2(n_1789),
.B(n_1787),
.Y(n_10901)
);

INVxp67_ASAP7_75t_L g10902 ( 
.A(n_10825),
.Y(n_10902)
);

OAI22xp5_ASAP7_75t_L g10903 ( 
.A1(n_10738),
.A2(n_1789),
.B1(n_1784),
.B2(n_1787),
.Y(n_10903)
);

OR2x2_ASAP7_75t_L g10904 ( 
.A(n_10761),
.B(n_1790),
.Y(n_10904)
);

AOI221x1_ASAP7_75t_SL g10905 ( 
.A1(n_10822),
.A2(n_1792),
.B1(n_1790),
.B2(n_1791),
.C(n_1793),
.Y(n_10905)
);

OAI21xp5_ASAP7_75t_L g10906 ( 
.A1(n_10833),
.A2(n_1793),
.B(n_1792),
.Y(n_10906)
);

NAND2xp5_ASAP7_75t_L g10907 ( 
.A(n_10721),
.B(n_1791),
.Y(n_10907)
);

INVx2_ASAP7_75t_SL g10908 ( 
.A(n_10756),
.Y(n_10908)
);

NAND4xp25_ASAP7_75t_SL g10909 ( 
.A(n_10792),
.B(n_1796),
.C(n_1794),
.D(n_1795),
.Y(n_10909)
);

NAND2xp5_ASAP7_75t_L g10910 ( 
.A(n_10735),
.B(n_1794),
.Y(n_10910)
);

AOI22xp33_ASAP7_75t_L g10911 ( 
.A1(n_10791),
.A2(n_1798),
.B1(n_1795),
.B2(n_1797),
.Y(n_10911)
);

INVx1_ASAP7_75t_L g10912 ( 
.A(n_10805),
.Y(n_10912)
);

XOR2xp5_ASAP7_75t_L g10913 ( 
.A(n_10730),
.B(n_10797),
.Y(n_10913)
);

OR2x2_ASAP7_75t_L g10914 ( 
.A(n_10776),
.B(n_10729),
.Y(n_10914)
);

INVx1_ASAP7_75t_L g10915 ( 
.A(n_10809),
.Y(n_10915)
);

OAI21xp5_ASAP7_75t_L g10916 ( 
.A1(n_10810),
.A2(n_1800),
.B(n_1799),
.Y(n_10916)
);

INVx1_ASAP7_75t_L g10917 ( 
.A(n_10798),
.Y(n_10917)
);

INVx1_ASAP7_75t_L g10918 ( 
.A(n_10832),
.Y(n_10918)
);

INVx1_ASAP7_75t_L g10919 ( 
.A(n_10816),
.Y(n_10919)
);

NAND3xp33_ASAP7_75t_L g10920 ( 
.A(n_10750),
.B(n_1798),
.C(n_1799),
.Y(n_10920)
);

INVx1_ASAP7_75t_L g10921 ( 
.A(n_10821),
.Y(n_10921)
);

NAND2xp5_ASAP7_75t_L g10922 ( 
.A(n_10763),
.B(n_1800),
.Y(n_10922)
);

NOR2xp67_ASAP7_75t_SL g10923 ( 
.A(n_10769),
.B(n_1801),
.Y(n_10923)
);

NAND2xp5_ASAP7_75t_L g10924 ( 
.A(n_10764),
.B(n_10815),
.Y(n_10924)
);

INVx1_ASAP7_75t_L g10925 ( 
.A(n_10802),
.Y(n_10925)
);

INVx1_ASAP7_75t_SL g10926 ( 
.A(n_10817),
.Y(n_10926)
);

INVx1_ASAP7_75t_L g10927 ( 
.A(n_10827),
.Y(n_10927)
);

INVx1_ASAP7_75t_SL g10928 ( 
.A(n_10804),
.Y(n_10928)
);

XNOR2xp5_ASAP7_75t_L g10929 ( 
.A(n_10812),
.B(n_1802),
.Y(n_10929)
);

XNOR2x1_ASAP7_75t_L g10930 ( 
.A(n_10814),
.B(n_10818),
.Y(n_10930)
);

O2A1O1Ixp33_ASAP7_75t_L g10931 ( 
.A1(n_10732),
.A2(n_1805),
.B(n_1803),
.C(n_1804),
.Y(n_10931)
);

AOI21xp33_ASAP7_75t_L g10932 ( 
.A1(n_10806),
.A2(n_1803),
.B(n_1806),
.Y(n_10932)
);

OAI21xp5_ASAP7_75t_SL g10933 ( 
.A1(n_10780),
.A2(n_1806),
.B(n_1807),
.Y(n_10933)
);

OAI22xp5_ASAP7_75t_L g10934 ( 
.A1(n_10789),
.A2(n_1810),
.B1(n_1807),
.B2(n_1808),
.Y(n_10934)
);

OAI221xp5_ASAP7_75t_L g10935 ( 
.A1(n_10800),
.A2(n_2255),
.B1(n_2256),
.B2(n_2254),
.C(n_2253),
.Y(n_10935)
);

AND2x2_ASAP7_75t_L g10936 ( 
.A(n_10788),
.B(n_1808),
.Y(n_10936)
);

OR2x2_ASAP7_75t_L g10937 ( 
.A(n_10778),
.B(n_1812),
.Y(n_10937)
);

AOI21xp5_ASAP7_75t_L g10938 ( 
.A1(n_10831),
.A2(n_10786),
.B(n_10807),
.Y(n_10938)
);

NAND2xp5_ASAP7_75t_L g10939 ( 
.A(n_10801),
.B(n_1812),
.Y(n_10939)
);

INVx1_ASAP7_75t_L g10940 ( 
.A(n_10796),
.Y(n_10940)
);

NAND2xp5_ASAP7_75t_L g10941 ( 
.A(n_10785),
.B(n_1814),
.Y(n_10941)
);

NAND3xp33_ASAP7_75t_L g10942 ( 
.A(n_10829),
.B(n_1815),
.C(n_1817),
.Y(n_10942)
);

INVxp67_ASAP7_75t_L g10943 ( 
.A(n_10823),
.Y(n_10943)
);

AOI22xp33_ASAP7_75t_L g10944 ( 
.A1(n_10820),
.A2(n_1819),
.B1(n_1815),
.B2(n_1818),
.Y(n_10944)
);

INVx1_ASAP7_75t_L g10945 ( 
.A(n_10835),
.Y(n_10945)
);

INVx1_ASAP7_75t_L g10946 ( 
.A(n_10838),
.Y(n_10946)
);

AOI22xp5_ASAP7_75t_L g10947 ( 
.A1(n_10858),
.A2(n_10771),
.B1(n_10782),
.B2(n_10768),
.Y(n_10947)
);

NAND3xp33_ASAP7_75t_L g10948 ( 
.A(n_10880),
.B(n_1818),
.C(n_1819),
.Y(n_10948)
);

CKINVDCx5p33_ASAP7_75t_R g10949 ( 
.A(n_10885),
.Y(n_10949)
);

XNOR2x1_ASAP7_75t_L g10950 ( 
.A(n_10930),
.B(n_1820),
.Y(n_10950)
);

NAND2xp5_ASAP7_75t_L g10951 ( 
.A(n_10905),
.B(n_1820),
.Y(n_10951)
);

AND2x2_ASAP7_75t_L g10952 ( 
.A(n_10839),
.B(n_1821),
.Y(n_10952)
);

NAND4xp25_ASAP7_75t_L g10953 ( 
.A(n_10859),
.B(n_10895),
.C(n_10888),
.D(n_10924),
.Y(n_10953)
);

INVx1_ASAP7_75t_L g10954 ( 
.A(n_10840),
.Y(n_10954)
);

XNOR2x2_ASAP7_75t_L g10955 ( 
.A(n_10837),
.B(n_1822),
.Y(n_10955)
);

INVx2_ASAP7_75t_L g10956 ( 
.A(n_10851),
.Y(n_10956)
);

AOI222xp33_ASAP7_75t_L g10957 ( 
.A1(n_10902),
.A2(n_1826),
.B1(n_1828),
.B2(n_1823),
.C1(n_1824),
.C2(n_1827),
.Y(n_10957)
);

NAND2xp5_ASAP7_75t_L g10958 ( 
.A(n_10853),
.B(n_1823),
.Y(n_10958)
);

OAI21xp5_ASAP7_75t_L g10959 ( 
.A1(n_10843),
.A2(n_1824),
.B(n_1826),
.Y(n_10959)
);

AOI22xp5_ASAP7_75t_L g10960 ( 
.A1(n_10852),
.A2(n_1829),
.B1(n_1827),
.B2(n_1828),
.Y(n_10960)
);

AND2x2_ASAP7_75t_L g10961 ( 
.A(n_10886),
.B(n_1829),
.Y(n_10961)
);

AOI221xp5_ASAP7_75t_L g10962 ( 
.A1(n_10868),
.A2(n_1834),
.B1(n_1830),
.B2(n_1831),
.C(n_1836),
.Y(n_10962)
);

INVx1_ASAP7_75t_L g10963 ( 
.A(n_10850),
.Y(n_10963)
);

INVx1_ASAP7_75t_L g10964 ( 
.A(n_10836),
.Y(n_10964)
);

OR2x2_ASAP7_75t_L g10965 ( 
.A(n_10846),
.B(n_1831),
.Y(n_10965)
);

AND2x2_ASAP7_75t_L g10966 ( 
.A(n_10856),
.B(n_1834),
.Y(n_10966)
);

XNOR2xp5_ASAP7_75t_L g10967 ( 
.A(n_10913),
.B(n_1836),
.Y(n_10967)
);

OAI21xp33_ASAP7_75t_SL g10968 ( 
.A1(n_10854),
.A2(n_1837),
.B(n_1838),
.Y(n_10968)
);

AO21x1_ASAP7_75t_L g10969 ( 
.A1(n_10841),
.A2(n_1839),
.B(n_1840),
.Y(n_10969)
);

OR2x2_ASAP7_75t_L g10970 ( 
.A(n_10874),
.B(n_1839),
.Y(n_10970)
);

NOR2x1_ASAP7_75t_L g10971 ( 
.A(n_10909),
.B(n_1840),
.Y(n_10971)
);

OAI211xp5_ASAP7_75t_L g10972 ( 
.A1(n_10861),
.A2(n_1843),
.B(n_1841),
.C(n_1842),
.Y(n_10972)
);

CKINVDCx5p33_ASAP7_75t_R g10973 ( 
.A(n_10860),
.Y(n_10973)
);

INVx1_ASAP7_75t_L g10974 ( 
.A(n_10929),
.Y(n_10974)
);

BUFx2_ASAP7_75t_L g10975 ( 
.A(n_10883),
.Y(n_10975)
);

INVx1_ASAP7_75t_L g10976 ( 
.A(n_10844),
.Y(n_10976)
);

NAND4xp25_ASAP7_75t_SL g10977 ( 
.A(n_10931),
.B(n_1844),
.C(n_1841),
.D(n_1843),
.Y(n_10977)
);

NAND2x1_ASAP7_75t_L g10978 ( 
.A(n_10923),
.B(n_1844),
.Y(n_10978)
);

A2O1A1Ixp33_ASAP7_75t_L g10979 ( 
.A1(n_10889),
.A2(n_1847),
.B(n_1845),
.C(n_1846),
.Y(n_10979)
);

XNOR2x1_ASAP7_75t_L g10980 ( 
.A(n_10891),
.B(n_1846),
.Y(n_10980)
);

INVx1_ASAP7_75t_L g10981 ( 
.A(n_10863),
.Y(n_10981)
);

INVx1_ASAP7_75t_L g10982 ( 
.A(n_10898),
.Y(n_10982)
);

NOR2x1_ASAP7_75t_L g10983 ( 
.A(n_10942),
.B(n_1848),
.Y(n_10983)
);

XNOR2xp5_ASAP7_75t_L g10984 ( 
.A(n_10928),
.B(n_1849),
.Y(n_10984)
);

NOR3xp33_ASAP7_75t_L g10985 ( 
.A(n_10908),
.B(n_1850),
.C(n_1851),
.Y(n_10985)
);

INVx1_ASAP7_75t_L g10986 ( 
.A(n_10896),
.Y(n_10986)
);

CKINVDCx14_ASAP7_75t_R g10987 ( 
.A(n_10914),
.Y(n_10987)
);

HB1xp67_ASAP7_75t_L g10988 ( 
.A(n_10855),
.Y(n_10988)
);

OR2x2_ASAP7_75t_L g10989 ( 
.A(n_10845),
.B(n_1850),
.Y(n_10989)
);

INVxp67_ASAP7_75t_SL g10990 ( 
.A(n_10882),
.Y(n_10990)
);

AOI21xp5_ASAP7_75t_L g10991 ( 
.A1(n_10890),
.A2(n_10938),
.B(n_10849),
.Y(n_10991)
);

NAND2xp5_ASAP7_75t_L g10992 ( 
.A(n_10897),
.B(n_10936),
.Y(n_10992)
);

CKINVDCx5p33_ASAP7_75t_R g10993 ( 
.A(n_10867),
.Y(n_10993)
);

INVx2_ASAP7_75t_L g10994 ( 
.A(n_10904),
.Y(n_10994)
);

OAI321xp33_ASAP7_75t_L g10995 ( 
.A1(n_10875),
.A2(n_1854),
.A3(n_1856),
.B1(n_1852),
.B2(n_1853),
.C(n_1855),
.Y(n_10995)
);

OAI31xp33_ASAP7_75t_L g10996 ( 
.A1(n_10876),
.A2(n_1862),
.A3(n_1871),
.B(n_1853),
.Y(n_10996)
);

INVx2_ASAP7_75t_L g10997 ( 
.A(n_10937),
.Y(n_10997)
);

AND2x2_ASAP7_75t_L g10998 ( 
.A(n_10869),
.B(n_1855),
.Y(n_10998)
);

AOI22xp5_ASAP7_75t_L g10999 ( 
.A1(n_10926),
.A2(n_1858),
.B1(n_1856),
.B2(n_1857),
.Y(n_10999)
);

INVx1_ASAP7_75t_L g11000 ( 
.A(n_10865),
.Y(n_11000)
);

INVxp67_ASAP7_75t_L g11001 ( 
.A(n_10878),
.Y(n_11001)
);

NAND2xp5_ASAP7_75t_SL g11002 ( 
.A(n_10870),
.B(n_1859),
.Y(n_11002)
);

A2O1A1Ixp33_ASAP7_75t_L g11003 ( 
.A1(n_10847),
.A2(n_1862),
.B(n_1860),
.C(n_1861),
.Y(n_11003)
);

INVx1_ASAP7_75t_L g11004 ( 
.A(n_10939),
.Y(n_11004)
);

XOR2x2_ASAP7_75t_L g11005 ( 
.A(n_10920),
.B(n_1860),
.Y(n_11005)
);

OR2x2_ASAP7_75t_L g11006 ( 
.A(n_10922),
.B(n_1861),
.Y(n_11006)
);

NAND2xp5_ASAP7_75t_L g11007 ( 
.A(n_10862),
.B(n_10864),
.Y(n_11007)
);

AOI22xp5_ASAP7_75t_L g11008 ( 
.A1(n_10943),
.A2(n_1865),
.B1(n_1863),
.B2(n_1864),
.Y(n_11008)
);

INVx1_ASAP7_75t_L g11009 ( 
.A(n_10907),
.Y(n_11009)
);

OAI22xp5_ASAP7_75t_L g11010 ( 
.A1(n_10899),
.A2(n_1865),
.B1(n_1863),
.B2(n_1864),
.Y(n_11010)
);

OAI211xp5_ASAP7_75t_L g11011 ( 
.A1(n_10933),
.A2(n_1868),
.B(n_1866),
.C(n_1867),
.Y(n_11011)
);

AOI211x1_ASAP7_75t_SL g11012 ( 
.A1(n_10893),
.A2(n_1870),
.B(n_1866),
.C(n_1867),
.Y(n_11012)
);

HB1xp67_ASAP7_75t_L g11013 ( 
.A(n_10848),
.Y(n_11013)
);

INVx1_ASAP7_75t_L g11014 ( 
.A(n_10877),
.Y(n_11014)
);

XOR2x2_ASAP7_75t_L g11015 ( 
.A(n_10916),
.B(n_10901),
.Y(n_11015)
);

INVx1_ASAP7_75t_L g11016 ( 
.A(n_10910),
.Y(n_11016)
);

OAI22xp5_ASAP7_75t_L g11017 ( 
.A1(n_10900),
.A2(n_1873),
.B1(n_1870),
.B2(n_1872),
.Y(n_11017)
);

XOR2x2_ASAP7_75t_L g11018 ( 
.A(n_10842),
.B(n_1873),
.Y(n_11018)
);

NAND2xp5_ASAP7_75t_SL g11019 ( 
.A(n_10857),
.B(n_1874),
.Y(n_11019)
);

AND2x2_ASAP7_75t_L g11020 ( 
.A(n_10884),
.B(n_1874),
.Y(n_11020)
);

AOI22xp33_ASAP7_75t_SL g11021 ( 
.A1(n_10940),
.A2(n_2261),
.B1(n_2249),
.B2(n_1877),
.Y(n_11021)
);

AOI211xp5_ASAP7_75t_L g11022 ( 
.A1(n_10879),
.A2(n_1877),
.B(n_1875),
.C(n_1876),
.Y(n_11022)
);

AOI22xp5_ASAP7_75t_L g11023 ( 
.A1(n_10881),
.A2(n_1880),
.B1(n_1876),
.B2(n_1878),
.Y(n_11023)
);

AOI211xp5_ASAP7_75t_SL g11024 ( 
.A1(n_10925),
.A2(n_1882),
.B(n_1880),
.C(n_1881),
.Y(n_11024)
);

NAND2xp5_ASAP7_75t_L g11025 ( 
.A(n_10944),
.B(n_1882),
.Y(n_11025)
);

INVx1_ASAP7_75t_L g11026 ( 
.A(n_10941),
.Y(n_11026)
);

INVx1_ASAP7_75t_L g11027 ( 
.A(n_10894),
.Y(n_11027)
);

INVx1_ASAP7_75t_L g11028 ( 
.A(n_10906),
.Y(n_11028)
);

OAI21xp33_ASAP7_75t_L g11029 ( 
.A1(n_10918),
.A2(n_2262),
.B(n_2257),
.Y(n_11029)
);

AOI21xp33_ASAP7_75t_L g11030 ( 
.A1(n_10915),
.A2(n_10912),
.B(n_10919),
.Y(n_11030)
);

AOI22xp33_ASAP7_75t_SL g11031 ( 
.A1(n_10871),
.A2(n_2263),
.B1(n_1885),
.B2(n_1883),
.Y(n_11031)
);

AND2x2_ASAP7_75t_L g11032 ( 
.A(n_10872),
.B(n_1883),
.Y(n_11032)
);

AOI311xp33_ASAP7_75t_L g11033 ( 
.A1(n_10892),
.A2(n_10927),
.A3(n_10873),
.B(n_10887),
.C(n_10921),
.Y(n_11033)
);

HB1xp67_ASAP7_75t_L g11034 ( 
.A(n_10903),
.Y(n_11034)
);

OAI22xp5_ASAP7_75t_L g11035 ( 
.A1(n_10911),
.A2(n_1887),
.B1(n_1884),
.B2(n_1886),
.Y(n_11035)
);

INVx1_ASAP7_75t_L g11036 ( 
.A(n_10934),
.Y(n_11036)
);

NAND3xp33_ASAP7_75t_L g11037 ( 
.A(n_10996),
.B(n_10932),
.C(n_10917),
.Y(n_11037)
);

NOR2x1_ASAP7_75t_L g11038 ( 
.A(n_10948),
.B(n_10866),
.Y(n_11038)
);

INVx2_ASAP7_75t_SL g11039 ( 
.A(n_10949),
.Y(n_11039)
);

OAI322xp33_ASAP7_75t_L g11040 ( 
.A1(n_10987),
.A2(n_10935),
.A3(n_1892),
.B1(n_1888),
.B2(n_1891),
.C1(n_1884),
.C2(n_1887),
.Y(n_11040)
);

NOR3xp33_ASAP7_75t_L g11041 ( 
.A(n_10953),
.B(n_1901),
.C(n_1888),
.Y(n_11041)
);

NOR2xp33_ASAP7_75t_L g11042 ( 
.A(n_10982),
.B(n_1889),
.Y(n_11042)
);

INVx1_ASAP7_75t_L g11043 ( 
.A(n_10961),
.Y(n_11043)
);

NOR2x1_ASAP7_75t_L g11044 ( 
.A(n_10978),
.B(n_1889),
.Y(n_11044)
);

NOR3xp33_ASAP7_75t_L g11045 ( 
.A(n_10954),
.B(n_1905),
.C(n_1892),
.Y(n_11045)
);

NAND3xp33_ASAP7_75t_L g11046 ( 
.A(n_10968),
.B(n_1895),
.C(n_1896),
.Y(n_11046)
);

NOR3x1_ASAP7_75t_L g11047 ( 
.A(n_10972),
.B(n_1895),
.C(n_1896),
.Y(n_11047)
);

NOR2x1_ASAP7_75t_SL g11048 ( 
.A(n_11011),
.B(n_1897),
.Y(n_11048)
);

OA211x2_ASAP7_75t_L g11049 ( 
.A1(n_10977),
.A2(n_1909),
.B(n_1917),
.C(n_1898),
.Y(n_11049)
);

NAND4xp75_ASAP7_75t_L g11050 ( 
.A(n_10983),
.B(n_1902),
.C(n_1898),
.D(n_1900),
.Y(n_11050)
);

AND4x1_ASAP7_75t_L g11051 ( 
.A(n_11033),
.B(n_11012),
.C(n_11024),
.D(n_10991),
.Y(n_11051)
);

NAND4xp25_ASAP7_75t_L g11052 ( 
.A(n_10947),
.B(n_1905),
.C(n_1902),
.D(n_1903),
.Y(n_11052)
);

NAND4xp75_ASAP7_75t_L g11053 ( 
.A(n_10969),
.B(n_1907),
.C(n_1903),
.D(n_1906),
.Y(n_11053)
);

AOI22x1_ASAP7_75t_L g11054 ( 
.A1(n_10975),
.A2(n_1908),
.B1(n_1906),
.B2(n_1907),
.Y(n_11054)
);

OA22x2_ASAP7_75t_L g11055 ( 
.A1(n_10967),
.A2(n_1912),
.B1(n_1910),
.B2(n_1911),
.Y(n_11055)
);

INVx1_ASAP7_75t_L g11056 ( 
.A(n_10984),
.Y(n_11056)
);

NOR4xp25_ASAP7_75t_L g11057 ( 
.A(n_11019),
.B(n_1913),
.C(n_1911),
.D(n_1912),
.Y(n_11057)
);

INVx1_ASAP7_75t_L g11058 ( 
.A(n_10952),
.Y(n_11058)
);

INVx1_ASAP7_75t_L g11059 ( 
.A(n_10988),
.Y(n_11059)
);

NOR3xp33_ASAP7_75t_L g11060 ( 
.A(n_11030),
.B(n_1921),
.C(n_1913),
.Y(n_11060)
);

NOR2xp33_ASAP7_75t_L g11061 ( 
.A(n_10946),
.B(n_11029),
.Y(n_11061)
);

AOI21xp5_ASAP7_75t_L g11062 ( 
.A1(n_11002),
.A2(n_11013),
.B(n_11007),
.Y(n_11062)
);

INVx1_ASAP7_75t_L g11063 ( 
.A(n_10966),
.Y(n_11063)
);

NOR2xp33_ASAP7_75t_L g11064 ( 
.A(n_10963),
.B(n_1914),
.Y(n_11064)
);

NAND3xp33_ASAP7_75t_L g11065 ( 
.A(n_11022),
.B(n_1914),
.C(n_1915),
.Y(n_11065)
);

AND2x4_ASAP7_75t_L g11066 ( 
.A(n_11020),
.B(n_1915),
.Y(n_11066)
);

NAND4xp25_ASAP7_75t_L g11067 ( 
.A(n_10945),
.B(n_1918),
.C(n_1916),
.D(n_1917),
.Y(n_11067)
);

AOI211xp5_ASAP7_75t_L g11068 ( 
.A1(n_11017),
.A2(n_1920),
.B(n_1918),
.C(n_1919),
.Y(n_11068)
);

OR2x2_ASAP7_75t_L g11069 ( 
.A(n_10951),
.B(n_1920),
.Y(n_11069)
);

NOR2x1_ASAP7_75t_L g11070 ( 
.A(n_10950),
.B(n_1921),
.Y(n_11070)
);

NOR3xp33_ASAP7_75t_SL g11071 ( 
.A(n_10993),
.B(n_1922),
.C(n_1923),
.Y(n_11071)
);

NAND2xp5_ASAP7_75t_L g11072 ( 
.A(n_11021),
.B(n_1924),
.Y(n_11072)
);

AOI22x1_ASAP7_75t_L g11073 ( 
.A1(n_10973),
.A2(n_11034),
.B1(n_10965),
.B2(n_10956),
.Y(n_11073)
);

NOR2xp33_ASAP7_75t_L g11074 ( 
.A(n_10981),
.B(n_1925),
.Y(n_11074)
);

NOR3xp33_ASAP7_75t_SL g11075 ( 
.A(n_10992),
.B(n_1926),
.C(n_1927),
.Y(n_11075)
);

NOR2x1_ASAP7_75t_L g11076 ( 
.A(n_10959),
.B(n_1926),
.Y(n_11076)
);

NOR3xp33_ASAP7_75t_L g11077 ( 
.A(n_11014),
.B(n_1937),
.C(n_1928),
.Y(n_11077)
);

AOI22xp5_ASAP7_75t_L g11078 ( 
.A1(n_10985),
.A2(n_1930),
.B1(n_1928),
.B2(n_1929),
.Y(n_11078)
);

NOR4xp25_ASAP7_75t_L g11079 ( 
.A(n_11027),
.B(n_11036),
.C(n_11028),
.D(n_10974),
.Y(n_11079)
);

AND2x2_ASAP7_75t_L g11080 ( 
.A(n_10971),
.B(n_1929),
.Y(n_11080)
);

NAND2xp5_ASAP7_75t_SL g11081 ( 
.A(n_10995),
.B(n_1930),
.Y(n_11081)
);

NAND2xp5_ASAP7_75t_L g11082 ( 
.A(n_10998),
.B(n_1931),
.Y(n_11082)
);

AOI22xp5_ASAP7_75t_L g11083 ( 
.A1(n_10986),
.A2(n_10976),
.B1(n_11035),
.B2(n_10997),
.Y(n_11083)
);

INVx1_ASAP7_75t_L g11084 ( 
.A(n_11032),
.Y(n_11084)
);

HB1xp67_ASAP7_75t_L g11085 ( 
.A(n_10955),
.Y(n_11085)
);

AOI22xp5_ASAP7_75t_L g11086 ( 
.A1(n_10990),
.A2(n_1933),
.B1(n_1931),
.B2(n_1932),
.Y(n_11086)
);

AND2x2_ASAP7_75t_L g11087 ( 
.A(n_10994),
.B(n_1932),
.Y(n_11087)
);

NAND2xp5_ASAP7_75t_L g11088 ( 
.A(n_11031),
.B(n_1933),
.Y(n_11088)
);

BUFx2_ASAP7_75t_L g11089 ( 
.A(n_10980),
.Y(n_11089)
);

INVx1_ASAP7_75t_L g11090 ( 
.A(n_10958),
.Y(n_11090)
);

AND2x4_ASAP7_75t_L g11091 ( 
.A(n_10964),
.B(n_1934),
.Y(n_11091)
);

NAND2xp5_ASAP7_75t_L g11092 ( 
.A(n_10957),
.B(n_1936),
.Y(n_11092)
);

OAI21xp33_ASAP7_75t_SL g11093 ( 
.A1(n_11009),
.A2(n_2249),
.B(n_2246),
.Y(n_11093)
);

INVx1_ASAP7_75t_L g11094 ( 
.A(n_10970),
.Y(n_11094)
);

AOI211xp5_ASAP7_75t_L g11095 ( 
.A1(n_10962),
.A2(n_1940),
.B(n_1938),
.C(n_1939),
.Y(n_11095)
);

AOI22xp5_ASAP7_75t_L g11096 ( 
.A1(n_11018),
.A2(n_1941),
.B1(n_1938),
.B2(n_1939),
.Y(n_11096)
);

HB1xp67_ASAP7_75t_L g11097 ( 
.A(n_11010),
.Y(n_11097)
);

NOR2x1_ASAP7_75t_L g11098 ( 
.A(n_11006),
.B(n_1943),
.Y(n_11098)
);

XNOR2xp5_ASAP7_75t_L g11099 ( 
.A(n_11015),
.B(n_11005),
.Y(n_11099)
);

NAND2xp5_ASAP7_75t_L g11100 ( 
.A(n_11003),
.B(n_1943),
.Y(n_11100)
);

NOR3xp33_ASAP7_75t_L g11101 ( 
.A(n_11001),
.B(n_1953),
.C(n_1944),
.Y(n_11101)
);

NOR2x1_ASAP7_75t_L g11102 ( 
.A(n_11044),
.B(n_10989),
.Y(n_11102)
);

AND2x2_ASAP7_75t_L g11103 ( 
.A(n_11059),
.B(n_11000),
.Y(n_11103)
);

NAND2x1p5_ASAP7_75t_L g11104 ( 
.A(n_11098),
.B(n_11004),
.Y(n_11104)
);

NAND4xp25_ASAP7_75t_SL g11105 ( 
.A(n_11041),
.B(n_11025),
.C(n_10979),
.D(n_11016),
.Y(n_11105)
);

AOI22xp5_ASAP7_75t_L g11106 ( 
.A1(n_11039),
.A2(n_11026),
.B1(n_10999),
.B2(n_11008),
.Y(n_11106)
);

AOI22xp5_ASAP7_75t_L g11107 ( 
.A1(n_11042),
.A2(n_10960),
.B1(n_11023),
.B2(n_1946),
.Y(n_11107)
);

BUFx3_ASAP7_75t_L g11108 ( 
.A(n_11043),
.Y(n_11108)
);

INVx1_ASAP7_75t_SL g11109 ( 
.A(n_11053),
.Y(n_11109)
);

INVx2_ASAP7_75t_L g11110 ( 
.A(n_11054),
.Y(n_11110)
);

INVx1_ASAP7_75t_L g11111 ( 
.A(n_11055),
.Y(n_11111)
);

NAND2xp33_ASAP7_75t_SL g11112 ( 
.A(n_11075),
.B(n_2248),
.Y(n_11112)
);

AOI22xp5_ASAP7_75t_L g11113 ( 
.A1(n_11061),
.A2(n_1946),
.B1(n_1944),
.B2(n_1945),
.Y(n_11113)
);

AOI22xp5_ASAP7_75t_L g11114 ( 
.A1(n_11038),
.A2(n_1949),
.B1(n_1945),
.B2(n_1947),
.Y(n_11114)
);

AOI22xp33_ASAP7_75t_L g11115 ( 
.A1(n_11085),
.A2(n_1950),
.B1(n_1951),
.B2(n_1949),
.Y(n_11115)
);

OAI211xp5_ASAP7_75t_L g11116 ( 
.A1(n_11093),
.A2(n_1951),
.B(n_1947),
.C(n_1950),
.Y(n_11116)
);

NAND4xp25_ASAP7_75t_L g11117 ( 
.A(n_11083),
.B(n_1955),
.C(n_1952),
.D(n_1954),
.Y(n_11117)
);

INVx2_ASAP7_75t_L g11118 ( 
.A(n_11091),
.Y(n_11118)
);

INVx2_ASAP7_75t_SL g11119 ( 
.A(n_11066),
.Y(n_11119)
);

AOI22xp5_ASAP7_75t_L g11120 ( 
.A1(n_11056),
.A2(n_1956),
.B1(n_1952),
.B2(n_1955),
.Y(n_11120)
);

BUFx2_ASAP7_75t_L g11121 ( 
.A(n_11066),
.Y(n_11121)
);

OAI22xp5_ASAP7_75t_SL g11122 ( 
.A1(n_11057),
.A2(n_1959),
.B1(n_1957),
.B2(n_1958),
.Y(n_11122)
);

AOI321xp33_ASAP7_75t_L g11123 ( 
.A1(n_11079),
.A2(n_1960),
.A3(n_1962),
.B1(n_1957),
.B2(n_1959),
.C(n_1961),
.Y(n_11123)
);

INVx3_ASAP7_75t_L g11124 ( 
.A(n_11091),
.Y(n_11124)
);

INVx1_ASAP7_75t_SL g11125 ( 
.A(n_11080),
.Y(n_11125)
);

AOI211xp5_ASAP7_75t_L g11126 ( 
.A1(n_11040),
.A2(n_11046),
.B(n_11060),
.C(n_11065),
.Y(n_11126)
);

INVx2_ASAP7_75t_L g11127 ( 
.A(n_11087),
.Y(n_11127)
);

INVx1_ASAP7_75t_SL g11128 ( 
.A(n_11050),
.Y(n_11128)
);

NOR3xp33_ASAP7_75t_L g11129 ( 
.A(n_11037),
.B(n_1964),
.C(n_1963),
.Y(n_11129)
);

CKINVDCx20_ASAP7_75t_R g11130 ( 
.A(n_11099),
.Y(n_11130)
);

OAI21xp5_ASAP7_75t_L g11131 ( 
.A1(n_11062),
.A2(n_1960),
.B(n_1964),
.Y(n_11131)
);

NOR3xp33_ASAP7_75t_L g11132 ( 
.A(n_11089),
.B(n_1967),
.C(n_1966),
.Y(n_11132)
);

INVx1_ASAP7_75t_L g11133 ( 
.A(n_11048),
.Y(n_11133)
);

AOI311xp33_ASAP7_75t_L g11134 ( 
.A1(n_11090),
.A2(n_1969),
.A3(n_1965),
.B(n_1968),
.C(n_1970),
.Y(n_11134)
);

INVxp67_ASAP7_75t_SL g11135 ( 
.A(n_11047),
.Y(n_11135)
);

AND2x2_ASAP7_75t_L g11136 ( 
.A(n_11071),
.B(n_1965),
.Y(n_11136)
);

A2O1A1Ixp33_ASAP7_75t_L g11137 ( 
.A1(n_11078),
.A2(n_1972),
.B(n_1969),
.C(n_1971),
.Y(n_11137)
);

NOR2x1_ASAP7_75t_L g11138 ( 
.A(n_11070),
.B(n_2246),
.Y(n_11138)
);

AOI31xp33_ASAP7_75t_L g11139 ( 
.A1(n_11076),
.A2(n_1975),
.A3(n_1971),
.B(n_1974),
.Y(n_11139)
);

OR2x2_ASAP7_75t_L g11140 ( 
.A(n_11052),
.B(n_1974),
.Y(n_11140)
);

AOI22xp5_ASAP7_75t_L g11141 ( 
.A1(n_11058),
.A2(n_1978),
.B1(n_1976),
.B2(n_1977),
.Y(n_11141)
);

NOR2xp33_ASAP7_75t_L g11142 ( 
.A(n_11117),
.B(n_11067),
.Y(n_11142)
);

AOI31xp33_ASAP7_75t_L g11143 ( 
.A1(n_11133),
.A2(n_11138),
.A3(n_11102),
.B(n_11104),
.Y(n_11143)
);

AND2x2_ASAP7_75t_L g11144 ( 
.A(n_11136),
.B(n_11097),
.Y(n_11144)
);

NOR3xp33_ASAP7_75t_L g11145 ( 
.A(n_11121),
.B(n_11063),
.C(n_11084),
.Y(n_11145)
);

NOR2xp33_ASAP7_75t_L g11146 ( 
.A(n_11124),
.B(n_11051),
.Y(n_11146)
);

NOR2xp33_ASAP7_75t_L g11147 ( 
.A(n_11139),
.B(n_11119),
.Y(n_11147)
);

INVx2_ASAP7_75t_L g11148 ( 
.A(n_11130),
.Y(n_11148)
);

NOR3xp33_ASAP7_75t_L g11149 ( 
.A(n_11105),
.B(n_11069),
.C(n_11094),
.Y(n_11149)
);

AND2x2_ASAP7_75t_L g11150 ( 
.A(n_11135),
.B(n_11111),
.Y(n_11150)
);

NOR2xp67_ASAP7_75t_L g11151 ( 
.A(n_11116),
.B(n_11096),
.Y(n_11151)
);

NAND3xp33_ASAP7_75t_SL g11152 ( 
.A(n_11123),
.B(n_11095),
.C(n_11068),
.Y(n_11152)
);

NAND2xp5_ASAP7_75t_L g11153 ( 
.A(n_11115),
.B(n_11064),
.Y(n_11153)
);

NAND2xp5_ASAP7_75t_SL g11154 ( 
.A(n_11134),
.B(n_11045),
.Y(n_11154)
);

NAND4xp25_ASAP7_75t_L g11155 ( 
.A(n_11126),
.B(n_11049),
.C(n_11092),
.D(n_11081),
.Y(n_11155)
);

NOR3xp33_ASAP7_75t_L g11156 ( 
.A(n_11131),
.B(n_11082),
.C(n_11072),
.Y(n_11156)
);

INVx4_ASAP7_75t_L g11157 ( 
.A(n_11118),
.Y(n_11157)
);

AND2x2_ASAP7_75t_L g11158 ( 
.A(n_11109),
.B(n_11088),
.Y(n_11158)
);

NOR3xp33_ASAP7_75t_L g11159 ( 
.A(n_11103),
.B(n_11100),
.C(n_11101),
.Y(n_11159)
);

NOR3xp33_ASAP7_75t_L g11160 ( 
.A(n_11129),
.B(n_11077),
.C(n_11074),
.Y(n_11160)
);

NOR3xp33_ASAP7_75t_L g11161 ( 
.A(n_11125),
.B(n_11073),
.C(n_11086),
.Y(n_11161)
);

HB1xp67_ASAP7_75t_L g11162 ( 
.A(n_11122),
.Y(n_11162)
);

NOR2xp33_ASAP7_75t_R g11163 ( 
.A(n_11112),
.B(n_1976),
.Y(n_11163)
);

INVx1_ASAP7_75t_L g11164 ( 
.A(n_11162),
.Y(n_11164)
);

AOI22xp5_ASAP7_75t_L g11165 ( 
.A1(n_11148),
.A2(n_11128),
.B1(n_11108),
.B2(n_11110),
.Y(n_11165)
);

INVx1_ASAP7_75t_SL g11166 ( 
.A(n_11163),
.Y(n_11166)
);

AOI221xp5_ASAP7_75t_L g11167 ( 
.A1(n_11143),
.A2(n_11127),
.B1(n_11106),
.B2(n_11107),
.C(n_11137),
.Y(n_11167)
);

AO22x2_ASAP7_75t_L g11168 ( 
.A1(n_11157),
.A2(n_11140),
.B1(n_11132),
.B2(n_11114),
.Y(n_11168)
);

AOI22xp5_ASAP7_75t_L g11169 ( 
.A1(n_11145),
.A2(n_11146),
.B1(n_11150),
.B2(n_11161),
.Y(n_11169)
);

NAND2xp5_ASAP7_75t_L g11170 ( 
.A(n_11147),
.B(n_11113),
.Y(n_11170)
);

AND2x2_ASAP7_75t_L g11171 ( 
.A(n_11144),
.B(n_11120),
.Y(n_11171)
);

AOI22xp33_ASAP7_75t_L g11172 ( 
.A1(n_11149),
.A2(n_11141),
.B1(n_1980),
.B2(n_1978),
.Y(n_11172)
);

NOR4xp25_ASAP7_75t_L g11173 ( 
.A(n_11155),
.B(n_2250),
.C(n_1981),
.D(n_1979),
.Y(n_11173)
);

AND2x4_ASAP7_75t_L g11174 ( 
.A(n_11158),
.B(n_1979),
.Y(n_11174)
);

NOR3xp33_ASAP7_75t_L g11175 ( 
.A(n_11159),
.B(n_1980),
.C(n_1981),
.Y(n_11175)
);

HB1xp67_ASAP7_75t_L g11176 ( 
.A(n_11151),
.Y(n_11176)
);

AND2x4_ASAP7_75t_L g11177 ( 
.A(n_11174),
.B(n_11156),
.Y(n_11177)
);

NOR2x1_ASAP7_75t_L g11178 ( 
.A(n_11164),
.B(n_11152),
.Y(n_11178)
);

INVx1_ASAP7_75t_L g11179 ( 
.A(n_11176),
.Y(n_11179)
);

NAND2xp5_ASAP7_75t_L g11180 ( 
.A(n_11173),
.B(n_11142),
.Y(n_11180)
);

OAI211xp5_ASAP7_75t_SL g11181 ( 
.A1(n_11169),
.A2(n_11153),
.B(n_11154),
.C(n_11160),
.Y(n_11181)
);

INVx2_ASAP7_75t_L g11182 ( 
.A(n_11168),
.Y(n_11182)
);

INVx1_ASAP7_75t_L g11183 ( 
.A(n_11168),
.Y(n_11183)
);

NAND3x2_ASAP7_75t_L g11184 ( 
.A(n_11171),
.B(n_1982),
.C(n_1983),
.Y(n_11184)
);

NOR4xp75_ASAP7_75t_L g11185 ( 
.A(n_11170),
.B(n_1985),
.C(n_1982),
.D(n_1984),
.Y(n_11185)
);

OAI22xp5_ASAP7_75t_SL g11186 ( 
.A1(n_11179),
.A2(n_11172),
.B1(n_11166),
.B2(n_11165),
.Y(n_11186)
);

AOI22xp5_ASAP7_75t_L g11187 ( 
.A1(n_11178),
.A2(n_11167),
.B1(n_11175),
.B2(n_1986),
.Y(n_11187)
);

NOR4xp25_ASAP7_75t_L g11188 ( 
.A(n_11181),
.B(n_1987),
.C(n_1984),
.D(n_1985),
.Y(n_11188)
);

NAND2x1p5_ASAP7_75t_L g11189 ( 
.A(n_11177),
.B(n_11183),
.Y(n_11189)
);

OAI222xp33_ASAP7_75t_R g11190 ( 
.A1(n_11182),
.A2(n_1989),
.B1(n_1991),
.B2(n_1987),
.C1(n_1988),
.C2(n_1990),
.Y(n_11190)
);

NAND5xp2_ASAP7_75t_L g11191 ( 
.A(n_11180),
.B(n_1992),
.C(n_1988),
.D(n_1990),
.E(n_1993),
.Y(n_11191)
);

NAND3xp33_ASAP7_75t_L g11192 ( 
.A(n_11187),
.B(n_11188),
.C(n_11184),
.Y(n_11192)
);

OAI21xp5_ASAP7_75t_L g11193 ( 
.A1(n_11189),
.A2(n_11185),
.B(n_1992),
.Y(n_11193)
);

INVx1_ASAP7_75t_L g11194 ( 
.A(n_11186),
.Y(n_11194)
);

INVxp67_ASAP7_75t_L g11195 ( 
.A(n_11193),
.Y(n_11195)
);

AND3x4_ASAP7_75t_L g11196 ( 
.A(n_11192),
.B(n_11190),
.C(n_11191),
.Y(n_11196)
);

OAI22xp5_ASAP7_75t_L g11197 ( 
.A1(n_11196),
.A2(n_11194),
.B1(n_11195),
.B2(n_1995),
.Y(n_11197)
);

OR4x1_ASAP7_75t_L g11198 ( 
.A(n_11196),
.B(n_1995),
.C(n_1993),
.D(n_1994),
.Y(n_11198)
);

NAND2xp5_ASAP7_75t_L g11199 ( 
.A(n_11197),
.B(n_1994),
.Y(n_11199)
);

XNOR2xp5_ASAP7_75t_L g11200 ( 
.A(n_11198),
.B(n_1996),
.Y(n_11200)
);

OAI22xp5_ASAP7_75t_L g11201 ( 
.A1(n_11200),
.A2(n_1998),
.B1(n_1996),
.B2(n_1997),
.Y(n_11201)
);

OAI31xp67_ASAP7_75t_SL g11202 ( 
.A1(n_11199),
.A2(n_2000),
.A3(n_1997),
.B(n_1999),
.Y(n_11202)
);

INVx1_ASAP7_75t_L g11203 ( 
.A(n_11201),
.Y(n_11203)
);

AOI21xp5_ASAP7_75t_L g11204 ( 
.A1(n_11202),
.A2(n_1999),
.B(n_2000),
.Y(n_11204)
);

INVx1_ASAP7_75t_L g11205 ( 
.A(n_11204),
.Y(n_11205)
);

AOI222xp33_ASAP7_75t_L g11206 ( 
.A1(n_11205),
.A2(n_11203),
.B1(n_2003),
.B2(n_2004),
.C1(n_2001),
.C2(n_2002),
.Y(n_11206)
);

OAI21x1_ASAP7_75t_SL g11207 ( 
.A1(n_11206),
.A2(n_2003),
.B(n_2002),
.Y(n_11207)
);

INVx1_ASAP7_75t_L g11208 ( 
.A(n_11207),
.Y(n_11208)
);

INVx1_ASAP7_75t_L g11209 ( 
.A(n_11207),
.Y(n_11209)
);

INVx1_ASAP7_75t_L g11210 ( 
.A(n_11207),
.Y(n_11210)
);

OR2x6_ASAP7_75t_L g11211 ( 
.A(n_11208),
.B(n_2004),
.Y(n_11211)
);

NAND2xp33_ASAP7_75t_SL g11212 ( 
.A(n_11209),
.B(n_11210),
.Y(n_11212)
);

AOI21xp5_ASAP7_75t_L g11213 ( 
.A1(n_11212),
.A2(n_2005),
.B(n_2007),
.Y(n_11213)
);

AOI211xp5_ASAP7_75t_L g11214 ( 
.A1(n_11213),
.A2(n_11211),
.B(n_2013),
.C(n_2009),
.Y(n_11214)
);


endmodule