module fake_jpeg_26830_n_332 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_332);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_332;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_145;
wire n_20;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_14),
.Y(n_26)
);

BUFx4f_ASAP7_75t_SL g27 ( 
.A(n_13),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g28 ( 
.A(n_13),
.B(n_10),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_13),
.B(n_0),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_10),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_11),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

INVx2_ASAP7_75t_SL g37 ( 
.A(n_19),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_41),
.Y(n_51)
);

BUFx10_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_28),
.B(n_7),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_42),
.B(n_25),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_46),
.B(n_57),
.Y(n_72)
);

AOI21xp33_ASAP7_75t_L g52 ( 
.A1(n_42),
.A2(n_29),
.B(n_28),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_52),
.B(n_26),
.C(n_30),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_53),
.B(n_25),
.Y(n_76)
);

BUFx12_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_56),
.Y(n_67)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_41),
.B(n_30),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_59),
.B(n_33),
.Y(n_85)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_60),
.Y(n_88)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_62),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_35),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_63),
.B(n_35),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_53),
.A2(n_44),
.B1(n_17),
.B2(n_32),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_64),
.A2(n_39),
.B1(n_23),
.B2(n_34),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_65),
.B(n_85),
.Y(n_100)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_61),
.Y(n_66)
);

INVx13_ASAP7_75t_L g97 ( 
.A(n_66),
.Y(n_97)
);

BUFx2_ASAP7_75t_L g68 ( 
.A(n_60),
.Y(n_68)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_68),
.Y(n_103)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_55),
.Y(n_69)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_69),
.Y(n_115)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_71),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_63),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_73),
.Y(n_96)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_74),
.Y(n_102)
);

OR2x2_ASAP7_75t_L g105 ( 
.A(n_75),
.B(n_76),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_61),
.A2(n_17),
.B1(n_44),
.B2(n_32),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_77),
.A2(n_81),
.B1(n_82),
.B2(n_50),
.Y(n_116)
);

HB1xp67_ASAP7_75t_L g78 ( 
.A(n_48),
.Y(n_78)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_78),
.Y(n_106)
);

HB1xp67_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_79),
.Y(n_120)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_48),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_80),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_61),
.A2(n_17),
.B1(n_32),
.B2(n_37),
.Y(n_81)
);

NAND2xp67_ASAP7_75t_SL g82 ( 
.A(n_52),
.B(n_27),
.Y(n_82)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_58),
.Y(n_83)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_83),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_55),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_84),
.Y(n_101)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_47),
.Y(n_86)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_86),
.Y(n_99)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_50),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_87),
.B(n_90),
.Y(n_121)
);

BUFx8_ASAP7_75t_L g89 ( 
.A(n_50),
.Y(n_89)
);

BUFx2_ASAP7_75t_L g122 ( 
.A(n_89),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_51),
.B(n_45),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_49),
.Y(n_91)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_91),
.Y(n_95)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_58),
.Y(n_92)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_92),
.Y(n_108)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_54),
.Y(n_93)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_93),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_90),
.B(n_51),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_104),
.B(n_107),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_82),
.B(n_62),
.C(n_54),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_87),
.A2(n_69),
.B1(n_74),
.B2(n_36),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_109),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_72),
.B(n_57),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_110),
.B(n_114),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_83),
.A2(n_45),
.B1(n_26),
.B2(n_33),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_112),
.A2(n_23),
.B1(n_18),
.B2(n_22),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_92),
.A2(n_39),
.B1(n_58),
.B2(n_49),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_113),
.A2(n_118),
.B1(n_60),
.B2(n_34),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_75),
.B(n_46),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_116),
.A2(n_76),
.B1(n_23),
.B2(n_18),
.Y(n_138)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_70),
.Y(n_117)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_117),
.Y(n_146)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_119),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_123),
.B(n_131),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_107),
.A2(n_77),
.B1(n_81),
.B2(n_80),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_124),
.A2(n_136),
.B1(n_145),
.B2(n_148),
.Y(n_171)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_122),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_125),
.B(n_129),
.Y(n_155)
);

INVx2_ASAP7_75t_SL g126 ( 
.A(n_95),
.Y(n_126)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_126),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_128),
.A2(n_138),
.B1(n_22),
.B2(n_20),
.Y(n_154)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_122),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_96),
.A2(n_101),
.B1(n_115),
.B2(n_98),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_130),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_100),
.B(n_59),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_110),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_132),
.B(n_141),
.Y(n_161)
);

INVxp33_ASAP7_75t_L g134 ( 
.A(n_119),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_134),
.B(n_140),
.Y(n_168)
);

INVx13_ASAP7_75t_L g135 ( 
.A(n_97),
.Y(n_135)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_135),
.Y(n_152)
);

NAND2xp33_ASAP7_75t_SL g137 ( 
.A(n_104),
.B(n_35),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_137),
.A2(n_139),
.B(n_38),
.Y(n_179)
);

XNOR2x1_ASAP7_75t_L g139 ( 
.A(n_114),
.B(n_27),
.Y(n_139)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_98),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_108),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_108),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_142),
.B(n_147),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_97),
.B(n_120),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_143),
.B(n_144),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_105),
.B(n_31),
.Y(n_144)
);

OAI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_105),
.A2(n_19),
.B1(n_21),
.B2(n_91),
.Y(n_145)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_106),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_118),
.A2(n_43),
.B1(n_40),
.B2(n_38),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_121),
.B(n_31),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_149),
.Y(n_175)
);

INVx1_ASAP7_75t_SL g151 ( 
.A(n_115),
.Y(n_151)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_151),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_154),
.A2(n_158),
.B1(n_165),
.B2(n_181),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_127),
.B(n_133),
.C(n_139),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_156),
.B(n_157),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_127),
.B(n_120),
.C(n_106),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_132),
.A2(n_95),
.B1(n_111),
.B2(n_94),
.Y(n_158)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_147),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_164),
.B(n_166),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_138),
.A2(n_103),
.B1(n_111),
.B2(n_117),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_141),
.Y(n_166)
);

OA21x2_ASAP7_75t_L g167 ( 
.A1(n_137),
.A2(n_103),
.B(n_34),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_167),
.A2(n_185),
.B(n_24),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_146),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_169),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_146),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_170),
.B(n_173),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_124),
.A2(n_99),
.B1(n_94),
.B2(n_102),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_172),
.A2(n_174),
.B1(n_182),
.B2(n_126),
.Y(n_186)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_142),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_136),
.A2(n_99),
.B1(n_102),
.B2(n_89),
.Y(n_174)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_148),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_176),
.B(n_177),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_135),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_133),
.B(n_56),
.C(n_43),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_SL g207 ( 
.A(n_178),
.B(n_179),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_150),
.A2(n_0),
.B(n_1),
.Y(n_180)
);

OAI21xp33_ASAP7_75t_L g192 ( 
.A1(n_180),
.A2(n_0),
.B(n_1),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_150),
.A2(n_40),
.B1(n_43),
.B2(n_20),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_140),
.A2(n_89),
.B1(n_40),
.B2(n_38),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_151),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_183),
.B(n_126),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_125),
.A2(n_129),
.B(n_24),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_186),
.A2(n_203),
.B1(n_153),
.B2(n_162),
.Y(n_227)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_187),
.Y(n_218)
);

OAI32xp33_ASAP7_75t_L g189 ( 
.A1(n_161),
.A2(n_19),
.A3(n_21),
.B1(n_38),
.B2(n_25),
.Y(n_189)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_189),
.Y(n_222)
);

BUFx3_ASAP7_75t_L g190 ( 
.A(n_152),
.Y(n_190)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_190),
.Y(n_241)
);

INVx13_ASAP7_75t_L g191 ( 
.A(n_152),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_191),
.B(n_194),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_192),
.B(n_195),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_193),
.A2(n_208),
.B1(n_182),
.B2(n_192),
.Y(n_238)
);

AND2x6_ASAP7_75t_L g194 ( 
.A(n_156),
.B(n_14),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_155),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_170),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_196),
.B(n_198),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_184),
.B(n_123),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_197),
.B(n_183),
.Y(n_223)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_163),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_163),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_199),
.B(n_200),
.Y(n_225)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_155),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_153),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_201),
.B(n_204),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_168),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_202),
.B(n_205),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_176),
.A2(n_68),
.B1(n_88),
.B2(n_21),
.Y(n_203)
);

INVx13_ASAP7_75t_L g204 ( 
.A(n_162),
.Y(n_204)
);

OR2x2_ASAP7_75t_L g205 ( 
.A(n_161),
.B(n_25),
.Y(n_205)
);

AO22x1_ASAP7_75t_SL g206 ( 
.A1(n_167),
.A2(n_88),
.B1(n_21),
.B2(n_16),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_206),
.B(n_181),
.Y(n_233)
);

OAI22x1_ASAP7_75t_SL g208 ( 
.A1(n_171),
.A2(n_24),
.B1(n_1),
.B2(n_2),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g211 ( 
.A(n_159),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_211),
.B(n_212),
.Y(n_242)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_158),
.Y(n_212)
);

HB1xp67_ASAP7_75t_L g215 ( 
.A(n_157),
.Y(n_215)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_215),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_216),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_SL g258 ( 
.A1(n_219),
.A2(n_233),
.B(n_237),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_209),
.B(n_178),
.C(n_179),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_221),
.B(n_207),
.C(n_205),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_223),
.B(n_226),
.Y(n_248)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_214),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_227),
.A2(n_213),
.B1(n_193),
.B2(n_202),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_186),
.A2(n_160),
.B1(n_171),
.B2(n_172),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_228),
.A2(n_206),
.B1(n_189),
.B2(n_207),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_210),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_229),
.Y(n_249)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_188),
.Y(n_231)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_231),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_209),
.B(n_185),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_232),
.B(n_175),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_208),
.A2(n_174),
.B1(n_160),
.B2(n_164),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_235),
.A2(n_236),
.B1(n_238),
.B2(n_206),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_213),
.A2(n_180),
.B1(n_167),
.B2(n_166),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_191),
.Y(n_237)
);

HB1xp67_ASAP7_75t_L g240 ( 
.A(n_190),
.Y(n_240)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_240),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_243),
.A2(n_252),
.B1(n_263),
.B2(n_241),
.Y(n_275)
);

INVx1_ASAP7_75t_SL g244 ( 
.A(n_230),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_244),
.B(n_256),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_246),
.A2(n_251),
.B1(n_260),
.B2(n_230),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_217),
.A2(n_222),
.B1(n_231),
.B2(n_228),
.Y(n_247)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_247),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_250),
.B(n_253),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_236),
.A2(n_203),
.B1(n_196),
.B2(n_201),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_221),
.B(n_194),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_222),
.A2(n_175),
.B1(n_204),
.B2(n_173),
.Y(n_254)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_254),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_SL g267 ( 
.A(n_255),
.B(n_257),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_232),
.B(n_67),
.C(n_56),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_224),
.B(n_56),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_233),
.A2(n_8),
.B1(n_15),
.B2(n_12),
.Y(n_259)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_259),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_235),
.A2(n_66),
.B1(n_67),
.B2(n_2),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_234),
.A2(n_7),
.B1(n_15),
.B2(n_12),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_262),
.B(n_242),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_227),
.A2(n_66),
.B1(n_1),
.B2(n_2),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_264),
.A2(n_266),
.B1(n_280),
.B2(n_263),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_246),
.A2(n_226),
.B1(n_219),
.B2(n_218),
.Y(n_266)
);

FAx1_ASAP7_75t_SL g268 ( 
.A(n_250),
.B(n_225),
.CI(n_252),
.CON(n_268),
.SN(n_268)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_268),
.Y(n_281)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_270),
.Y(n_285)
);

AOI22xp33_ASAP7_75t_L g271 ( 
.A1(n_244),
.A2(n_237),
.B1(n_241),
.B2(n_218),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_271),
.A2(n_275),
.B1(n_278),
.B2(n_261),
.Y(n_284)
);

AND2x2_ASAP7_75t_L g272 ( 
.A(n_251),
.B(n_220),
.Y(n_272)
);

AO21x1_ASAP7_75t_L g289 ( 
.A1(n_272),
.A2(n_258),
.B(n_245),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_249),
.B(n_229),
.Y(n_274)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_274),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_249),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_276),
.B(n_248),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_258),
.A2(n_224),
.B1(n_239),
.B2(n_16),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_260),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_280)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_282),
.Y(n_304)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_283),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_284),
.B(n_288),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_265),
.B(n_256),
.C(n_255),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_287),
.B(n_290),
.C(n_292),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_278),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_289),
.A2(n_294),
.B(n_295),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_269),
.B(n_253),
.C(n_257),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_269),
.B(n_245),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_291),
.B(n_267),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_273),
.B(n_261),
.C(n_8),
.Y(n_292)
);

OAI21xp33_ASAP7_75t_L g293 ( 
.A1(n_277),
.A2(n_9),
.B(n_11),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_293),
.B(n_280),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_272),
.A2(n_9),
.B(n_4),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_272),
.A2(n_279),
.B(n_268),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_288),
.A2(n_275),
.B1(n_268),
.B2(n_266),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_297),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_287),
.B(n_267),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_298),
.B(n_299),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_290),
.B(n_264),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_301),
.B(n_305),
.C(n_307),
.Y(n_309)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_303),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_291),
.B(n_3),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_281),
.B(n_3),
.C(n_4),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_307),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_311),
.B(n_315),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_304),
.A2(n_289),
.B(n_286),
.Y(n_312)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_312),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_300),
.A2(n_285),
.B(n_292),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_SL g317 ( 
.A(n_313),
.B(n_305),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g315 ( 
.A1(n_302),
.A2(n_283),
.B(n_293),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_306),
.B(n_3),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_316),
.B(n_4),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_317),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_318),
.B(n_319),
.C(n_320),
.Y(n_325)
);

NOR2x1_ASAP7_75t_L g319 ( 
.A(n_308),
.B(n_296),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_314),
.A2(n_301),
.B1(n_296),
.B2(n_299),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_321),
.B(n_309),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_323),
.B(n_321),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_326),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_327),
.B(n_325),
.C(n_323),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_328),
.B(n_324),
.C(n_322),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_329),
.A2(n_316),
.B1(n_310),
.B2(n_6),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_L g331 ( 
.A1(n_330),
.A2(n_4),
.B(n_5),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_331),
.B(n_6),
.Y(n_332)
);


endmodule