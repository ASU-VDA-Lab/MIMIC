module fake_jpeg_12638_n_595 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_595);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_595;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_393;
wire n_288;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_18;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx1_ASAP7_75t_SL g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx8_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

BUFx12_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_9),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_12),
.Y(n_35)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_4),
.Y(n_38)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_0),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_11),
.B(n_12),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_5),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

INVx2_ASAP7_75t_SL g44 ( 
.A(n_5),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_1),
.Y(n_45)
);

CKINVDCx5p33_ASAP7_75t_R g46 ( 
.A(n_3),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_11),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_7),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_14),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_12),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_1),
.Y(n_51)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_9),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_16),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_13),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_1),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_4),
.B(n_2),
.Y(n_56)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_5),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_13),
.Y(n_58)
);

BUFx24_ASAP7_75t_L g59 ( 
.A(n_15),
.Y(n_59)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_59),
.Y(n_60)
);

INVx11_ASAP7_75t_L g129 ( 
.A(n_60),
.Y(n_129)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_59),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g179 ( 
.A(n_61),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_30),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_62),
.B(n_63),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_30),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_31),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g137 ( 
.A(n_64),
.Y(n_137)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_27),
.Y(n_65)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_65),
.Y(n_134)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_27),
.Y(n_66)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_66),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_19),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_67),
.Y(n_125)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_54),
.Y(n_68)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_68),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_19),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_69),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_19),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_70),
.Y(n_130)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_59),
.Y(n_71)
);

INVx5_ASAP7_75t_L g153 ( 
.A(n_71),
.Y(n_153)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_54),
.Y(n_72)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_72),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_53),
.B(n_58),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_73),
.B(n_79),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_41),
.A2(n_17),
.B1(n_16),
.B2(n_15),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g145 ( 
.A1(n_74),
.A2(n_25),
.B1(n_44),
.B2(n_28),
.Y(n_145)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_31),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g161 ( 
.A(n_75),
.Y(n_161)
);

INVx3_ASAP7_75t_SL g76 ( 
.A(n_59),
.Y(n_76)
);

CKINVDCx6p67_ASAP7_75t_R g183 ( 
.A(n_76),
.Y(n_183)
);

INVx8_ASAP7_75t_SL g77 ( 
.A(n_46),
.Y(n_77)
);

INVx4_ASAP7_75t_SL g157 ( 
.A(n_77),
.Y(n_157)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_50),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g166 ( 
.A(n_78),
.Y(n_166)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_20),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_29),
.Y(n_80)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_80),
.Y(n_126)
);

AND2x2_ASAP7_75t_SL g81 ( 
.A(n_46),
.B(n_0),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_81),
.B(n_82),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_30),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_22),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_83),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_50),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g188 ( 
.A(n_84),
.Y(n_188)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_49),
.Y(n_85)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_85),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_32),
.Y(n_86)
);

INVx5_ASAP7_75t_L g164 ( 
.A(n_86),
.Y(n_164)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_22),
.Y(n_87)
);

INVx5_ASAP7_75t_L g170 ( 
.A(n_87),
.Y(n_170)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_32),
.Y(n_88)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_88),
.Y(n_141)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_29),
.Y(n_89)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_89),
.Y(n_140)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_20),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_90),
.B(n_93),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_22),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_91),
.Y(n_144)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_39),
.Y(n_92)
);

INVx6_ASAP7_75t_L g201 ( 
.A(n_92),
.Y(n_201)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_21),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_36),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_94),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_36),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_95),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_36),
.Y(n_96)
);

INVx8_ASAP7_75t_L g174 ( 
.A(n_96),
.Y(n_174)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_49),
.Y(n_97)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_97),
.Y(n_159)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_32),
.Y(n_98)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_98),
.Y(n_148)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_49),
.Y(n_99)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_99),
.Y(n_136)
);

BUFx10_ASAP7_75t_L g100 ( 
.A(n_26),
.Y(n_100)
);

INVx2_ASAP7_75t_SL g163 ( 
.A(n_100),
.Y(n_163)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_32),
.Y(n_101)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_101),
.Y(n_151)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_49),
.Y(n_102)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_102),
.Y(n_162)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_49),
.Y(n_103)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_103),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_52),
.Y(n_104)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_104),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_41),
.B(n_56),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_105),
.B(n_110),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_52),
.Y(n_106)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_106),
.Y(n_152)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_32),
.Y(n_107)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_107),
.Y(n_177)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_52),
.Y(n_108)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_108),
.Y(n_167)
);

BUFx5_ASAP7_75t_L g109 ( 
.A(n_39),
.Y(n_109)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_109),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_56),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_34),
.Y(n_111)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_111),
.Y(n_180)
);

AND2x6_ASAP7_75t_L g112 ( 
.A(n_53),
.B(n_14),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_112),
.B(n_116),
.Y(n_173)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_57),
.Y(n_113)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_113),
.Y(n_194)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_34),
.Y(n_114)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_114),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_57),
.Y(n_115)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_115),
.Y(n_185)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_21),
.Y(n_116)
);

INVx1_ASAP7_75t_SL g117 ( 
.A(n_25),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_117),
.B(n_118),
.Y(n_176)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_23),
.Y(n_118)
);

INVx8_ASAP7_75t_L g119 ( 
.A(n_39),
.Y(n_119)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_119),
.Y(n_186)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_23),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_120),
.B(n_55),
.Y(n_181)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_34),
.Y(n_121)
);

HB1xp67_ASAP7_75t_L g146 ( 
.A(n_121),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_57),
.Y(n_122)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_122),
.Y(n_187)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_26),
.Y(n_123)
);

INVx2_ASAP7_75t_SL g168 ( 
.A(n_123),
.Y(n_168)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_26),
.Y(n_124)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_124),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_81),
.B(n_58),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_127),
.B(n_133),
.Y(n_227)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_114),
.B(n_25),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g244 ( 
.A(n_131),
.B(n_149),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_60),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_132),
.B(n_156),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_121),
.B(n_35),
.Y(n_133)
);

INVx6_ASAP7_75t_SL g142 ( 
.A(n_100),
.Y(n_142)
);

CKINVDCx9p33_ASAP7_75t_R g272 ( 
.A(n_142),
.Y(n_272)
);

INVx11_ASAP7_75t_L g143 ( 
.A(n_100),
.Y(n_143)
);

CKINVDCx6p67_ASAP7_75t_R g232 ( 
.A(n_143),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_145),
.A2(n_44),
.B1(n_34),
.B2(n_47),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_76),
.B(n_26),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_64),
.A2(n_44),
.B1(n_34),
.B2(n_28),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_154),
.A2(n_38),
.B(n_33),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_119),
.Y(n_156)
);

NAND3xp33_ASAP7_75t_L g160 ( 
.A(n_112),
.B(n_37),
.C(n_51),
.Y(n_160)
);

NOR3xp33_ASAP7_75t_L g275 ( 
.A(n_160),
.B(n_6),
.C(n_7),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_87),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_165),
.B(n_175),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_92),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_181),
.B(n_193),
.Y(n_254)
);

INVx4_ASAP7_75t_SL g182 ( 
.A(n_94),
.Y(n_182)
);

INVx4_ASAP7_75t_SL g249 ( 
.A(n_182),
.Y(n_249)
);

OAI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_67),
.A2(n_28),
.B1(n_51),
.B2(n_48),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_184),
.A2(n_30),
.B1(n_2),
.B2(n_3),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_86),
.B(n_18),
.Y(n_193)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_69),
.Y(n_195)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_195),
.Y(n_206)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_70),
.Y(n_197)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_197),
.Y(n_208)
);

INVx4_ASAP7_75t_SL g198 ( 
.A(n_122),
.Y(n_198)
);

INVx4_ASAP7_75t_L g209 ( 
.A(n_198),
.Y(n_209)
);

BUFx10_ASAP7_75t_L g199 ( 
.A(n_75),
.Y(n_199)
);

BUFx2_ASAP7_75t_L g219 ( 
.A(n_199),
.Y(n_219)
);

INVx4_ASAP7_75t_SL g200 ( 
.A(n_115),
.Y(n_200)
);

INVx1_ASAP7_75t_SL g224 ( 
.A(n_200),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_88),
.B(n_18),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_202),
.B(n_203),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_111),
.B(n_33),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_169),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_207),
.B(n_213),
.Y(n_278)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_177),
.Y(n_210)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_210),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_211),
.A2(n_217),
.B1(n_238),
.B2(n_274),
.Y(n_279)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_170),
.Y(n_212)
);

INVx4_ASAP7_75t_L g283 ( 
.A(n_212),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_169),
.Y(n_213)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_159),
.Y(n_215)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_215),
.Y(n_282)
);

AOI22xp33_ASAP7_75t_L g216 ( 
.A1(n_184),
.A2(n_91),
.B1(n_83),
.B2(n_96),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_216),
.A2(n_261),
.B1(n_154),
.B2(n_193),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_173),
.A2(n_106),
.B1(n_104),
.B2(n_95),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_137),
.A2(n_84),
.B1(n_78),
.B2(n_101),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_SL g294 ( 
.A1(n_218),
.A2(n_226),
.B1(n_255),
.B2(n_256),
.Y(n_294)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_134),
.Y(n_220)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_220),
.Y(n_286)
);

OR2x4_ASAP7_75t_L g221 ( 
.A(n_158),
.B(n_98),
.Y(n_221)
);

AO22x1_ASAP7_75t_L g290 ( 
.A1(n_221),
.A2(n_264),
.B1(n_269),
.B2(n_163),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_149),
.Y(n_222)
);

HB1xp67_ASAP7_75t_L g296 ( 
.A(n_222),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_147),
.B(n_55),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_223),
.B(n_231),
.Y(n_312)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_186),
.Y(n_225)
);

INVx4_ASAP7_75t_L g295 ( 
.A(n_225),
.Y(n_295)
);

AOI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_161),
.A2(n_166),
.B1(n_188),
.B2(n_174),
.Y(n_226)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_164),
.Y(n_228)
);

INVx3_ASAP7_75t_L g323 ( 
.A(n_228),
.Y(n_323)
);

INVx6_ASAP7_75t_L g229 ( 
.A(n_125),
.Y(n_229)
);

INVx5_ASAP7_75t_L g314 ( 
.A(n_229),
.Y(n_314)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_155),
.Y(n_230)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_230),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_147),
.B(n_24),
.Y(n_231)
);

BUFx3_ASAP7_75t_L g233 ( 
.A(n_179),
.Y(n_233)
);

BUFx3_ASAP7_75t_L g288 ( 
.A(n_233),
.Y(n_288)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_125),
.Y(n_234)
);

INVx5_ASAP7_75t_L g318 ( 
.A(n_234),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_172),
.B(n_24),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_235),
.B(n_239),
.Y(n_287)
);

INVx6_ASAP7_75t_L g236 ( 
.A(n_128),
.Y(n_236)
);

INVx5_ASAP7_75t_L g324 ( 
.A(n_236),
.Y(n_324)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_162),
.Y(n_237)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_237),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_173),
.A2(n_38),
.B1(n_35),
.B2(n_45),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_172),
.B(n_48),
.Y(n_239)
);

INVx6_ASAP7_75t_L g240 ( 
.A(n_128),
.Y(n_240)
);

INVx3_ASAP7_75t_L g334 ( 
.A(n_240),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_139),
.B(n_47),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_241),
.B(n_243),
.Y(n_289)
);

CKINVDCx12_ASAP7_75t_R g242 ( 
.A(n_157),
.Y(n_242)
);

INVx4_ASAP7_75t_SL g297 ( 
.A(n_242),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_139),
.B(n_43),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_181),
.B(n_43),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_245),
.B(n_266),
.Y(n_316)
);

HB1xp67_ASAP7_75t_L g246 ( 
.A(n_146),
.Y(n_246)
);

HB1xp67_ASAP7_75t_L g327 ( 
.A(n_246),
.Y(n_327)
);

HB1xp67_ASAP7_75t_L g247 ( 
.A(n_146),
.Y(n_247)
);

CKINVDCx16_ASAP7_75t_R g299 ( 
.A(n_247),
.Y(n_299)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_171),
.Y(n_248)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_248),
.Y(n_304)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_191),
.Y(n_250)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_250),
.Y(n_308)
);

INVx6_ASAP7_75t_L g251 ( 
.A(n_130),
.Y(n_251)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_251),
.Y(n_305)
);

BUFx12f_ASAP7_75t_L g252 ( 
.A(n_199),
.Y(n_252)
);

BUFx3_ASAP7_75t_L g302 ( 
.A(n_252),
.Y(n_302)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_196),
.Y(n_253)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_253),
.Y(n_306)
);

AOI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_199),
.A2(n_37),
.B1(n_42),
.B2(n_40),
.Y(n_255)
);

AOI22xp33_ASAP7_75t_SL g256 ( 
.A1(n_150),
.A2(n_45),
.B1(n_42),
.B2(n_40),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g313 ( 
.A1(n_257),
.A2(n_129),
.B(n_183),
.Y(n_313)
);

CKINVDCx12_ASAP7_75t_R g258 ( 
.A(n_157),
.Y(n_258)
);

NAND2x1_ASAP7_75t_SL g333 ( 
.A(n_258),
.B(n_228),
.Y(n_333)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_185),
.Y(n_259)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_259),
.Y(n_310)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_204),
.Y(n_260)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_260),
.Y(n_329)
);

A2O1A1Ixp33_ASAP7_75t_L g262 ( 
.A1(n_158),
.A2(n_17),
.B(n_14),
.C(n_13),
.Y(n_262)
);

O2A1O1Ixp33_ASAP7_75t_L g315 ( 
.A1(n_262),
.A2(n_183),
.B(n_8),
.C(n_9),
.Y(n_315)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_187),
.Y(n_263)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_263),
.Y(n_317)
);

OR2x4_ASAP7_75t_L g264 ( 
.A(n_160),
.B(n_17),
.Y(n_264)
);

INVx3_ASAP7_75t_L g265 ( 
.A(n_152),
.Y(n_265)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_265),
.Y(n_277)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_135),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_126),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_267),
.B(n_268),
.Y(n_320)
);

INVx6_ASAP7_75t_L g268 ( 
.A(n_130),
.Y(n_268)
);

NOR2x1_ASAP7_75t_L g269 ( 
.A(n_131),
.B(n_0),
.Y(n_269)
);

INVx5_ASAP7_75t_L g270 ( 
.A(n_141),
.Y(n_270)
);

AND2x2_ASAP7_75t_L g301 ( 
.A(n_270),
.B(n_271),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_176),
.B(n_3),
.Y(n_271)
);

INVx6_ASAP7_75t_L g273 ( 
.A(n_138),
.Y(n_273)
);

AOI22xp33_ASAP7_75t_SL g298 ( 
.A1(n_273),
.A2(n_163),
.B1(n_179),
.B2(n_153),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_145),
.A2(n_3),
.B1(n_6),
.B2(n_7),
.Y(n_274)
);

AND2x2_ASAP7_75t_L g309 ( 
.A(n_275),
.B(n_272),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_216),
.A2(n_201),
.B1(n_140),
.B2(n_144),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_280),
.A2(n_321),
.B1(n_330),
.B2(n_331),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_276),
.B(n_176),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_284),
.B(n_325),
.Y(n_335)
);

AND2x2_ASAP7_75t_L g347 ( 
.A(n_285),
.B(n_313),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_290),
.B(n_309),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_214),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_291),
.B(n_309),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_222),
.A2(n_194),
.B1(n_167),
.B2(n_178),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g343 ( 
.A(n_292),
.Y(n_343)
);

AOI22xp33_ASAP7_75t_L g293 ( 
.A1(n_244),
.A2(n_192),
.B1(n_189),
.B2(n_168),
.Y(n_293)
);

OA22x2_ASAP7_75t_L g378 ( 
.A1(n_293),
.A2(n_300),
.B1(n_280),
.B2(n_321),
.Y(n_378)
);

INVxp67_ASAP7_75t_L g362 ( 
.A(n_298),
.Y(n_362)
);

AOI22xp33_ASAP7_75t_L g300 ( 
.A1(n_244),
.A2(n_168),
.B1(n_190),
.B2(n_202),
.Y(n_300)
);

AOI22xp33_ASAP7_75t_SL g311 ( 
.A1(n_224),
.A2(n_148),
.B1(n_180),
.B2(n_151),
.Y(n_311)
);

OAI22xp33_ASAP7_75t_SL g358 ( 
.A1(n_311),
.A2(n_328),
.B1(n_233),
.B2(n_219),
.Y(n_358)
);

AND2x2_ASAP7_75t_L g357 ( 
.A(n_315),
.B(n_322),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_227),
.B(n_254),
.C(n_221),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_319),
.B(n_255),
.C(n_219),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_205),
.A2(n_136),
.B1(n_200),
.B2(n_182),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_256),
.A2(n_198),
.B1(n_183),
.B2(n_11),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_262),
.B(n_6),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_L g326 ( 
.A1(n_226),
.A2(n_8),
.B(n_218),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_L g359 ( 
.A1(n_326),
.A2(n_232),
.B(n_234),
.Y(n_359)
);

AOI22xp33_ASAP7_75t_SL g328 ( 
.A1(n_224),
.A2(n_272),
.B1(n_265),
.B2(n_212),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_264),
.A2(n_206),
.B1(n_208),
.B2(n_225),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_229),
.A2(n_268),
.B1(n_251),
.B2(n_240),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_249),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_332),
.B(n_232),
.Y(n_354)
);

INVx1_ASAP7_75t_SL g376 ( 
.A(n_333),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_327),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_336),
.B(n_342),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_284),
.B(n_269),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_338),
.B(n_350),
.Y(n_384)
);

INVx3_ASAP7_75t_L g339 ( 
.A(n_283),
.Y(n_339)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_339),
.Y(n_388)
);

INVx2_ASAP7_75t_SL g340 ( 
.A(n_314),
.Y(n_340)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_340),
.Y(n_392)
);

BUFx6f_ASAP7_75t_L g341 ( 
.A(n_318),
.Y(n_341)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_341),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_333),
.Y(n_342)
);

INVx13_ASAP7_75t_L g344 ( 
.A(n_297),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_344),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_345),
.B(n_299),
.C(n_329),
.Y(n_393)
);

AOI22xp33_ASAP7_75t_L g346 ( 
.A1(n_296),
.A2(n_209),
.B1(n_273),
.B2(n_236),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_L g390 ( 
.A1(n_346),
.A2(n_378),
.B1(n_331),
.B2(n_277),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_SL g349 ( 
.A(n_278),
.B(n_249),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_SL g396 ( 
.A(n_349),
.B(n_366),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_301),
.B(n_270),
.Y(n_350)
);

INVx8_ASAP7_75t_L g351 ( 
.A(n_318),
.Y(n_351)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_351),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_301),
.B(n_209),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_352),
.B(n_361),
.Y(n_387)
);

AND2x6_ASAP7_75t_L g353 ( 
.A(n_319),
.B(n_232),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_SL g389 ( 
.A(n_353),
.B(n_367),
.C(n_277),
.Y(n_389)
);

NAND3xp33_ASAP7_75t_L g409 ( 
.A(n_354),
.B(n_371),
.C(n_373),
.Y(n_409)
);

INVx3_ASAP7_75t_L g355 ( 
.A(n_283),
.Y(n_355)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_355),
.Y(n_402)
);

INVx3_ASAP7_75t_L g356 ( 
.A(n_314),
.Y(n_356)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_356),
.Y(n_407)
);

AOI22xp33_ASAP7_75t_SL g410 ( 
.A1(n_358),
.A2(n_369),
.B1(n_370),
.B2(n_377),
.Y(n_410)
);

AOI21xp5_ASAP7_75t_L g385 ( 
.A1(n_359),
.A2(n_376),
.B(n_362),
.Y(n_385)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_286),
.Y(n_360)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_360),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_301),
.B(n_252),
.Y(n_361)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_323),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_363),
.B(n_372),
.Y(n_394)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_307),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_364),
.B(n_365),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_320),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_312),
.B(n_252),
.Y(n_366)
);

AND2x6_ASAP7_75t_L g367 ( 
.A(n_290),
.B(n_313),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_316),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_368),
.Y(n_405)
);

BUFx6f_ASAP7_75t_L g369 ( 
.A(n_324),
.Y(n_369)
);

INVx8_ASAP7_75t_L g370 ( 
.A(n_324),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_SL g371 ( 
.A(n_287),
.B(n_289),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_325),
.B(n_279),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_308),
.B(n_309),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_374),
.Y(n_386)
);

INVx13_ASAP7_75t_L g375 ( 
.A(n_297),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_375),
.Y(n_391)
);

INVx6_ASAP7_75t_L g377 ( 
.A(n_334),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_SL g379 ( 
.A1(n_372),
.A2(n_279),
.B1(n_294),
.B2(n_326),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_379),
.B(n_397),
.Y(n_429)
);

NAND2x1_ASAP7_75t_SL g380 ( 
.A(n_345),
.B(n_323),
.Y(n_380)
);

AND2x2_ASAP7_75t_L g431 ( 
.A(n_380),
.B(n_355),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_SL g381 ( 
.A(n_338),
.B(n_330),
.Y(n_381)
);

XOR2x2_ASAP7_75t_L g417 ( 
.A(n_381),
.B(n_357),
.Y(n_417)
);

AOI21xp5_ASAP7_75t_SL g382 ( 
.A1(n_347),
.A2(n_315),
.B(n_292),
.Y(n_382)
);

INVxp67_ASAP7_75t_L g423 ( 
.A(n_382),
.Y(n_423)
);

INVxp67_ASAP7_75t_L g435 ( 
.A(n_385),
.Y(n_435)
);

AND2x6_ASAP7_75t_L g428 ( 
.A(n_389),
.B(n_357),
.Y(n_428)
);

BUFx2_ASAP7_75t_L g420 ( 
.A(n_390),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_393),
.B(n_413),
.C(n_414),
.Y(n_418)
);

OAI22xp33_ASAP7_75t_SL g397 ( 
.A1(n_343),
.A2(n_334),
.B1(n_305),
.B2(n_295),
.Y(n_397)
);

OAI21xp5_ASAP7_75t_SL g398 ( 
.A1(n_347),
.A2(n_376),
.B(n_343),
.Y(n_398)
);

OR2x2_ASAP7_75t_L g439 ( 
.A(n_398),
.B(n_415),
.Y(n_439)
);

AO22x1_ASAP7_75t_SL g403 ( 
.A1(n_347),
.A2(n_367),
.B1(n_337),
.B2(n_378),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_403),
.B(n_411),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_344),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_404),
.B(n_406),
.Y(n_419)
);

FAx1_ASAP7_75t_SL g406 ( 
.A(n_335),
.B(n_317),
.CI(n_310),
.CON(n_406),
.SN(n_406)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_337),
.A2(n_357),
.B1(n_335),
.B2(n_359),
.Y(n_411)
);

FAx1_ASAP7_75t_SL g412 ( 
.A(n_353),
.B(n_306),
.CI(n_282),
.CON(n_412),
.SN(n_412)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_412),
.B(n_378),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_L g413 ( 
.A(n_352),
.B(n_281),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_350),
.B(n_281),
.C(n_282),
.Y(n_414)
);

OAI21xp5_ASAP7_75t_SL g415 ( 
.A1(n_361),
.A2(n_329),
.B(n_304),
.Y(n_415)
);

CKINVDCx14_ASAP7_75t_R g416 ( 
.A(n_396),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_416),
.B(n_428),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_L g466 ( 
.A(n_417),
.B(n_380),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_SL g421 ( 
.A(n_386),
.B(n_348),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_SL g467 ( 
.A(n_421),
.B(n_427),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_L g450 ( 
.A1(n_422),
.A2(n_449),
.B1(n_384),
.B2(n_394),
.Y(n_450)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_408),
.Y(n_424)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_424),
.Y(n_477)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_408),
.Y(n_425)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_425),
.Y(n_452)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_399),
.Y(n_426)
);

INVx1_ASAP7_75t_SL g478 ( 
.A(n_426),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_405),
.B(n_288),
.Y(n_427)
);

AND2x2_ASAP7_75t_L g472 ( 
.A(n_431),
.B(n_442),
.Y(n_472)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_407),
.Y(n_432)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_432),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_393),
.B(n_363),
.C(n_378),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_433),
.B(n_379),
.C(n_414),
.Y(n_453)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_401),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_434),
.B(n_438),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g436 ( 
.A(n_386),
.B(n_339),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_SL g469 ( 
.A(n_436),
.B(n_437),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_395),
.B(n_288),
.Y(n_437)
);

AND2x6_ASAP7_75t_L g438 ( 
.A(n_389),
.B(n_375),
.Y(n_438)
);

AND2x2_ASAP7_75t_L g440 ( 
.A(n_398),
.B(n_356),
.Y(n_440)
);

INVxp67_ASAP7_75t_L g463 ( 
.A(n_440),
.Y(n_463)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_407),
.Y(n_441)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_441),
.Y(n_468)
);

INVx4_ASAP7_75t_SL g442 ( 
.A(n_383),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_392),
.Y(n_443)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_443),
.Y(n_470)
);

OR2x2_ASAP7_75t_L g444 ( 
.A(n_411),
.B(n_295),
.Y(n_444)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_444),
.Y(n_471)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_392),
.Y(n_445)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_445),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_406),
.B(n_369),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_SL g479 ( 
.A(n_446),
.B(n_448),
.Y(n_479)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_388),
.Y(n_447)
);

INVx2_ASAP7_75t_SL g461 ( 
.A(n_447),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_406),
.B(n_302),
.Y(n_448)
);

CKINVDCx14_ASAP7_75t_R g449 ( 
.A(n_384),
.Y(n_449)
);

OR2x2_ASAP7_75t_L g480 ( 
.A(n_450),
.B(n_456),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_453),
.B(n_457),
.C(n_476),
.Y(n_487)
);

AOI22xp5_ASAP7_75t_L g454 ( 
.A1(n_420),
.A2(n_394),
.B1(n_412),
.B2(n_403),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_SL g493 ( 
.A1(n_454),
.A2(n_444),
.B1(n_439),
.B2(n_429),
.Y(n_493)
);

OAI21xp33_ASAP7_75t_L g456 ( 
.A1(n_434),
.A2(n_409),
.B(n_387),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_418),
.B(n_381),
.C(n_413),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g459 ( 
.A(n_442),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_459),
.B(n_462),
.Y(n_502)
);

XNOR2xp5_ASAP7_75t_SL g460 ( 
.A(n_418),
.B(n_417),
.Y(n_460)
);

XNOR2xp5_ASAP7_75t_SL g497 ( 
.A(n_460),
.B(n_466),
.Y(n_497)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_442),
.Y(n_462)
);

XOR2xp5_ASAP7_75t_L g464 ( 
.A(n_433),
.B(n_387),
.Y(n_464)
);

XOR2xp5_ASAP7_75t_L g481 ( 
.A(n_464),
.B(n_430),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_443),
.B(n_415),
.Y(n_465)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_465),
.Y(n_499)
);

OAI21xp5_ASAP7_75t_L g474 ( 
.A1(n_435),
.A2(n_385),
.B(n_380),
.Y(n_474)
);

INVxp67_ASAP7_75t_L g485 ( 
.A(n_474),
.Y(n_485)
);

OAI21xp5_ASAP7_75t_L g475 ( 
.A1(n_435),
.A2(n_382),
.B(n_403),
.Y(n_475)
);

OAI21xp5_ASAP7_75t_L g490 ( 
.A1(n_475),
.A2(n_439),
.B(n_423),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_431),
.B(n_412),
.C(n_400),
.Y(n_476)
);

XOR2xp5_ASAP7_75t_L g512 ( 
.A(n_481),
.B(n_483),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_461),
.B(n_445),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g516 ( 
.A(n_482),
.Y(n_516)
);

XOR2xp5_ASAP7_75t_L g483 ( 
.A(n_464),
.B(n_430),
.Y(n_483)
);

AOI22xp5_ASAP7_75t_SL g484 ( 
.A1(n_476),
.A2(n_423),
.B1(n_431),
.B2(n_429),
.Y(n_484)
);

OAI22xp5_ASAP7_75t_SL g513 ( 
.A1(n_484),
.A2(n_501),
.B1(n_505),
.B2(n_463),
.Y(n_513)
);

CKINVDCx20_ASAP7_75t_R g486 ( 
.A(n_472),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_486),
.B(n_488),
.Y(n_510)
);

CKINVDCx16_ASAP7_75t_R g488 ( 
.A(n_469),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_460),
.B(n_440),
.C(n_444),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_489),
.B(n_495),
.C(n_496),
.Y(n_507)
);

AOI21xp5_ASAP7_75t_L g515 ( 
.A1(n_490),
.A2(n_458),
.B(n_470),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_461),
.B(n_441),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_491),
.B(n_498),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_SL g492 ( 
.A(n_467),
.B(n_421),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_SL g527 ( 
.A(n_492),
.B(n_494),
.Y(n_527)
);

AOI22xp5_ASAP7_75t_SL g514 ( 
.A1(n_493),
.A2(n_503),
.B1(n_463),
.B2(n_465),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_SL g494 ( 
.A(n_451),
.B(n_419),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_457),
.B(n_440),
.C(n_439),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_453),
.B(n_432),
.C(n_447),
.Y(n_496)
);

CKINVDCx16_ASAP7_75t_R g498 ( 
.A(n_472),
.Y(n_498)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_455),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_500),
.B(n_504),
.Y(n_525)
);

AOI22xp5_ASAP7_75t_SL g501 ( 
.A1(n_471),
.A2(n_420),
.B1(n_362),
.B2(n_438),
.Y(n_501)
);

OAI22xp5_ASAP7_75t_SL g503 ( 
.A1(n_454),
.A2(n_420),
.B1(n_428),
.B2(n_410),
.Y(n_503)
);

CKINVDCx20_ASAP7_75t_R g504 ( 
.A(n_472),
.Y(n_504)
);

AOI22xp5_ASAP7_75t_SL g505 ( 
.A1(n_471),
.A2(n_426),
.B1(n_400),
.B2(n_424),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_496),
.B(n_479),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_SL g533 ( 
.A(n_506),
.B(n_521),
.Y(n_533)
);

INVxp33_ASAP7_75t_L g508 ( 
.A(n_502),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_508),
.B(n_523),
.Y(n_530)
);

MAJIxp5_ASAP7_75t_L g509 ( 
.A(n_487),
.B(n_466),
.C(n_474),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_SL g528 ( 
.A(n_509),
.B(n_519),
.Y(n_528)
);

XNOR2xp5_ASAP7_75t_L g511 ( 
.A(n_487),
.B(n_475),
.Y(n_511)
);

XOR2xp5_ASAP7_75t_L g531 ( 
.A(n_511),
.B(n_513),
.Y(n_531)
);

OAI22xp5_ASAP7_75t_L g529 ( 
.A1(n_514),
.A2(n_501),
.B1(n_485),
.B2(n_505),
.Y(n_529)
);

OAI21xp5_ASAP7_75t_SL g534 ( 
.A1(n_515),
.A2(n_485),
.B(n_480),
.Y(n_534)
);

XNOR2xp5_ASAP7_75t_L g517 ( 
.A(n_495),
.B(n_489),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g542 ( 
.A(n_517),
.B(n_520),
.C(n_522),
.Y(n_542)
);

XNOR2xp5_ASAP7_75t_L g519 ( 
.A(n_481),
.B(n_458),
.Y(n_519)
);

XNOR2xp5_ASAP7_75t_L g520 ( 
.A(n_483),
.B(n_461),
.Y(n_520)
);

CKINVDCx16_ASAP7_75t_R g521 ( 
.A(n_482),
.Y(n_521)
);

XOR2xp5_ASAP7_75t_L g522 ( 
.A(n_497),
.B(n_473),
.Y(n_522)
);

XOR2xp5_ASAP7_75t_L g523 ( 
.A(n_497),
.B(n_473),
.Y(n_523)
);

XOR2xp5_ASAP7_75t_L g524 ( 
.A(n_484),
.B(n_470),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_524),
.B(n_468),
.Y(n_540)
);

XNOR2xp5_ASAP7_75t_SL g526 ( 
.A(n_493),
.B(n_499),
.Y(n_526)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_526),
.Y(n_535)
);

XOR2xp5_ASAP7_75t_L g549 ( 
.A(n_529),
.B(n_512),
.Y(n_549)
);

OAI321xp33_ASAP7_75t_L g532 ( 
.A1(n_510),
.A2(n_499),
.A3(n_491),
.B1(n_480),
.B2(n_500),
.C(n_503),
.Y(n_532)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_532),
.Y(n_559)
);

AOI21xp5_ASAP7_75t_L g560 ( 
.A1(n_534),
.A2(n_543),
.B(n_545),
.Y(n_560)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_518),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_536),
.B(n_537),
.Y(n_556)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_525),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_526),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_L g551 ( 
.A(n_538),
.B(n_383),
.Y(n_551)
);

AOI22xp5_ASAP7_75t_L g539 ( 
.A1(n_516),
.A2(n_490),
.B1(n_478),
.B2(n_455),
.Y(n_539)
);

OAI22xp5_ASAP7_75t_L g555 ( 
.A1(n_539),
.A2(n_544),
.B1(n_404),
.B2(n_391),
.Y(n_555)
);

XNOR2xp5_ASAP7_75t_L g547 ( 
.A(n_540),
.B(n_512),
.Y(n_547)
);

CKINVDCx16_ASAP7_75t_R g541 ( 
.A(n_514),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_SL g553 ( 
.A(n_541),
.B(n_452),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_508),
.B(n_478),
.Y(n_543)
);

AOI22xp5_ASAP7_75t_L g544 ( 
.A1(n_524),
.A2(n_523),
.B1(n_522),
.B2(n_507),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_520),
.B(n_468),
.Y(n_545)
);

FAx1_ASAP7_75t_SL g546 ( 
.A(n_540),
.B(n_509),
.CI(n_507),
.CON(n_546),
.SN(n_546)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_546),
.B(n_548),
.Y(n_567)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_547),
.Y(n_563)
);

MAJIxp5_ASAP7_75t_L g548 ( 
.A(n_542),
.B(n_517),
.C(n_511),
.Y(n_548)
);

XNOR2xp5_ASAP7_75t_L g566 ( 
.A(n_549),
.B(n_553),
.Y(n_566)
);

MAJIxp5_ASAP7_75t_L g550 ( 
.A(n_542),
.B(n_388),
.C(n_402),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_550),
.B(n_551),
.Y(n_569)
);

NOR2xp33_ASAP7_75t_L g552 ( 
.A(n_533),
.B(n_527),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_SL g571 ( 
.A(n_552),
.B(n_554),
.Y(n_571)
);

NOR2xp33_ASAP7_75t_L g554 ( 
.A(n_537),
.B(n_399),
.Y(n_554)
);

XOR2xp5_ASAP7_75t_L g564 ( 
.A(n_555),
.B(n_543),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_SL g557 ( 
.A(n_528),
.B(n_391),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_L g562 ( 
.A(n_557),
.B(n_530),
.Y(n_562)
);

MAJIxp5_ASAP7_75t_L g558 ( 
.A(n_531),
.B(n_402),
.C(n_452),
.Y(n_558)
);

MAJIxp5_ASAP7_75t_L g565 ( 
.A(n_558),
.B(n_550),
.C(n_548),
.Y(n_565)
);

OAI21xp5_ASAP7_75t_L g561 ( 
.A1(n_559),
.A2(n_534),
.B(n_535),
.Y(n_561)
);

NOR3xp33_ASAP7_75t_L g576 ( 
.A(n_561),
.B(n_538),
.C(n_535),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_562),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_564),
.B(n_565),
.Y(n_574)
);

OAI21xp5_ASAP7_75t_SL g568 ( 
.A1(n_560),
.A2(n_530),
.B(n_544),
.Y(n_568)
);

AOI21xp5_ASAP7_75t_L g572 ( 
.A1(n_568),
.A2(n_570),
.B(n_558),
.Y(n_572)
);

AOI21xp5_ASAP7_75t_L g570 ( 
.A1(n_556),
.A2(n_539),
.B(n_536),
.Y(n_570)
);

OAI21xp5_ASAP7_75t_L g582 ( 
.A1(n_572),
.A2(n_576),
.B(n_570),
.Y(n_582)
);

AND2x2_ASAP7_75t_L g573 ( 
.A(n_567),
.B(n_549),
.Y(n_573)
);

AOI21xp5_ASAP7_75t_L g584 ( 
.A1(n_573),
.A2(n_575),
.B(n_569),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_L g575 ( 
.A(n_571),
.B(n_546),
.Y(n_575)
);

AOI22xp5_ASAP7_75t_SL g578 ( 
.A1(n_563),
.A2(n_546),
.B1(n_545),
.B2(n_531),
.Y(n_578)
);

XNOR2xp5_ASAP7_75t_L g580 ( 
.A(n_578),
.B(n_561),
.Y(n_580)
);

INVx6_ASAP7_75t_L g579 ( 
.A(n_565),
.Y(n_579)
);

NOR2xp33_ASAP7_75t_L g581 ( 
.A(n_579),
.B(n_566),
.Y(n_581)
);

AOI21xp5_ASAP7_75t_L g588 ( 
.A1(n_580),
.A2(n_582),
.B(n_584),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_SL g586 ( 
.A(n_581),
.B(n_583),
.Y(n_586)
);

XNOR2xp5_ASAP7_75t_L g583 ( 
.A(n_574),
.B(n_566),
.Y(n_583)
);

OAI21xp5_ASAP7_75t_SL g585 ( 
.A1(n_575),
.A2(n_564),
.B(n_547),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_SL g587 ( 
.A(n_585),
.B(n_577),
.Y(n_587)
);

OAI22xp5_ASAP7_75t_L g589 ( 
.A1(n_587),
.A2(n_581),
.B1(n_586),
.B2(n_588),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_589),
.B(n_590),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_L g590 ( 
.A(n_587),
.B(n_477),
.Y(n_590)
);

A2O1A1O1Ixp25_ASAP7_75t_L g592 ( 
.A1(n_591),
.A2(n_425),
.B(n_340),
.C(n_370),
.D(n_377),
.Y(n_592)
);

FAx1_ASAP7_75t_SL g593 ( 
.A(n_592),
.B(n_340),
.CI(n_351),
.CON(n_593),
.SN(n_593)
);

AOI332xp33_ASAP7_75t_L g594 ( 
.A1(n_593),
.A2(n_302),
.A3(n_303),
.B1(n_304),
.B2(n_305),
.B3(n_306),
.C1(n_341),
.C2(n_587),
.Y(n_594)
);

BUFx24_ASAP7_75t_SL g595 ( 
.A(n_594),
.Y(n_595)
);


endmodule