module real_jpeg_15143_n_17 (n_8, n_0, n_2, n_69, n_10, n_9, n_12, n_68, n_6, n_11, n_14, n_7, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_17);

input n_8;
input n_0;
input n_2;
input n_69;
input n_10;
input n_9;
input n_12;
input n_68;
input n_6;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_17;

wire n_43;
wire n_54;
wire n_57;
wire n_21;
wire n_37;
wire n_65;
wire n_33;
wire n_38;
wire n_50;
wire n_35;
wire n_29;
wire n_55;
wire n_49;
wire n_52;
wire n_58;
wire n_31;
wire n_63;
wire n_24;
wire n_66;
wire n_34;
wire n_44;
wire n_60;
wire n_28;
wire n_46;
wire n_62;
wire n_59;
wire n_64;
wire n_23;
wire n_51;
wire n_47;
wire n_45;
wire n_25;
wire n_61;
wire n_42;
wire n_53;
wire n_18;
wire n_22;
wire n_40;
wire n_39;
wire n_36;
wire n_41;
wire n_27;
wire n_56;
wire n_20;
wire n_19;
wire n_48;
wire n_26;
wire n_30;
wire n_32;

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_0),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_0),
.B(n_63),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_1),
.B(n_52),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_1),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_2),
.B(n_7),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_2),
.B(n_7),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_3),
.B(n_15),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_3),
.B(n_15),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_4),
.B(n_8),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_4),
.B(n_8),
.Y(n_48)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_9),
.B(n_12),
.C(n_25),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_10),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_11),
.B(n_69),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_13),
.A2(n_50),
.B1(n_53),
.B2(n_54),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_13),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_13),
.B(n_60),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_14),
.B(n_51),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_14),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_SL g26 ( 
.A1(n_16),
.A2(n_27),
.B(n_30),
.Y(n_26)
);

AOI221xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_49),
.B1(n_55),
.B2(n_58),
.C(n_66),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_SL g18 ( 
.A1(n_19),
.A2(n_43),
.B1(n_44),
.B2(n_48),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_19),
.A2(n_44),
.B1(n_56),
.B2(n_57),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_22),
.B1(n_33),
.B2(n_41),
.Y(n_19)
);

CKINVDCx16_ASAP7_75t_R g20 ( 
.A(n_21),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_21),
.A2(n_33),
.B1(n_42),
.B2(n_45),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_37),
.B1(n_38),
.B2(n_40),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_23),
.A2(n_38),
.B1(n_46),
.B2(n_47),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_33),
.Y(n_23)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_31),
.C(n_32),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_29),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_28),
.B(n_29),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_33),
.B(n_39),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_33),
.B(n_63),
.Y(n_66)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx16f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_43),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_48),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_50),
.Y(n_54)
);

OAI21xp33_ASAP7_75t_L g58 ( 
.A1(n_53),
.A2(n_59),
.B(n_64),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_62),
.Y(n_60)
);

INVxp33_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_68),
.Y(n_28)
);


endmodule