module real_aes_8437_n_382 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_357, n_64, n_254, n_207, n_10, n_83, n_181, n_362, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_355, n_239, n_100, n_54, n_112, n_319, n_364, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_376, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_353, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_379, n_374, n_26, n_235, n_378, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_356, n_184, n_28, n_372, n_202, n_56, n_370, n_34, n_98, n_121, n_352, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_369, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_381, n_311, n_324, n_25, n_278, n_236, n_367, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_363, n_323, n_199, n_350, n_142, n_223, n_67, n_368, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_360, n_58, n_165, n_361, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_351, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_366, n_346, n_193, n_293, n_162, n_358, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_377, n_273, n_114, n_276, n_295, n_265, n_354, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_373, n_60, n_233, n_290, n_365, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_359, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_371, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_375, n_340, n_13, n_380, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_382);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_357;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_362;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_355;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_364;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_376;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_353;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_379;
input n_374;
input n_26;
input n_235;
input n_378;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_356;
input n_184;
input n_28;
input n_372;
input n_202;
input n_56;
input n_370;
input n_34;
input n_98;
input n_121;
input n_352;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_369;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_381;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_367;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_363;
input n_323;
input n_199;
input n_350;
input n_142;
input n_223;
input n_67;
input n_368;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_360;
input n_58;
input n_165;
input n_361;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_351;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_366;
input n_346;
input n_193;
input n_293;
input n_162;
input n_358;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_377;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_354;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_373;
input n_60;
input n_233;
input n_290;
input n_365;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_359;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_371;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_375;
input n_340;
input n_13;
input n_380;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_382;
wire n_480;
wire n_1073;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_887;
wire n_684;
wire n_1066;
wire n_390;
wire n_1096;
wire n_821;
wire n_830;
wire n_624;
wire n_1018;
wire n_980;
wire n_618;
wire n_778;
wire n_800;
wire n_1106;
wire n_522;
wire n_1092;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_943;
wire n_977;
wire n_503;
wire n_635;
wire n_673;
wire n_386;
wire n_792;
wire n_518;
wire n_905;
wire n_1067;
wire n_878;
wire n_665;
wire n_667;
wire n_991;
wire n_1114;
wire n_577;
wire n_580;
wire n_1004;
wire n_469;
wire n_987;
wire n_979;
wire n_759;
wire n_445;
wire n_1065;
wire n_596;
wire n_592;
wire n_540;
wire n_1064;
wire n_1075;
wire n_657;
wire n_900;
wire n_718;
wire n_841;
wire n_669;
wire n_1091;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_1014;
wire n_421;
wire n_555;
wire n_766;
wire n_852;
wire n_1113;
wire n_974;
wire n_857;
wire n_1089;
wire n_919;
wire n_1122;
wire n_461;
wire n_1047;
wire n_1016;
wire n_908;
wire n_571;
wire n_1123;
wire n_549;
wire n_491;
wire n_694;
wire n_894;
wire n_923;
wire n_1034;
wire n_952;
wire n_429;
wire n_1110;
wire n_752;
wire n_448;
wire n_556;
wire n_545;
wire n_593;
wire n_460;
wire n_742;
wire n_937;
wire n_773;
wire n_989;
wire n_401;
wire n_538;
wire n_431;
wire n_1044;
wire n_963;
wire n_865;
wire n_537;
wire n_666;
wire n_551;
wire n_884;
wire n_560;
wire n_660;
wire n_1094;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_983;
wire n_767;
wire n_696;
wire n_955;
wire n_889;
wire n_975;
wire n_704;
wire n_941;
wire n_453;
wire n_932;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_1046;
wire n_677;
wire n_958;
wire n_1021;
wire n_591;
wire n_775;
wire n_763;
wire n_1093;
wire n_1109;
wire n_870;
wire n_961;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_415;
wire n_572;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_1116;
wire n_573;
wire n_510;
wire n_1099;
wire n_709;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_626;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_953;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_550;
wire n_966;
wire n_1108;
wire n_670;
wire n_818;
wire n_716;
wire n_918;
wire n_478;
wire n_883;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_578;
wire n_528;
wire n_892;
wire n_495;
wire n_994;
wire n_1078;
wire n_1072;
wire n_384;
wire n_744;
wire n_938;
wire n_935;
wire n_1098;
wire n_824;
wire n_467;
wire n_875;
wire n_951;
wire n_774;
wire n_992;
wire n_813;
wire n_791;
wire n_981;
wire n_559;
wire n_976;
wire n_636;
wire n_1053;
wire n_1049;
wire n_466;
wire n_872;
wire n_477;
wire n_906;
wire n_515;
wire n_984;
wire n_1019;
wire n_680;
wire n_595;
wire n_1086;
wire n_726;
wire n_1070;
wire n_517;
wire n_683;
wire n_931;
wire n_904;
wire n_780;
wire n_570;
wire n_675;
wire n_840;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_1117;
wire n_834;
wire n_882;
wire n_784;
wire n_496;
wire n_693;
wire n_962;
wire n_1082;
wire n_468;
wire n_746;
wire n_532;
wire n_656;
wire n_755;
wire n_1025;
wire n_409;
wire n_781;
wire n_748;
wire n_909;
wire n_523;
wire n_860;
wire n_996;
wire n_439;
wire n_1062;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_801;
wire n_1126;
wire n_383;
wire n_529;
wire n_1115;
wire n_504;
wire n_455;
wire n_725;
wire n_960;
wire n_1081;
wire n_671;
wire n_973;
wire n_1084;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_1029;
wire n_1020;
wire n_457;
wire n_1121;
wire n_885;
wire n_1059;
wire n_950;
wire n_993;
wire n_493;
wire n_664;
wire n_819;
wire n_737;
wire n_1013;
wire n_1017;
wire n_581;
wire n_610;
wire n_936;
wire n_1035;
wire n_620;
wire n_582;
wire n_641;
wire n_1063;
wire n_828;
wire n_808;
wire n_770;
wire n_940;
wire n_722;
wire n_745;
wire n_867;
wire n_398;
wire n_1100;
wire n_688;
wire n_425;
wire n_609;
wire n_1042;
wire n_879;
wire n_417;
wire n_1006;
wire n_607;
wire n_449;
wire n_754;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_706;
wire n_901;
wire n_561;
wire n_947;
wire n_970;
wire n_876;
wire n_437;
wire n_1112;
wire n_428;
wire n_405;
wire n_621;
wire n_783;
wire n_1107;
wire n_1012;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1054;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_1050;
wire n_426;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_658;
wire n_676;
wire n_986;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_1037;
wire n_1031;
wire n_1103;
wire n_1008;
wire n_807;
wire n_1011;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_913;
wire n_999;
wire n_619;
wire n_391;
wire n_1095;
wire n_1060;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_1080;
wire n_917;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_985;
wire n_777;
wire n_1077;
wire n_501;
wire n_1041;
wire n_488;
wire n_1111;
wire n_910;
wire n_642;
wire n_613;
wire n_869;
wire n_387;
wire n_1125;
wire n_957;
wire n_995;
wire n_1124;
wire n_702;
wire n_954;
wire n_969;
wire n_912;
wire n_1009;
wire n_1007;
wire n_464;
wire n_945;
wire n_604;
wire n_734;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_1022;
wire n_404;
wire n_598;
wire n_756;
wire n_713;
wire n_735;
wire n_728;
wire n_569;
wire n_997;
wire n_785;
wire n_563;
wire n_891;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_1105;
wire n_853;
wire n_810;
wire n_1079;
wire n_843;
wire n_579;
wire n_1033;
wire n_699;
wire n_533;
wire n_1000;
wire n_1003;
wire n_1028;
wire n_727;
wire n_1083;
wire n_397;
wire n_385;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_536;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_915;
wire n_1002;
wire n_934;
wire n_494;
wire n_1001;
wire n_711;
wire n_864;
wire n_1027;
wire n_1058;
wire n_927;
wire n_1038;
wire n_965;
wire n_723;
wire n_662;
wire n_1085;
wire n_845;
wire n_1043;
wire n_850;
wire n_720;
wire n_968;
wire n_972;
wire n_435;
wire n_1127;
wire n_1026;
wire n_511;
wire n_484;
wire n_893;
wire n_492;
wire n_1068;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_1023;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_1057;
wire n_411;
wire n_697;
wire n_978;
wire n_847;
wire n_907;
wire n_779;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_648;
wire n_589;
wire n_628;
wire n_939;
wire n_1005;
wire n_487;
wire n_831;
wire n_653;
wire n_637;
wire n_526;
wire n_899;
wire n_928;
wire n_692;
wire n_544;
wire n_789;
wire n_1087;
wire n_1051;
wire n_389;
wire n_738;
wire n_701;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_926;
wire n_922;
wire n_942;
wire n_1048;
wire n_472;
wire n_1120;
wire n_971;
wire n_866;
wire n_452;
wire n_1071;
wire n_787;
wire n_1052;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_1097;
wire n_715;
wire n_959;
wire n_946;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_741;
wire n_753;
wire n_623;
wire n_1032;
wire n_446;
wire n_721;
wire n_681;
wire n_982;
wire n_456;
wire n_717;
wire n_1090;
wire n_712;
wire n_433;
wire n_516;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_575;
wire n_762;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_740;
wire n_541;
wire n_839;
wire n_639;
wire n_546;
wire n_587;
wire n_1010;
wire n_811;
wire n_1015;
wire n_459;
wire n_558;
wire n_863;
wire n_998;
wire n_724;
wire n_440;
wire n_525;
wire n_1074;
wire n_644;
wire n_674;
wire n_836;
wire n_888;
wire n_793;
wire n_1056;
wire n_583;
wire n_833;
wire n_414;
wire n_757;
wire n_929;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_949;
wire n_614;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_719;
wire n_465;
wire n_473;
wire n_566;
wire n_1045;
wire n_837;
wire n_967;
wire n_871;
wire n_474;
wire n_829;
wire n_1030;
wire n_988;
wire n_1055;
wire n_1088;
wire n_921;
wire n_597;
wire n_640;
wire n_483;
wire n_611;
wire n_1036;
wire n_394;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_710;
wire n_650;
wire n_743;
wire n_823;
wire n_393;
wire n_1040;
wire n_652;
wire n_703;
wire n_601;
wire n_500;
wire n_1102;
wire n_661;
wire n_1076;
wire n_463;
wire n_396;
wire n_804;
wire n_1101;
wire n_447;
wire n_603;
wire n_403;
wire n_854;
wire n_1119;
wire n_424;
wire n_802;
wire n_868;
wire n_877;
wire n_1039;
wire n_574;
wire n_1069;
wire n_1024;
wire n_842;
wire n_1104;
wire n_849;
wire n_1061;
wire n_475;
wire n_554;
wire n_897;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
AOI22xp33_ASAP7_75t_L g600 ( .A1(n_0), .A2(n_190), .B1(n_477), .B2(n_601), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g967 ( .A(n_1), .B(n_593), .Y(n_967) );
INVx1_ASAP7_75t_L g1024 ( .A(n_2), .Y(n_1024) );
AOI22xp33_ASAP7_75t_SL g643 ( .A1(n_3), .A2(n_243), .B1(n_608), .B2(n_644), .Y(n_643) );
AOI222xp33_ASAP7_75t_L g784 ( .A1(n_4), .A2(n_183), .B1(n_340), .B2(n_427), .C1(n_561), .C2(n_785), .Y(n_784) );
AOI22xp33_ASAP7_75t_L g656 ( .A1(n_5), .A2(n_115), .B1(n_533), .B2(n_607), .Y(n_656) );
AOI22xp33_ASAP7_75t_SL g802 ( .A1(n_6), .A2(n_166), .B1(n_571), .B2(n_803), .Y(n_802) );
AOI22xp33_ASAP7_75t_L g753 ( .A1(n_7), .A2(n_236), .B1(n_610), .B2(n_639), .Y(n_753) );
NAND2xp5_ASAP7_75t_SL g797 ( .A(n_8), .B(n_798), .Y(n_797) );
AO22x2_ASAP7_75t_L g409 ( .A1(n_9), .A2(n_224), .B1(n_410), .B2(n_411), .Y(n_409) );
INVx1_ASAP7_75t_L g1061 ( .A(n_9), .Y(n_1061) );
CKINVDCx20_ASAP7_75t_R g819 ( .A(n_10), .Y(n_819) );
AOI22xp33_ASAP7_75t_L g776 ( .A1(n_11), .A2(n_175), .B1(n_481), .B2(n_719), .Y(n_776) );
AOI22xp33_ASAP7_75t_SL g881 ( .A1(n_12), .A2(n_363), .B1(n_436), .B2(n_783), .Y(n_881) );
CKINVDCx20_ASAP7_75t_R g763 ( .A(n_13), .Y(n_763) );
AOI22xp5_ASAP7_75t_L g567 ( .A1(n_14), .A2(n_163), .B1(n_535), .B2(n_568), .Y(n_567) );
INVx1_ASAP7_75t_L g979 ( .A(n_15), .Y(n_979) );
AOI22xp33_ASAP7_75t_L g935 ( .A1(n_16), .A2(n_197), .B1(n_516), .B2(n_519), .Y(n_935) );
AOI22xp33_ASAP7_75t_L g874 ( .A1(n_17), .A2(n_254), .B1(n_535), .B2(n_731), .Y(n_874) );
AOI22xp33_ASAP7_75t_L g660 ( .A1(n_18), .A2(n_328), .B1(n_486), .B2(n_661), .Y(n_660) );
CKINVDCx20_ASAP7_75t_R g1081 ( .A(n_19), .Y(n_1081) );
AOI22xp33_ASAP7_75t_L g492 ( .A1(n_20), .A2(n_230), .B1(n_493), .B2(n_497), .Y(n_492) );
AOI222xp33_ASAP7_75t_L g733 ( .A1(n_21), .A2(n_71), .B1(n_288), .B2(n_436), .C1(n_559), .C2(n_734), .Y(n_733) );
AOI22xp33_ASAP7_75t_SL g541 ( .A1(n_22), .A2(n_315), .B1(n_470), .B2(n_490), .Y(n_541) );
CKINVDCx20_ASAP7_75t_R g830 ( .A(n_23), .Y(n_830) );
AOI22xp5_ASAP7_75t_SL g869 ( .A1(n_24), .A2(n_251), .B1(n_568), .B2(n_870), .Y(n_869) );
CKINVDCx20_ASAP7_75t_R g548 ( .A(n_25), .Y(n_548) );
AOI22xp33_ASAP7_75t_SL g531 ( .A1(n_26), .A2(n_312), .B1(n_532), .B2(n_533), .Y(n_531) );
AOI22xp33_ASAP7_75t_L g647 ( .A1(n_27), .A2(n_257), .B1(n_481), .B2(n_648), .Y(n_647) );
AOI22xp33_ASAP7_75t_L g569 ( .A1(n_28), .A2(n_367), .B1(n_570), .B2(n_571), .Y(n_569) );
CKINVDCx20_ASAP7_75t_R g765 ( .A(n_29), .Y(n_765) );
AOI22xp33_ASAP7_75t_L g938 ( .A1(n_30), .A2(n_249), .B1(n_719), .B2(n_806), .Y(n_938) );
AO22x2_ASAP7_75t_L g413 ( .A1(n_31), .A2(n_130), .B1(n_410), .B2(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g420 ( .A(n_32), .Y(n_420) );
AOI22xp33_ASAP7_75t_L g942 ( .A1(n_33), .A2(n_179), .B1(n_491), .B2(n_498), .Y(n_942) );
CKINVDCx20_ASAP7_75t_R g735 ( .A(n_34), .Y(n_735) );
AOI22xp5_ASAP7_75t_L g581 ( .A1(n_35), .A2(n_582), .B1(n_611), .B2(n_612), .Y(n_581) );
INVx1_ASAP7_75t_L g612 ( .A(n_35), .Y(n_612) );
AOI22xp33_ASAP7_75t_L g1084 ( .A1(n_36), .A2(n_63), .B1(n_464), .B2(n_806), .Y(n_1084) );
AOI22xp33_ASAP7_75t_SL g941 ( .A1(n_37), .A2(n_65), .B1(n_481), .B2(n_494), .Y(n_941) );
AOI22xp33_ASAP7_75t_L g962 ( .A1(n_38), .A2(n_70), .B1(n_803), .B2(n_963), .Y(n_962) );
INVx1_ASAP7_75t_L g1003 ( .A(n_39), .Y(n_1003) );
AOI22xp5_ASAP7_75t_L g931 ( .A1(n_40), .A2(n_298), .B1(n_561), .B2(n_932), .Y(n_931) );
CKINVDCx20_ASAP7_75t_R g814 ( .A(n_41), .Y(n_814) );
AOI22xp5_ASAP7_75t_L g1031 ( .A1(n_42), .A2(n_66), .B1(n_483), .B2(n_573), .Y(n_1031) );
AOI22xp33_ASAP7_75t_L g899 ( .A1(n_43), .A2(n_169), .B1(n_577), .B2(n_719), .Y(n_899) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_44), .B(n_704), .Y(n_703) );
AOI22xp33_ASAP7_75t_L g606 ( .A1(n_45), .A2(n_308), .B1(n_607), .B2(n_608), .Y(n_606) );
AOI22xp33_ASAP7_75t_L g682 ( .A1(n_46), .A2(n_135), .B1(n_658), .B2(n_683), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_47), .B(n_516), .Y(n_702) );
INVx1_ASAP7_75t_L g895 ( .A(n_48), .Y(n_895) );
AOI22xp33_ASAP7_75t_L g924 ( .A1(n_49), .A2(n_369), .B1(n_528), .B2(n_596), .Y(n_924) );
CKINVDCx20_ASAP7_75t_R g820 ( .A(n_50), .Y(n_820) );
AOI22xp5_ASAP7_75t_L g1001 ( .A1(n_51), .A2(n_212), .B1(n_446), .B2(n_529), .Y(n_1001) );
AOI22xp33_ASAP7_75t_L g817 ( .A1(n_52), .A2(n_329), .B1(n_672), .B2(n_700), .Y(n_817) );
AOI222xp33_ASAP7_75t_L g671 ( .A1(n_53), .A2(n_306), .B1(n_327), .B2(n_556), .C1(n_590), .C2(n_672), .Y(n_671) );
AOI22xp5_ASAP7_75t_SL g867 ( .A1(n_54), .A2(n_322), .B1(n_721), .B2(n_868), .Y(n_867) );
AOI22xp33_ASAP7_75t_L g923 ( .A1(n_55), .A2(n_305), .B1(n_781), .B2(n_891), .Y(n_923) );
CKINVDCx20_ASAP7_75t_R g686 ( .A(n_56), .Y(n_686) );
CKINVDCx20_ASAP7_75t_R g786 ( .A(n_57), .Y(n_786) );
AOI22xp33_ASAP7_75t_L g745 ( .A1(n_58), .A2(n_131), .B1(n_464), .B2(n_746), .Y(n_745) );
AOI222xp33_ASAP7_75t_L g1122 ( .A1(n_59), .A2(n_180), .B1(n_351), .B2(n_428), .C1(n_558), .C2(n_1123), .Y(n_1122) );
AOI22xp5_ASAP7_75t_SL g1030 ( .A1(n_60), .A2(n_222), .B1(n_535), .B2(n_868), .Y(n_1030) );
AOI22xp33_ASAP7_75t_SL g510 ( .A1(n_61), .A2(n_85), .B1(n_434), .B2(n_511), .Y(n_510) );
INVx1_ASAP7_75t_L g985 ( .A(n_62), .Y(n_985) );
AOI22xp33_ASAP7_75t_L g725 ( .A1(n_64), .A2(n_337), .B1(n_726), .B2(n_727), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g1077 ( .A(n_67), .B(n_590), .Y(n_1077) );
CKINVDCx20_ASAP7_75t_R g943 ( .A(n_68), .Y(n_943) );
AOI22xp33_ASAP7_75t_SL g860 ( .A1(n_69), .A2(n_250), .B1(n_610), .B2(n_639), .Y(n_860) );
AOI22xp33_ASAP7_75t_L g983 ( .A1(n_72), .A2(n_276), .B1(n_511), .B2(n_528), .Y(n_983) );
AOI22xp33_ASAP7_75t_L g991 ( .A1(n_73), .A2(n_365), .B1(n_472), .B2(n_603), .Y(n_991) );
AOI22xp5_ASAP7_75t_L g896 ( .A1(n_74), .A2(n_105), .B1(n_561), .B2(n_727), .Y(n_896) );
CKINVDCx20_ASAP7_75t_R g828 ( .A(n_75), .Y(n_828) );
INVx1_ASAP7_75t_L g442 ( .A(n_76), .Y(n_442) );
AOI22xp33_ASAP7_75t_SL g801 ( .A1(n_77), .A2(n_139), .B1(n_575), .B2(n_730), .Y(n_801) );
AOI22xp33_ASAP7_75t_L g1115 ( .A1(n_78), .A2(n_345), .B1(n_644), .B2(n_859), .Y(n_1115) );
AOI22xp33_ASAP7_75t_L g476 ( .A1(n_79), .A2(n_358), .B1(n_477), .B2(n_481), .Y(n_476) );
INVx1_ASAP7_75t_L g1022 ( .A(n_80), .Y(n_1022) );
AOI22xp33_ASAP7_75t_L g1088 ( .A1(n_81), .A2(n_157), .B1(n_490), .B2(n_1089), .Y(n_1088) );
NAND2xp5_ASAP7_75t_SL g1011 ( .A(n_82), .B(n_873), .Y(n_1011) );
CKINVDCx20_ASAP7_75t_R g586 ( .A(n_83), .Y(n_586) );
AOI22xp33_ASAP7_75t_SL g638 ( .A1(n_84), .A2(n_208), .B1(n_639), .B2(n_641), .Y(n_638) );
CKINVDCx20_ASAP7_75t_R g565 ( .A(n_86), .Y(n_565) );
AOI22xp33_ASAP7_75t_L g882 ( .A1(n_87), .A2(n_221), .B1(n_517), .B2(n_519), .Y(n_882) );
INVx1_ASAP7_75t_L g628 ( .A(n_88), .Y(n_628) );
INVx1_ASAP7_75t_L g982 ( .A(n_89), .Y(n_982) );
AOI22xp33_ASAP7_75t_L g1085 ( .A1(n_90), .A2(n_108), .B1(n_648), .B2(n_1086), .Y(n_1085) );
AOI22xp33_ASAP7_75t_SL g862 ( .A1(n_91), .A2(n_227), .B1(n_722), .B2(n_863), .Y(n_862) );
AOI22xp5_ASAP7_75t_SL g1033 ( .A1(n_92), .A2(n_109), .B1(n_806), .B2(n_863), .Y(n_1033) );
CKINVDCx20_ASAP7_75t_R g1107 ( .A(n_93), .Y(n_1107) );
AO22x2_ASAP7_75t_L g417 ( .A1(n_94), .A2(n_265), .B1(n_410), .B2(n_411), .Y(n_417) );
INVx1_ASAP7_75t_L g1058 ( .A(n_94), .Y(n_1058) );
AOI22xp33_ASAP7_75t_SL g635 ( .A1(n_95), .A2(n_96), .B1(n_636), .B2(n_637), .Y(n_635) );
AOI22xp33_ASAP7_75t_L g732 ( .A1(n_97), .A2(n_275), .B1(n_498), .B2(n_570), .Y(n_732) );
AOI22xp33_ASAP7_75t_L g557 ( .A1(n_98), .A2(n_360), .B1(n_558), .B2(n_559), .Y(n_557) );
AOI22xp33_ASAP7_75t_L g576 ( .A1(n_99), .A2(n_359), .B1(n_577), .B2(n_578), .Y(n_576) );
AOI22xp33_ASAP7_75t_L g1091 ( .A1(n_100), .A2(n_375), .B1(n_963), .B2(n_1092), .Y(n_1091) );
AOI22xp33_ASAP7_75t_L g592 ( .A1(n_101), .A2(n_302), .B1(n_593), .B2(n_594), .Y(n_592) );
AOI22xp33_ASAP7_75t_L g911 ( .A1(n_102), .A2(n_377), .B1(n_912), .B2(n_913), .Y(n_911) );
AOI22xp5_ASAP7_75t_L g587 ( .A1(n_103), .A2(n_218), .B1(n_588), .B2(n_590), .Y(n_587) );
CKINVDCx20_ASAP7_75t_R g509 ( .A(n_104), .Y(n_509) );
AOI22xp33_ASAP7_75t_L g572 ( .A1(n_106), .A2(n_317), .B1(n_573), .B2(n_575), .Y(n_572) );
OA22x2_ASAP7_75t_L g652 ( .A1(n_107), .A2(n_653), .B1(n_654), .B2(n_673), .Y(n_652) );
INVx1_ASAP7_75t_L g653 ( .A(n_107), .Y(n_653) );
AOI22xp5_ASAP7_75t_L g900 ( .A1(n_110), .A2(n_126), .B1(n_730), .B2(n_806), .Y(n_900) );
AOI22xp33_ASAP7_75t_SL g1034 ( .A1(n_111), .A2(n_209), .B1(n_608), .B2(n_873), .Y(n_1034) );
CKINVDCx16_ASAP7_75t_R g1099 ( .A(n_112), .Y(n_1099) );
AOI22xp5_ASAP7_75t_L g1101 ( .A1(n_112), .A2(n_1099), .B1(n_1102), .B2(n_1124), .Y(n_1101) );
AOI22xp33_ASAP7_75t_SL g934 ( .A1(n_113), .A2(n_119), .B1(n_672), .B2(n_783), .Y(n_934) );
INVx1_ASAP7_75t_L g1027 ( .A(n_114), .Y(n_1027) );
AOI22xp33_ASAP7_75t_L g602 ( .A1(n_116), .A2(n_138), .B1(n_603), .B2(n_604), .Y(n_602) );
AOI22xp33_ASAP7_75t_L g705 ( .A1(n_117), .A2(n_355), .B1(n_523), .B2(n_528), .Y(n_705) );
AOI22xp33_ASAP7_75t_SL g851 ( .A1(n_118), .A2(n_165), .B1(n_523), .B2(n_526), .Y(n_851) );
CKINVDCx20_ASAP7_75t_R g877 ( .A(n_120), .Y(n_877) );
CKINVDCx20_ASAP7_75t_R g1010 ( .A(n_121), .Y(n_1010) );
NAND2xp5_ASAP7_75t_L g890 ( .A(n_122), .B(n_891), .Y(n_890) );
AOI22xp33_ASAP7_75t_L g485 ( .A1(n_123), .A2(n_152), .B1(n_486), .B2(n_489), .Y(n_485) );
CKINVDCx20_ASAP7_75t_R g1004 ( .A(n_124), .Y(n_1004) );
AOI22xp5_ASAP7_75t_L g993 ( .A1(n_125), .A2(n_247), .B1(n_570), .B2(n_918), .Y(n_993) );
CKINVDCx20_ASAP7_75t_R g689 ( .A(n_127), .Y(n_689) );
AOI22xp33_ASAP7_75t_L g959 ( .A1(n_128), .A2(n_286), .B1(n_608), .B2(n_637), .Y(n_959) );
XOR2xp5_ASAP7_75t_L g1064 ( .A(n_129), .B(n_1065), .Y(n_1064) );
INVx1_ASAP7_75t_L g1062 ( .A(n_130), .Y(n_1062) );
AOI22xp33_ASAP7_75t_SL g536 ( .A1(n_132), .A2(n_155), .B1(n_497), .B2(n_537), .Y(n_536) );
CKINVDCx20_ASAP7_75t_R g793 ( .A(n_133), .Y(n_793) );
CKINVDCx20_ASAP7_75t_R g750 ( .A(n_134), .Y(n_750) );
AOI22xp33_ASAP7_75t_L g903 ( .A1(n_136), .A2(n_141), .B1(n_608), .B2(n_904), .Y(n_903) );
OAI22xp5_ASAP7_75t_L g616 ( .A1(n_137), .A2(n_617), .B1(n_618), .B2(n_619), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_137), .Y(n_617) );
CKINVDCx20_ASAP7_75t_R g1119 ( .A(n_140), .Y(n_1119) );
AOI22xp33_ASAP7_75t_L g758 ( .A1(n_142), .A2(n_266), .B1(n_526), .B2(n_596), .Y(n_758) );
CKINVDCx20_ASAP7_75t_R g1037 ( .A(n_143), .Y(n_1037) );
XNOR2x2_ASAP7_75t_L g955 ( .A(n_144), .B(n_956), .Y(n_955) );
CKINVDCx20_ASAP7_75t_R g1007 ( .A(n_145), .Y(n_1007) );
AOI22xp33_ASAP7_75t_L g917 ( .A1(n_146), .A2(n_198), .B1(n_870), .B2(n_918), .Y(n_917) );
CKINVDCx20_ASAP7_75t_R g744 ( .A(n_147), .Y(n_744) );
INVx1_ASAP7_75t_L g905 ( .A(n_148), .Y(n_905) );
AOI22xp33_ASAP7_75t_L g921 ( .A1(n_149), .A2(n_196), .B1(n_639), .B2(n_641), .Y(n_921) );
AOI22xp33_ASAP7_75t_L g663 ( .A1(n_150), .A2(n_344), .B1(n_664), .B2(n_666), .Y(n_663) );
AOI22xp5_ASAP7_75t_L g939 ( .A1(n_151), .A2(n_178), .B1(n_646), .B2(n_730), .Y(n_939) );
AOI22xp5_ASAP7_75t_L g1041 ( .A1(n_153), .A2(n_264), .B1(n_511), .B2(n_528), .Y(n_1041) );
AOI22xp33_ASAP7_75t_SL g463 ( .A1(n_154), .A2(n_245), .B1(n_464), .B2(n_470), .Y(n_463) );
AOI22xp33_ASAP7_75t_L g893 ( .A1(n_156), .A2(n_364), .B1(n_436), .B2(n_783), .Y(n_893) );
AOI22xp33_ASAP7_75t_L g774 ( .A1(n_158), .A2(n_188), .B1(n_494), .B2(n_498), .Y(n_774) );
AOI22xp33_ASAP7_75t_L g1121 ( .A1(n_159), .A2(n_207), .B1(n_727), .B2(n_783), .Y(n_1121) );
AOI22xp33_ASAP7_75t_L g670 ( .A1(n_160), .A2(n_281), .B1(n_523), .B2(n_529), .Y(n_670) );
AOI22xp33_ASAP7_75t_L g609 ( .A1(n_161), .A2(n_232), .B1(n_493), .B2(n_610), .Y(n_609) );
CKINVDCx20_ASAP7_75t_R g813 ( .A(n_162), .Y(n_813) );
AND2x6_ASAP7_75t_L g385 ( .A(n_164), .B(n_386), .Y(n_385) );
HB1xp67_ASAP7_75t_L g1055 ( .A(n_164), .Y(n_1055) );
CKINVDCx20_ASAP7_75t_R g1006 ( .A(n_167), .Y(n_1006) );
CKINVDCx20_ASAP7_75t_R g1043 ( .A(n_168), .Y(n_1043) );
AOI22xp33_ASAP7_75t_SL g902 ( .A1(n_170), .A2(n_361), .B1(n_494), .B2(n_532), .Y(n_902) );
AOI22xp5_ASAP7_75t_L g879 ( .A1(n_171), .A2(n_242), .B1(n_529), .B2(n_561), .Y(n_879) );
AOI22xp33_ASAP7_75t_SL g805 ( .A1(n_172), .A2(n_376), .B1(n_719), .B2(n_806), .Y(n_805) );
CKINVDCx20_ASAP7_75t_R g808 ( .A(n_173), .Y(n_808) );
AOI222xp33_ASAP7_75t_L g925 ( .A1(n_174), .A2(n_191), .B1(n_210), .B2(n_511), .C1(n_734), .C2(n_785), .Y(n_925) );
CKINVDCx20_ASAP7_75t_R g691 ( .A(n_176), .Y(n_691) );
AOI22xp33_ASAP7_75t_L g657 ( .A1(n_177), .A2(n_273), .B1(n_537), .B2(n_658), .Y(n_657) );
CKINVDCx20_ASAP7_75t_R g831 ( .A(n_181), .Y(n_831) );
INVx1_ASAP7_75t_L g632 ( .A(n_182), .Y(n_632) );
CKINVDCx20_ASAP7_75t_R g816 ( .A(n_184), .Y(n_816) );
CKINVDCx20_ASAP7_75t_R g1079 ( .A(n_185), .Y(n_1079) );
AOI22xp33_ASAP7_75t_SL g539 ( .A1(n_186), .A2(n_272), .B1(n_486), .B2(n_540), .Y(n_539) );
AO22x2_ASAP7_75t_L g419 ( .A1(n_187), .A2(n_252), .B1(n_410), .B2(n_414), .Y(n_419) );
NOR2xp33_ASAP7_75t_L g1059 ( .A(n_187), .B(n_1060), .Y(n_1059) );
CKINVDCx20_ASAP7_75t_R g551 ( .A(n_189), .Y(n_551) );
AOI22xp33_ASAP7_75t_SL g807 ( .A1(n_192), .A2(n_271), .B1(n_568), .B2(n_721), .Y(n_807) );
AOI22xp33_ASAP7_75t_L g773 ( .A1(n_193), .A2(n_255), .B1(n_573), .B2(n_646), .Y(n_773) );
AOI22xp33_ASAP7_75t_L g848 ( .A1(n_194), .A2(n_313), .B1(n_511), .B2(n_849), .Y(n_848) );
AOI222xp33_ASAP7_75t_L g969 ( .A1(n_195), .A2(n_223), .B1(n_299), .B2(n_436), .C1(n_511), .C2(n_734), .Y(n_969) );
AOI22xp33_ASAP7_75t_L g629 ( .A1(n_199), .A2(n_381), .B1(n_436), .B2(n_511), .Y(n_629) );
INVx1_ASAP7_75t_L g622 ( .A(n_200), .Y(n_622) );
AOI22xp33_ASAP7_75t_SL g990 ( .A1(n_201), .A2(n_343), .B1(n_636), .B2(n_646), .Y(n_990) );
INVx1_ASAP7_75t_L g631 ( .A(n_202), .Y(n_631) );
AOI22xp5_ASAP7_75t_SL g872 ( .A1(n_203), .A2(n_283), .B1(n_859), .B2(n_873), .Y(n_872) );
AOI22xp33_ASAP7_75t_L g718 ( .A1(n_204), .A2(n_239), .B1(n_578), .B2(n_719), .Y(n_718) );
CKINVDCx20_ASAP7_75t_R g1069 ( .A(n_205), .Y(n_1069) );
CKINVDCx20_ASAP7_75t_R g1120 ( .A(n_206), .Y(n_1120) );
NAND2xp5_ASAP7_75t_L g780 ( .A(n_211), .B(n_781), .Y(n_780) );
CKINVDCx20_ASAP7_75t_R g756 ( .A(n_213), .Y(n_756) );
AOI22xp33_ASAP7_75t_SL g522 ( .A1(n_214), .A2(n_253), .B1(n_523), .B2(n_526), .Y(n_522) );
CKINVDCx20_ASAP7_75t_R g1075 ( .A(n_215), .Y(n_1075) );
AOI211xp5_ASAP7_75t_L g382 ( .A1(n_216), .A2(n_383), .B(n_391), .C(n_1063), .Y(n_382) );
CKINVDCx20_ASAP7_75t_R g1105 ( .A(n_217), .Y(n_1105) );
CKINVDCx20_ASAP7_75t_R g554 ( .A(n_219), .Y(n_554) );
INVx1_ASAP7_75t_L g432 ( .A(n_220), .Y(n_432) );
CKINVDCx20_ASAP7_75t_R g757 ( .A(n_225), .Y(n_757) );
CKINVDCx20_ASAP7_75t_R g742 ( .A(n_226), .Y(n_742) );
AOI22xp33_ASAP7_75t_L g595 ( .A1(n_228), .A2(n_304), .B1(n_526), .B2(n_596), .Y(n_595) );
AOI22xp33_ASAP7_75t_L g777 ( .A1(n_229), .A2(n_373), .B1(n_490), .B2(n_578), .Y(n_777) );
CKINVDCx20_ASAP7_75t_R g883 ( .A(n_231), .Y(n_883) );
CKINVDCx20_ASAP7_75t_R g1110 ( .A(n_233), .Y(n_1110) );
AOI22xp33_ASAP7_75t_L g823 ( .A1(n_234), .A2(n_303), .B1(n_472), .B2(n_664), .Y(n_823) );
XNOR2xp5_ASAP7_75t_L g504 ( .A(n_235), .B(n_505), .Y(n_504) );
CKINVDCx20_ASAP7_75t_R g698 ( .A(n_237), .Y(n_698) );
AOI22xp33_ASAP7_75t_SL g856 ( .A1(n_238), .A2(n_277), .B1(n_857), .B2(n_859), .Y(n_856) );
AOI22xp5_ASAP7_75t_SL g400 ( .A1(n_240), .A2(n_401), .B1(n_501), .B2(n_502), .Y(n_400) );
INVx1_ASAP7_75t_L g502 ( .A(n_240), .Y(n_502) );
AOI22xp33_ASAP7_75t_L g1116 ( .A1(n_241), .A2(n_267), .B1(n_498), .B2(n_570), .Y(n_1116) );
AOI22xp33_ASAP7_75t_L g824 ( .A1(n_244), .A2(n_378), .B1(n_639), .B2(n_658), .Y(n_824) );
INVx2_ASAP7_75t_L g390 ( .A(n_246), .Y(n_390) );
AOI22xp33_ASAP7_75t_SL g794 ( .A1(n_248), .A2(n_335), .B1(n_436), .B2(n_446), .Y(n_794) );
INVx1_ASAP7_75t_L g404 ( .A(n_256), .Y(n_404) );
AOI22xp33_ASAP7_75t_L g720 ( .A1(n_258), .A2(n_270), .B1(n_721), .B2(n_722), .Y(n_720) );
OA22x2_ASAP7_75t_L g973 ( .A1(n_259), .A2(n_974), .B1(n_975), .B2(n_976), .Y(n_973) );
INVx1_ASAP7_75t_L g974 ( .A(n_259), .Y(n_974) );
AOI22xp33_ASAP7_75t_SL g994 ( .A1(n_260), .A2(n_294), .B1(n_575), .B2(n_963), .Y(n_994) );
AOI22xp5_ASAP7_75t_L g736 ( .A1(n_261), .A2(n_737), .B1(n_766), .B2(n_767), .Y(n_736) );
INVx1_ASAP7_75t_L g766 ( .A(n_261), .Y(n_766) );
INVx1_ASAP7_75t_L g454 ( .A(n_262), .Y(n_454) );
AOI22xp33_ASAP7_75t_L g729 ( .A1(n_263), .A2(n_320), .B1(n_730), .B2(n_731), .Y(n_729) );
INVx1_ASAP7_75t_L g1000 ( .A(n_268), .Y(n_1000) );
CKINVDCx20_ASAP7_75t_R g847 ( .A(n_269), .Y(n_847) );
CKINVDCx20_ASAP7_75t_R g1076 ( .A(n_274), .Y(n_1076) );
AOI22xp33_ASAP7_75t_L g958 ( .A1(n_278), .A2(n_318), .B1(n_741), .B2(n_920), .Y(n_958) );
AOI22xp33_ASAP7_75t_L g668 ( .A1(n_279), .A2(n_326), .B1(n_594), .B2(n_669), .Y(n_668) );
AOI22xp33_ASAP7_75t_L g915 ( .A1(n_280), .A2(n_297), .B1(n_472), .B2(n_575), .Y(n_915) );
NAND2xp5_ASAP7_75t_SL g796 ( .A(n_282), .B(n_516), .Y(n_796) );
AOI22xp33_ASAP7_75t_L g680 ( .A1(n_284), .A2(n_325), .B1(n_470), .B2(n_681), .Y(n_680) );
CKINVDCx20_ASAP7_75t_R g1019 ( .A(n_285), .Y(n_1019) );
AOI22xp33_ASAP7_75t_L g724 ( .A1(n_287), .A2(n_370), .B1(n_516), .B2(n_593), .Y(n_724) );
AOI22xp33_ASAP7_75t_SL g864 ( .A1(n_289), .A2(n_380), .B1(n_636), .B2(n_648), .Y(n_864) );
CKINVDCx20_ASAP7_75t_R g1038 ( .A(n_290), .Y(n_1038) );
INVx1_ASAP7_75t_L g410 ( .A(n_291), .Y(n_410) );
INVx1_ASAP7_75t_L g412 ( .A(n_291), .Y(n_412) );
AOI22xp33_ASAP7_75t_L g852 ( .A1(n_292), .A2(n_296), .B1(n_669), .B2(n_853), .Y(n_852) );
INVx1_ASAP7_75t_L g624 ( .A(n_293), .Y(n_624) );
CKINVDCx20_ASAP7_75t_R g1070 ( .A(n_295), .Y(n_1070) );
CKINVDCx20_ASAP7_75t_R g1013 ( .A(n_300), .Y(n_1013) );
CKINVDCx20_ASAP7_75t_R g1017 ( .A(n_301), .Y(n_1017) );
CKINVDCx20_ASAP7_75t_R g1045 ( .A(n_307), .Y(n_1045) );
CKINVDCx20_ASAP7_75t_R g761 ( .A(n_309), .Y(n_761) );
AOI22xp33_ASAP7_75t_SL g799 ( .A1(n_310), .A2(n_357), .B1(n_524), .B2(n_727), .Y(n_799) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_311), .B(n_444), .Y(n_443) );
CKINVDCx20_ASAP7_75t_R g1112 ( .A(n_314), .Y(n_1112) );
CKINVDCx20_ASAP7_75t_R g563 ( .A(n_316), .Y(n_563) );
AOI22xp33_ASAP7_75t_L g782 ( .A1(n_319), .A2(n_347), .B1(n_528), .B2(n_783), .Y(n_782) );
NAND2xp5_ASAP7_75t_SL g518 ( .A(n_321), .B(n_519), .Y(n_518) );
AO22x2_ASAP7_75t_L g544 ( .A1(n_323), .A2(n_545), .B1(n_579), .B2(n_580), .Y(n_544) );
CKINVDCx20_ASAP7_75t_R g580 ( .A(n_323), .Y(n_580) );
AOI22xp33_ASAP7_75t_SL g699 ( .A1(n_324), .A2(n_350), .B1(n_434), .B2(n_700), .Y(n_699) );
CKINVDCx20_ASAP7_75t_R g843 ( .A(n_330), .Y(n_843) );
INVx1_ASAP7_75t_L g389 ( .A(n_331), .Y(n_389) );
AOI22xp33_ASAP7_75t_L g961 ( .A1(n_332), .A2(n_341), .B1(n_487), .B2(n_636), .Y(n_961) );
CKINVDCx20_ASAP7_75t_R g685 ( .A(n_333), .Y(n_685) );
INVx1_ASAP7_75t_L g386 ( .A(n_334), .Y(n_386) );
XOR2x2_ASAP7_75t_L g908 ( .A(n_336), .B(n_909), .Y(n_908) );
NAND2xp5_ASAP7_75t_L g892 ( .A(n_338), .B(n_781), .Y(n_892) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_339), .B(n_514), .Y(n_513) );
INVx1_ASAP7_75t_L g1025 ( .A(n_342), .Y(n_1025) );
AOI22xp5_ASAP7_75t_SL g809 ( .A1(n_346), .A2(n_810), .B1(n_832), .B2(n_833), .Y(n_809) );
INVx1_ASAP7_75t_L g833 ( .A(n_346), .Y(n_833) );
AOI22xp33_ASAP7_75t_L g968 ( .A1(n_348), .A2(n_362), .B1(n_596), .B2(n_932), .Y(n_968) );
INVx1_ASAP7_75t_L g987 ( .A(n_349), .Y(n_987) );
CKINVDCx20_ASAP7_75t_R g752 ( .A(n_352), .Y(n_752) );
CKINVDCx20_ASAP7_75t_R g1014 ( .A(n_353), .Y(n_1014) );
CKINVDCx20_ASAP7_75t_R g1040 ( .A(n_354), .Y(n_1040) );
CKINVDCx20_ASAP7_75t_R g779 ( .A(n_356), .Y(n_779) );
CKINVDCx20_ASAP7_75t_R g965 ( .A(n_366), .Y(n_965) );
CKINVDCx20_ASAP7_75t_R g826 ( .A(n_368), .Y(n_826) );
OAI22xp5_ASAP7_75t_L g675 ( .A1(n_371), .A2(n_676), .B1(n_677), .B2(n_706), .Y(n_675) );
INVx1_ASAP7_75t_L g706 ( .A(n_371), .Y(n_706) );
INVx1_ASAP7_75t_L g449 ( .A(n_372), .Y(n_449) );
INVx1_ASAP7_75t_L g980 ( .A(n_374), .Y(n_980) );
CKINVDCx20_ASAP7_75t_R g930 ( .A(n_379), .Y(n_930) );
INVx2_ASAP7_75t_SL g383 ( .A(n_384), .Y(n_383) );
NAND2xp5_ASAP7_75t_SL g384 ( .A(n_385), .B(n_387), .Y(n_384) );
HB1xp67_ASAP7_75t_L g1054 ( .A(n_386), .Y(n_1054) );
OA21x2_ASAP7_75t_L g1097 ( .A1(n_387), .A2(n_1053), .B(n_1098), .Y(n_1097) );
NOR2xp33_ASAP7_75t_L g387 ( .A(n_388), .B(n_390), .Y(n_387) );
HB1xp67_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
AOI221xp5_ASAP7_75t_L g391 ( .A1(n_392), .A2(n_838), .B1(n_1048), .B2(n_1049), .C(n_1050), .Y(n_391) );
INVx1_ASAP7_75t_L g1048 ( .A(n_392), .Y(n_1048) );
AOI22xp5_ASAP7_75t_SL g392 ( .A1(n_393), .A2(n_711), .B1(n_712), .B2(n_837), .Y(n_392) );
INVx1_ASAP7_75t_L g837 ( .A(n_393), .Y(n_837) );
AOI22xp5_ASAP7_75t_L g393 ( .A1(n_394), .A2(n_613), .B1(n_709), .B2(n_710), .Y(n_393) );
INVx1_ASAP7_75t_L g709 ( .A(n_394), .Y(n_709) );
OAI22xp5_ASAP7_75t_L g394 ( .A1(n_395), .A2(n_396), .B1(n_542), .B2(n_543), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
OAI22xp5_ASAP7_75t_L g396 ( .A1(n_397), .A2(n_398), .B1(n_503), .B2(n_504), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
HB1xp67_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx2_ASAP7_75t_SL g501 ( .A(n_401), .Y(n_501) );
AND2x2_ASAP7_75t_L g401 ( .A(n_402), .B(n_461), .Y(n_401) );
NOR3xp33_ASAP7_75t_L g402 ( .A(n_403), .B(n_425), .C(n_448), .Y(n_402) );
OAI22xp5_ASAP7_75t_L g403 ( .A1(n_404), .A2(n_405), .B1(n_420), .B2(n_421), .Y(n_403) );
OAI22xp5_ASAP7_75t_L g978 ( .A1(n_405), .A2(n_625), .B1(n_979), .B2(n_980), .Y(n_978) );
OAI21xp5_ASAP7_75t_SL g1039 ( .A1(n_405), .A2(n_1040), .B(n_1041), .Y(n_1039) );
OAI221xp5_ASAP7_75t_SL g1118 ( .A1(n_405), .A2(n_1071), .B1(n_1119), .B2(n_1120), .C(n_1121), .Y(n_1118) );
BUFx6f_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx2_ASAP7_75t_L g550 ( .A(n_406), .Y(n_550) );
OAI22xp5_ASAP7_75t_SL g812 ( .A1(n_406), .A2(n_626), .B1(n_813), .B2(n_814), .Y(n_812) );
OAI21xp5_ASAP7_75t_L g999 ( .A1(n_406), .A2(n_1000), .B(n_1001), .Y(n_999) );
OR2x2_ASAP7_75t_L g406 ( .A(n_407), .B(n_415), .Y(n_406) );
INVx2_ASAP7_75t_L g480 ( .A(n_407), .Y(n_480) );
OR2x2_ASAP7_75t_L g407 ( .A(n_408), .B(n_413), .Y(n_407) );
AND2x2_ASAP7_75t_L g424 ( .A(n_408), .B(n_413), .Y(n_424) );
AND2x2_ASAP7_75t_L g469 ( .A(n_408), .B(n_440), .Y(n_469) );
INVx2_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
AND2x2_ASAP7_75t_L g429 ( .A(n_409), .B(n_413), .Y(n_429) );
AND2x2_ASAP7_75t_L g441 ( .A(n_409), .B(n_419), .Y(n_441) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g414 ( .A(n_412), .Y(n_414) );
INVx2_ASAP7_75t_L g440 ( .A(n_413), .Y(n_440) );
INVx1_ASAP7_75t_L g500 ( .A(n_413), .Y(n_500) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
NAND2x1p5_ASAP7_75t_L g423 ( .A(n_416), .B(n_424), .Y(n_423) );
AND2x4_ASAP7_75t_L g491 ( .A(n_416), .B(n_469), .Y(n_491) );
AND2x6_ASAP7_75t_L g517 ( .A(n_416), .B(n_424), .Y(n_517) );
AND2x4_ASAP7_75t_L g521 ( .A(n_416), .B(n_480), .Y(n_521) );
AND2x2_ASAP7_75t_L g416 ( .A(n_417), .B(n_418), .Y(n_416) );
INVx1_ASAP7_75t_L g431 ( .A(n_417), .Y(n_431) );
INVx1_ASAP7_75t_L g439 ( .A(n_417), .Y(n_439) );
INVx1_ASAP7_75t_L g460 ( .A(n_417), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_417), .B(n_419), .Y(n_475) );
AND2x2_ASAP7_75t_L g430 ( .A(n_418), .B(n_431), .Y(n_430) );
INVx2_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
AND2x2_ASAP7_75t_L g468 ( .A(n_419), .B(n_460), .Y(n_468) );
INVx1_ASAP7_75t_SL g421 ( .A(n_422), .Y(n_421) );
INVx2_ASAP7_75t_L g552 ( .A(n_422), .Y(n_552) );
INVx1_ASAP7_75t_L g966 ( .A(n_422), .Y(n_966) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
BUFx3_ASAP7_75t_L g626 ( .A(n_423), .Y(n_626) );
AND2x4_ASAP7_75t_L g483 ( .A(n_424), .B(n_430), .Y(n_483) );
AND2x2_ASAP7_75t_L g496 ( .A(n_424), .B(n_468), .Y(n_496) );
NAND2xp5_ASAP7_75t_SL g1020 ( .A(n_424), .B(n_468), .Y(n_1020) );
OAI221xp5_ASAP7_75t_L g425 ( .A1(n_426), .A2(n_432), .B1(n_433), .B2(n_442), .C(n_443), .Y(n_425) );
OAI21xp33_ASAP7_75t_SL g627 ( .A1(n_426), .A2(n_628), .B(n_629), .Y(n_627) );
OAI21xp33_ASAP7_75t_L g981 ( .A1(n_426), .A2(n_982), .B(n_983), .Y(n_981) );
INVx2_ASAP7_75t_SL g426 ( .A(n_427), .Y(n_426) );
INVx2_ASAP7_75t_L g508 ( .A(n_427), .Y(n_508) );
BUFx6f_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
BUFx3_ASAP7_75t_L g556 ( .A(n_428), .Y(n_556) );
INVx2_ASAP7_75t_L g585 ( .A(n_428), .Y(n_585) );
INVx4_ASAP7_75t_L g697 ( .A(n_428), .Y(n_697) );
INVx2_ASAP7_75t_SL g762 ( .A(n_428), .Y(n_762) );
INVx2_ASAP7_75t_L g878 ( .A(n_428), .Y(n_878) );
AND2x6_ASAP7_75t_L g428 ( .A(n_429), .B(n_430), .Y(n_428) );
INVx1_ASAP7_75t_L g457 ( .A(n_429), .Y(n_457) );
AND2x4_ASAP7_75t_L g529 ( .A(n_429), .B(n_459), .Y(n_529) );
AND2x6_ASAP7_75t_L g479 ( .A(n_430), .B(n_480), .Y(n_479) );
AND2x2_ASAP7_75t_L g488 ( .A(n_430), .B(n_469), .Y(n_488) );
OAI221xp5_ASAP7_75t_L g1073 ( .A1(n_433), .A2(n_1074), .B1(n_1075), .B2(n_1076), .C(n_1077), .Y(n_1073) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx3_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
OAI22xp5_ASAP7_75t_L g1005 ( .A1(n_435), .A2(n_762), .B1(n_1006), .B2(n_1007), .Y(n_1005) );
INVx4_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
BUFx2_ASAP7_75t_L g849 ( .A(n_436), .Y(n_849) );
INVx2_ASAP7_75t_L g1044 ( .A(n_436), .Y(n_1044) );
BUFx6f_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
BUFx2_ASAP7_75t_L g558 ( .A(n_437), .Y(n_558) );
BUFx6f_ASAP7_75t_L g589 ( .A(n_437), .Y(n_589) );
BUFx4f_ASAP7_75t_SL g672 ( .A(n_437), .Y(n_672) );
BUFx6f_ASAP7_75t_L g785 ( .A(n_437), .Y(n_785) );
AND2x4_ASAP7_75t_L g437 ( .A(n_438), .B(n_441), .Y(n_437) );
AND2x2_ASAP7_75t_L g438 ( .A(n_439), .B(n_440), .Y(n_438) );
INVx1_ASAP7_75t_L g447 ( .A(n_439), .Y(n_447) );
INVx1_ASAP7_75t_L g453 ( .A(n_440), .Y(n_453) );
AND2x4_ASAP7_75t_L g446 ( .A(n_441), .B(n_447), .Y(n_446) );
NAND2x1p5_ASAP7_75t_L g452 ( .A(n_441), .B(n_453), .Y(n_452) );
AND2x4_ASAP7_75t_L g524 ( .A(n_441), .B(n_525), .Y(n_524) );
BUFx3_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx2_ASAP7_75t_L g764 ( .A(n_445), .Y(n_764) );
BUFx2_ASAP7_75t_L g1123 ( .A(n_445), .Y(n_1123) );
BUFx6f_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
BUFx6f_ASAP7_75t_L g511 ( .A(n_446), .Y(n_511) );
BUFx12f_ASAP7_75t_L g561 ( .A(n_446), .Y(n_561) );
OAI22xp5_ASAP7_75t_L g448 ( .A1(n_449), .A2(n_450), .B1(n_454), .B2(n_455), .Y(n_448) );
OAI22xp5_ASAP7_75t_SL g818 ( .A1(n_450), .A2(n_455), .B1(n_819), .B2(n_820), .Y(n_818) );
OAI22xp5_ASAP7_75t_SL g1036 ( .A1(n_450), .A2(n_552), .B1(n_1037), .B2(n_1038), .Y(n_1036) );
INVx3_ASAP7_75t_SL g450 ( .A(n_451), .Y(n_450) );
INVx2_ASAP7_75t_L g564 ( .A(n_451), .Y(n_564) );
INVx4_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
OAI22xp5_ASAP7_75t_L g630 ( .A1(n_452), .A2(n_455), .B1(n_631), .B2(n_632), .Y(n_630) );
OAI22xp5_ASAP7_75t_L g984 ( .A1(n_452), .A2(n_985), .B1(n_986), .B2(n_987), .Y(n_984) );
OAI22xp5_ASAP7_75t_L g1002 ( .A1(n_452), .A2(n_626), .B1(n_1003), .B2(n_1004), .Y(n_1002) );
BUFx3_ASAP7_75t_L g1080 ( .A(n_452), .Y(n_1080) );
AND2x2_ASAP7_75t_L g873 ( .A(n_453), .B(n_474), .Y(n_873) );
OAI22xp5_ASAP7_75t_L g1078 ( .A1(n_455), .A2(n_1079), .B1(n_1080), .B2(n_1081), .Y(n_1078) );
BUFx2_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
OAI22xp5_ASAP7_75t_L g562 ( .A1(n_456), .A2(n_563), .B1(n_564), .B2(n_565), .Y(n_562) );
OR2x6_ASAP7_75t_L g456 ( .A(n_457), .B(n_458), .Y(n_456) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
NOR2xp33_ASAP7_75t_L g461 ( .A(n_462), .B(n_484), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_463), .B(n_476), .Y(n_462) );
INVx1_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
BUFx4f_ASAP7_75t_SL g636 ( .A(n_466), .Y(n_636) );
BUFx3_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
BUFx3_ASAP7_75t_L g535 ( .A(n_467), .Y(n_535) );
BUFx3_ASAP7_75t_L g604 ( .A(n_467), .Y(n_604) );
BUFx3_ASAP7_75t_L g719 ( .A(n_467), .Y(n_719) );
AND2x2_ASAP7_75t_L g467 ( .A(n_468), .B(n_469), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_468), .B(n_469), .Y(n_694) );
AND2x4_ASAP7_75t_L g473 ( .A(n_469), .B(n_474), .Y(n_473) );
INVx2_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
INVx2_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
BUFx3_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
BUFx3_ASAP7_75t_L g578 ( .A(n_473), .Y(n_578) );
BUFx2_ASAP7_75t_SL g601 ( .A(n_473), .Y(n_601) );
BUFx2_ASAP7_75t_SL g637 ( .A(n_473), .Y(n_637) );
BUFx2_ASAP7_75t_L g666 ( .A(n_473), .Y(n_666) );
BUFx3_ASAP7_75t_L g806 ( .A(n_473), .Y(n_806) );
BUFx3_ASAP7_75t_L g859 ( .A(n_473), .Y(n_859) );
INVx1_ASAP7_75t_L g1018 ( .A(n_473), .Y(n_1018) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
OR2x6_ASAP7_75t_L g499 ( .A(n_475), .B(n_500), .Y(n_499) );
INVx2_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
INVx4_ASAP7_75t_L g540 ( .A(n_478), .Y(n_540) );
INVx2_ASAP7_75t_SL g577 ( .A(n_478), .Y(n_577) );
INVx5_ASAP7_75t_SL g646 ( .A(n_478), .Y(n_646) );
INVx1_ASAP7_75t_L g741 ( .A(n_478), .Y(n_741) );
NOR2xp33_ASAP7_75t_L g1023 ( .A(n_478), .B(n_1024), .Y(n_1023) );
INVx11_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
INVx11_ASAP7_75t_L g662 ( .A(n_479), .Y(n_662) );
INVx3_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx2_ASAP7_75t_L g607 ( .A(n_482), .Y(n_607) );
INVx2_ASAP7_75t_L g722 ( .A(n_482), .Y(n_722) );
OAI22xp5_ASAP7_75t_L g825 ( .A1(n_482), .A2(n_826), .B1(n_827), .B2(n_828), .Y(n_825) );
OAI22xp5_ASAP7_75t_SL g1012 ( .A1(n_482), .A2(n_574), .B1(n_1013), .B2(n_1014), .Y(n_1012) );
INVx6_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
BUFx3_ASAP7_75t_L g532 ( .A(n_483), .Y(n_532) );
BUFx3_ASAP7_75t_L g568 ( .A(n_483), .Y(n_568) );
BUFx3_ASAP7_75t_L g920 ( .A(n_483), .Y(n_920) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_485), .B(n_492), .Y(n_484) );
BUFx3_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
BUFx6f_ASAP7_75t_L g648 ( .A(n_487), .Y(n_648) );
BUFx3_ASAP7_75t_L g746 ( .A(n_487), .Y(n_746) );
BUFx6f_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
INVx2_ASAP7_75t_L g574 ( .A(n_488), .Y(n_574) );
BUFx2_ASAP7_75t_SL g603 ( .A(n_488), .Y(n_603) );
BUFx2_ASAP7_75t_SL g870 ( .A(n_488), .Y(n_870) );
BUFx2_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
BUFx3_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
BUFx3_ASAP7_75t_L g575 ( .A(n_491), .Y(n_575) );
BUFx6f_ASAP7_75t_L g608 ( .A(n_491), .Y(n_608) );
BUFx3_ASAP7_75t_L g731 ( .A(n_491), .Y(n_731) );
INVx2_ASAP7_75t_L g858 ( .A(n_491), .Y(n_858) );
BUFx6f_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
BUFx2_ASAP7_75t_L g1092 ( .A(n_494), .Y(n_1092) );
INVx5_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
INVx4_ASAP7_75t_L g538 ( .A(n_495), .Y(n_538) );
INVx2_ASAP7_75t_L g570 ( .A(n_495), .Y(n_570) );
INVx1_ASAP7_75t_L g803 ( .A(n_495), .Y(n_803) );
INVx3_ASAP7_75t_L g868 ( .A(n_495), .Y(n_868) );
INVx8_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
BUFx4f_ASAP7_75t_SL g497 ( .A(n_498), .Y(n_497) );
BUFx2_ASAP7_75t_L g571 ( .A(n_498), .Y(n_571) );
BUFx2_ASAP7_75t_L g641 ( .A(n_498), .Y(n_641) );
BUFx2_ASAP7_75t_L g658 ( .A(n_498), .Y(n_658) );
INVx6_ASAP7_75t_SL g498 ( .A(n_499), .Y(n_498) );
INVx1_ASAP7_75t_SL g610 ( .A(n_499), .Y(n_610) );
INVx1_ASAP7_75t_SL g904 ( .A(n_499), .Y(n_904) );
INVx1_ASAP7_75t_L g963 ( .A(n_499), .Y(n_963) );
INVx1_ASAP7_75t_L g525 ( .A(n_500), .Y(n_525) );
INVx1_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
NAND4xp75_ASAP7_75t_SL g505 ( .A(n_506), .B(n_530), .C(n_539), .D(n_541), .Y(n_505) );
NOR2xp67_ASAP7_75t_L g506 ( .A(n_507), .B(n_512), .Y(n_506) );
OAI21xp5_ASAP7_75t_SL g507 ( .A1(n_508), .A2(n_509), .B(n_510), .Y(n_507) );
OAI21xp5_ASAP7_75t_SL g846 ( .A1(n_508), .A2(n_847), .B(n_848), .Y(n_846) );
BUFx4f_ASAP7_75t_L g700 ( .A(n_511), .Y(n_700) );
NAND3xp33_ASAP7_75t_L g512 ( .A(n_513), .B(n_518), .C(n_522), .Y(n_512) );
INVx1_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
BUFx4f_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
BUFx2_ASAP7_75t_L g594 ( .A(n_517), .Y(n_594) );
INVx1_ASAP7_75t_SL g854 ( .A(n_517), .Y(n_854) );
BUFx2_ASAP7_75t_L g891 ( .A(n_517), .Y(n_891) );
BUFx6f_ASAP7_75t_L g669 ( .A(n_519), .Y(n_669) );
HB1xp67_ASAP7_75t_L g704 ( .A(n_519), .Y(n_704) );
INVx5_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
INVx2_ASAP7_75t_L g593 ( .A(n_520), .Y(n_593) );
INVx2_ASAP7_75t_L g781 ( .A(n_520), .Y(n_781) );
INVx2_ASAP7_75t_L g798 ( .A(n_520), .Y(n_798) );
INVx4_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
BUFx2_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
INVx1_ASAP7_75t_L g597 ( .A(n_524), .Y(n_597) );
BUFx2_ASAP7_75t_L g726 ( .A(n_524), .Y(n_726) );
BUFx3_ASAP7_75t_L g783 ( .A(n_524), .Y(n_783) );
INVx2_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
INVx1_ASAP7_75t_SL g527 ( .A(n_528), .Y(n_527) );
BUFx6f_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
BUFx3_ASAP7_75t_L g727 ( .A(n_529), .Y(n_727) );
BUFx2_ASAP7_75t_SL g932 ( .A(n_529), .Y(n_932) );
AND2x2_ASAP7_75t_L g530 ( .A(n_531), .B(n_536), .Y(n_530) );
INVx1_ASAP7_75t_L g687 ( .A(n_532), .Y(n_687) );
INVx2_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
BUFx2_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
INVx2_ASAP7_75t_L g640 ( .A(n_538), .Y(n_640) );
BUFx6f_ASAP7_75t_L g683 ( .A(n_538), .Y(n_683) );
INVx1_ASAP7_75t_SL g827 ( .A(n_540), .Y(n_827) );
INVx2_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
XNOR2x2_ASAP7_75t_L g543 ( .A(n_544), .B(n_581), .Y(n_543) );
XNOR2xp5_ASAP7_75t_L g674 ( .A(n_544), .B(n_675), .Y(n_674) );
INVx1_ASAP7_75t_SL g579 ( .A(n_545), .Y(n_579) );
AND2x2_ASAP7_75t_SL g545 ( .A(n_546), .B(n_566), .Y(n_545) );
NOR3xp33_ASAP7_75t_L g546 ( .A(n_547), .B(n_553), .C(n_562), .Y(n_546) );
OAI22xp5_ASAP7_75t_L g547 ( .A1(n_548), .A2(n_549), .B1(n_551), .B2(n_552), .Y(n_547) );
INVx2_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
INVx2_ASAP7_75t_L g623 ( .A(n_550), .Y(n_623) );
OAI21xp33_ASAP7_75t_L g553 ( .A1(n_554), .A2(n_555), .B(n_557), .Y(n_553) );
INVx3_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
INVx3_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
INVx2_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
BUFx4f_ASAP7_75t_SL g590 ( .A(n_561), .Y(n_590) );
AND4x1_ASAP7_75t_L g566 ( .A(n_567), .B(n_569), .C(n_572), .D(n_576), .Y(n_566) );
INVx1_ASAP7_75t_L g743 ( .A(n_568), .Y(n_743) );
INVx3_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
INVx3_ASAP7_75t_L g730 ( .A(n_574), .Y(n_730) );
BUFx2_ASAP7_75t_L g749 ( .A(n_575), .Y(n_749) );
INVxp67_ASAP7_75t_L g1113 ( .A(n_575), .Y(n_1113) );
INVx1_ASAP7_75t_L g1090 ( .A(n_577), .Y(n_1090) );
INVx2_ASAP7_75t_SL g611 ( .A(n_582), .Y(n_611) );
AND2x2_ASAP7_75t_L g582 ( .A(n_583), .B(n_598), .Y(n_582) );
NOR2xp33_ASAP7_75t_L g583 ( .A(n_584), .B(n_591), .Y(n_583) );
OAI21xp5_ASAP7_75t_SL g584 ( .A1(n_585), .A2(n_586), .B(n_587), .Y(n_584) );
OAI21xp5_ASAP7_75t_SL g792 ( .A1(n_585), .A2(n_793), .B(n_794), .Y(n_792) );
OAI21xp5_ASAP7_75t_SL g894 ( .A1(n_585), .A2(n_895), .B(n_896), .Y(n_894) );
OAI21xp5_ASAP7_75t_L g929 ( .A1(n_585), .A2(n_930), .B(n_931), .Y(n_929) );
BUFx6f_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
INVx1_ASAP7_75t_L g986 ( .A(n_589), .Y(n_986) );
NAND2xp5_ASAP7_75t_SL g591 ( .A(n_592), .B(n_595), .Y(n_591) );
INVx1_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
NOR2xp33_ASAP7_75t_L g598 ( .A(n_599), .B(n_605), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_600), .B(n_602), .Y(n_599) );
INVx1_ASAP7_75t_L g690 ( .A(n_603), .Y(n_690) );
INVx1_ASAP7_75t_L g914 ( .A(n_604), .Y(n_914) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_606), .B(n_609), .Y(n_605) );
INVx2_ASAP7_75t_L g1106 ( .A(n_607), .Y(n_1106) );
INVx4_ASAP7_75t_L g665 ( .A(n_608), .Y(n_665) );
INVx1_ASAP7_75t_L g710 ( .A(n_613), .Y(n_710) );
AOI22xp5_ASAP7_75t_L g613 ( .A1(n_614), .A2(n_649), .B1(n_650), .B2(n_708), .Y(n_613) );
INVx1_ASAP7_75t_L g708 ( .A(n_614), .Y(n_708) );
HB1xp67_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
INVx1_ASAP7_75t_SL g618 ( .A(n_619), .Y(n_618) );
AND2x2_ASAP7_75t_L g619 ( .A(n_620), .B(n_633), .Y(n_619) );
NOR3xp33_ASAP7_75t_L g620 ( .A(n_621), .B(n_627), .C(n_630), .Y(n_620) );
OAI22xp5_ASAP7_75t_L g621 ( .A1(n_622), .A2(n_623), .B1(n_624), .B2(n_625), .Y(n_621) );
OAI221xp5_ASAP7_75t_SL g755 ( .A1(n_623), .A2(n_625), .B1(n_756), .B2(n_757), .C(n_758), .Y(n_755) );
OAI22xp5_ASAP7_75t_L g1068 ( .A1(n_623), .A2(n_1069), .B1(n_1070), .B2(n_1071), .Y(n_1068) );
BUFx3_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
OA211x2_ASAP7_75t_L g778 ( .A1(n_626), .A2(n_779), .B(n_780), .C(n_782), .Y(n_778) );
INVx2_ASAP7_75t_L g1072 ( .A(n_626), .Y(n_1072) );
NOR2xp33_ASAP7_75t_L g633 ( .A(n_634), .B(n_642), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_635), .B(n_638), .Y(n_634) );
INVx1_ASAP7_75t_L g751 ( .A(n_637), .Y(n_751) );
INVx3_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_643), .B(n_647), .Y(n_642) );
INVx2_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
OAI22xp5_ASAP7_75t_L g684 ( .A1(n_645), .A2(n_685), .B1(n_686), .B2(n_687), .Y(n_684) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
INVx1_ASAP7_75t_SL g1111 ( .A(n_648), .Y(n_1111) );
INVx2_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
AO22x1_ASAP7_75t_L g650 ( .A1(n_651), .A2(n_652), .B1(n_674), .B2(n_707), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
INVx1_ASAP7_75t_SL g673 ( .A(n_654), .Y(n_673) );
NAND4xp75_ASAP7_75t_L g654 ( .A(n_655), .B(n_659), .C(n_667), .D(n_671), .Y(n_654) );
AND2x2_ASAP7_75t_L g655 ( .A(n_656), .B(n_657), .Y(n_655) );
AND2x2_ASAP7_75t_L g659 ( .A(n_660), .B(n_663), .Y(n_659) );
INVx2_ASAP7_75t_SL g661 ( .A(n_662), .Y(n_661) );
INVx3_ASAP7_75t_L g721 ( .A(n_662), .Y(n_721) );
INVx4_ASAP7_75t_L g863 ( .A(n_662), .Y(n_863) );
INVx4_ASAP7_75t_L g912 ( .A(n_662), .Y(n_912) );
INVx3_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
INVx4_ASAP7_75t_L g681 ( .A(n_665), .Y(n_681) );
AND2x2_ASAP7_75t_SL g667 ( .A(n_668), .B(n_670), .Y(n_667) );
INVx1_ASAP7_75t_L g760 ( .A(n_672), .Y(n_760) );
INVx1_ASAP7_75t_L g707 ( .A(n_674), .Y(n_707) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
AND2x2_ASAP7_75t_SL g677 ( .A(n_678), .B(n_695), .Y(n_677) );
NOR3xp33_ASAP7_75t_L g678 ( .A(n_679), .B(n_684), .C(n_688), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_680), .B(n_682), .Y(n_679) );
INVx1_ASAP7_75t_L g1086 ( .A(n_687), .Y(n_1086) );
OAI22xp5_ASAP7_75t_L g688 ( .A1(n_689), .A2(n_690), .B1(n_691), .B2(n_692), .Y(n_688) );
OAI22xp5_ASAP7_75t_L g829 ( .A1(n_690), .A2(n_692), .B1(n_830), .B2(n_831), .Y(n_829) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
INVx1_ASAP7_75t_L g1108 ( .A(n_693), .Y(n_1108) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
NOR2xp33_ASAP7_75t_L g1021 ( .A(n_694), .B(n_1022), .Y(n_1021) );
NOR2xp33_ASAP7_75t_L g695 ( .A(n_696), .B(n_701), .Y(n_695) );
OAI21xp5_ASAP7_75t_SL g696 ( .A1(n_697), .A2(n_698), .B(n_699), .Y(n_696) );
INVx4_ASAP7_75t_L g734 ( .A(n_697), .Y(n_734) );
OAI21xp5_ASAP7_75t_SL g815 ( .A1(n_697), .A2(n_816), .B(n_817), .Y(n_815) );
OAI22xp5_ASAP7_75t_SL g1042 ( .A1(n_697), .A2(n_1043), .B1(n_1044), .B2(n_1045), .Y(n_1042) );
BUFx2_ASAP7_75t_L g1074 ( .A(n_697), .Y(n_1074) );
NAND3xp33_ASAP7_75t_L g701 ( .A(n_702), .B(n_703), .C(n_705), .Y(n_701) );
INVx1_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
XOR2x2_ASAP7_75t_L g712 ( .A(n_713), .B(n_769), .Y(n_712) );
AOI22xp5_ASAP7_75t_L g713 ( .A1(n_714), .A2(n_715), .B1(n_736), .B2(n_768), .Y(n_713) );
INVx2_ASAP7_75t_SL g714 ( .A(n_715), .Y(n_714) );
XOR2x2_ASAP7_75t_L g715 ( .A(n_716), .B(n_735), .Y(n_715) );
NAND4xp75_ASAP7_75t_L g716 ( .A(n_717), .B(n_723), .C(n_728), .D(n_733), .Y(n_716) );
AND2x2_ASAP7_75t_L g717 ( .A(n_718), .B(n_720), .Y(n_717) );
AND2x2_ASAP7_75t_SL g723 ( .A(n_724), .B(n_725), .Y(n_723) );
AND2x2_ASAP7_75t_L g728 ( .A(n_729), .B(n_732), .Y(n_728) );
INVx1_ASAP7_75t_L g768 ( .A(n_736), .Y(n_768) );
INVx1_ASAP7_75t_L g767 ( .A(n_737), .Y(n_767) );
AND2x2_ASAP7_75t_L g737 ( .A(n_738), .B(n_754), .Y(n_737) );
NOR2xp33_ASAP7_75t_L g738 ( .A(n_739), .B(n_747), .Y(n_738) );
OAI221xp5_ASAP7_75t_SL g739 ( .A1(n_740), .A2(n_742), .B1(n_743), .B2(n_744), .C(n_745), .Y(n_739) );
INVx2_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
OAI221xp5_ASAP7_75t_SL g747 ( .A1(n_748), .A2(n_750), .B1(n_751), .B2(n_752), .C(n_753), .Y(n_747) );
INVx1_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
NOR2xp33_ASAP7_75t_SL g754 ( .A(n_755), .B(n_759), .Y(n_754) );
OAI222xp33_ASAP7_75t_L g759 ( .A1(n_760), .A2(n_761), .B1(n_762), .B2(n_763), .C1(n_764), .C2(n_765), .Y(n_759) );
AO22x1_ASAP7_75t_L g769 ( .A1(n_770), .A2(n_787), .B1(n_788), .B2(n_836), .Y(n_769) );
INVx2_ASAP7_75t_SL g836 ( .A(n_770), .Y(n_836) );
XOR2x2_ASAP7_75t_L g770 ( .A(n_771), .B(n_786), .Y(n_770) );
NAND4xp75_ASAP7_75t_L g771 ( .A(n_772), .B(n_775), .C(n_778), .D(n_784), .Y(n_771) );
AND2x2_ASAP7_75t_L g772 ( .A(n_773), .B(n_774), .Y(n_772) );
AND2x2_ASAP7_75t_L g775 ( .A(n_776), .B(n_777), .Y(n_775) );
INVx1_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
AO22x2_ASAP7_75t_SL g788 ( .A1(n_789), .A2(n_809), .B1(n_834), .B2(n_835), .Y(n_788) );
INVx4_ASAP7_75t_SL g834 ( .A(n_789), .Y(n_834) );
XOR2x2_ASAP7_75t_L g789 ( .A(n_790), .B(n_808), .Y(n_789) );
NAND3x1_ASAP7_75t_L g790 ( .A(n_791), .B(n_800), .C(n_804), .Y(n_790) );
NOR2xp33_ASAP7_75t_L g791 ( .A(n_792), .B(n_795), .Y(n_791) );
NAND3xp33_ASAP7_75t_L g795 ( .A(n_796), .B(n_797), .C(n_799), .Y(n_795) );
AND2x2_ASAP7_75t_L g800 ( .A(n_801), .B(n_802), .Y(n_800) );
AND2x2_ASAP7_75t_L g804 ( .A(n_805), .B(n_807), .Y(n_804) );
INVx1_ASAP7_75t_L g835 ( .A(n_809), .Y(n_835) );
INVx1_ASAP7_75t_L g832 ( .A(n_810), .Y(n_832) );
AND2x2_ASAP7_75t_L g810 ( .A(n_811), .B(n_821), .Y(n_810) );
NOR3xp33_ASAP7_75t_L g811 ( .A(n_812), .B(n_815), .C(n_818), .Y(n_811) );
NOR3xp33_ASAP7_75t_L g821 ( .A(n_822), .B(n_825), .C(n_829), .Y(n_821) );
NAND2xp5_ASAP7_75t_L g822 ( .A(n_823), .B(n_824), .Y(n_822) );
INVx1_ASAP7_75t_L g1049 ( .A(n_838), .Y(n_1049) );
AOI22xp5_ASAP7_75t_SL g838 ( .A1(n_839), .A2(n_948), .B1(n_949), .B2(n_1047), .Y(n_838) );
INVx1_ASAP7_75t_L g1047 ( .A(n_839), .Y(n_1047) );
AOI22xp33_ASAP7_75t_L g839 ( .A1(n_840), .A2(n_841), .B1(n_884), .B2(n_947), .Y(n_839) );
INVx1_ASAP7_75t_L g840 ( .A(n_841), .Y(n_840) );
XOR2x2_ASAP7_75t_L g841 ( .A(n_842), .B(n_865), .Y(n_841) );
XNOR2xp5_ASAP7_75t_L g842 ( .A(n_843), .B(n_844), .Y(n_842) );
NAND3xp33_ASAP7_75t_L g844 ( .A(n_845), .B(n_855), .C(n_861), .Y(n_844) );
NOR2xp33_ASAP7_75t_L g845 ( .A(n_846), .B(n_850), .Y(n_845) );
NAND2xp5_ASAP7_75t_L g850 ( .A(n_851), .B(n_852), .Y(n_850) );
INVx1_ASAP7_75t_SL g853 ( .A(n_854), .Y(n_853) );
AND2x2_ASAP7_75t_L g855 ( .A(n_856), .B(n_860), .Y(n_855) );
INVx2_ASAP7_75t_L g857 ( .A(n_858), .Y(n_857) );
OAI21xp5_ASAP7_75t_SL g1009 ( .A1(n_858), .A2(n_1010), .B(n_1011), .Y(n_1009) );
AND2x2_ASAP7_75t_L g861 ( .A(n_862), .B(n_864), .Y(n_861) );
OAI22xp5_ASAP7_75t_L g952 ( .A1(n_865), .A2(n_953), .B1(n_954), .B2(n_955), .Y(n_952) );
INVx2_ASAP7_75t_L g953 ( .A(n_865), .Y(n_953) );
XOR2x2_ASAP7_75t_L g865 ( .A(n_866), .B(n_883), .Y(n_865) );
NAND4xp75_ASAP7_75t_SL g866 ( .A(n_867), .B(n_869), .C(n_871), .D(n_875), .Y(n_866) );
AND2x2_ASAP7_75t_L g871 ( .A(n_872), .B(n_874), .Y(n_871) );
NOR2xp33_ASAP7_75t_L g875 ( .A(n_876), .B(n_880), .Y(n_875) );
OAI21xp5_ASAP7_75t_L g876 ( .A1(n_877), .A2(n_878), .B(n_879), .Y(n_876) );
NAND2xp5_ASAP7_75t_L g880 ( .A(n_881), .B(n_882), .Y(n_880) );
INVx1_ASAP7_75t_L g947 ( .A(n_884), .Y(n_947) );
AOI22xp5_ASAP7_75t_L g884 ( .A1(n_885), .A2(n_906), .B1(n_907), .B2(n_946), .Y(n_884) );
INVx1_ASAP7_75t_SL g946 ( .A(n_885), .Y(n_946) );
INVx1_ASAP7_75t_L g885 ( .A(n_886), .Y(n_885) );
XOR2x2_ASAP7_75t_SL g886 ( .A(n_887), .B(n_905), .Y(n_886) );
NAND2x1p5_ASAP7_75t_L g887 ( .A(n_888), .B(n_897), .Y(n_887) );
NOR2xp33_ASAP7_75t_L g888 ( .A(n_889), .B(n_894), .Y(n_888) );
NAND3xp33_ASAP7_75t_L g889 ( .A(n_890), .B(n_892), .C(n_893), .Y(n_889) );
NOR2x1_ASAP7_75t_L g897 ( .A(n_898), .B(n_901), .Y(n_897) );
NAND2xp5_ASAP7_75t_L g898 ( .A(n_899), .B(n_900), .Y(n_898) );
NAND2xp5_ASAP7_75t_L g901 ( .A(n_902), .B(n_903), .Y(n_901) );
INVx1_ASAP7_75t_L g906 ( .A(n_907), .Y(n_906) );
AO22x1_ASAP7_75t_SL g907 ( .A1(n_908), .A2(n_926), .B1(n_944), .B2(n_945), .Y(n_907) );
INVx1_ASAP7_75t_L g944 ( .A(n_908), .Y(n_944) );
NAND4xp75_ASAP7_75t_L g909 ( .A(n_910), .B(n_916), .C(n_922), .D(n_925), .Y(n_909) );
AND2x2_ASAP7_75t_L g910 ( .A(n_911), .B(n_915), .Y(n_910) );
INVx1_ASAP7_75t_L g913 ( .A(n_914), .Y(n_913) );
AND2x2_ASAP7_75t_L g916 ( .A(n_917), .B(n_921), .Y(n_916) );
INVx2_ASAP7_75t_L g918 ( .A(n_919), .Y(n_918) );
INVx3_ASAP7_75t_L g919 ( .A(n_920), .Y(n_919) );
AND2x2_ASAP7_75t_SL g922 ( .A(n_923), .B(n_924), .Y(n_922) );
INVx3_ASAP7_75t_SL g945 ( .A(n_926), .Y(n_945) );
XOR2x2_ASAP7_75t_L g926 ( .A(n_927), .B(n_943), .Y(n_926) );
NAND2xp5_ASAP7_75t_SL g927 ( .A(n_928), .B(n_936), .Y(n_927) );
NOR2xp33_ASAP7_75t_L g928 ( .A(n_929), .B(n_933), .Y(n_928) );
NAND2xp5_ASAP7_75t_L g933 ( .A(n_934), .B(n_935), .Y(n_933) );
NOR2xp33_ASAP7_75t_L g936 ( .A(n_937), .B(n_940), .Y(n_936) );
NAND2xp5_ASAP7_75t_L g937 ( .A(n_938), .B(n_939), .Y(n_937) );
NAND2xp5_ASAP7_75t_L g940 ( .A(n_941), .B(n_942), .Y(n_940) );
INVx1_ASAP7_75t_L g948 ( .A(n_949), .Y(n_948) );
XOR2xp5_ASAP7_75t_L g949 ( .A(n_950), .B(n_970), .Y(n_949) );
HB1xp67_ASAP7_75t_L g950 ( .A(n_951), .Y(n_950) );
INVx1_ASAP7_75t_L g951 ( .A(n_952), .Y(n_951) );
INVx1_ASAP7_75t_L g954 ( .A(n_955), .Y(n_954) );
NAND4xp75_ASAP7_75t_L g956 ( .A(n_957), .B(n_960), .C(n_964), .D(n_969), .Y(n_956) );
AND2x2_ASAP7_75t_L g957 ( .A(n_958), .B(n_959), .Y(n_957) );
AND2x2_ASAP7_75t_L g960 ( .A(n_961), .B(n_962), .Y(n_960) );
OA211x2_ASAP7_75t_L g964 ( .A1(n_965), .A2(n_966), .B(n_967), .C(n_968), .Y(n_964) );
INVx1_ASAP7_75t_L g970 ( .A(n_971), .Y(n_970) );
AO22x2_ASAP7_75t_L g971 ( .A1(n_972), .A2(n_973), .B1(n_995), .B2(n_1046), .Y(n_971) );
INVx1_ASAP7_75t_L g972 ( .A(n_973), .Y(n_972) );
INVx1_ASAP7_75t_L g975 ( .A(n_976), .Y(n_975) );
AND2x2_ASAP7_75t_L g976 ( .A(n_977), .B(n_988), .Y(n_976) );
NOR3xp33_ASAP7_75t_L g977 ( .A(n_978), .B(n_981), .C(n_984), .Y(n_977) );
NOR2xp33_ASAP7_75t_L g988 ( .A(n_989), .B(n_992), .Y(n_988) );
NAND2xp5_ASAP7_75t_L g989 ( .A(n_990), .B(n_991), .Y(n_989) );
NAND2xp5_ASAP7_75t_L g992 ( .A(n_993), .B(n_994), .Y(n_992) );
INVx2_ASAP7_75t_L g1046 ( .A(n_995), .Y(n_1046) );
XOR2x2_ASAP7_75t_L g995 ( .A(n_996), .B(n_1026), .Y(n_995) );
XNOR2x1_ASAP7_75t_L g996 ( .A(n_997), .B(n_1025), .Y(n_996) );
AND3x2_ASAP7_75t_L g997 ( .A(n_998), .B(n_1008), .C(n_1015), .Y(n_997) );
NOR3xp33_ASAP7_75t_L g998 ( .A(n_999), .B(n_1002), .C(n_1005), .Y(n_998) );
NOR2xp33_ASAP7_75t_L g1008 ( .A(n_1009), .B(n_1012), .Y(n_1008) );
NOR3xp33_ASAP7_75t_L g1015 ( .A(n_1016), .B(n_1021), .C(n_1023), .Y(n_1015) );
OAI22xp5_ASAP7_75t_L g1016 ( .A1(n_1017), .A2(n_1018), .B1(n_1019), .B2(n_1020), .Y(n_1016) );
XNOR2xp5_ASAP7_75t_L g1026 ( .A(n_1027), .B(n_1028), .Y(n_1026) );
NAND3x1_ASAP7_75t_SL g1028 ( .A(n_1029), .B(n_1032), .C(n_1035), .Y(n_1028) );
AND2x2_ASAP7_75t_L g1029 ( .A(n_1030), .B(n_1031), .Y(n_1029) );
AND2x2_ASAP7_75t_L g1032 ( .A(n_1033), .B(n_1034), .Y(n_1032) );
NOR3xp33_ASAP7_75t_L g1035 ( .A(n_1036), .B(n_1039), .C(n_1042), .Y(n_1035) );
INVx1_ASAP7_75t_SL g1050 ( .A(n_1051), .Y(n_1050) );
NOR2x1_ASAP7_75t_L g1051 ( .A(n_1052), .B(n_1056), .Y(n_1051) );
OR2x2_ASAP7_75t_SL g1127 ( .A(n_1052), .B(n_1057), .Y(n_1127) );
NAND2xp5_ASAP7_75t_L g1052 ( .A(n_1053), .B(n_1055), .Y(n_1052) );
INVx1_ASAP7_75t_L g1053 ( .A(n_1054), .Y(n_1053) );
OAI322xp33_ASAP7_75t_L g1063 ( .A1(n_1054), .A2(n_1064), .A3(n_1093), .B1(n_1095), .B2(n_1099), .C1(n_1100), .C2(n_1125), .Y(n_1063) );
NAND2xp5_ASAP7_75t_L g1098 ( .A(n_1054), .B(n_1094), .Y(n_1098) );
CKINVDCx16_ASAP7_75t_R g1094 ( .A(n_1055), .Y(n_1094) );
CKINVDCx20_ASAP7_75t_R g1056 ( .A(n_1057), .Y(n_1056) );
NAND2xp5_ASAP7_75t_L g1057 ( .A(n_1058), .B(n_1059), .Y(n_1057) );
NAND2xp5_ASAP7_75t_L g1060 ( .A(n_1061), .B(n_1062), .Y(n_1060) );
INVx1_ASAP7_75t_L g1065 ( .A(n_1066), .Y(n_1065) );
NAND2xp5_ASAP7_75t_L g1066 ( .A(n_1067), .B(n_1082), .Y(n_1066) );
NOR3xp33_ASAP7_75t_L g1067 ( .A(n_1068), .B(n_1073), .C(n_1078), .Y(n_1067) );
INVx2_ASAP7_75t_L g1071 ( .A(n_1072), .Y(n_1071) );
NOR2xp67_ASAP7_75t_L g1082 ( .A(n_1083), .B(n_1087), .Y(n_1082) );
NAND2xp5_ASAP7_75t_L g1083 ( .A(n_1084), .B(n_1085), .Y(n_1083) );
NAND2xp5_ASAP7_75t_L g1087 ( .A(n_1088), .B(n_1091), .Y(n_1087) );
INVx1_ASAP7_75t_L g1089 ( .A(n_1090), .Y(n_1089) );
INVx1_ASAP7_75t_L g1093 ( .A(n_1094), .Y(n_1093) );
INVx1_ASAP7_75t_L g1095 ( .A(n_1096), .Y(n_1095) );
CKINVDCx20_ASAP7_75t_R g1096 ( .A(n_1097), .Y(n_1096) );
HB1xp67_ASAP7_75t_L g1100 ( .A(n_1101), .Y(n_1100) );
INVx2_ASAP7_75t_SL g1124 ( .A(n_1102), .Y(n_1124) );
AND4x1_ASAP7_75t_L g1102 ( .A(n_1103), .B(n_1114), .C(n_1117), .D(n_1122), .Y(n_1102) );
NOR2xp33_ASAP7_75t_L g1103 ( .A(n_1104), .B(n_1109), .Y(n_1103) );
OAI22xp5_ASAP7_75t_L g1104 ( .A1(n_1105), .A2(n_1106), .B1(n_1107), .B2(n_1108), .Y(n_1104) );
OAI22xp5_ASAP7_75t_L g1109 ( .A1(n_1110), .A2(n_1111), .B1(n_1112), .B2(n_1113), .Y(n_1109) );
AND2x2_ASAP7_75t_L g1114 ( .A(n_1115), .B(n_1116), .Y(n_1114) );
INVx1_ASAP7_75t_L g1117 ( .A(n_1118), .Y(n_1117) );
CKINVDCx20_ASAP7_75t_R g1125 ( .A(n_1126), .Y(n_1125) );
CKINVDCx20_ASAP7_75t_R g1126 ( .A(n_1127), .Y(n_1126) );
endmodule