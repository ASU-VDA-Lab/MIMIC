module fake_netlist_1_12093_n_38 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_38);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_38;
wire n_20;
wire n_36;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
AND2x4_ASAP7_75t_L g11 ( .A(n_5), .B(n_10), .Y(n_11) );
NOR2x1_ASAP7_75t_L g12 ( .A(n_5), .B(n_2), .Y(n_12) );
NAND2xp5_ASAP7_75t_SL g13 ( .A(n_2), .B(n_4), .Y(n_13) );
BUFx6f_ASAP7_75t_L g14 ( .A(n_4), .Y(n_14) );
AND2x4_ASAP7_75t_L g15 ( .A(n_8), .B(n_7), .Y(n_15) );
INVx2_ASAP7_75t_L g16 ( .A(n_1), .Y(n_16) );
NAND2xp5_ASAP7_75t_L g17 ( .A(n_15), .B(n_0), .Y(n_17) );
HB1xp67_ASAP7_75t_L g18 ( .A(n_16), .Y(n_18) );
NAND2xp5_ASAP7_75t_L g19 ( .A(n_15), .B(n_0), .Y(n_19) );
INVx1_ASAP7_75t_L g20 ( .A(n_16), .Y(n_20) );
HB1xp67_ASAP7_75t_L g21 ( .A(n_18), .Y(n_21) );
AND2x2_ASAP7_75t_L g22 ( .A(n_20), .B(n_11), .Y(n_22) );
AND2x2_ASAP7_75t_L g23 ( .A(n_21), .B(n_19), .Y(n_23) );
OR2x6_ASAP7_75t_SL g24 ( .A(n_22), .B(n_17), .Y(n_24) );
NAND2xp5_ASAP7_75t_L g25 ( .A(n_23), .B(n_22), .Y(n_25) );
CKINVDCx5p33_ASAP7_75t_R g26 ( .A(n_24), .Y(n_26) );
OAI22xp33_ASAP7_75t_L g27 ( .A1(n_26), .A2(n_24), .B1(n_23), .B2(n_13), .Y(n_27) );
INVx1_ASAP7_75t_L g28 ( .A(n_25), .Y(n_28) );
OA22x2_ASAP7_75t_L g29 ( .A1(n_28), .A2(n_25), .B1(n_13), .B2(n_11), .Y(n_29) );
OAI21xp5_ASAP7_75t_L g30 ( .A1(n_27), .A2(n_11), .B(n_12), .Y(n_30) );
NOR2x1_ASAP7_75t_L g31 ( .A(n_27), .B(n_20), .Y(n_31) );
NAND2xp5_ASAP7_75t_L g32 ( .A(n_31), .B(n_14), .Y(n_32) );
NAND2xp5_ASAP7_75t_L g33 ( .A(n_30), .B(n_14), .Y(n_33) );
OR5x1_ASAP7_75t_L g34 ( .A(n_29), .B(n_1), .C(n_3), .D(n_6), .E(n_7), .Y(n_34) );
AND3x2_ASAP7_75t_L g35 ( .A(n_32), .B(n_3), .C(n_6), .Y(n_35) );
NAND4xp25_ASAP7_75t_L g36 ( .A(n_33), .B(n_8), .C(n_9), .D(n_14), .Y(n_36) );
NAND2xp5_ASAP7_75t_L g37 ( .A(n_35), .B(n_14), .Y(n_37) );
AOI22xp5_ASAP7_75t_SL g38 ( .A1(n_37), .A2(n_36), .B1(n_34), .B2(n_9), .Y(n_38) );
endmodule