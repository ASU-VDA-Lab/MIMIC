module real_jpeg_30976_n_30 (n_17, n_8, n_0, n_21, n_212, n_2, n_29, n_209, n_201, n_10, n_9, n_12, n_24, n_6, n_28, n_208, n_207, n_202, n_203, n_23, n_11, n_14, n_211, n_25, n_205, n_7, n_22, n_18, n_3, n_206, n_210, n_5, n_4, n_1, n_26, n_27, n_20, n_19, n_200, n_204, n_16, n_15, n_13, n_30);

input n_17;
input n_8;
input n_0;
input n_21;
input n_212;
input n_2;
input n_29;
input n_209;
input n_201;
input n_10;
input n_9;
input n_12;
input n_24;
input n_6;
input n_28;
input n_208;
input n_207;
input n_202;
input n_203;
input n_23;
input n_11;
input n_14;
input n_211;
input n_25;
input n_205;
input n_7;
input n_22;
input n_18;
input n_3;
input n_206;
input n_210;
input n_5;
input n_4;
input n_1;
input n_26;
input n_27;
input n_20;
input n_19;
input n_200;
input n_204;
input n_16;
input n_15;
input n_13;

output n_30;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_166;
wire n_176;
wire n_194;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_173;
wire n_105;
wire n_115;
wire n_98;
wire n_56;
wire n_184;
wire n_164;
wire n_48;
wire n_140;
wire n_126;
wire n_113;
wire n_120;
wire n_155;
wire n_93;
wire n_141;
wire n_95;
wire n_139;
wire n_33;
wire n_65;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_172;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_148;
wire n_118;
wire n_123;
wire n_116;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_198;
wire n_192;
wire n_100;
wire n_51;
wire n_71;
wire n_90;
wire n_195;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_150;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_92;
wire n_75;
wire n_187;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_179;
wire n_133;
wire n_138;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_0),
.Y(n_70)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_1),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g190 ( 
.A(n_1),
.B(n_98),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_2),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_3),
.B(n_126),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_3),
.B(n_126),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_4),
.B(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_4),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_5),
.B(n_92),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_5),
.B(n_92),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_6),
.Y(n_59)
);

AOI221xp5_ASAP7_75t_L g138 ( 
.A1(n_7),
.A2(n_13),
.B1(n_139),
.B2(n_144),
.C(n_147),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_7),
.B(n_139),
.C(n_144),
.Y(n_150)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_8),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_9),
.B(n_76),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_10),
.B(n_54),
.C(n_195),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_11),
.B(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_12),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_12),
.B(n_164),
.Y(n_175)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_13),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_14),
.B(n_82),
.Y(n_81)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_14),
.Y(n_193)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_16),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_16),
.A2(n_56),
.B1(n_58),
.B2(n_180),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_17),
.B(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_17),
.Y(n_177)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_18),
.Y(n_156)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_19),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_20),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_21),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_22),
.A2(n_32),
.B1(n_42),
.B2(n_43),
.Y(n_31)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_22),
.B(n_47),
.Y(n_198)
);

NOR2x1_ASAP7_75t_L g85 ( 
.A(n_23),
.B(n_86),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_23),
.B(n_86),
.Y(n_191)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_24),
.Y(n_117)
);

AOI322xp5_ASAP7_75t_L g173 ( 
.A1(n_24),
.A2(n_111),
.A3(n_113),
.B1(n_119),
.B2(n_174),
.C1(n_176),
.C2(n_210),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_25),
.B(n_141),
.Y(n_140)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_26),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_26),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_27),
.B(n_87),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_28),
.B(n_99),
.Y(n_98)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_29),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_29),
.B(n_121),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_44),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_41),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_SL g34 ( 
.A(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_38),
.Y(n_137)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_40),
.Y(n_84)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_40),
.Y(n_89)
);

A2O1A1Ixp33_ASAP7_75t_L g45 ( 
.A1(n_42),
.A2(n_46),
.B(n_53),
.C(n_198),
.Y(n_45)
);

HB1xp67_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_52),
.Y(n_47)
);

BUFx2_ASAP7_75t_L g197 ( 
.A(n_48),
.Y(n_197)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_49),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_51),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_51),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_51),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_101),
.B(n_179),
.Y(n_54)
);

NAND4xp25_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_65),
.C(n_90),
.D(n_96),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_64),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_60),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_62),
.Y(n_146)
);

INVx6_ASAP7_75t_L g167 ( 
.A(n_62),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_63),
.Y(n_72)
);

NOR3xp33_ASAP7_75t_SL g65 ( 
.A(n_66),
.B(n_74),
.C(n_79),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

NAND3xp33_ASAP7_75t_L g188 ( 
.A(n_67),
.B(n_189),
.C(n_190),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_68),
.B(n_73),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_68),
.B(n_73),
.Y(n_183)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_71),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_74),
.Y(n_182)
);

OAI322xp33_ASAP7_75t_L g187 ( 
.A1(n_74),
.A2(n_81),
.A3(n_188),
.B1(n_191),
.B2(n_192),
.C1(n_193),
.C2(n_212),
.Y(n_187)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_75),
.Y(n_186)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_77),
.Y(n_99)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

AOI321xp33_ASAP7_75t_L g181 ( 
.A1(n_80),
.A2(n_182),
.A3(n_183),
.B1(n_184),
.B2(n_187),
.C(n_211),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_85),
.Y(n_80)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_82),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_85),
.Y(n_189)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_91),
.A2(n_181),
.B(n_194),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_94),
.Y(n_92)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_97),
.B(n_100),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

AOI31xp67_ASAP7_75t_L g101 ( 
.A1(n_102),
.A2(n_129),
.A3(n_162),
.B(n_169),
.Y(n_101)
);

NOR3xp33_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_118),
.C(n_125),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_103),
.A2(n_170),
.B(n_173),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_111),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

NOR3xp33_ASAP7_75t_L g174 ( 
.A(n_105),
.B(n_125),
.C(n_175),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_106),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_108),
.Y(n_106)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_SL g123 ( 
.A(n_109),
.Y(n_123)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_109),
.Y(n_128)
);

BUFx12f_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_112),
.B(n_117),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_201),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_115),
.B(n_161),
.Y(n_160)
);

BUFx2_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

OA21x2_ASAP7_75t_SL g170 ( 
.A1(n_118),
.A2(n_171),
.B(n_172),
.Y(n_170)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_120),
.B(n_124),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_123),
.Y(n_121)
);

NOR2x1_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_128),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_158),
.C(n_159),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_131),
.A2(n_151),
.B(n_157),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_132),
.A2(n_138),
.B1(n_149),
.B2(n_150),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_135),
.Y(n_133)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_140),
.B(n_148),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_143),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_143),
.Y(n_155)
);

INVx2_ASAP7_75t_SL g148 ( 
.A(n_144),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_206),
.Y(n_144)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_152),
.B(n_156),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_152),
.B(n_156),
.Y(n_157)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_155),
.Y(n_153)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_163),
.B(n_168),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_166),
.Y(n_164)
);

INVx8_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_178),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_186),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_197),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_200),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_202),
.Y(n_122)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_203),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_204),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_205),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_207),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_208),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_209),
.Y(n_165)
);


endmodule