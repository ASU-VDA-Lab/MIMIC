module fake_netlist_6_2592_n_109 (n_16, n_1, n_9, n_8, n_18, n_10, n_6, n_15, n_3, n_14, n_0, n_4, n_13, n_11, n_17, n_12, n_7, n_2, n_5, n_109);

input n_16;
input n_1;
input n_9;
input n_8;
input n_18;
input n_10;
input n_6;
input n_15;
input n_3;
input n_14;
input n_0;
input n_4;
input n_13;
input n_11;
input n_17;
input n_12;
input n_7;
input n_2;
input n_5;

output n_109;

wire n_52;
wire n_91;
wire n_46;
wire n_21;
wire n_88;
wire n_98;
wire n_39;
wire n_63;
wire n_73;
wire n_22;
wire n_68;
wire n_28;
wire n_50;
wire n_49;
wire n_83;
wire n_101;
wire n_77;
wire n_106;
wire n_92;
wire n_42;
wire n_96;
wire n_90;
wire n_24;
wire n_105;
wire n_54;
wire n_102;
wire n_87;
wire n_32;
wire n_66;
wire n_85;
wire n_99;
wire n_78;
wire n_84;
wire n_100;
wire n_23;
wire n_20;
wire n_19;
wire n_47;
wire n_62;
wire n_29;
wire n_75;
wire n_45;
wire n_34;
wire n_70;
wire n_67;
wire n_37;
wire n_33;
wire n_82;
wire n_27;
wire n_38;
wire n_61;
wire n_81;
wire n_59;
wire n_76;
wire n_36;
wire n_26;
wire n_55;
wire n_97;
wire n_94;
wire n_108;
wire n_58;
wire n_64;
wire n_48;
wire n_65;
wire n_25;
wire n_40;
wire n_93;
wire n_80;
wire n_41;
wire n_86;
wire n_104;
wire n_95;
wire n_107;
wire n_71;
wire n_74;
wire n_72;
wire n_89;
wire n_103;
wire n_60;
wire n_35;
wire n_69;
wire n_30;
wire n_79;
wire n_43;
wire n_31;
wire n_57;
wire n_53;
wire n_51;
wire n_44;
wire n_56;

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

CKINVDCx16_ASAP7_75t_R g26 ( 
.A(n_8),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

CKINVDCx5p33_ASAP7_75t_R g29 ( 
.A(n_0),
.Y(n_29)
);

CKINVDCx5p33_ASAP7_75t_R g30 ( 
.A(n_3),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

HB1xp67_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_26),
.B(n_2),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_25),
.Y(n_45)
);

AND2x4_ASAP7_75t_L g46 ( 
.A(n_32),
.B(n_2),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

INVx1_ASAP7_75t_SL g48 ( 
.A(n_41),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

OR2x6_ASAP7_75t_L g51 ( 
.A(n_36),
.B(n_32),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_34),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

AO22x2_ASAP7_75t_L g54 ( 
.A1(n_46),
.A2(n_28),
.B1(n_31),
.B2(n_30),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

AO22x2_ASAP7_75t_L g56 ( 
.A1(n_46),
.A2(n_10),
.B1(n_11),
.B2(n_14),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_49),
.Y(n_57)
);

CKINVDCx5p33_ASAP7_75t_R g58 ( 
.A(n_48),
.Y(n_58)
);

CKINVDCx5p33_ASAP7_75t_R g59 ( 
.A(n_51),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_52),
.B(n_45),
.Y(n_60)
);

AND2x6_ASAP7_75t_SL g61 ( 
.A(n_51),
.B(n_38),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_50),
.Y(n_62)
);

OR2x2_ASAP7_75t_L g63 ( 
.A(n_58),
.B(n_60),
.Y(n_63)
);

A2O1A1Ixp33_ASAP7_75t_L g64 ( 
.A1(n_57),
.A2(n_36),
.B(n_47),
.C(n_44),
.Y(n_64)
);

AOI21xp5_ASAP7_75t_L g65 ( 
.A1(n_62),
.A2(n_57),
.B(n_55),
.Y(n_65)
);

AND2x2_ASAP7_75t_SL g66 ( 
.A(n_61),
.B(n_56),
.Y(n_66)
);

AND2x4_ASAP7_75t_L g67 ( 
.A(n_59),
.B(n_39),
.Y(n_67)
);

HB1xp67_ASAP7_75t_L g68 ( 
.A(n_58),
.Y(n_68)
);

A2O1A1Ixp33_ASAP7_75t_L g69 ( 
.A1(n_64),
.A2(n_63),
.B(n_65),
.C(n_68),
.Y(n_69)
);

AND2x4_ASAP7_75t_L g70 ( 
.A(n_67),
.B(n_37),
.Y(n_70)
);

AO32x2_ASAP7_75t_L g71 ( 
.A1(n_66),
.A2(n_56),
.A3(n_54),
.B1(n_47),
.B2(n_42),
.Y(n_71)
);

NAND2xp33_ASAP7_75t_L g72 ( 
.A(n_67),
.B(n_54),
.Y(n_72)
);

NOR2x1_ASAP7_75t_SL g73 ( 
.A(n_63),
.B(n_53),
.Y(n_73)
);

AO21x2_ASAP7_75t_L g74 ( 
.A1(n_69),
.A2(n_37),
.B(n_43),
.Y(n_74)
);

OA21x2_ASAP7_75t_L g75 ( 
.A1(n_70),
.A2(n_43),
.B(n_35),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_73),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_71),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_L g78 ( 
.A1(n_72),
.A2(n_35),
.B(n_43),
.Y(n_78)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_76),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_74),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_77),
.Y(n_81)
);

AND2x4_ASAP7_75t_SL g82 ( 
.A(n_77),
.B(n_71),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_81),
.Y(n_83)
);

BUFx2_ASAP7_75t_L g84 ( 
.A(n_79),
.Y(n_84)
);

HB1xp67_ASAP7_75t_L g85 ( 
.A(n_79),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_82),
.B(n_75),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_82),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_80),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_83),
.Y(n_89)
);

INVx1_ASAP7_75t_SL g90 ( 
.A(n_84),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_85),
.B(n_76),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_88),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_90),
.Y(n_93)
);

NOR2x1_ASAP7_75t_L g94 ( 
.A(n_92),
.B(n_84),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_89),
.B(n_87),
.Y(n_95)
);

INVx1_ASAP7_75t_SL g96 ( 
.A(n_91),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_89),
.Y(n_97)
);

AND2x4_ASAP7_75t_L g98 ( 
.A(n_93),
.B(n_86),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_97),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_95),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_96),
.A2(n_76),
.B1(n_78),
.B2(n_74),
.Y(n_101)
);

HB1xp67_ASAP7_75t_L g102 ( 
.A(n_100),
.Y(n_102)
);

NOR3xp33_ASAP7_75t_SL g103 ( 
.A(n_99),
.B(n_78),
.C(n_94),
.Y(n_103)
);

OR2x2_ASAP7_75t_L g104 ( 
.A(n_98),
.B(n_80),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_102),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_105),
.A2(n_101),
.B1(n_103),
.B2(n_104),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_106),
.A2(n_74),
.B(n_86),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_107),
.B(n_17),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_108),
.A2(n_74),
.B1(n_75),
.B2(n_18),
.Y(n_109)
);


endmodule