module fake_jpeg_3445_n_690 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_690);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_690;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_686;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_678;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_543;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_672;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_688;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_689;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_195;
wire n_450;
wire n_557;
wire n_681;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_668;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_682;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_679;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_676;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_670;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_683;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_674;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_684;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_680;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_687;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_673;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_665;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_677;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_671;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_669;
wire n_524;
wire n_402;
wire n_563;
wire n_685;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_675;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_19),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_18),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_19),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_18),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_18),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

BUFx16f_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_14),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_7),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_2),
.B(n_16),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_5),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_8),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_1),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_8),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g50 ( 
.A(n_19),
.Y(n_50)
);

BUFx4f_ASAP7_75t_L g51 ( 
.A(n_8),
.Y(n_51)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_2),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_8),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_1),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_15),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_5),
.Y(n_56)
);

INVx13_ASAP7_75t_L g57 ( 
.A(n_2),
.Y(n_57)
);

BUFx2_ASAP7_75t_L g58 ( 
.A(n_19),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_20),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_59),
.Y(n_151)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_60),
.Y(n_138)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_61),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_36),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_62),
.B(n_65),
.Y(n_136)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_63),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_20),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_64),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_42),
.B(n_10),
.Y(n_65)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_66),
.Y(n_148)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_36),
.Y(n_67)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_67),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_42),
.B(n_23),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_68),
.B(n_92),
.Y(n_135)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_53),
.Y(n_69)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_69),
.Y(n_149)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_36),
.Y(n_70)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_70),
.Y(n_142)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_53),
.Y(n_71)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_71),
.Y(n_153)
);

INVx6_ASAP7_75t_SL g72 ( 
.A(n_57),
.Y(n_72)
);

CKINVDCx6p67_ASAP7_75t_R g216 ( 
.A(n_72),
.Y(n_216)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_41),
.Y(n_73)
);

BUFx2_ASAP7_75t_L g150 ( 
.A(n_73),
.Y(n_150)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_21),
.Y(n_74)
);

INVx4_ASAP7_75t_SL g202 ( 
.A(n_74),
.Y(n_202)
);

BUFx5_ASAP7_75t_L g75 ( 
.A(n_23),
.Y(n_75)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_75),
.Y(n_170)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_21),
.Y(n_76)
);

INVx4_ASAP7_75t_SL g222 ( 
.A(n_76),
.Y(n_222)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_51),
.Y(n_77)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_77),
.Y(n_159)
);

BUFx2_ASAP7_75t_L g78 ( 
.A(n_58),
.Y(n_78)
);

BUFx2_ASAP7_75t_L g161 ( 
.A(n_78),
.Y(n_161)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_51),
.Y(n_79)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_79),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_20),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_80),
.Y(n_160)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_45),
.Y(n_81)
);

INVx5_ASAP7_75t_L g171 ( 
.A(n_81),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_20),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_82),
.Y(n_180)
);

BUFx5_ASAP7_75t_L g83 ( 
.A(n_29),
.Y(n_83)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_83),
.Y(n_185)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_51),
.Y(n_84)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_84),
.Y(n_187)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_54),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g232 ( 
.A(n_85),
.Y(n_232)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_24),
.Y(n_86)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_86),
.Y(n_158)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_45),
.Y(n_87)
);

INVx5_ASAP7_75t_L g183 ( 
.A(n_87),
.Y(n_183)
);

INVx4_ASAP7_75t_SL g88 ( 
.A(n_28),
.Y(n_88)
);

OR2x2_ASAP7_75t_L g174 ( 
.A(n_88),
.B(n_128),
.Y(n_174)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_32),
.Y(n_89)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_89),
.Y(n_178)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_24),
.Y(n_90)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_90),
.Y(n_206)
);

BUFx12f_ASAP7_75t_L g91 ( 
.A(n_21),
.Y(n_91)
);

INVx8_ASAP7_75t_L g168 ( 
.A(n_91),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_50),
.B(n_10),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_44),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_93),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_33),
.B(n_10),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_94),
.B(n_100),
.Y(n_144)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_45),
.Y(n_95)
);

INVx5_ASAP7_75t_L g199 ( 
.A(n_95),
.Y(n_199)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_24),
.Y(n_96)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_96),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_44),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_97),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_44),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_98),
.Y(n_205)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_54),
.Y(n_99)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_99),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_33),
.B(n_10),
.Y(n_100)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_32),
.Y(n_101)
);

INVx4_ASAP7_75t_L g215 ( 
.A(n_101),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_56),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_102),
.Y(n_226)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_22),
.Y(n_103)
);

INVx5_ASAP7_75t_L g214 ( 
.A(n_103),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_56),
.Y(n_104)
);

INVx6_ASAP7_75t_L g154 ( 
.A(n_104),
.Y(n_154)
);

INVx13_ASAP7_75t_L g105 ( 
.A(n_57),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_105),
.Y(n_207)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_58),
.Y(n_106)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_106),
.Y(n_137)
);

INVx11_ASAP7_75t_L g107 ( 
.A(n_45),
.Y(n_107)
);

INVx11_ASAP7_75t_L g217 ( 
.A(n_107),
.Y(n_217)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_32),
.Y(n_108)
);

INVx4_ASAP7_75t_L g223 ( 
.A(n_108),
.Y(n_223)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_30),
.Y(n_109)
);

INVx4_ASAP7_75t_L g231 ( 
.A(n_109),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_56),
.Y(n_110)
);

INVx6_ASAP7_75t_L g203 ( 
.A(n_110),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_54),
.Y(n_111)
);

INVx6_ASAP7_75t_L g221 ( 
.A(n_111),
.Y(n_221)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_58),
.Y(n_112)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_112),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_25),
.B(n_17),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_113),
.B(n_129),
.Y(n_169)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_22),
.Y(n_114)
);

INVx5_ASAP7_75t_L g224 ( 
.A(n_114),
.Y(n_224)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_30),
.Y(n_115)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_115),
.Y(n_195)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_22),
.Y(n_116)
);

INVx6_ASAP7_75t_L g227 ( 
.A(n_116),
.Y(n_227)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_58),
.Y(n_117)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_117),
.Y(n_189)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_51),
.Y(n_118)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_118),
.Y(n_218)
);

BUFx12_ASAP7_75t_L g119 ( 
.A(n_57),
.Y(n_119)
);

BUFx12_ASAP7_75t_L g220 ( 
.A(n_119),
.Y(n_220)
);

BUFx5_ASAP7_75t_L g120 ( 
.A(n_29),
.Y(n_120)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_120),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_30),
.A2(n_17),
.B1(n_16),
.B2(n_15),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_121),
.A2(n_31),
.B1(n_38),
.B2(n_48),
.Y(n_140)
);

BUFx5_ASAP7_75t_L g122 ( 
.A(n_29),
.Y(n_122)
);

NAND2xp33_ASAP7_75t_SL g164 ( 
.A(n_122),
.B(n_126),
.Y(n_164)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_41),
.Y(n_123)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_123),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_34),
.Y(n_124)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_124),
.Y(n_210)
);

INVx8_ASAP7_75t_L g125 ( 
.A(n_28),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_125),
.B(n_127),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g126 ( 
.A(n_34),
.Y(n_126)
);

INVx6_ASAP7_75t_L g127 ( 
.A(n_41),
.Y(n_127)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_35),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_34),
.Y(n_129)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_28),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_130),
.B(n_131),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_28),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_28),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_132),
.B(n_0),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_88),
.A2(n_52),
.B1(n_38),
.B2(n_31),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_134),
.A2(n_139),
.B1(n_143),
.B2(n_145),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_93),
.A2(n_55),
.B1(n_26),
.B2(n_37),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_140),
.A2(n_198),
.B1(n_211),
.B2(n_137),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_70),
.B(n_55),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_141),
.B(n_147),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_97),
.A2(n_25),
.B1(n_26),
.B2(n_37),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_98),
.A2(n_48),
.B1(n_52),
.B2(n_49),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_78),
.B(n_46),
.Y(n_147)
);

OA22x2_ASAP7_75t_L g152 ( 
.A1(n_123),
.A2(n_127),
.B1(n_99),
.B2(n_85),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_152),
.B(n_208),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_74),
.B(n_76),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_157),
.B(n_165),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_102),
.A2(n_52),
.B1(n_49),
.B2(n_47),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_162),
.A2(n_163),
.B1(n_173),
.B2(n_175),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_89),
.A2(n_101),
.B1(n_128),
.B2(n_108),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_74),
.B(n_47),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_76),
.B(n_40),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_172),
.B(n_177),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_104),
.A2(n_46),
.B1(n_40),
.B2(n_27),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_107),
.A2(n_27),
.B1(n_35),
.B2(n_43),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_103),
.A2(n_43),
.B1(n_35),
.B2(n_21),
.Y(n_176)
);

OAI22xp33_ASAP7_75t_SL g313 ( 
.A1(n_176),
.A2(n_229),
.B1(n_181),
.B2(n_204),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_114),
.B(n_11),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_116),
.A2(n_43),
.B1(n_21),
.B2(n_11),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_181),
.A2(n_182),
.B1(n_190),
.B2(n_191),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_110),
.A2(n_17),
.B1(n_16),
.B2(n_15),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_91),
.B(n_17),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_184),
.B(n_194),
.Y(n_293)
);

AND2x2_ASAP7_75t_SL g186 ( 
.A(n_91),
.B(n_0),
.Y(n_186)
);

NAND2x1_ASAP7_75t_SL g310 ( 
.A(n_186),
.B(n_148),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_59),
.A2(n_15),
.B1(n_14),
.B2(n_13),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_126),
.A2(n_13),
.B1(n_12),
.B2(n_11),
.Y(n_191)
);

CKINVDCx14_ASAP7_75t_SL g193 ( 
.A(n_105),
.Y(n_193)
);

INVx11_ASAP7_75t_L g279 ( 
.A(n_193),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_125),
.B(n_13),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_60),
.B(n_12),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_197),
.B(n_212),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_64),
.A2(n_12),
.B1(n_1),
.B2(n_2),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_81),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g252 ( 
.A1(n_204),
.A2(n_129),
.B1(n_132),
.B2(n_6),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_80),
.B(n_3),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_209),
.B(n_6),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_82),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_87),
.B(n_3),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_95),
.B(n_3),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_213),
.B(n_219),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_131),
.B(n_4),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_124),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_229)
);

OA22x2_ASAP7_75t_L g230 ( 
.A1(n_111),
.A2(n_4),
.B1(n_6),
.B2(n_9),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_230),
.A2(n_202),
.B1(n_222),
.B2(n_191),
.Y(n_305)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_159),
.Y(n_233)
);

BUFx2_ASAP7_75t_L g365 ( 
.A(n_233),
.Y(n_365)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_166),
.Y(n_234)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_234),
.Y(n_321)
);

INVx13_ASAP7_75t_L g235 ( 
.A(n_216),
.Y(n_235)
);

INVx1_ASAP7_75t_SL g324 ( 
.A(n_235),
.Y(n_324)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_188),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g338 ( 
.A(n_236),
.Y(n_338)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_187),
.Y(n_237)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_237),
.Y(n_322)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_161),
.Y(n_238)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_238),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_L g323 ( 
.A1(n_239),
.A2(n_271),
.B1(n_301),
.B2(n_305),
.Y(n_323)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_218),
.Y(n_240)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_240),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_193),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_241),
.B(n_251),
.Y(n_343)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_179),
.Y(n_242)
);

HB1xp67_ASAP7_75t_L g326 ( 
.A(n_242),
.Y(n_326)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_189),
.Y(n_243)
);

HB1xp67_ASAP7_75t_L g344 ( 
.A(n_243),
.Y(n_344)
);

AND2x2_ASAP7_75t_SL g244 ( 
.A(n_186),
.B(n_169),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_244),
.B(n_222),
.C(n_202),
.Y(n_325)
);

INVx6_ASAP7_75t_L g247 ( 
.A(n_188),
.Y(n_247)
);

INVx4_ASAP7_75t_L g320 ( 
.A(n_247),
.Y(n_320)
);

INVx3_ASAP7_75t_L g248 ( 
.A(n_138),
.Y(n_248)
);

INVx4_ASAP7_75t_L g348 ( 
.A(n_248),
.Y(n_348)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_200),
.Y(n_249)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_249),
.Y(n_355)
);

INVx2_ASAP7_75t_SL g250 ( 
.A(n_161),
.Y(n_250)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_250),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_216),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g331 ( 
.A(n_252),
.Y(n_331)
);

INVx3_ASAP7_75t_L g253 ( 
.A(n_138),
.Y(n_253)
);

INVx3_ASAP7_75t_L g334 ( 
.A(n_253),
.Y(n_334)
);

INVx3_ASAP7_75t_L g254 ( 
.A(n_171),
.Y(n_254)
);

BUFx3_ASAP7_75t_L g340 ( 
.A(n_254),
.Y(n_340)
);

AOI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_155),
.A2(n_119),
.B1(n_6),
.B2(n_9),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g342 ( 
.A(n_255),
.Y(n_342)
);

INVx13_ASAP7_75t_L g256 ( 
.A(n_216),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g370 ( 
.A(n_256),
.Y(n_370)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_174),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_257),
.B(n_280),
.Y(n_349)
);

INVx3_ASAP7_75t_L g258 ( 
.A(n_171),
.Y(n_258)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_258),
.Y(n_366)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_142),
.Y(n_259)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_259),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_SL g363 ( 
.A(n_260),
.B(n_265),
.Y(n_363)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_196),
.Y(n_261)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_261),
.Y(n_380)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_210),
.Y(n_262)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_262),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_174),
.Y(n_265)
);

BUFx2_ASAP7_75t_L g266 ( 
.A(n_142),
.Y(n_266)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_266),
.Y(n_367)
);

NAND2x1p5_ASAP7_75t_L g267 ( 
.A(n_186),
.B(n_119),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_L g381 ( 
.A1(n_267),
.A2(n_278),
.B(n_299),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_155),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g374 ( 
.A(n_268),
.B(n_274),
.Y(n_374)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_201),
.Y(n_269)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_269),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_230),
.A2(n_9),
.B1(n_135),
.B2(n_152),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_144),
.B(n_136),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_272),
.B(n_278),
.Y(n_352)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_192),
.Y(n_273)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_273),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_221),
.Y(n_274)
);

BUFx6f_ASAP7_75t_L g275 ( 
.A(n_196),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_275),
.Y(n_329)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_192),
.Y(n_276)
);

AND2x2_ASAP7_75t_L g328 ( 
.A(n_276),
.B(n_285),
.Y(n_328)
);

AOI22xp33_ASAP7_75t_SL g277 ( 
.A1(n_185),
.A2(n_9),
.B1(n_152),
.B2(n_225),
.Y(n_277)
);

AOI22xp33_ASAP7_75t_SL g337 ( 
.A1(n_277),
.A2(n_284),
.B1(n_295),
.B2(n_300),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_133),
.B(n_9),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_221),
.Y(n_280)
);

CKINVDCx16_ASAP7_75t_R g281 ( 
.A(n_207),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_281),
.B(n_283),
.Y(n_354)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_195),
.Y(n_283)
);

AOI22xp33_ASAP7_75t_SL g284 ( 
.A1(n_185),
.A2(n_150),
.B1(n_178),
.B2(n_176),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_146),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_149),
.Y(n_286)
);

AND2x2_ASAP7_75t_L g336 ( 
.A(n_286),
.B(n_287),
.Y(n_336)
);

INVx4_ASAP7_75t_L g287 ( 
.A(n_183),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_153),
.Y(n_288)
);

OR2x2_ASAP7_75t_L g347 ( 
.A(n_288),
.B(n_289),
.Y(n_347)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_178),
.Y(n_289)
);

FAx1_ASAP7_75t_SL g290 ( 
.A(n_164),
.B(n_229),
.CI(n_230),
.CON(n_290),
.SN(n_290)
);

NOR2xp33_ASAP7_75t_SL g335 ( 
.A(n_290),
.B(n_312),
.Y(n_335)
);

BUFx6f_ASAP7_75t_L g292 ( 
.A(n_205),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_292),
.Y(n_369)
);

INVx8_ASAP7_75t_L g295 ( 
.A(n_227),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_158),
.Y(n_296)
);

OR2x2_ASAP7_75t_L g382 ( 
.A(n_296),
.B(n_304),
.Y(n_382)
);

BUFx2_ASAP7_75t_L g297 ( 
.A(n_148),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_297),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_134),
.B(n_206),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_298),
.B(n_299),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_158),
.B(n_206),
.Y(n_299)
);

BUFx6f_ASAP7_75t_L g300 ( 
.A(n_205),
.Y(n_300)
);

AOI22xp33_ASAP7_75t_L g301 ( 
.A1(n_228),
.A2(n_226),
.B1(n_156),
.B2(n_151),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_154),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_302),
.B(n_303),
.Y(n_373)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_228),
.Y(n_303)
);

INVx4_ASAP7_75t_SL g304 ( 
.A(n_220),
.Y(n_304)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_154),
.Y(n_306)
);

AOI22xp33_ASAP7_75t_SL g357 ( 
.A1(n_306),
.A2(n_307),
.B1(n_309),
.B2(n_314),
.Y(n_357)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_203),
.Y(n_307)
);

CKINVDCx16_ASAP7_75t_R g308 ( 
.A(n_150),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_308),
.B(n_310),
.Y(n_372)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_203),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_183),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_313),
.A2(n_318),
.B1(n_214),
.B2(n_224),
.Y(n_332)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_215),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_231),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_SL g378 ( 
.A(n_315),
.B(n_316),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_199),
.Y(n_316)
);

INVx3_ASAP7_75t_L g317 ( 
.A(n_199),
.Y(n_317)
);

AOI22xp33_ASAP7_75t_L g364 ( 
.A1(n_317),
.A2(n_319),
.B1(n_217),
.B2(n_250),
.Y(n_364)
);

OAI22xp33_ASAP7_75t_L g318 ( 
.A1(n_175),
.A2(n_163),
.B1(n_226),
.B2(n_160),
.Y(n_318)
);

BUFx2_ASAP7_75t_L g319 ( 
.A(n_167),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_325),
.B(n_288),
.Y(n_392)
);

AOI21xp5_ASAP7_75t_L g327 ( 
.A1(n_298),
.A2(n_167),
.B(n_215),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_L g431 ( 
.A1(n_327),
.A2(n_368),
.B(n_372),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_244),
.B(n_223),
.C(n_231),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_330),
.B(n_339),
.C(n_371),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_332),
.A2(n_345),
.B1(n_359),
.B2(n_361),
.Y(n_385)
);

MAJx2_ASAP7_75t_L g339 ( 
.A(n_244),
.B(n_220),
.C(n_223),
.Y(n_339)
);

AO22x2_ASAP7_75t_L g341 ( 
.A1(n_263),
.A2(n_214),
.B1(n_224),
.B2(n_170),
.Y(n_341)
);

AND2x2_ASAP7_75t_L g412 ( 
.A(n_341),
.B(n_381),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_271),
.A2(n_151),
.B1(n_156),
.B2(n_160),
.Y(n_345)
);

AOI32xp33_ASAP7_75t_L g346 ( 
.A1(n_311),
.A2(n_294),
.A3(n_293),
.B1(n_257),
.B2(n_310),
.Y(n_346)
);

A2O1A1Ixp33_ASAP7_75t_L g406 ( 
.A1(n_346),
.A2(n_235),
.B(n_256),
.C(n_237),
.Y(n_406)
);

AND2x4_ASAP7_75t_L g356 ( 
.A(n_267),
.B(n_170),
.Y(n_356)
);

INVx1_ASAP7_75t_SL g432 ( 
.A(n_356),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_L g359 ( 
.A1(n_239),
.A2(n_180),
.B1(n_227),
.B2(n_232),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_L g361 ( 
.A1(n_291),
.A2(n_180),
.B1(n_232),
.B2(n_168),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_291),
.A2(n_168),
.B1(n_217),
.B2(n_220),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_362),
.A2(n_375),
.B1(n_304),
.B2(n_317),
.Y(n_390)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_364),
.Y(n_388)
);

AOI21xp5_ASAP7_75t_L g368 ( 
.A1(n_267),
.A2(n_291),
.B(n_318),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g371 ( 
.A(n_269),
.B(n_245),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_L g375 ( 
.A1(n_282),
.A2(n_246),
.B1(n_305),
.B2(n_264),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_352),
.B(n_260),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_383),
.B(n_396),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_368),
.A2(n_290),
.B1(n_270),
.B2(n_272),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g433 ( 
.A1(n_384),
.A2(n_386),
.B1(n_387),
.B2(n_418),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_L g386 ( 
.A1(n_360),
.A2(n_290),
.B1(n_306),
.B2(n_302),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_L g387 ( 
.A1(n_360),
.A2(n_307),
.B1(n_309),
.B2(n_247),
.Y(n_387)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_351),
.Y(n_389)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_389),
.Y(n_449)
);

AND2x2_ASAP7_75t_L g460 ( 
.A(n_390),
.B(n_429),
.Y(n_460)
);

BUFx3_ASAP7_75t_L g391 ( 
.A(n_370),
.Y(n_391)
);

INVx4_ASAP7_75t_L g442 ( 
.A(n_391),
.Y(n_442)
);

XOR2xp5_ASAP7_75t_L g445 ( 
.A(n_392),
.B(n_420),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_371),
.B(n_289),
.Y(n_393)
);

INVxp67_ASAP7_75t_L g454 ( 
.A(n_393),
.Y(n_454)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_358),
.Y(n_394)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_394),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_346),
.B(n_266),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_395),
.B(n_398),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_352),
.B(n_262),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_SL g397 ( 
.A1(n_342),
.A2(n_248),
.B1(n_258),
.B2(n_253),
.Y(n_397)
);

OAI21xp5_ASAP7_75t_SL g436 ( 
.A1(n_397),
.A2(n_324),
.B(n_382),
.Y(n_436)
);

AOI32xp33_ASAP7_75t_L g398 ( 
.A1(n_381),
.A2(n_287),
.A3(n_296),
.B1(n_273),
.B2(n_276),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_SL g399 ( 
.A(n_363),
.B(n_285),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_399),
.B(n_401),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_326),
.B(n_314),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_358),
.Y(n_402)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_402),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_377),
.B(n_286),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_403),
.B(n_409),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_344),
.B(n_319),
.Y(n_404)
);

INVxp67_ASAP7_75t_SL g472 ( 
.A(n_404),
.Y(n_472)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_323),
.A2(n_249),
.B1(n_234),
.B2(n_233),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_L g438 ( 
.A1(n_405),
.A2(n_416),
.B1(n_423),
.B2(n_425),
.Y(n_438)
);

OAI21xp5_ASAP7_75t_L g453 ( 
.A1(n_406),
.A2(n_336),
.B(n_324),
.Y(n_453)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_351),
.Y(n_407)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_407),
.Y(n_446)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_350),
.Y(n_408)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_408),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_377),
.B(n_240),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_350),
.Y(n_410)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_410),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_339),
.B(n_254),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_411),
.B(n_413),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_330),
.B(n_238),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_353),
.Y(n_414)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_414),
.Y(n_452)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_353),
.Y(n_415)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_415),
.Y(n_468)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_345),
.A2(n_236),
.B1(n_292),
.B2(n_261),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_373),
.Y(n_417)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_417),
.Y(n_469)
);

OAI22xp5_ASAP7_75t_SL g418 ( 
.A1(n_332),
.A2(n_275),
.B1(n_300),
.B2(n_295),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_SL g419 ( 
.A(n_335),
.B(n_250),
.Y(n_419)
);

MAJx2_ASAP7_75t_L g470 ( 
.A(n_419),
.B(n_421),
.C(n_376),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_349),
.B(n_297),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_335),
.B(n_279),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_328),
.Y(n_422)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_422),
.Y(n_465)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_356),
.A2(n_279),
.B1(n_327),
.B2(n_362),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_328),
.Y(n_424)
);

INVx1_ASAP7_75t_SL g443 ( 
.A(n_424),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_356),
.A2(n_342),
.B1(n_331),
.B2(n_341),
.Y(n_425)
);

INVx3_ASAP7_75t_L g426 ( 
.A(n_320),
.Y(n_426)
);

BUFx2_ASAP7_75t_L g473 ( 
.A(n_426),
.Y(n_473)
);

OAI22xp5_ASAP7_75t_SL g427 ( 
.A1(n_337),
.A2(n_341),
.B1(n_331),
.B2(n_372),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_L g435 ( 
.A1(n_427),
.A2(n_341),
.B1(n_382),
.B2(n_378),
.Y(n_435)
);

CKINVDCx14_ASAP7_75t_R g428 ( 
.A(n_356),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_428),
.Y(n_444)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_328),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_SL g430 ( 
.A(n_374),
.B(n_325),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_430),
.Y(n_462)
);

NAND2xp33_ASAP7_75t_SL g455 ( 
.A(n_431),
.B(n_336),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_L g492 ( 
.A1(n_435),
.A2(n_459),
.B1(n_464),
.B2(n_471),
.Y(n_492)
);

INVxp67_ASAP7_75t_L g496 ( 
.A(n_436),
.Y(n_496)
);

OAI21xp5_ASAP7_75t_SL g437 ( 
.A1(n_431),
.A2(n_343),
.B(n_354),
.Y(n_437)
);

AOI21xp5_ASAP7_75t_L g494 ( 
.A1(n_437),
.A2(n_450),
.B(n_455),
.Y(n_494)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_412),
.A2(n_341),
.B1(n_378),
.B2(n_369),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_L g487 ( 
.A1(n_440),
.A2(n_441),
.B1(n_451),
.B2(n_466),
.Y(n_487)
);

OAI22xp5_ASAP7_75t_L g441 ( 
.A1(n_412),
.A2(n_347),
.B1(n_369),
.B2(n_329),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_SL g447 ( 
.A1(n_427),
.A2(n_329),
.B1(n_334),
.B2(n_366),
.Y(n_447)
);

INVx1_ASAP7_75t_SL g507 ( 
.A(n_447),
.Y(n_507)
);

OAI21xp5_ASAP7_75t_SL g450 ( 
.A1(n_432),
.A2(n_347),
.B(n_357),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_L g451 ( 
.A1(n_412),
.A2(n_320),
.B1(n_380),
.B2(n_334),
.Y(n_451)
);

HB1xp67_ASAP7_75t_L g503 ( 
.A(n_453),
.Y(n_503)
);

OAI22xp5_ASAP7_75t_SL g459 ( 
.A1(n_385),
.A2(n_380),
.B1(n_366),
.B2(n_338),
.Y(n_459)
);

OAI22xp5_ASAP7_75t_SL g464 ( 
.A1(n_385),
.A2(n_338),
.B1(n_348),
.B2(n_336),
.Y(n_464)
);

AOI22xp5_ASAP7_75t_L g466 ( 
.A1(n_386),
.A2(n_348),
.B1(n_376),
.B2(n_338),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_470),
.B(n_475),
.Y(n_479)
);

OAI22xp5_ASAP7_75t_SL g471 ( 
.A1(n_390),
.A2(n_425),
.B1(n_411),
.B2(n_423),
.Y(n_471)
);

MAJx2_ASAP7_75t_L g474 ( 
.A(n_400),
.B(n_379),
.C(n_355),
.Y(n_474)
);

XOR2xp5_ASAP7_75t_L g501 ( 
.A(n_474),
.B(n_398),
.Y(n_501)
);

AOI21xp5_ASAP7_75t_L g475 ( 
.A1(n_432),
.A2(n_370),
.B(n_367),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_446),
.Y(n_476)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_476),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_SL g477 ( 
.A(n_462),
.B(n_396),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_477),
.B(n_481),
.Y(n_537)
);

XNOR2xp5_ASAP7_75t_L g478 ( 
.A(n_445),
.B(n_400),
.Y(n_478)
);

XOR2xp5_ASAP7_75t_L g544 ( 
.A(n_478),
.B(n_486),
.Y(n_544)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_456),
.Y(n_480)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_480),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_SL g481 ( 
.A(n_462),
.B(n_399),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_454),
.B(n_417),
.Y(n_482)
);

CKINVDCx16_ASAP7_75t_R g523 ( 
.A(n_482),
.Y(n_523)
);

CKINVDCx20_ASAP7_75t_R g483 ( 
.A(n_467),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g529 ( 
.A(n_483),
.Y(n_529)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_474),
.B(n_392),
.C(n_413),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_484),
.B(n_485),
.C(n_489),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_474),
.B(n_384),
.C(n_383),
.Y(n_485)
);

XNOR2xp5_ASAP7_75t_L g486 ( 
.A(n_445),
.B(n_430),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_458),
.B(n_409),
.Y(n_488)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_488),
.Y(n_549)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_463),
.B(n_406),
.C(n_420),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_463),
.B(n_458),
.C(n_437),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_490),
.B(n_509),
.C(n_443),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_SL g491 ( 
.A(n_461),
.B(n_419),
.Y(n_491)
);

CKINVDCx20_ASAP7_75t_R g517 ( 
.A(n_491),
.Y(n_517)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_446),
.Y(n_493)
);

INVxp67_ASAP7_75t_L g533 ( 
.A(n_493),
.Y(n_533)
);

CKINVDCx20_ASAP7_75t_R g495 ( 
.A(n_467),
.Y(n_495)
);

CKINVDCx20_ASAP7_75t_R g536 ( 
.A(n_495),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_461),
.B(n_403),
.Y(n_497)
);

CKINVDCx20_ASAP7_75t_R g538 ( 
.A(n_497),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_465),
.B(n_402),
.Y(n_498)
);

CKINVDCx20_ASAP7_75t_R g542 ( 
.A(n_498),
.Y(n_542)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_434),
.Y(n_499)
);

HB1xp67_ASAP7_75t_L g520 ( 
.A(n_499),
.Y(n_520)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_434),
.Y(n_500)
);

OAI22xp5_ASAP7_75t_L g519 ( 
.A1(n_500),
.A2(n_502),
.B1(n_504),
.B2(n_505),
.Y(n_519)
);

XNOR2xp5_ASAP7_75t_SL g518 ( 
.A(n_501),
.B(n_457),
.Y(n_518)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_456),
.Y(n_502)
);

AOI22xp5_ASAP7_75t_L g504 ( 
.A1(n_471),
.A2(n_418),
.B1(n_405),
.B2(n_387),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_439),
.Y(n_505)
);

CKINVDCx20_ASAP7_75t_R g506 ( 
.A(n_473),
.Y(n_506)
);

OAI21xp5_ASAP7_75t_SL g551 ( 
.A1(n_506),
.A2(n_449),
.B(n_389),
.Y(n_551)
);

AOI22xp5_ASAP7_75t_L g508 ( 
.A1(n_438),
.A2(n_421),
.B1(n_416),
.B2(n_394),
.Y(n_508)
);

OAI22xp5_ASAP7_75t_L g524 ( 
.A1(n_508),
.A2(n_510),
.B1(n_511),
.B2(n_513),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g509 ( 
.A(n_457),
.B(n_429),
.C(n_424),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_469),
.B(n_391),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_469),
.B(n_340),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_439),
.Y(n_512)
);

OAI22xp5_ASAP7_75t_L g553 ( 
.A1(n_512),
.A2(n_410),
.B1(n_365),
.B2(n_426),
.Y(n_553)
);

CKINVDCx16_ASAP7_75t_R g513 ( 
.A(n_473),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_448),
.Y(n_514)
);

OAI22xp5_ASAP7_75t_L g528 ( 
.A1(n_514),
.A2(n_515),
.B1(n_443),
.B2(n_448),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_SL g515 ( 
.A(n_472),
.B(n_415),
.Y(n_515)
);

XNOR2xp5_ASAP7_75t_L g516 ( 
.A(n_478),
.B(n_470),
.Y(n_516)
);

XOR2xp5_ASAP7_75t_L g562 ( 
.A(n_516),
.B(n_518),
.Y(n_562)
);

AOI22xp5_ASAP7_75t_L g522 ( 
.A1(n_487),
.A2(n_438),
.B1(n_435),
.B2(n_460),
.Y(n_522)
);

OAI22xp5_ASAP7_75t_L g563 ( 
.A1(n_522),
.A2(n_525),
.B1(n_532),
.B2(n_508),
.Y(n_563)
);

AOI22xp5_ASAP7_75t_L g525 ( 
.A1(n_487),
.A2(n_460),
.B1(n_440),
.B2(n_433),
.Y(n_525)
);

XNOR2xp5_ASAP7_75t_L g555 ( 
.A(n_526),
.B(n_544),
.Y(n_555)
);

INVxp67_ASAP7_75t_SL g559 ( 
.A(n_528),
.Y(n_559)
);

OAI22xp5_ASAP7_75t_SL g530 ( 
.A1(n_492),
.A2(n_433),
.B1(n_447),
.B2(n_460),
.Y(n_530)
);

AOI22xp5_ASAP7_75t_L g560 ( 
.A1(n_530),
.A2(n_540),
.B1(n_550),
.B2(n_519),
.Y(n_560)
);

MAJIxp5_ASAP7_75t_L g531 ( 
.A(n_484),
.B(n_444),
.C(n_465),
.Y(n_531)
);

MAJIxp5_ASAP7_75t_L g565 ( 
.A(n_531),
.B(n_535),
.C(n_546),
.Y(n_565)
);

AOI22xp5_ASAP7_75t_L g532 ( 
.A1(n_492),
.A2(n_453),
.B1(n_441),
.B2(n_464),
.Y(n_532)
);

MAJIxp5_ASAP7_75t_L g535 ( 
.A(n_486),
.B(n_444),
.C(n_470),
.Y(n_535)
);

XNOR2xp5_ASAP7_75t_L g539 ( 
.A(n_485),
.B(n_455),
.Y(n_539)
);

XOR2xp5_ASAP7_75t_L g568 ( 
.A(n_539),
.B(n_541),
.Y(n_568)
);

OAI22xp5_ASAP7_75t_SL g540 ( 
.A1(n_483),
.A2(n_466),
.B1(n_475),
.B2(n_468),
.Y(n_540)
);

XNOR2xp5_ASAP7_75t_SL g541 ( 
.A(n_490),
.B(n_450),
.Y(n_541)
);

XNOR2xp5_ASAP7_75t_L g543 ( 
.A(n_489),
.B(n_422),
.Y(n_543)
);

XOR2xp5_ASAP7_75t_L g574 ( 
.A(n_543),
.B(n_545),
.Y(n_574)
);

XNOR2x1_ASAP7_75t_SL g545 ( 
.A(n_509),
.B(n_451),
.Y(n_545)
);

MAJIxp5_ASAP7_75t_L g546 ( 
.A(n_501),
.B(n_468),
.C(n_452),
.Y(n_546)
);

MAJIxp5_ASAP7_75t_L g547 ( 
.A(n_503),
.B(n_452),
.C(n_408),
.Y(n_547)
);

MAJIxp5_ASAP7_75t_L g569 ( 
.A(n_547),
.B(n_548),
.C(n_514),
.Y(n_569)
);

MAJIxp5_ASAP7_75t_L g548 ( 
.A(n_494),
.B(n_414),
.C(n_407),
.Y(n_548)
);

OAI22xp5_ASAP7_75t_SL g550 ( 
.A1(n_495),
.A2(n_459),
.B1(n_449),
.B2(n_388),
.Y(n_550)
);

OAI21xp5_ASAP7_75t_SL g564 ( 
.A1(n_551),
.A2(n_552),
.B(n_479),
.Y(n_564)
);

OAI21xp5_ASAP7_75t_SL g552 ( 
.A1(n_494),
.A2(n_436),
.B(n_397),
.Y(n_552)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_553),
.Y(n_554)
);

XNOR2xp5_ASAP7_75t_L g588 ( 
.A(n_555),
.B(n_569),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_537),
.B(n_477),
.Y(n_556)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_556),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_533),
.B(n_498),
.Y(n_557)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_557),
.Y(n_605)
);

INVxp67_ASAP7_75t_L g558 ( 
.A(n_551),
.Y(n_558)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_558),
.Y(n_608)
);

OAI22xp5_ASAP7_75t_SL g586 ( 
.A1(n_560),
.A2(n_561),
.B1(n_567),
.B2(n_571),
.Y(n_586)
);

AOI22xp5_ASAP7_75t_L g561 ( 
.A1(n_530),
.A2(n_496),
.B1(n_479),
.B2(n_507),
.Y(n_561)
);

AOI22xp5_ASAP7_75t_SL g597 ( 
.A1(n_563),
.A2(n_540),
.B1(n_524),
.B2(n_542),
.Y(n_597)
);

AOI21xp5_ASAP7_75t_L g595 ( 
.A1(n_564),
.A2(n_575),
.B(n_552),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_517),
.B(n_497),
.Y(n_566)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_566),
.Y(n_609)
);

AOI22xp5_ASAP7_75t_L g567 ( 
.A1(n_522),
.A2(n_496),
.B1(n_507),
.B2(n_504),
.Y(n_567)
);

MAJIxp5_ASAP7_75t_L g570 ( 
.A(n_544),
.B(n_488),
.C(n_512),
.Y(n_570)
);

MAJIxp5_ASAP7_75t_L g589 ( 
.A(n_570),
.B(n_573),
.C(n_584),
.Y(n_589)
);

AOI22xp5_ASAP7_75t_L g571 ( 
.A1(n_525),
.A2(n_481),
.B1(n_491),
.B2(n_476),
.Y(n_571)
);

AOI22xp5_ASAP7_75t_L g572 ( 
.A1(n_529),
.A2(n_536),
.B1(n_532),
.B2(n_542),
.Y(n_572)
);

OAI22xp5_ASAP7_75t_SL g610 ( 
.A1(n_572),
.A2(n_579),
.B1(n_560),
.B2(n_557),
.Y(n_610)
);

MAJIxp5_ASAP7_75t_L g573 ( 
.A(n_521),
.B(n_499),
.C(n_505),
.Y(n_573)
);

OAI21xp5_ASAP7_75t_L g575 ( 
.A1(n_529),
.A2(n_500),
.B(n_493),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_520),
.Y(n_576)
);

HB1xp67_ASAP7_75t_L g591 ( 
.A(n_576),
.Y(n_591)
);

XNOR2xp5_ASAP7_75t_L g577 ( 
.A(n_543),
.B(n_502),
.Y(n_577)
);

XNOR2xp5_ASAP7_75t_L g602 ( 
.A(n_577),
.B(n_550),
.Y(n_602)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_533),
.Y(n_578)
);

HB1xp67_ASAP7_75t_L g603 ( 
.A(n_578),
.Y(n_603)
);

AOI22xp5_ASAP7_75t_L g579 ( 
.A1(n_536),
.A2(n_506),
.B1(n_480),
.B2(n_388),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_527),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_SL g606 ( 
.A(n_580),
.B(n_583),
.Y(n_606)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_534),
.Y(n_581)
);

INVx4_ASAP7_75t_L g590 ( 
.A(n_581),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_SL g582 ( 
.A(n_523),
.B(n_442),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_SL g594 ( 
.A(n_582),
.B(n_571),
.Y(n_594)
);

CKINVDCx16_ASAP7_75t_R g583 ( 
.A(n_547),
.Y(n_583)
);

MAJIxp5_ASAP7_75t_L g584 ( 
.A(n_521),
.B(n_526),
.C(n_546),
.Y(n_584)
);

XOR2xp5_ASAP7_75t_L g585 ( 
.A(n_539),
.B(n_473),
.Y(n_585)
);

XOR2xp5_ASAP7_75t_L g598 ( 
.A(n_585),
.B(n_516),
.Y(n_598)
);

CKINVDCx20_ASAP7_75t_R g587 ( 
.A(n_575),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_587),
.B(n_592),
.Y(n_617)
);

MAJIxp5_ASAP7_75t_L g592 ( 
.A(n_573),
.B(n_531),
.C(n_545),
.Y(n_592)
);

XNOR2xp5_ASAP7_75t_SL g593 ( 
.A(n_568),
.B(n_541),
.Y(n_593)
);

XOR2xp5_ASAP7_75t_L g616 ( 
.A(n_593),
.B(n_596),
.Y(n_616)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_594),
.Y(n_632)
);

AOI21xp5_ASAP7_75t_L g626 ( 
.A1(n_595),
.A2(n_579),
.B(n_367),
.Y(n_626)
);

XNOR2x1_ASAP7_75t_L g596 ( 
.A(n_585),
.B(n_535),
.Y(n_596)
);

OAI22xp5_ASAP7_75t_L g629 ( 
.A1(n_597),
.A2(n_365),
.B1(n_379),
.B2(n_333),
.Y(n_629)
);

XOR2xp5_ASAP7_75t_L g627 ( 
.A(n_598),
.B(n_611),
.Y(n_627)
);

A2O1A1Ixp33_ASAP7_75t_L g599 ( 
.A1(n_564),
.A2(n_538),
.B(n_549),
.C(n_548),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_599),
.B(n_572),
.Y(n_612)
);

MAJIxp5_ASAP7_75t_L g600 ( 
.A(n_584),
.B(n_518),
.C(n_549),
.Y(n_600)
);

MAJIxp5_ASAP7_75t_L g613 ( 
.A(n_600),
.B(n_565),
.C(n_569),
.Y(n_613)
);

XNOR2xp5_ASAP7_75t_L g615 ( 
.A(n_602),
.B(n_604),
.Y(n_615)
);

XNOR2xp5_ASAP7_75t_L g604 ( 
.A(n_555),
.B(n_538),
.Y(n_604)
);

XNOR2xp5_ASAP7_75t_L g607 ( 
.A(n_565),
.B(n_527),
.Y(n_607)
);

XNOR2xp5_ASAP7_75t_L g619 ( 
.A(n_607),
.B(n_574),
.Y(n_619)
);

AOI22xp33_ASAP7_75t_SL g622 ( 
.A1(n_610),
.A2(n_554),
.B1(n_567),
.B2(n_581),
.Y(n_622)
);

XOR2xp5_ASAP7_75t_L g611 ( 
.A(n_570),
.B(n_534),
.Y(n_611)
);

AOI21xp5_ASAP7_75t_L g636 ( 
.A1(n_612),
.A2(n_626),
.B(n_608),
.Y(n_636)
);

XNOR2xp5_ASAP7_75t_L g639 ( 
.A(n_613),
.B(n_619),
.Y(n_639)
);

MAJIxp5_ASAP7_75t_L g614 ( 
.A(n_588),
.B(n_577),
.C(n_559),
.Y(n_614)
);

MAJIxp5_ASAP7_75t_L g642 ( 
.A(n_614),
.B(n_620),
.C(n_621),
.Y(n_642)
);

BUFx24_ASAP7_75t_SL g618 ( 
.A(n_601),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_L g640 ( 
.A(n_618),
.B(n_631),
.Y(n_640)
);

MAJIxp5_ASAP7_75t_L g620 ( 
.A(n_588),
.B(n_574),
.C(n_568),
.Y(n_620)
);

MAJIxp5_ASAP7_75t_L g621 ( 
.A(n_589),
.B(n_562),
.C(n_558),
.Y(n_621)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_622),
.Y(n_637)
);

MAJIxp5_ASAP7_75t_L g623 ( 
.A(n_589),
.B(n_562),
.C(n_561),
.Y(n_623)
);

MAJIxp5_ASAP7_75t_L g643 ( 
.A(n_623),
.B(n_611),
.C(n_592),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_L g624 ( 
.A(n_607),
.B(n_442),
.Y(n_624)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_624),
.Y(n_641)
);

CKINVDCx20_ASAP7_75t_R g625 ( 
.A(n_591),
.Y(n_625)
);

AOI22xp33_ASAP7_75t_SL g638 ( 
.A1(n_625),
.A2(n_603),
.B1(n_605),
.B2(n_590),
.Y(n_638)
);

NOR2xp33_ASAP7_75t_L g628 ( 
.A(n_609),
.B(n_340),
.Y(n_628)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_628),
.Y(n_644)
);

AOI22xp5_ASAP7_75t_L g647 ( 
.A1(n_629),
.A2(n_630),
.B1(n_633),
.B2(n_590),
.Y(n_647)
);

AOI22xp5_ASAP7_75t_L g630 ( 
.A1(n_586),
.A2(n_365),
.B1(n_322),
.B2(n_333),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_SL g631 ( 
.A(n_606),
.B(n_355),
.Y(n_631)
);

AOI22xp5_ASAP7_75t_L g633 ( 
.A1(n_586),
.A2(n_321),
.B1(n_322),
.B2(n_610),
.Y(n_633)
);

XOR2xp5_ASAP7_75t_L g634 ( 
.A(n_619),
.B(n_596),
.Y(n_634)
);

AND2x2_ASAP7_75t_L g661 ( 
.A(n_634),
.B(n_635),
.Y(n_661)
);

XOR2xp5_ASAP7_75t_L g635 ( 
.A(n_615),
.B(n_604),
.Y(n_635)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_636),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_638),
.B(n_643),
.Y(n_653)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_612),
.Y(n_645)
);

NOR2xp33_ASAP7_75t_L g652 ( 
.A(n_645),
.B(n_646),
.Y(n_652)
);

NOR2xp33_ASAP7_75t_L g646 ( 
.A(n_617),
.B(n_600),
.Y(n_646)
);

XNOR2xp5_ASAP7_75t_L g658 ( 
.A(n_647),
.B(n_648),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_632),
.B(n_602),
.Y(n_648)
);

MAJIxp5_ASAP7_75t_L g649 ( 
.A(n_613),
.B(n_614),
.C(n_621),
.Y(n_649)
);

MAJIxp5_ASAP7_75t_L g655 ( 
.A(n_649),
.B(n_651),
.C(n_627),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_615),
.B(n_599),
.Y(n_650)
);

XNOR2xp5_ASAP7_75t_L g660 ( 
.A(n_650),
.B(n_616),
.Y(n_660)
);

MAJIxp5_ASAP7_75t_L g651 ( 
.A(n_623),
.B(n_598),
.C(n_597),
.Y(n_651)
);

OAI21xp5_ASAP7_75t_SL g654 ( 
.A1(n_650),
.A2(n_626),
.B(n_633),
.Y(n_654)
);

AOI21xp5_ASAP7_75t_L g668 ( 
.A1(n_654),
.A2(n_662),
.B(n_664),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_655),
.B(n_656),
.Y(n_673)
);

MAJIxp5_ASAP7_75t_L g656 ( 
.A(n_639),
.B(n_627),
.C(n_620),
.Y(n_656)
);

NOR2xp33_ASAP7_75t_L g657 ( 
.A(n_644),
.B(n_630),
.Y(n_657)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_657),
.Y(n_667)
);

MAJIxp5_ASAP7_75t_L g659 ( 
.A(n_639),
.B(n_616),
.C(n_593),
.Y(n_659)
);

MAJIxp5_ASAP7_75t_L g666 ( 
.A(n_659),
.B(n_665),
.C(n_642),
.Y(n_666)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_660),
.Y(n_675)
);

OAI21xp5_ASAP7_75t_SL g662 ( 
.A1(n_636),
.A2(n_321),
.B(n_637),
.Y(n_662)
);

NOR2xp33_ASAP7_75t_L g664 ( 
.A(n_649),
.B(n_640),
.Y(n_664)
);

MAJIxp5_ASAP7_75t_L g665 ( 
.A(n_643),
.B(n_642),
.C(n_635),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_SL g680 ( 
.A(n_666),
.B(n_672),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_L g669 ( 
.A(n_665),
.B(n_648),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_669),
.B(n_670),
.Y(n_681)
);

NOR2xp33_ASAP7_75t_L g670 ( 
.A(n_663),
.B(n_641),
.Y(n_670)
);

INVxp67_ASAP7_75t_L g671 ( 
.A(n_653),
.Y(n_671)
);

NOR2xp33_ASAP7_75t_L g677 ( 
.A(n_671),
.B(n_655),
.Y(n_677)
);

NOR2xp33_ASAP7_75t_L g672 ( 
.A(n_658),
.B(n_651),
.Y(n_672)
);

OAI21xp5_ASAP7_75t_L g674 ( 
.A1(n_658),
.A2(n_647),
.B(n_634),
.Y(n_674)
);

AOI21xp5_ASAP7_75t_L g676 ( 
.A1(n_674),
.A2(n_652),
.B(n_660),
.Y(n_676)
);

AOI22xp5_ASAP7_75t_L g682 ( 
.A1(n_676),
.A2(n_677),
.B1(n_679),
.B2(n_667),
.Y(n_682)
);

AND2x2_ASAP7_75t_L g678 ( 
.A(n_673),
.B(n_656),
.Y(n_678)
);

CKINVDCx20_ASAP7_75t_R g684 ( 
.A(n_678),
.Y(n_684)
);

AOI21xp5_ASAP7_75t_L g679 ( 
.A1(n_666),
.A2(n_661),
.B(n_659),
.Y(n_679)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_682),
.Y(n_685)
);

NOR2xp33_ASAP7_75t_SL g683 ( 
.A(n_681),
.B(n_675),
.Y(n_683)
);

MAJx2_ASAP7_75t_L g686 ( 
.A(n_683),
.B(n_680),
.C(n_668),
.Y(n_686)
);

MAJIxp5_ASAP7_75t_L g687 ( 
.A(n_686),
.B(n_684),
.C(n_671),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_687),
.B(n_685),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_SL g689 ( 
.A(n_688),
.B(n_674),
.Y(n_689)
);

XNOR2xp5_ASAP7_75t_L g690 ( 
.A(n_689),
.B(n_661),
.Y(n_690)
);


endmodule