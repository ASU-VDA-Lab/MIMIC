module fake_jpeg_16507_n_55 (n_13, n_21, n_1, n_10, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_55);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_55;

wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_27;
wire n_47;
wire n_51;
wire n_40;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_31;
wire n_25;
wire n_29;
wire n_43;
wire n_37;
wire n_50;
wire n_32;

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_22),
.B(n_14),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

AOI21xp33_ASAP7_75t_L g28 ( 
.A1(n_10),
.A2(n_2),
.B(n_18),
.Y(n_28)
);

OR2x2_ASAP7_75t_L g29 ( 
.A(n_3),
.B(n_13),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

AOI21xp5_ASAP7_75t_L g31 ( 
.A1(n_28),
.A2(n_20),
.B(n_9),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_31),
.A2(n_23),
.B1(n_8),
.B2(n_15),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_29),
.B(n_26),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_32),
.B(n_35),
.Y(n_37)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_25),
.Y(n_33)
);

OR2x2_ASAP7_75t_L g41 ( 
.A(n_33),
.B(n_36),
.Y(n_41)
);

CKINVDCx12_ASAP7_75t_R g34 ( 
.A(n_24),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g35 ( 
.A(n_29),
.B(n_0),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

OAI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_33),
.A2(n_11),
.B1(n_19),
.B2(n_16),
.Y(n_38)
);

NOR3xp33_ASAP7_75t_L g45 ( 
.A(n_38),
.B(n_39),
.C(n_5),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_35),
.B(n_30),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_42),
.B(n_43),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_35),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_43)
);

INVx5_ASAP7_75t_SL g44 ( 
.A(n_40),
.Y(n_44)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_45),
.Y(n_48)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

AOI221xp5_ASAP7_75t_L g50 ( 
.A1(n_48),
.A2(n_46),
.B1(n_47),
.B2(n_45),
.C(n_37),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_50),
.A2(n_41),
.B1(n_49),
.B2(n_27),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_51),
.B(n_41),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_52),
.Y(n_53)
);

AO21x1_ASAP7_75t_L g54 ( 
.A1(n_53),
.A2(n_6),
.B(n_7),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_54),
.Y(n_55)
);


endmodule