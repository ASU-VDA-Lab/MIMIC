module fake_ariane_3007_n_2168 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_195, n_38, n_213, n_47, n_110, n_153, n_18, n_197, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_203, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_205, n_71, n_24, n_7, n_109, n_208, n_96, n_156, n_209, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_210, n_147, n_204, n_200, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_199, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_201, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_212, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_198, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_206, n_13, n_27, n_207, n_29, n_41, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_211, n_194, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_202, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_2168);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_195;
input n_38;
input n_213;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_203;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_205;
input n_71;
input n_24;
input n_7;
input n_109;
input n_208;
input n_96;
input n_156;
input n_209;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_210;
input n_147;
input n_204;
input n_200;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_199;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_201;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_198;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_206;
input n_13;
input n_27;
input n_207;
input n_29;
input n_41;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_211;
input n_194;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_202;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_2168;

wire n_913;
wire n_1681;
wire n_2163;
wire n_1486;
wire n_1507;
wire n_1938;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_2131;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_2135;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_2002;
wire n_1463;
wire n_1238;
wire n_2011;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_2013;
wire n_1566;
wire n_717;
wire n_2006;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_214;
wire n_2042;
wire n_2123;
wire n_1853;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_2084;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_1985;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1909;
wire n_2156;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1979;
wire n_1277;
wire n_2107;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_2109;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_1944;
wire n_331;
wire n_559;
wire n_495;
wire n_267;
wire n_1988;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_2149;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_2078;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_2162;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_1977;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_2060;
wire n_1850;
wire n_238;
wire n_365;
wire n_2004;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_661;
wire n_2098;
wire n_1751;
wire n_300;
wire n_533;
wire n_1917;
wire n_1924;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_2045;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_2061;
wire n_2094;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_2043;
wire n_780;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_2077;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_225;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_2038;
wire n_2116;
wire n_2145;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_2134;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_2166;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_2015;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_2072;
wire n_306;
wire n_436;
wire n_324;
wire n_2087;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_2161;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_2155;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_1880;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_2100;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_2147;
wire n_1226;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1970;
wire n_1920;
wire n_2083;
wire n_815;
wire n_542;
wire n_2167;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1911;
wire n_1908;
wire n_1825;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_2066;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_1914;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_2019;
wire n_698;
wire n_2130;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_2160;
wire n_1992;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_2142;
wire n_1633;
wire n_404;
wire n_1913;
wire n_2069;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_2144;
wire n_564;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_2120;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_2041;
wire n_2113;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_552;
wire n_348;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1951;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_2132;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_720;
wire n_926;
wire n_1943;
wire n_1802;
wire n_2112;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_2146;
wire n_1868;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_2099;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_1413;
wire n_2129;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_2059;
wire n_1439;
wire n_814;
wire n_578;
wire n_2074;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_2122;
wire n_320;
wire n_1414;
wire n_1134;
wire n_2067;
wire n_1484;
wire n_1901;
wire n_647;
wire n_2055;
wire n_2027;
wire n_1423;
wire n_2117;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_1939;
wire n_1906;
wire n_529;
wire n_1899;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1828;
wire n_2159;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_2102;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_2023;
wire n_1278;
wire n_707;
wire n_983;
wire n_699;
wire n_590;
wire n_727;
wire n_301;
wire n_1726;
wire n_2075;
wire n_1945;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_2031;
wire n_2118;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_1963;
wire n_729;
wire n_887;
wire n_2057;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_2125;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_2033;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_1883;
wire n_1969;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1927;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_1957;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_534;
wire n_1791;
wire n_2124;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_2119;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_2008;
wire n_454;
wire n_298;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_2127;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_2071;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_2082;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_2140;
wire n_873;
wire n_1301;
wire n_1748;
wire n_2157;
wire n_1966;
wire n_1243;
wire n_1400;
wire n_342;
wire n_2035;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_2128;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1993;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1897;
wire n_2137;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_2026;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_642;
wire n_1804;
wire n_2106;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_2091;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_1929;
wire n_1950;
wire n_805;
wire n_2032;
wire n_2090;
wire n_295;
wire n_1658;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1997;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_463;
wire n_1524;
wire n_1476;
wire n_1733;
wire n_1856;
wire n_2016;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_1971;
wire n_586;
wire n_1429;
wire n_1324;
wire n_2064;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_2022;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_2143;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_2076;
wire n_2133;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_2001;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_2158;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_2070;
wire n_2136;
wire n_426;
wire n_433;
wire n_398;
wire n_1090;
wire n_1367;
wire n_2044;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_2020;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_1881;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_1958;
wire n_467;
wire n_1511;
wire n_1422;
wire n_1965;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_2036;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_2003;
wire n_1307;
wire n_1128;
wire n_2053;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1955;
wire n_2110;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_2121;
wire n_601;
wire n_683;
wire n_236;
wire n_565;
wire n_628;
wire n_1300;
wire n_1960;
wire n_2068;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_1978;
wire n_571;
wire n_414;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_526;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_2154;
wire n_1789;
wire n_763;
wire n_1986;
wire n_540;
wire n_216;
wire n_692;
wire n_2054;
wire n_1857;
wire n_984;
wire n_1687;
wire n_2073;
wire n_223;
wire n_2150;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_2046;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_2093;
wire n_2018;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_493;
wire n_1311;
wire n_1956;
wire n_1589;
wire n_2151;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_2114;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_2014;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_2141;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_508;
wire n_1679;
wire n_2126;
wire n_1952;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_1834;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_2050;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_1980;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_1998;
wire n_2165;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_2028;
wire n_919;
wire n_1663;
wire n_2092;
wire n_1625;
wire n_2086;
wire n_1926;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_2138;
wire n_2065;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1904;
wire n_2000;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_2096;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1937;
wire n_2012;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_2111;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_2103;
wire n_1710;
wire n_1865;
wire n_309;
wire n_1344;
wire n_1390;
wire n_485;
wire n_401;
wire n_1792;
wire n_504;
wire n_2062;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_2153;
wire n_1510;
wire n_2139;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1727;
wire n_1991;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_2034;
wire n_1845;
wire n_2101;
wire n_1934;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_2104;
wire n_1265;
wire n_1576;
wire n_2105;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_2088;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_2005;
wire n_2048;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_2108;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_1866;
wire n_2056;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_838;
wire n_383;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_2085;
wire n_1686;
wire n_1964;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_1982;
wire n_2097;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_2115;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_2148;
wire n_1946;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_2051;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_2164;
wire n_1732;
wire n_415;
wire n_1967;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_2052;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_2080;
wire n_2058;
wire n_1126;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_2047;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_2081;
wire n_265;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_925;
wire n_246;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1905;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_2063;
wire n_1925;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_2079;
wire n_1228;
wire n_2152;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_484;
wire n_411;
wire n_849;
wire n_2095;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_1989;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2037;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_2089;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_53),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_34),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_147),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_81),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_23),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_11),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_2),
.Y(n_220)
);

INVx1_ASAP7_75t_SL g221 ( 
.A(n_44),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_117),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_104),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_76),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_94),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_185),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_9),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_5),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_65),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_102),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_99),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_34),
.Y(n_232)
);

BUFx3_ASAP7_75t_L g233 ( 
.A(n_26),
.Y(n_233)
);

INVx2_ASAP7_75t_SL g234 ( 
.A(n_49),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_53),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_90),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_56),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_161),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_183),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_154),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_52),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_23),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_148),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_64),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_51),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_212),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_58),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_136),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_129),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_1),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_137),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_78),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_46),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_143),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_206),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_72),
.Y(n_256)
);

CKINVDCx16_ASAP7_75t_R g257 ( 
.A(n_68),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_41),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_157),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_74),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_85),
.Y(n_261)
);

BUFx2_ASAP7_75t_L g262 ( 
.A(n_114),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_1),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_25),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_79),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_139),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_142),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_155),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_165),
.Y(n_269)
);

HB1xp67_ASAP7_75t_L g270 ( 
.A(n_188),
.Y(n_270)
);

BUFx10_ASAP7_75t_L g271 ( 
.A(n_130),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_182),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_13),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_207),
.Y(n_274)
);

BUFx3_ASAP7_75t_L g275 ( 
.A(n_51),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_59),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_44),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_208),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_45),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_83),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_171),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_169),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_79),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_69),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_87),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_209),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_10),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_164),
.Y(n_288)
);

BUFx8_ASAP7_75t_SL g289 ( 
.A(n_69),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_178),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_55),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_5),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_187),
.Y(n_293)
);

INVx2_ASAP7_75t_SL g294 ( 
.A(n_176),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_158),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_111),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_50),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_36),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_201),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_122),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_106),
.Y(n_301)
);

BUFx2_ASAP7_75t_L g302 ( 
.A(n_61),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_193),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_105),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_199),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_177),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_135),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_167),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_174),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_73),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_77),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_31),
.Y(n_312)
);

BUFx6f_ASAP7_75t_L g313 ( 
.A(n_190),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_192),
.Y(n_314)
);

CKINVDCx14_ASAP7_75t_R g315 ( 
.A(n_82),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_92),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_49),
.Y(n_317)
);

BUFx2_ASAP7_75t_L g318 ( 
.A(n_153),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_113),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_71),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_112),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_3),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_156),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_30),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_39),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_57),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_180),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_110),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_11),
.Y(n_329)
);

INVxp67_ASAP7_75t_L g330 ( 
.A(n_131),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_9),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_78),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_172),
.Y(n_333)
);

INVx1_ASAP7_75t_SL g334 ( 
.A(n_36),
.Y(n_334)
);

INVx1_ASAP7_75t_SL g335 ( 
.A(n_162),
.Y(n_335)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_71),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_66),
.Y(n_337)
);

INVx1_ASAP7_75t_SL g338 ( 
.A(n_186),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_144),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_195),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_21),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_55),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_73),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_57),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_152),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_47),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_108),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_159),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_63),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_109),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_91),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_80),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_202),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_37),
.Y(n_354)
);

BUFx6f_ASAP7_75t_L g355 ( 
.A(n_7),
.Y(n_355)
);

BUFx2_ASAP7_75t_L g356 ( 
.A(n_7),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_37),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_120),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_133),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_25),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_118),
.Y(n_361)
);

BUFx3_ASAP7_75t_L g362 ( 
.A(n_198),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_181),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_18),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_68),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_138),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_46),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_67),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_2),
.Y(n_369)
);

INVx1_ASAP7_75t_SL g370 ( 
.A(n_116),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_141),
.Y(n_371)
);

BUFx10_ASAP7_75t_L g372 ( 
.A(n_134),
.Y(n_372)
);

HB1xp67_ASAP7_75t_L g373 ( 
.A(n_197),
.Y(n_373)
);

BUFx2_ASAP7_75t_L g374 ( 
.A(n_163),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_74),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_128),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_62),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_29),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_30),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_59),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_124),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_150),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_205),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_196),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_89),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_15),
.Y(n_386)
);

BUFx10_ASAP7_75t_L g387 ( 
.A(n_56),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_35),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_121),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_66),
.Y(n_390)
);

INVx1_ASAP7_75t_SL g391 ( 
.A(n_38),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_43),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_6),
.Y(n_393)
);

INVx2_ASAP7_75t_SL g394 ( 
.A(n_119),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_184),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_61),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_168),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_132),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_19),
.Y(n_399)
);

BUFx6f_ASAP7_75t_L g400 ( 
.A(n_8),
.Y(n_400)
);

INVx1_ASAP7_75t_SL g401 ( 
.A(n_145),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_127),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_45),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_33),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_13),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_203),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_191),
.Y(n_407)
);

BUFx6f_ASAP7_75t_L g408 ( 
.A(n_67),
.Y(n_408)
);

INVx1_ASAP7_75t_SL g409 ( 
.A(n_126),
.Y(n_409)
);

INVx1_ASAP7_75t_SL g410 ( 
.A(n_194),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_95),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_21),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_60),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_52),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_170),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_97),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_70),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_64),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_75),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_81),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_189),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_166),
.Y(n_422)
);

INVxp67_ASAP7_75t_SL g423 ( 
.A(n_233),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_289),
.Y(n_424)
);

INVxp67_ASAP7_75t_L g425 ( 
.A(n_302),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_257),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_216),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_355),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_222),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_299),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_363),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_222),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_223),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_395),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_223),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_220),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_226),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_226),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_228),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_235),
.Y(n_440)
);

INVxp67_ASAP7_75t_SL g441 ( 
.A(n_233),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_238),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_214),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_R g444 ( 
.A(n_315),
.B(n_84),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_215),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_283),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_218),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_238),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_239),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_219),
.Y(n_450)
);

HB1xp67_ASAP7_75t_L g451 ( 
.A(n_302),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_224),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_291),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_227),
.Y(n_454)
);

AND2x2_ASAP7_75t_L g455 ( 
.A(n_356),
.B(n_0),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_325),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_239),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_332),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_262),
.B(n_0),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_229),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_232),
.Y(n_461)
);

HB1xp67_ASAP7_75t_L g462 ( 
.A(n_356),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_262),
.B(n_318),
.Y(n_463)
);

BUFx2_ASAP7_75t_L g464 ( 
.A(n_275),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_318),
.B(n_3),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_241),
.Y(n_466)
);

AND2x2_ASAP7_75t_L g467 ( 
.A(n_374),
.B(n_387),
.Y(n_467)
);

NOR2xp67_ASAP7_75t_L g468 ( 
.A(n_234),
.B(n_4),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_240),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_244),
.Y(n_470)
);

INVxp33_ASAP7_75t_SL g471 ( 
.A(n_245),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_240),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g473 ( 
.A(n_337),
.Y(n_473)
);

INVxp67_ASAP7_75t_SL g474 ( 
.A(n_275),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_247),
.Y(n_475)
);

CKINVDCx20_ASAP7_75t_R g476 ( 
.A(n_368),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_252),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_243),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_243),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_403),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_254),
.Y(n_481)
);

NOR2xp67_ASAP7_75t_L g482 ( 
.A(n_234),
.B(n_4),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_355),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_253),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_254),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_355),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_256),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_255),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_255),
.Y(n_489)
);

CKINVDCx20_ASAP7_75t_R g490 ( 
.A(n_404),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_258),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_259),
.Y(n_492)
);

INVxp67_ASAP7_75t_L g493 ( 
.A(n_217),
.Y(n_493)
);

CKINVDCx20_ASAP7_75t_R g494 ( 
.A(n_412),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_259),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_261),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_260),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_261),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_263),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_264),
.Y(n_500)
);

CKINVDCx20_ASAP7_75t_R g501 ( 
.A(n_418),
.Y(n_501)
);

NOR2xp67_ASAP7_75t_L g502 ( 
.A(n_336),
.B(n_6),
.Y(n_502)
);

BUFx10_ASAP7_75t_L g503 ( 
.A(n_294),
.Y(n_503)
);

HB1xp67_ASAP7_75t_L g504 ( 
.A(n_273),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_374),
.B(n_8),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_272),
.Y(n_506)
);

INVxp67_ASAP7_75t_SL g507 ( 
.A(n_355),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_272),
.Y(n_508)
);

INVx3_ASAP7_75t_L g509 ( 
.A(n_355),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_274),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_279),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_274),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_285),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_285),
.Y(n_514)
);

INVxp67_ASAP7_75t_L g515 ( 
.A(n_217),
.Y(n_515)
);

INVxp67_ASAP7_75t_L g516 ( 
.A(n_237),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_293),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_284),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_292),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_293),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_301),
.Y(n_521)
);

INVxp33_ASAP7_75t_L g522 ( 
.A(n_237),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_301),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_297),
.Y(n_524)
);

CKINVDCx20_ASAP7_75t_R g525 ( 
.A(n_271),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_329),
.Y(n_526)
);

CKINVDCx20_ASAP7_75t_R g527 ( 
.A(n_271),
.Y(n_527)
);

BUFx3_ASAP7_75t_L g528 ( 
.A(n_362),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_331),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_307),
.Y(n_530)
);

CKINVDCx20_ASAP7_75t_R g531 ( 
.A(n_271),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_509),
.Y(n_532)
);

AND2x2_ASAP7_75t_L g533 ( 
.A(n_467),
.B(n_429),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_463),
.B(n_270),
.Y(n_534)
);

AND2x2_ASAP7_75t_L g535 ( 
.A(n_467),
.B(n_360),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_509),
.Y(n_536)
);

BUFx6f_ASAP7_75t_L g537 ( 
.A(n_509),
.Y(n_537)
);

BUFx6f_ASAP7_75t_L g538 ( 
.A(n_509),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_428),
.Y(n_539)
);

XNOR2x2_ASAP7_75t_R g540 ( 
.A(n_424),
.B(n_387),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_428),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_483),
.Y(n_542)
);

BUFx2_ASAP7_75t_L g543 ( 
.A(n_426),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_483),
.Y(n_544)
);

BUFx6f_ASAP7_75t_L g545 ( 
.A(n_486),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_507),
.Y(n_546)
);

AND2x4_ASAP7_75t_L g547 ( 
.A(n_429),
.B(n_400),
.Y(n_547)
);

HB1xp67_ASAP7_75t_L g548 ( 
.A(n_451),
.Y(n_548)
);

BUFx6f_ASAP7_75t_L g549 ( 
.A(n_486),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_432),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_432),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_433),
.B(n_373),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_433),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_435),
.Y(n_554)
);

INVx3_ASAP7_75t_L g555 ( 
.A(n_435),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_437),
.B(n_438),
.Y(n_556)
);

AND2x2_ASAP7_75t_L g557 ( 
.A(n_437),
.B(n_360),
.Y(n_557)
);

BUFx2_ASAP7_75t_L g558 ( 
.A(n_443),
.Y(n_558)
);

NAND2xp33_ASAP7_75t_L g559 ( 
.A(n_455),
.B(n_400),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_438),
.Y(n_560)
);

BUFx6f_ASAP7_75t_L g561 ( 
.A(n_442),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_442),
.Y(n_562)
);

INVx3_ASAP7_75t_L g563 ( 
.A(n_448),
.Y(n_563)
);

BUFx6f_ASAP7_75t_L g564 ( 
.A(n_448),
.Y(n_564)
);

BUFx6f_ASAP7_75t_L g565 ( 
.A(n_449),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_449),
.B(n_457),
.Y(n_566)
);

NAND2xp33_ASAP7_75t_L g567 ( 
.A(n_455),
.B(n_400),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_457),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_469),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_469),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_472),
.Y(n_571)
);

AND2x6_ASAP7_75t_L g572 ( 
.A(n_472),
.B(n_313),
.Y(n_572)
);

CKINVDCx6p67_ASAP7_75t_R g573 ( 
.A(n_525),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_478),
.Y(n_574)
);

AND2x2_ASAP7_75t_L g575 ( 
.A(n_478),
.B(n_271),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_479),
.Y(n_576)
);

BUFx6f_ASAP7_75t_L g577 ( 
.A(n_479),
.Y(n_577)
);

AND2x6_ASAP7_75t_L g578 ( 
.A(n_481),
.B(n_313),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_481),
.Y(n_579)
);

AND2x2_ASAP7_75t_L g580 ( 
.A(n_485),
.B(n_372),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_485),
.Y(n_581)
);

BUFx6f_ASAP7_75t_L g582 ( 
.A(n_488),
.Y(n_582)
);

AOI22xp5_ASAP7_75t_L g583 ( 
.A1(n_425),
.A2(n_334),
.B1(n_391),
.B2(n_221),
.Y(n_583)
);

HB1xp67_ASAP7_75t_L g584 ( 
.A(n_462),
.Y(n_584)
);

AND2x2_ASAP7_75t_L g585 ( 
.A(n_488),
.B(n_372),
.Y(n_585)
);

BUFx6f_ASAP7_75t_L g586 ( 
.A(n_489),
.Y(n_586)
);

BUFx6f_ASAP7_75t_L g587 ( 
.A(n_489),
.Y(n_587)
);

AND2x2_ASAP7_75t_L g588 ( 
.A(n_492),
.B(n_372),
.Y(n_588)
);

INVx3_ASAP7_75t_L g589 ( 
.A(n_492),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_495),
.Y(n_590)
);

BUFx6f_ASAP7_75t_L g591 ( 
.A(n_495),
.Y(n_591)
);

INVx6_ASAP7_75t_L g592 ( 
.A(n_503),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_496),
.Y(n_593)
);

INVx3_ASAP7_75t_L g594 ( 
.A(n_496),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_498),
.Y(n_595)
);

INVx4_ASAP7_75t_L g596 ( 
.A(n_503),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_498),
.Y(n_597)
);

BUFx2_ASAP7_75t_L g598 ( 
.A(n_445),
.Y(n_598)
);

BUFx6f_ASAP7_75t_L g599 ( 
.A(n_506),
.Y(n_599)
);

BUFx6f_ASAP7_75t_L g600 ( 
.A(n_506),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_508),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_508),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_510),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_510),
.Y(n_604)
);

INVx3_ASAP7_75t_L g605 ( 
.A(n_512),
.Y(n_605)
);

OA21x2_ASAP7_75t_L g606 ( 
.A1(n_512),
.A2(n_514),
.B(n_513),
.Y(n_606)
);

AND2x4_ASAP7_75t_L g607 ( 
.A(n_513),
.B(n_400),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_514),
.Y(n_608)
);

AND2x2_ASAP7_75t_L g609 ( 
.A(n_517),
.B(n_372),
.Y(n_609)
);

OAI22xp5_ASAP7_75t_SL g610 ( 
.A1(n_436),
.A2(n_250),
.B1(n_265),
.B2(n_242),
.Y(n_610)
);

BUFx2_ASAP7_75t_L g611 ( 
.A(n_447),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_517),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_SL g613 ( 
.A(n_459),
.B(n_400),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_520),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_520),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_521),
.B(n_307),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_521),
.Y(n_617)
);

AND2x4_ASAP7_75t_L g618 ( 
.A(n_523),
.B(n_408),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_532),
.Y(n_619)
);

CKINVDCx20_ASAP7_75t_R g620 ( 
.A(n_558),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_561),
.Y(n_621)
);

BUFx3_ASAP7_75t_L g622 ( 
.A(n_546),
.Y(n_622)
);

OAI22xp5_ASAP7_75t_L g623 ( 
.A1(n_534),
.A2(n_505),
.B1(n_465),
.B2(n_471),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_L g624 ( 
.A(n_534),
.B(n_450),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_SL g625 ( 
.A(n_558),
.B(n_452),
.Y(n_625)
);

AOI22xp33_ASAP7_75t_L g626 ( 
.A1(n_575),
.A2(n_468),
.B1(n_482),
.B2(n_522),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_561),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_561),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_561),
.Y(n_629)
);

BUFx6f_ASAP7_75t_L g630 ( 
.A(n_561),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_561),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_532),
.Y(n_632)
);

NOR2xp33_ASAP7_75t_L g633 ( 
.A(n_546),
.B(n_454),
.Y(n_633)
);

INVx5_ASAP7_75t_L g634 ( 
.A(n_572),
.Y(n_634)
);

INVx1_ASAP7_75t_SL g635 ( 
.A(n_543),
.Y(n_635)
);

INVx3_ASAP7_75t_L g636 ( 
.A(n_606),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_575),
.B(n_503),
.Y(n_637)
);

NOR2xp33_ASAP7_75t_L g638 ( 
.A(n_596),
.B(n_460),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_532),
.Y(n_639)
);

AND2x2_ASAP7_75t_L g640 ( 
.A(n_533),
.B(n_423),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_532),
.Y(n_641)
);

AND3x1_ASAP7_75t_L g642 ( 
.A(n_583),
.B(n_250),
.C(n_242),
.Y(n_642)
);

CKINVDCx20_ASAP7_75t_R g643 ( 
.A(n_558),
.Y(n_643)
);

AOI22xp33_ASAP7_75t_L g644 ( 
.A1(n_575),
.A2(n_468),
.B1(n_482),
.B2(n_444),
.Y(n_644)
);

NAND3xp33_ASAP7_75t_L g645 ( 
.A(n_533),
.B(n_466),
.C(n_461),
.Y(n_645)
);

INVx1_ASAP7_75t_SL g646 ( 
.A(n_543),
.Y(n_646)
);

OAI22xp33_ASAP7_75t_L g647 ( 
.A1(n_583),
.A2(n_502),
.B1(n_475),
.B2(n_477),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_580),
.B(n_503),
.Y(n_648)
);

BUFx6f_ASAP7_75t_L g649 ( 
.A(n_561),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_561),
.Y(n_650)
);

INVxp67_ASAP7_75t_SL g651 ( 
.A(n_556),
.Y(n_651)
);

INVx2_ASAP7_75t_SL g652 ( 
.A(n_580),
.Y(n_652)
);

OAI21xp33_ASAP7_75t_SL g653 ( 
.A1(n_533),
.A2(n_585),
.B(n_580),
.Y(n_653)
);

NOR2xp33_ASAP7_75t_L g654 ( 
.A(n_596),
.B(n_470),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_564),
.Y(n_655)
);

BUFx8_ASAP7_75t_SL g656 ( 
.A(n_543),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_564),
.Y(n_657)
);

INVx3_ASAP7_75t_L g658 ( 
.A(n_606),
.Y(n_658)
);

NOR2xp33_ASAP7_75t_L g659 ( 
.A(n_596),
.B(n_484),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_539),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_539),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_SL g662 ( 
.A(n_598),
.B(n_487),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_539),
.Y(n_663)
);

NOR2xp33_ASAP7_75t_L g664 ( 
.A(n_596),
.B(n_491),
.Y(n_664)
);

BUFx3_ASAP7_75t_L g665 ( 
.A(n_555),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_539),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_542),
.Y(n_667)
);

OR2x2_ASAP7_75t_L g668 ( 
.A(n_548),
.B(n_430),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_SL g669 ( 
.A(n_598),
.B(n_497),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_564),
.Y(n_670)
);

AOI22xp5_ASAP7_75t_L g671 ( 
.A1(n_585),
.A2(n_500),
.B1(n_511),
.B2(n_499),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_542),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_564),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_542),
.Y(n_674)
);

INVxp33_ASAP7_75t_L g675 ( 
.A(n_548),
.Y(n_675)
);

AND2x2_ASAP7_75t_SL g676 ( 
.A(n_559),
.B(n_267),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_542),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_564),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_564),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_585),
.B(n_528),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_564),
.Y(n_681)
);

NOR3xp33_ASAP7_75t_L g682 ( 
.A(n_598),
.B(n_519),
.C(n_518),
.Y(n_682)
);

HB1xp67_ASAP7_75t_L g683 ( 
.A(n_584),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_588),
.B(n_528),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_564),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_565),
.Y(n_686)
);

CKINVDCx20_ASAP7_75t_R g687 ( 
.A(n_611),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_565),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_565),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_573),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_588),
.B(n_528),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_565),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_565),
.Y(n_693)
);

BUFx3_ASAP7_75t_L g694 ( 
.A(n_555),
.Y(n_694)
);

AND2x2_ASAP7_75t_L g695 ( 
.A(n_588),
.B(n_609),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_565),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_SL g697 ( 
.A(n_611),
.B(n_524),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_565),
.Y(n_698)
);

AOI22xp5_ASAP7_75t_L g699 ( 
.A1(n_609),
.A2(n_526),
.B1(n_529),
.B2(n_502),
.Y(n_699)
);

NAND2xp33_ASAP7_75t_L g700 ( 
.A(n_565),
.B(n_408),
.Y(n_700)
);

NAND2xp33_ASAP7_75t_L g701 ( 
.A(n_577),
.B(n_408),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_SL g702 ( 
.A(n_611),
.B(n_504),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_609),
.B(n_523),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_577),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_SL g705 ( 
.A(n_596),
.B(n_431),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_592),
.B(n_530),
.Y(n_706)
);

NOR2xp33_ASAP7_75t_L g707 ( 
.A(n_592),
.B(n_441),
.Y(n_707)
);

OAI22xp33_ASAP7_75t_SL g708 ( 
.A1(n_552),
.A2(n_493),
.B1(n_516),
.B2(n_515),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_577),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_L g710 ( 
.A(n_592),
.B(n_474),
.Y(n_710)
);

INVx3_ASAP7_75t_L g711 ( 
.A(n_606),
.Y(n_711)
);

BUFx6f_ASAP7_75t_L g712 ( 
.A(n_577),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_577),
.Y(n_713)
);

NOR2x1p5_ASAP7_75t_L g714 ( 
.A(n_573),
.B(n_434),
.Y(n_714)
);

XNOR2x2_ASAP7_75t_L g715 ( 
.A(n_610),
.B(n_531),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_577),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_592),
.B(n_530),
.Y(n_717)
);

INVx3_ASAP7_75t_L g718 ( 
.A(n_606),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_577),
.Y(n_719)
);

CKINVDCx20_ASAP7_75t_R g720 ( 
.A(n_573),
.Y(n_720)
);

AND2x6_ASAP7_75t_L g721 ( 
.A(n_547),
.B(n_314),
.Y(n_721)
);

BUFx8_ASAP7_75t_SL g722 ( 
.A(n_540),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_SL g723 ( 
.A(n_552),
.B(n_527),
.Y(n_723)
);

INVx5_ASAP7_75t_L g724 ( 
.A(n_572),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_577),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_582),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_582),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_592),
.B(n_464),
.Y(n_728)
);

NOR2xp33_ASAP7_75t_L g729 ( 
.A(n_592),
.B(n_464),
.Y(n_729)
);

INVx1_ASAP7_75t_SL g730 ( 
.A(n_584),
.Y(n_730)
);

OAI22xp5_ASAP7_75t_L g731 ( 
.A1(n_556),
.A2(n_342),
.B1(n_343),
.B2(n_341),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_582),
.Y(n_732)
);

BUFx2_ASAP7_75t_L g733 ( 
.A(n_535),
.Y(n_733)
);

BUFx6f_ASAP7_75t_L g734 ( 
.A(n_582),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_582),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_582),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_SL g737 ( 
.A(n_535),
.B(n_387),
.Y(n_737)
);

AND2x2_ASAP7_75t_L g738 ( 
.A(n_557),
.B(n_387),
.Y(n_738)
);

INVx4_ASAP7_75t_L g739 ( 
.A(n_555),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_582),
.Y(n_740)
);

INVx6_ASAP7_75t_L g741 ( 
.A(n_547),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_582),
.Y(n_742)
);

INVx2_ASAP7_75t_SL g743 ( 
.A(n_535),
.Y(n_743)
);

INVxp67_ASAP7_75t_SL g744 ( 
.A(n_566),
.Y(n_744)
);

INVx2_ASAP7_75t_SL g745 ( 
.A(n_606),
.Y(n_745)
);

AND2x2_ASAP7_75t_L g746 ( 
.A(n_557),
.B(n_265),
.Y(n_746)
);

NAND2xp33_ASAP7_75t_L g747 ( 
.A(n_586),
.B(n_587),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_555),
.B(n_335),
.Y(n_748)
);

INVx4_ASAP7_75t_L g749 ( 
.A(n_555),
.Y(n_749)
);

NOR2xp33_ASAP7_75t_L g750 ( 
.A(n_579),
.B(n_248),
.Y(n_750)
);

INVx3_ASAP7_75t_L g751 ( 
.A(n_606),
.Y(n_751)
);

NOR2xp33_ASAP7_75t_L g752 ( 
.A(n_581),
.B(n_330),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_563),
.B(n_338),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_586),
.Y(n_754)
);

BUFx10_ASAP7_75t_L g755 ( 
.A(n_547),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_586),
.Y(n_756)
);

INVx3_ASAP7_75t_L g757 ( 
.A(n_586),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_586),
.Y(n_758)
);

NOR3xp33_ASAP7_75t_L g759 ( 
.A(n_610),
.B(n_277),
.C(n_276),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_586),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_586),
.Y(n_761)
);

INVx5_ASAP7_75t_L g762 ( 
.A(n_572),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_586),
.Y(n_763)
);

BUFx4f_ASAP7_75t_L g764 ( 
.A(n_587),
.Y(n_764)
);

AND2x2_ASAP7_75t_L g765 ( 
.A(n_557),
.B(n_276),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_SL g766 ( 
.A(n_563),
.B(n_346),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_587),
.Y(n_767)
);

BUFx6f_ASAP7_75t_L g768 ( 
.A(n_587),
.Y(n_768)
);

INVx1_ASAP7_75t_SL g769 ( 
.A(n_616),
.Y(n_769)
);

INVx3_ASAP7_75t_L g770 ( 
.A(n_587),
.Y(n_770)
);

OAI221xp5_ASAP7_75t_L g771 ( 
.A1(n_623),
.A2(n_317),
.B1(n_320),
.B2(n_379),
.C(n_312),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_769),
.B(n_563),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_SL g773 ( 
.A(n_739),
.B(n_587),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_619),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_622),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_SL g776 ( 
.A(n_739),
.B(n_587),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_624),
.B(n_563),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_622),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_651),
.B(n_563),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_SL g780 ( 
.A(n_671),
.B(n_589),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_619),
.Y(n_781)
);

INVx1_ASAP7_75t_SL g782 ( 
.A(n_635),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_665),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_632),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_744),
.B(n_589),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_632),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_SL g787 ( 
.A(n_652),
.B(n_589),
.Y(n_787)
);

INVx2_ASAP7_75t_SL g788 ( 
.A(n_646),
.Y(n_788)
);

AO221x1_ASAP7_75t_L g789 ( 
.A1(n_647),
.A2(n_408),
.B1(n_399),
.B2(n_324),
.C(n_312),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_695),
.B(n_589),
.Y(n_790)
);

INVx2_ASAP7_75t_SL g791 ( 
.A(n_730),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_695),
.B(n_589),
.Y(n_792)
);

OAI22xp33_ASAP7_75t_L g793 ( 
.A1(n_652),
.A2(n_616),
.B1(n_566),
.B2(n_593),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_665),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_SL g795 ( 
.A(n_739),
.B(n_587),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_SL g796 ( 
.A(n_729),
.B(n_633),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_639),
.Y(n_797)
);

NOR2xp33_ASAP7_75t_L g798 ( 
.A(n_653),
.B(n_613),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_638),
.B(n_594),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_SL g800 ( 
.A(n_699),
.B(n_594),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_654),
.B(n_594),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_694),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_659),
.B(n_594),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_664),
.B(n_594),
.Y(n_804)
);

AOI22xp5_ASAP7_75t_L g805 ( 
.A1(n_676),
.A2(n_567),
.B1(n_559),
.B2(n_613),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_694),
.Y(n_806)
);

NOR2xp33_ASAP7_75t_L g807 ( 
.A(n_645),
.B(n_605),
.Y(n_807)
);

NAND2xp33_ASAP7_75t_L g808 ( 
.A(n_630),
.B(n_591),
.Y(n_808)
);

BUFx5_ASAP7_75t_L g809 ( 
.A(n_621),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_703),
.B(n_605),
.Y(n_810)
);

INVx8_ASAP7_75t_L g811 ( 
.A(n_721),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_707),
.B(n_605),
.Y(n_812)
);

NOR2xp33_ASAP7_75t_L g813 ( 
.A(n_637),
.B(n_605),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_639),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_SL g815 ( 
.A(n_749),
.B(n_591),
.Y(n_815)
);

NOR2xp33_ASAP7_75t_L g816 ( 
.A(n_648),
.B(n_605),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_641),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_SL g818 ( 
.A(n_749),
.B(n_591),
.Y(n_818)
);

AND2x2_ASAP7_75t_L g819 ( 
.A(n_738),
.B(n_427),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_SL g820 ( 
.A(n_749),
.B(n_591),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_710),
.B(n_550),
.Y(n_821)
);

AND2x2_ASAP7_75t_L g822 ( 
.A(n_738),
.B(n_439),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_641),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_741),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_741),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_SL g826 ( 
.A(n_745),
.B(n_591),
.Y(n_826)
);

INVx2_ASAP7_75t_SL g827 ( 
.A(n_668),
.Y(n_827)
);

NOR2xp33_ASAP7_75t_L g828 ( 
.A(n_743),
.B(n_733),
.Y(n_828)
);

OR2x2_ASAP7_75t_L g829 ( 
.A(n_668),
.B(n_581),
.Y(n_829)
);

INVx2_ASAP7_75t_SL g830 ( 
.A(n_683),
.Y(n_830)
);

INVx3_ASAP7_75t_L g831 ( 
.A(n_755),
.Y(n_831)
);

AOI22xp33_ASAP7_75t_L g832 ( 
.A1(n_759),
.A2(n_567),
.B1(n_595),
.B2(n_593),
.Y(n_832)
);

OAI22xp5_ASAP7_75t_L g833 ( 
.A1(n_676),
.A2(n_554),
.B1(n_562),
.B2(n_550),
.Y(n_833)
);

BUFx5_ASAP7_75t_L g834 ( 
.A(n_621),
.Y(n_834)
);

INVxp67_ASAP7_75t_L g835 ( 
.A(n_656),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_680),
.B(n_554),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_684),
.B(n_562),
.Y(n_837)
);

AOI22xp5_ASAP7_75t_L g838 ( 
.A1(n_743),
.A2(n_597),
.B1(n_604),
.B2(n_595),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_SL g839 ( 
.A(n_682),
.B(n_562),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_691),
.B(n_568),
.Y(n_840)
);

AND2x2_ASAP7_75t_L g841 ( 
.A(n_675),
.B(n_440),
.Y(n_841)
);

CKINVDCx20_ASAP7_75t_R g842 ( 
.A(n_620),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_660),
.Y(n_843)
);

INVxp67_ASAP7_75t_L g844 ( 
.A(n_723),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_750),
.B(n_568),
.Y(n_845)
);

NAND3xp33_ASAP7_75t_SL g846 ( 
.A(n_643),
.B(n_453),
.C(n_446),
.Y(n_846)
);

AOI22xp33_ASAP7_75t_L g847 ( 
.A1(n_626),
.A2(n_604),
.B1(n_614),
.B2(n_597),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_752),
.B(n_568),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_661),
.Y(n_849)
);

O2A1O1Ixp5_ASAP7_75t_L g850 ( 
.A1(n_766),
.A2(n_614),
.B(n_590),
.C(n_603),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_741),
.Y(n_851)
);

NOR2xp33_ASAP7_75t_L g852 ( 
.A(n_733),
.B(n_569),
.Y(n_852)
);

BUFx3_ASAP7_75t_L g853 ( 
.A(n_755),
.Y(n_853)
);

NOR2xp67_ASAP7_75t_L g854 ( 
.A(n_625),
.B(n_551),
.Y(n_854)
);

NOR2xp33_ASAP7_75t_L g855 ( 
.A(n_640),
.B(n_569),
.Y(n_855)
);

INVx2_ASAP7_75t_SL g856 ( 
.A(n_640),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_SL g857 ( 
.A(n_644),
.B(n_728),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_661),
.Y(n_858)
);

AOI22xp5_ASAP7_75t_L g859 ( 
.A1(n_721),
.A2(n_590),
.B1(n_603),
.B2(n_569),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_748),
.B(n_590),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_663),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_753),
.B(n_603),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_741),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_746),
.B(n_615),
.Y(n_864)
);

BUFx6f_ASAP7_75t_L g865 ( 
.A(n_630),
.Y(n_865)
);

AND2x6_ASAP7_75t_L g866 ( 
.A(n_636),
.B(n_615),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_746),
.B(n_765),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_SL g868 ( 
.A(n_745),
.B(n_591),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_663),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_755),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_765),
.B(n_615),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_SL g872 ( 
.A(n_636),
.B(n_591),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_666),
.Y(n_873)
);

NOR2xp33_ASAP7_75t_L g874 ( 
.A(n_705),
.B(n_617),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_721),
.B(n_617),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_SL g876 ( 
.A(n_708),
.B(n_617),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_721),
.B(n_551),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_721),
.B(n_551),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_666),
.Y(n_879)
);

NOR2xp33_ASAP7_75t_L g880 ( 
.A(n_737),
.B(n_551),
.Y(n_880)
);

BUFx6f_ASAP7_75t_L g881 ( 
.A(n_630),
.Y(n_881)
);

AND2x2_ASAP7_75t_L g882 ( 
.A(n_702),
.B(n_456),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_721),
.B(n_553),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_667),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_SL g885 ( 
.A(n_662),
.B(n_591),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_667),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_672),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_721),
.B(n_553),
.Y(n_888)
);

INVx2_ASAP7_75t_L g889 ( 
.A(n_672),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_674),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_636),
.B(n_553),
.Y(n_891)
);

NAND3xp33_ASAP7_75t_L g892 ( 
.A(n_669),
.B(n_600),
.C(n_599),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_674),
.Y(n_893)
);

NOR2xp33_ASAP7_75t_L g894 ( 
.A(n_697),
.B(n_553),
.Y(n_894)
);

AOI22xp33_ASAP7_75t_L g895 ( 
.A1(n_658),
.A2(n_547),
.B1(n_618),
.B2(n_607),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_SL g896 ( 
.A(n_731),
.B(n_599),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_658),
.B(n_560),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_677),
.Y(n_898)
);

INVx3_ASAP7_75t_L g899 ( 
.A(n_658),
.Y(n_899)
);

OR2x6_ASAP7_75t_L g900 ( 
.A(n_714),
.B(n_547),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_677),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_711),
.B(n_560),
.Y(n_902)
);

BUFx6f_ASAP7_75t_SL g903 ( 
.A(n_722),
.Y(n_903)
);

OAI221xp5_ASAP7_75t_L g904 ( 
.A1(n_642),
.A2(n_320),
.B1(n_354),
.B2(n_352),
.C(n_344),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_711),
.Y(n_905)
);

AO221x1_ASAP7_75t_L g906 ( 
.A1(n_715),
.A2(n_408),
.B1(n_364),
.B2(n_277),
.C(n_413),
.Y(n_906)
);

NOR2xp33_ASAP7_75t_L g907 ( 
.A(n_711),
.B(n_560),
.Y(n_907)
);

NOR2xp33_ASAP7_75t_L g908 ( 
.A(n_718),
.B(n_560),
.Y(n_908)
);

NOR2xp33_ASAP7_75t_L g909 ( 
.A(n_718),
.B(n_570),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_718),
.Y(n_910)
);

NOR2xp33_ASAP7_75t_L g911 ( 
.A(n_751),
.B(n_570),
.Y(n_911)
);

NOR2xp33_ASAP7_75t_L g912 ( 
.A(n_751),
.B(n_570),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_751),
.Y(n_913)
);

AND2x4_ASAP7_75t_L g914 ( 
.A(n_714),
.B(n_547),
.Y(n_914)
);

BUFx3_ASAP7_75t_L g915 ( 
.A(n_630),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_706),
.B(n_570),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_717),
.B(n_571),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_757),
.B(n_571),
.Y(n_918)
);

NOR2xp33_ASAP7_75t_L g919 ( 
.A(n_757),
.B(n_571),
.Y(n_919)
);

INVx4_ASAP7_75t_L g920 ( 
.A(n_630),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_757),
.B(n_571),
.Y(n_921)
);

INVx4_ASAP7_75t_L g922 ( 
.A(n_649),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_SL g923 ( 
.A(n_649),
.B(n_599),
.Y(n_923)
);

NOR2xp33_ASAP7_75t_L g924 ( 
.A(n_770),
.B(n_574),
.Y(n_924)
);

AOI22xp33_ASAP7_75t_L g925 ( 
.A1(n_715),
.A2(n_618),
.B1(n_607),
.B2(n_600),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_627),
.Y(n_926)
);

NOR2xp33_ASAP7_75t_L g927 ( 
.A(n_770),
.B(n_574),
.Y(n_927)
);

NOR2xp33_ASAP7_75t_L g928 ( 
.A(n_770),
.B(n_574),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_627),
.Y(n_929)
);

AOI21xp5_ASAP7_75t_L g930 ( 
.A1(n_764),
.A2(n_576),
.B(n_574),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_689),
.B(n_576),
.Y(n_931)
);

NOR2xp33_ASAP7_75t_L g932 ( 
.A(n_628),
.B(n_629),
.Y(n_932)
);

AND2x2_ASAP7_75t_L g933 ( 
.A(n_687),
.B(n_690),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_689),
.Y(n_934)
);

INVx2_ASAP7_75t_SL g935 ( 
.A(n_690),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_SL g936 ( 
.A(n_649),
.B(n_599),
.Y(n_936)
);

OAI22xp5_ASAP7_75t_L g937 ( 
.A1(n_764),
.A2(n_601),
.B1(n_602),
.B2(n_576),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_698),
.B(n_576),
.Y(n_938)
);

INVx2_ASAP7_75t_L g939 ( 
.A(n_698),
.Y(n_939)
);

OAI22xp5_ASAP7_75t_L g940 ( 
.A1(n_764),
.A2(n_602),
.B1(n_608),
.B2(n_601),
.Y(n_940)
);

AOI21xp5_ASAP7_75t_L g941 ( 
.A1(n_872),
.A2(n_747),
.B(n_629),
.Y(n_941)
);

INVx3_ASAP7_75t_L g942 ( 
.A(n_853),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_SL g943 ( 
.A(n_853),
.B(n_649),
.Y(n_943)
);

CKINVDCx20_ASAP7_75t_R g944 ( 
.A(n_842),
.Y(n_944)
);

INVx4_ASAP7_75t_L g945 ( 
.A(n_811),
.Y(n_945)
);

AOI22xp33_ASAP7_75t_L g946 ( 
.A1(n_925),
.A2(n_473),
.B1(n_476),
.B2(n_458),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_SL g947 ( 
.A(n_782),
.B(n_768),
.Y(n_947)
);

AOI21xp5_ASAP7_75t_L g948 ( 
.A1(n_872),
.A2(n_747),
.B(n_631),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_855),
.B(n_601),
.Y(n_949)
);

O2A1O1Ixp33_ASAP7_75t_L g950 ( 
.A1(n_867),
.A2(n_602),
.B(n_608),
.C(n_601),
.Y(n_950)
);

NOR2xp33_ASAP7_75t_L g951 ( 
.A(n_788),
.B(n_480),
.Y(n_951)
);

O2A1O1Ixp33_ASAP7_75t_L g952 ( 
.A1(n_771),
.A2(n_608),
.B(n_612),
.C(n_602),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_843),
.Y(n_953)
);

NAND2xp33_ASAP7_75t_L g954 ( 
.A(n_866),
.B(n_649),
.Y(n_954)
);

OAI22xp5_ASAP7_75t_L g955 ( 
.A1(n_777),
.A2(n_631),
.B1(n_650),
.B2(n_628),
.Y(n_955)
);

OR2x6_ASAP7_75t_L g956 ( 
.A(n_811),
.B(n_720),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_855),
.B(n_852),
.Y(n_957)
);

INVx3_ASAP7_75t_L g958 ( 
.A(n_831),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_852),
.B(n_608),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_796),
.B(n_612),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_828),
.B(n_612),
.Y(n_961)
);

OAI22xp5_ASAP7_75t_L g962 ( 
.A1(n_828),
.A2(n_650),
.B1(n_657),
.B2(n_655),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_772),
.B(n_612),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_856),
.B(n_599),
.Y(n_964)
);

AOI22xp33_ASAP7_75t_L g965 ( 
.A1(n_906),
.A2(n_494),
.B1(n_501),
.B2(n_490),
.Y(n_965)
);

AOI21x1_ASAP7_75t_L g966 ( 
.A1(n_773),
.A2(n_657),
.B(n_655),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_845),
.B(n_848),
.Y(n_967)
);

NAND2xp33_ASAP7_75t_L g968 ( 
.A(n_866),
.B(n_712),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_864),
.B(n_599),
.Y(n_969)
);

AOI21xp5_ASAP7_75t_L g970 ( 
.A1(n_826),
.A2(n_673),
.B(n_670),
.Y(n_970)
);

A2O1A1Ixp33_ASAP7_75t_L g971 ( 
.A1(n_798),
.A2(n_716),
.B(n_726),
.C(n_713),
.Y(n_971)
);

AND2x2_ASAP7_75t_L g972 ( 
.A(n_791),
.B(n_607),
.Y(n_972)
);

INVx2_ASAP7_75t_L g973 ( 
.A(n_843),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_871),
.B(n_599),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_894),
.B(n_599),
.Y(n_975)
);

AOI21xp5_ASAP7_75t_L g976 ( 
.A1(n_826),
.A2(n_868),
.B(n_891),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_894),
.B(n_600),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_793),
.B(n_600),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_790),
.B(n_600),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_775),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_SL g981 ( 
.A(n_831),
.B(n_870),
.Y(n_981)
);

INVx3_ASAP7_75t_L g982 ( 
.A(n_811),
.Y(n_982)
);

OAI21xp5_ASAP7_75t_L g983 ( 
.A1(n_907),
.A2(n_673),
.B(n_670),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_792),
.B(n_600),
.Y(n_984)
);

AND2x2_ASAP7_75t_L g985 ( 
.A(n_819),
.B(n_607),
.Y(n_985)
);

AND3x1_ASAP7_75t_SL g986 ( 
.A(n_904),
.B(n_298),
.C(n_287),
.Y(n_986)
);

AOI21xp5_ASAP7_75t_L g987 ( 
.A1(n_868),
.A2(n_679),
.B(n_678),
.Y(n_987)
);

OAI21xp33_ASAP7_75t_L g988 ( 
.A1(n_874),
.A2(n_829),
.B(n_838),
.Y(n_988)
);

INVx3_ASAP7_75t_L g989 ( 
.A(n_920),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_778),
.Y(n_990)
);

AOI22xp5_ASAP7_75t_L g991 ( 
.A1(n_827),
.A2(n_679),
.B1(n_681),
.B2(n_678),
.Y(n_991)
);

AOI21xp5_ASAP7_75t_L g992 ( 
.A1(n_897),
.A2(n_685),
.B(n_681),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_832),
.B(n_600),
.Y(n_993)
);

O2A1O1Ixp33_ASAP7_75t_L g994 ( 
.A1(n_836),
.A2(n_298),
.B(n_310),
.C(n_287),
.Y(n_994)
);

OR2x6_ASAP7_75t_SL g995 ( 
.A(n_903),
.B(n_349),
.Y(n_995)
);

OAI21xp5_ASAP7_75t_L g996 ( 
.A1(n_907),
.A2(n_686),
.B(n_685),
.Y(n_996)
);

AOI21xp5_ASAP7_75t_L g997 ( 
.A1(n_902),
.A2(n_688),
.B(n_686),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_813),
.B(n_600),
.Y(n_998)
);

A2O1A1Ixp33_ASAP7_75t_L g999 ( 
.A1(n_798),
.A2(n_716),
.B(n_726),
.C(n_713),
.Y(n_999)
);

A2O1A1Ixp33_ASAP7_75t_L g1000 ( 
.A1(n_807),
.A2(n_742),
.B(n_763),
.C(n_732),
.Y(n_1000)
);

INVx2_ASAP7_75t_L g1001 ( 
.A(n_849),
.Y(n_1001)
);

BUFx6f_ASAP7_75t_L g1002 ( 
.A(n_865),
.Y(n_1002)
);

NAND2x1_ASAP7_75t_L g1003 ( 
.A(n_866),
.B(n_688),
.Y(n_1003)
);

OAI21xp5_ASAP7_75t_L g1004 ( 
.A1(n_908),
.A2(n_693),
.B(n_692),
.Y(n_1004)
);

O2A1O1Ixp33_ASAP7_75t_L g1005 ( 
.A1(n_787),
.A2(n_311),
.B(n_317),
.C(n_310),
.Y(n_1005)
);

NOR2x2_ASAP7_75t_L g1006 ( 
.A(n_900),
.B(n_732),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_813),
.B(n_607),
.Y(n_1007)
);

AO21x1_ASAP7_75t_L g1008 ( 
.A1(n_807),
.A2(n_693),
.B(n_692),
.Y(n_1008)
);

CKINVDCx5p33_ASAP7_75t_R g1009 ( 
.A(n_903),
.Y(n_1009)
);

AND2x2_ASAP7_75t_L g1010 ( 
.A(n_822),
.B(n_607),
.Y(n_1010)
);

AOI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_908),
.A2(n_704),
.B(n_696),
.Y(n_1011)
);

AOI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_909),
.A2(n_704),
.B(n_696),
.Y(n_1012)
);

NOR2xp33_ASAP7_75t_L g1013 ( 
.A(n_844),
.B(n_709),
.Y(n_1013)
);

NOR3xp33_ASAP7_75t_L g1014 ( 
.A(n_830),
.B(n_322),
.C(n_311),
.Y(n_1014)
);

AOI21xp5_ASAP7_75t_L g1015 ( 
.A1(n_909),
.A2(n_719),
.B(n_709),
.Y(n_1015)
);

BUFx6f_ASAP7_75t_L g1016 ( 
.A(n_865),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_816),
.B(n_618),
.Y(n_1017)
);

OAI21xp5_ASAP7_75t_L g1018 ( 
.A1(n_911),
.A2(n_725),
.B(n_719),
.Y(n_1018)
);

OAI321xp33_ASAP7_75t_L g1019 ( 
.A1(n_805),
.A2(n_399),
.A3(n_322),
.B1(n_324),
.B2(n_326),
.C(n_344),
.Y(n_1019)
);

OAI22xp5_ASAP7_75t_L g1020 ( 
.A1(n_779),
.A2(n_725),
.B1(n_735),
.B2(n_727),
.Y(n_1020)
);

AOI21x1_ASAP7_75t_L g1021 ( 
.A1(n_773),
.A2(n_735),
.B(n_727),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_816),
.B(n_618),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_847),
.B(n_618),
.Y(n_1023)
);

AOI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_911),
.A2(n_740),
.B(n_736),
.Y(n_1024)
);

BUFx6f_ASAP7_75t_L g1025 ( 
.A(n_865),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_785),
.B(n_618),
.Y(n_1026)
);

INVx1_ASAP7_75t_SL g1027 ( 
.A(n_841),
.Y(n_1027)
);

AOI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_912),
.A2(n_740),
.B(n_736),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_817),
.Y(n_1029)
);

AOI21x1_ASAP7_75t_L g1030 ( 
.A1(n_776),
.A2(n_756),
.B(n_754),
.Y(n_1030)
);

NOR2x1_ASAP7_75t_L g1031 ( 
.A(n_900),
.B(n_754),
.Y(n_1031)
);

OAI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_912),
.A2(n_758),
.B(n_756),
.Y(n_1032)
);

AOI21xp33_ASAP7_75t_L g1033 ( 
.A1(n_880),
.A2(n_760),
.B(n_758),
.Y(n_1033)
);

AOI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_812),
.A2(n_761),
.B(n_760),
.Y(n_1034)
);

OAI22xp5_ASAP7_75t_L g1035 ( 
.A1(n_859),
.A2(n_799),
.B1(n_803),
.B2(n_801),
.Y(n_1035)
);

BUFx2_ASAP7_75t_L g1036 ( 
.A(n_933),
.Y(n_1036)
);

INVx2_ASAP7_75t_SL g1037 ( 
.A(n_914),
.Y(n_1037)
);

BUFx6f_ASAP7_75t_L g1038 ( 
.A(n_865),
.Y(n_1038)
);

AOI21xp5_ASAP7_75t_L g1039 ( 
.A1(n_804),
.A2(n_767),
.B(n_761),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_SL g1040 ( 
.A(n_935),
.B(n_768),
.Y(n_1040)
);

INVx2_ASAP7_75t_L g1041 ( 
.A(n_849),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_873),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_879),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_SL g1044 ( 
.A(n_914),
.B(n_768),
.Y(n_1044)
);

NOR2xp67_ASAP7_75t_L g1045 ( 
.A(n_835),
.B(n_742),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_886),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_810),
.B(n_763),
.Y(n_1047)
);

NOR2xp33_ASAP7_75t_L g1048 ( 
.A(n_882),
.B(n_767),
.Y(n_1048)
);

BUFx4f_ASAP7_75t_L g1049 ( 
.A(n_900),
.Y(n_1049)
);

HB1xp67_ASAP7_75t_L g1050 ( 
.A(n_914),
.Y(n_1050)
);

NOR3xp33_ASAP7_75t_L g1051 ( 
.A(n_839),
.B(n_846),
.C(n_885),
.Y(n_1051)
);

AOI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_918),
.A2(n_734),
.B(n_712),
.Y(n_1052)
);

OAI21xp5_ASAP7_75t_L g1053 ( 
.A1(n_905),
.A2(n_701),
.B(n_700),
.Y(n_1053)
);

OAI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_905),
.A2(n_701),
.B(n_700),
.Y(n_1054)
);

O2A1O1Ixp33_ASAP7_75t_SL g1055 ( 
.A1(n_776),
.A2(n_389),
.B(n_381),
.C(n_385),
.Y(n_1055)
);

AOI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_921),
.A2(n_734),
.B(n_712),
.Y(n_1056)
);

BUFx3_ASAP7_75t_L g1057 ( 
.A(n_824),
.Y(n_1057)
);

AOI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_931),
.A2(n_734),
.B(n_712),
.Y(n_1058)
);

A2O1A1Ixp33_ASAP7_75t_L g1059 ( 
.A1(n_874),
.A2(n_389),
.B(n_314),
.C(n_321),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_893),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_821),
.B(n_712),
.Y(n_1061)
);

BUFx12f_ASAP7_75t_L g1062 ( 
.A(n_881),
.Y(n_1062)
);

AND2x4_ASAP7_75t_L g1063 ( 
.A(n_825),
.B(n_734),
.Y(n_1063)
);

AOI22xp5_ASAP7_75t_L g1064 ( 
.A1(n_857),
.A2(n_768),
.B1(n_734),
.B2(n_394),
.Y(n_1064)
);

OAI21xp33_ASAP7_75t_L g1065 ( 
.A1(n_860),
.A2(n_365),
.B(n_357),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_901),
.Y(n_1066)
);

AND2x2_ASAP7_75t_L g1067 ( 
.A(n_876),
.B(n_326),
.Y(n_1067)
);

BUFx12f_ASAP7_75t_L g1068 ( 
.A(n_881),
.Y(n_1068)
);

A2O1A1Ixp33_ASAP7_75t_L g1069 ( 
.A1(n_880),
.A2(n_397),
.B(n_321),
.C(n_323),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_774),
.Y(n_1070)
);

OAI22xp5_ASAP7_75t_L g1071 ( 
.A1(n_833),
.A2(n_768),
.B1(n_367),
.B2(n_369),
.Y(n_1071)
);

AND2x2_ASAP7_75t_SL g1072 ( 
.A(n_895),
.B(n_352),
.Y(n_1072)
);

INVx11_ASAP7_75t_L g1073 ( 
.A(n_866),
.Y(n_1073)
);

NOR2xp33_ASAP7_75t_L g1074 ( 
.A(n_851),
.B(n_375),
.Y(n_1074)
);

AOI22xp33_ASAP7_75t_L g1075 ( 
.A1(n_789),
.A2(n_390),
.B1(n_392),
.B2(n_393),
.Y(n_1075)
);

INVx2_ASAP7_75t_L g1076 ( 
.A(n_858),
.Y(n_1076)
);

AOI21xp5_ASAP7_75t_L g1077 ( 
.A1(n_938),
.A2(n_536),
.B(n_537),
.Y(n_1077)
);

O2A1O1Ixp33_ASAP7_75t_L g1078 ( 
.A1(n_837),
.A2(n_392),
.B(n_414),
.C(n_413),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_862),
.B(n_840),
.Y(n_1079)
);

A2O1A1Ixp33_ASAP7_75t_L g1080 ( 
.A1(n_780),
.A2(n_323),
.B(n_381),
.C(n_385),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_781),
.Y(n_1081)
);

O2A1O1Ixp33_ASAP7_75t_L g1082 ( 
.A1(n_800),
.A2(n_393),
.B(n_390),
.C(n_414),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_SL g1083 ( 
.A(n_863),
.B(n_854),
.Y(n_1083)
);

OAI22xp5_ASAP7_75t_L g1084 ( 
.A1(n_899),
.A2(n_396),
.B1(n_386),
.B2(n_388),
.Y(n_1084)
);

AND2x2_ASAP7_75t_L g1085 ( 
.A(n_783),
.B(n_354),
.Y(n_1085)
);

AO21x2_ASAP7_75t_L g1086 ( 
.A1(n_896),
.A2(n_544),
.B(n_541),
.Y(n_1086)
);

BUFx3_ASAP7_75t_L g1087 ( 
.A(n_794),
.Y(n_1087)
);

A2O1A1Ixp33_ASAP7_75t_L g1088 ( 
.A1(n_932),
.A2(n_351),
.B(n_416),
.C(n_397),
.Y(n_1088)
);

BUFx3_ASAP7_75t_L g1089 ( 
.A(n_802),
.Y(n_1089)
);

AO21x1_ASAP7_75t_L g1090 ( 
.A1(n_930),
.A2(n_415),
.B(n_351),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_806),
.B(n_536),
.Y(n_1091)
);

AO21x1_ASAP7_75t_L g1092 ( 
.A1(n_937),
.A2(n_940),
.B(n_932),
.Y(n_1092)
);

O2A1O1Ixp33_ASAP7_75t_L g1093 ( 
.A1(n_926),
.A2(n_364),
.B(n_378),
.C(n_379),
.Y(n_1093)
);

BUFx5_ASAP7_75t_L g1094 ( 
.A(n_866),
.Y(n_1094)
);

NOR2xp33_ASAP7_75t_SL g1095 ( 
.A(n_875),
.B(n_920),
.Y(n_1095)
);

AOI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_795),
.A2(n_538),
.B(n_537),
.Y(n_1096)
);

INVx11_ASAP7_75t_L g1097 ( 
.A(n_892),
.Y(n_1097)
);

AOI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_795),
.A2(n_538),
.B(n_537),
.Y(n_1098)
);

OAI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_910),
.A2(n_416),
.B(n_415),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_SL g1100 ( 
.A(n_881),
.B(n_809),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_910),
.B(n_378),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_913),
.B(n_377),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_SL g1103 ( 
.A(n_881),
.B(n_380),
.Y(n_1103)
);

AND2x6_ASAP7_75t_L g1104 ( 
.A(n_913),
.B(n_422),
.Y(n_1104)
);

BUFx6f_ASAP7_75t_L g1105 ( 
.A(n_915),
.Y(n_1105)
);

AOI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_815),
.A2(n_538),
.B(n_537),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_919),
.B(n_405),
.Y(n_1107)
);

NOR2xp33_ASAP7_75t_L g1108 ( 
.A(n_899),
.B(n_417),
.Y(n_1108)
);

A2O1A1Ixp33_ASAP7_75t_L g1109 ( 
.A1(n_919),
.A2(n_924),
.B(n_927),
.C(n_928),
.Y(n_1109)
);

AND2x2_ASAP7_75t_L g1110 ( 
.A(n_784),
.B(n_419),
.Y(n_1110)
);

AOI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_815),
.A2(n_538),
.B(n_537),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_924),
.B(n_420),
.Y(n_1112)
);

BUFx6f_ASAP7_75t_L g1113 ( 
.A(n_915),
.Y(n_1113)
);

AND2x2_ASAP7_75t_L g1114 ( 
.A(n_784),
.B(n_541),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_927),
.B(n_370),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_928),
.B(n_401),
.Y(n_1116)
);

AOI22xp33_ASAP7_75t_L g1117 ( 
.A1(n_858),
.A2(n_362),
.B1(n_422),
.B2(n_394),
.Y(n_1117)
);

AOI21xp5_ASAP7_75t_L g1118 ( 
.A1(n_818),
.A2(n_538),
.B(n_537),
.Y(n_1118)
);

AOI22xp5_ASAP7_75t_L g1119 ( 
.A1(n_877),
.A2(n_294),
.B1(n_281),
.B2(n_280),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_SL g1120 ( 
.A(n_809),
.B(n_724),
.Y(n_1120)
);

BUFx2_ASAP7_75t_L g1121 ( 
.A(n_878),
.Y(n_1121)
);

NOR2xp33_ASAP7_75t_L g1122 ( 
.A(n_818),
.B(n_820),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_786),
.B(n_409),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_797),
.B(n_410),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_814),
.Y(n_1125)
);

A2O1A1Ixp33_ASAP7_75t_L g1126 ( 
.A1(n_883),
.A2(n_384),
.B(n_544),
.C(n_538),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_814),
.B(n_537),
.Y(n_1127)
);

NOR2x1_ASAP7_75t_L g1128 ( 
.A(n_944),
.B(n_922),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_957),
.B(n_823),
.Y(n_1129)
);

CKINVDCx20_ASAP7_75t_R g1130 ( 
.A(n_1009),
.Y(n_1130)
);

A2O1A1Ixp33_ASAP7_75t_L g1131 ( 
.A1(n_988),
.A2(n_850),
.B(n_888),
.C(n_929),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_1029),
.Y(n_1132)
);

NOR2xp33_ASAP7_75t_L g1133 ( 
.A(n_951),
.B(n_823),
.Y(n_1133)
);

OAI22xp5_ASAP7_75t_SL g1134 ( 
.A1(n_946),
.A2(n_251),
.B1(n_225),
.B2(n_421),
.Y(n_1134)
);

INVx2_ASAP7_75t_L g1135 ( 
.A(n_953),
.Y(n_1135)
);

O2A1O1Ixp33_ASAP7_75t_L g1136 ( 
.A1(n_967),
.A2(n_820),
.B(n_917),
.C(n_916),
.Y(n_1136)
);

NOR2xp33_ASAP7_75t_R g1137 ( 
.A(n_1062),
.B(n_808),
.Y(n_1137)
);

AOI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_1079),
.A2(n_936),
.B(n_923),
.Y(n_1138)
);

BUFx2_ASAP7_75t_L g1139 ( 
.A(n_1036),
.Y(n_1139)
);

AOI21xp5_ASAP7_75t_L g1140 ( 
.A1(n_954),
.A2(n_936),
.B(n_922),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_1042),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_1072),
.B(n_861),
.Y(n_1142)
);

OAI22x1_ASAP7_75t_L g1143 ( 
.A1(n_1048),
.A2(n_939),
.B1(n_934),
.B2(n_898),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_1043),
.Y(n_1144)
);

BUFx2_ASAP7_75t_L g1145 ( 
.A(n_956),
.Y(n_1145)
);

NOR2xp33_ASAP7_75t_L g1146 ( 
.A(n_1027),
.B(n_934),
.Y(n_1146)
);

OR2x6_ASAP7_75t_SL g1147 ( 
.A(n_1084),
.B(n_230),
.Y(n_1147)
);

O2A1O1Ixp33_ASAP7_75t_L g1148 ( 
.A1(n_1059),
.A2(n_939),
.B(n_898),
.C(n_890),
.Y(n_1148)
);

AOI21xp5_ASAP7_75t_L g1149 ( 
.A1(n_968),
.A2(n_890),
.B(n_869),
.Y(n_1149)
);

AOI21xp5_ASAP7_75t_L g1150 ( 
.A1(n_1035),
.A2(n_869),
.B(n_861),
.Y(n_1150)
);

NOR2xp67_ASAP7_75t_L g1151 ( 
.A(n_1068),
.B(n_884),
.Y(n_1151)
);

OAI21x1_ASAP7_75t_L g1152 ( 
.A1(n_992),
.A2(n_889),
.B(n_887),
.Y(n_1152)
);

CKINVDCx14_ASAP7_75t_R g1153 ( 
.A(n_995),
.Y(n_1153)
);

AOI21xp5_ASAP7_75t_L g1154 ( 
.A1(n_1109),
.A2(n_889),
.B(n_887),
.Y(n_1154)
);

INVx3_ASAP7_75t_SL g1155 ( 
.A(n_956),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_SL g1156 ( 
.A(n_1049),
.B(n_809),
.Y(n_1156)
);

AOI22xp33_ASAP7_75t_L g1157 ( 
.A1(n_965),
.A2(n_884),
.B1(n_834),
.B2(n_809),
.Y(n_1157)
);

AOI22xp5_ASAP7_75t_L g1158 ( 
.A1(n_1037),
.A2(n_809),
.B1(n_834),
.B2(n_340),
.Y(n_1158)
);

OA21x2_ASAP7_75t_L g1159 ( 
.A1(n_1008),
.A2(n_834),
.B(n_809),
.Y(n_1159)
);

INVxp67_ASAP7_75t_L g1160 ( 
.A(n_1067),
.Y(n_1160)
);

AOI21xp5_ASAP7_75t_L g1161 ( 
.A1(n_1061),
.A2(n_834),
.B(n_333),
.Y(n_1161)
);

INVx2_ASAP7_75t_L g1162 ( 
.A(n_973),
.Y(n_1162)
);

AOI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_949),
.A2(n_834),
.B(n_339),
.Y(n_1163)
);

BUFx3_ASAP7_75t_L g1164 ( 
.A(n_956),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_959),
.B(n_834),
.Y(n_1165)
);

BUFx6f_ASAP7_75t_L g1166 ( 
.A(n_1105),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_961),
.B(n_537),
.Y(n_1167)
);

BUFx12f_ASAP7_75t_L g1168 ( 
.A(n_1105),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_1122),
.B(n_538),
.Y(n_1169)
);

A2O1A1Ixp33_ASAP7_75t_SL g1170 ( 
.A1(n_1108),
.A2(n_10),
.B(n_12),
.C(n_14),
.Y(n_1170)
);

AND2x4_ASAP7_75t_L g1171 ( 
.A(n_945),
.B(n_634),
.Y(n_1171)
);

OR2x6_ASAP7_75t_L g1172 ( 
.A(n_945),
.B(n_545),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_1046),
.Y(n_1173)
);

AND2x4_ASAP7_75t_L g1174 ( 
.A(n_1050),
.B(n_1031),
.Y(n_1174)
);

NAND2x1_ASAP7_75t_L g1175 ( 
.A(n_982),
.B(n_538),
.Y(n_1175)
);

AOI22xp5_ASAP7_75t_L g1176 ( 
.A1(n_1051),
.A2(n_328),
.B1(n_236),
.B2(n_246),
.Y(n_1176)
);

A2O1A1Ixp33_ASAP7_75t_L g1177 ( 
.A1(n_1082),
.A2(n_545),
.B(n_549),
.C(n_231),
.Y(n_1177)
);

BUFx12f_ASAP7_75t_L g1178 ( 
.A(n_1105),
.Y(n_1178)
);

AOI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_998),
.A2(n_545),
.B(n_549),
.Y(n_1179)
);

HAxp5_ASAP7_75t_L g1180 ( 
.A(n_986),
.B(n_12),
.CON(n_1180),
.SN(n_1180)
);

O2A1O1Ixp5_ASAP7_75t_L g1181 ( 
.A1(n_1092),
.A2(n_14),
.B(n_15),
.C(n_16),
.Y(n_1181)
);

OAI22xp5_ASAP7_75t_L g1182 ( 
.A1(n_1073),
.A2(n_411),
.B1(n_308),
.B2(n_306),
.Y(n_1182)
);

OAI21xp33_ASAP7_75t_L g1183 ( 
.A1(n_1065),
.A2(n_319),
.B(n_309),
.Y(n_1183)
);

AND2x2_ASAP7_75t_L g1184 ( 
.A(n_985),
.B(n_1010),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_1060),
.Y(n_1185)
);

NOR2xp33_ASAP7_75t_L g1186 ( 
.A(n_1087),
.B(n_1089),
.Y(n_1186)
);

NOR2x1p5_ASAP7_75t_SL g1187 ( 
.A(n_1094),
.B(n_572),
.Y(n_1187)
);

CKINVDCx5p33_ASAP7_75t_R g1188 ( 
.A(n_1057),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_1066),
.Y(n_1189)
);

NAND3xp33_ASAP7_75t_SL g1190 ( 
.A(n_1014),
.B(n_300),
.C(n_296),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_SL g1191 ( 
.A(n_1049),
.B(n_249),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_960),
.B(n_545),
.Y(n_1192)
);

NOR3xp33_ASAP7_75t_SL g1193 ( 
.A(n_1103),
.B(n_1074),
.C(n_1040),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_SL g1194 ( 
.A(n_942),
.B(n_266),
.Y(n_1194)
);

O2A1O1Ixp33_ASAP7_75t_L g1195 ( 
.A1(n_1088),
.A2(n_1069),
.B(n_1078),
.C(n_994),
.Y(n_1195)
);

INVx8_ASAP7_75t_L g1196 ( 
.A(n_1104),
.Y(n_1196)
);

AOI21xp5_ASAP7_75t_L g1197 ( 
.A1(n_1047),
.A2(n_350),
.B(n_269),
.Y(n_1197)
);

AND2x4_ASAP7_75t_L g1198 ( 
.A(n_982),
.B(n_762),
.Y(n_1198)
);

AOI221xp5_ASAP7_75t_SL g1199 ( 
.A1(n_1093),
.A2(n_545),
.B1(n_549),
.B2(n_18),
.C(n_19),
.Y(n_1199)
);

NOR2xp33_ASAP7_75t_L g1200 ( 
.A(n_980),
.B(n_268),
.Y(n_1200)
);

AOI21xp5_ASAP7_75t_L g1201 ( 
.A1(n_1011),
.A2(n_358),
.B(n_282),
.Y(n_1201)
);

CKINVDCx5p33_ASAP7_75t_R g1202 ( 
.A(n_1113),
.Y(n_1202)
);

OAI22xp5_ASAP7_75t_L g1203 ( 
.A1(n_1007),
.A2(n_290),
.B1(n_288),
.B2(n_286),
.Y(n_1203)
);

AOI21xp5_ASAP7_75t_L g1204 ( 
.A1(n_1011),
.A2(n_361),
.B(n_295),
.Y(n_1204)
);

OR2x6_ASAP7_75t_L g1205 ( 
.A(n_1044),
.B(n_545),
.Y(n_1205)
);

AO32x2_ASAP7_75t_L g1206 ( 
.A1(n_962),
.A2(n_545),
.A3(n_549),
.B1(n_20),
.B2(n_22),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_1070),
.B(n_545),
.Y(n_1207)
);

BUFx8_ASAP7_75t_L g1208 ( 
.A(n_1085),
.Y(n_1208)
);

CKINVDCx5p33_ASAP7_75t_R g1209 ( 
.A(n_1113),
.Y(n_1209)
);

BUFx2_ASAP7_75t_L g1210 ( 
.A(n_972),
.Y(n_1210)
);

NOR2xp33_ASAP7_75t_L g1211 ( 
.A(n_990),
.B(n_278),
.Y(n_1211)
);

AOI21xp5_ASAP7_75t_L g1212 ( 
.A1(n_1012),
.A2(n_366),
.B(n_304),
.Y(n_1212)
);

OAI22xp5_ASAP7_75t_L g1213 ( 
.A1(n_1017),
.A2(n_1022),
.B1(n_1026),
.B2(n_978),
.Y(n_1213)
);

A2O1A1Ixp33_ASAP7_75t_SL g1214 ( 
.A1(n_950),
.A2(n_16),
.B(n_17),
.C(n_20),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_1101),
.Y(n_1215)
);

NOR2xp33_ASAP7_75t_R g1216 ( 
.A(n_942),
.B(n_303),
.Y(n_1216)
);

A2O1A1Ixp33_ASAP7_75t_SL g1217 ( 
.A1(n_950),
.A2(n_17),
.B(n_22),
.C(n_24),
.Y(n_1217)
);

OAI21xp33_ASAP7_75t_L g1218 ( 
.A1(n_1107),
.A2(n_305),
.B(n_407),
.Y(n_1218)
);

A2O1A1Ixp33_ASAP7_75t_L g1219 ( 
.A1(n_1082),
.A2(n_549),
.B(n_316),
.C(n_327),
.Y(n_1219)
);

BUFx2_ASAP7_75t_L g1220 ( 
.A(n_1006),
.Y(n_1220)
);

INVx2_ASAP7_75t_L g1221 ( 
.A(n_1001),
.Y(n_1221)
);

AOI21xp5_ASAP7_75t_L g1222 ( 
.A1(n_1012),
.A2(n_382),
.B(n_353),
.Y(n_1222)
);

OAI21xp5_ASAP7_75t_L g1223 ( 
.A1(n_976),
.A2(n_572),
.B(n_578),
.Y(n_1223)
);

INVx2_ASAP7_75t_L g1224 ( 
.A(n_1041),
.Y(n_1224)
);

O2A1O1Ixp33_ASAP7_75t_SL g1225 ( 
.A1(n_1100),
.A2(n_24),
.B(n_26),
.C(n_27),
.Y(n_1225)
);

BUFx6f_ASAP7_75t_L g1226 ( 
.A(n_1113),
.Y(n_1226)
);

INVx2_ASAP7_75t_L g1227 ( 
.A(n_1076),
.Y(n_1227)
);

AOI21xp5_ASAP7_75t_L g1228 ( 
.A1(n_1015),
.A2(n_383),
.B(n_359),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_L g1229 ( 
.A(n_1081),
.B(n_549),
.Y(n_1229)
);

AOI21xp5_ASAP7_75t_L g1230 ( 
.A1(n_1015),
.A2(n_398),
.B(n_371),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_SL g1231 ( 
.A(n_1094),
.B(n_345),
.Y(n_1231)
);

AOI21xp5_ASAP7_75t_L g1232 ( 
.A1(n_1024),
.A2(n_402),
.B(n_347),
.Y(n_1232)
);

INVx4_ASAP7_75t_L g1233 ( 
.A(n_1002),
.Y(n_1233)
);

CKINVDCx16_ASAP7_75t_R g1234 ( 
.A(n_1110),
.Y(n_1234)
);

OR2x6_ASAP7_75t_L g1235 ( 
.A(n_1045),
.B(n_549),
.Y(n_1235)
);

OAI22xp5_ASAP7_75t_L g1236 ( 
.A1(n_1099),
.A2(n_348),
.B1(n_376),
.B2(n_406),
.Y(n_1236)
);

AOI21xp5_ASAP7_75t_L g1237 ( 
.A1(n_1024),
.A2(n_724),
.B(n_762),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_1125),
.B(n_1121),
.Y(n_1238)
);

AOI21xp5_ASAP7_75t_L g1239 ( 
.A1(n_1028),
.A2(n_724),
.B(n_762),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1091),
.Y(n_1240)
);

O2A1O1Ixp33_ASAP7_75t_L g1241 ( 
.A1(n_994),
.A2(n_27),
.B(n_28),
.C(n_29),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_L g1242 ( 
.A(n_963),
.B(n_549),
.Y(n_1242)
);

O2A1O1Ixp33_ASAP7_75t_SL g1243 ( 
.A1(n_1003),
.A2(n_28),
.B(n_31),
.C(n_32),
.Y(n_1243)
);

INVx2_ASAP7_75t_L g1244 ( 
.A(n_1114),
.Y(n_1244)
);

NOR2xp33_ASAP7_75t_L g1245 ( 
.A(n_1013),
.B(n_32),
.Y(n_1245)
);

INVx2_ASAP7_75t_L g1246 ( 
.A(n_1127),
.Y(n_1246)
);

NAND3xp33_ASAP7_75t_SL g1247 ( 
.A(n_1078),
.B(n_33),
.C(n_35),
.Y(n_1247)
);

BUFx3_ASAP7_75t_L g1248 ( 
.A(n_1063),
.Y(n_1248)
);

BUFx3_ASAP7_75t_L g1249 ( 
.A(n_1063),
.Y(n_1249)
);

BUFx2_ASAP7_75t_L g1250 ( 
.A(n_1104),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_SL g1251 ( 
.A(n_1094),
.B(n_724),
.Y(n_1251)
);

BUFx2_ASAP7_75t_L g1252 ( 
.A(n_1104),
.Y(n_1252)
);

CKINVDCx14_ASAP7_75t_R g1253 ( 
.A(n_1002),
.Y(n_1253)
);

CKINVDCx6p67_ASAP7_75t_R g1254 ( 
.A(n_1104),
.Y(n_1254)
);

INVx6_ASAP7_75t_L g1255 ( 
.A(n_1002),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_L g1256 ( 
.A(n_969),
.B(n_578),
.Y(n_1256)
);

A2O1A1Ixp33_ASAP7_75t_L g1257 ( 
.A1(n_1019),
.A2(n_313),
.B(n_724),
.C(n_634),
.Y(n_1257)
);

NOR2xp33_ASAP7_75t_SL g1258 ( 
.A(n_1094),
.B(n_724),
.Y(n_1258)
);

AOI21xp5_ASAP7_75t_L g1259 ( 
.A1(n_1028),
.A2(n_762),
.B(n_634),
.Y(n_1259)
);

INVx3_ASAP7_75t_L g1260 ( 
.A(n_1016),
.Y(n_1260)
);

OAI21x1_ASAP7_75t_L g1261 ( 
.A1(n_992),
.A2(n_578),
.B(n_572),
.Y(n_1261)
);

AND2x4_ASAP7_75t_L g1262 ( 
.A(n_958),
.B(n_762),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_952),
.Y(n_1263)
);

NAND3xp33_ASAP7_75t_L g1264 ( 
.A(n_1080),
.B(n_313),
.C(n_634),
.Y(n_1264)
);

BUFx6f_ASAP7_75t_L g1265 ( 
.A(n_1016),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_952),
.Y(n_1266)
);

INVx2_ASAP7_75t_L g1267 ( 
.A(n_964),
.Y(n_1267)
);

BUFx2_ASAP7_75t_L g1268 ( 
.A(n_1104),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_L g1269 ( 
.A(n_974),
.B(n_578),
.Y(n_1269)
);

AOI21xp5_ASAP7_75t_L g1270 ( 
.A1(n_976),
.A2(n_634),
.B(n_313),
.Y(n_1270)
);

INVxp67_ASAP7_75t_L g1271 ( 
.A(n_1102),
.Y(n_1271)
);

AOI21xp5_ASAP7_75t_L g1272 ( 
.A1(n_1058),
.A2(n_96),
.B(n_213),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1123),
.Y(n_1273)
);

OAI22xp5_ASAP7_75t_SL g1274 ( 
.A1(n_1075),
.A2(n_1115),
.B1(n_1116),
.B2(n_1119),
.Y(n_1274)
);

AOI22xp33_ASAP7_75t_L g1275 ( 
.A1(n_1023),
.A2(n_578),
.B1(n_572),
.B2(n_40),
.Y(n_1275)
);

O2A1O1Ixp33_ASAP7_75t_SL g1276 ( 
.A1(n_943),
.A2(n_38),
.B(n_39),
.C(n_40),
.Y(n_1276)
);

BUFx3_ASAP7_75t_L g1277 ( 
.A(n_1016),
.Y(n_1277)
);

A2O1A1Ixp33_ASAP7_75t_L g1278 ( 
.A1(n_1005),
.A2(n_578),
.B(n_572),
.C(n_43),
.Y(n_1278)
);

AOI21xp5_ASAP7_75t_L g1279 ( 
.A1(n_1058),
.A2(n_100),
.B(n_211),
.Y(n_1279)
);

INVx2_ASAP7_75t_L g1280 ( 
.A(n_1086),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1124),
.Y(n_1281)
);

NOR3xp33_ASAP7_75t_SL g1282 ( 
.A(n_1071),
.B(n_41),
.C(n_42),
.Y(n_1282)
);

INVx2_ASAP7_75t_L g1283 ( 
.A(n_1086),
.Y(n_1283)
);

CKINVDCx5p33_ASAP7_75t_R g1284 ( 
.A(n_1097),
.Y(n_1284)
);

OR2x6_ASAP7_75t_L g1285 ( 
.A(n_947),
.B(n_42),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_958),
.B(n_578),
.Y(n_1286)
);

CKINVDCx8_ASAP7_75t_R g1287 ( 
.A(n_1025),
.Y(n_1287)
);

INVx3_ASAP7_75t_L g1288 ( 
.A(n_1287),
.Y(n_1288)
);

O2A1O1Ixp5_ASAP7_75t_L g1289 ( 
.A1(n_1245),
.A2(n_1090),
.B(n_955),
.C(n_999),
.Y(n_1289)
);

INVx1_ASAP7_75t_SL g1290 ( 
.A(n_1139),
.Y(n_1290)
);

INVx1_ASAP7_75t_SL g1291 ( 
.A(n_1248),
.Y(n_1291)
);

BUFx6f_ASAP7_75t_L g1292 ( 
.A(n_1168),
.Y(n_1292)
);

AND2x2_ASAP7_75t_L g1293 ( 
.A(n_1234),
.B(n_1112),
.Y(n_1293)
);

A2O1A1Ixp33_ASAP7_75t_L g1294 ( 
.A1(n_1195),
.A2(n_1064),
.B(n_991),
.C(n_1095),
.Y(n_1294)
);

NOR2xp33_ASAP7_75t_L g1295 ( 
.A(n_1284),
.B(n_1083),
.Y(n_1295)
);

AND2x2_ASAP7_75t_L g1296 ( 
.A(n_1160),
.B(n_1117),
.Y(n_1296)
);

INVx3_ASAP7_75t_L g1297 ( 
.A(n_1233),
.Y(n_1297)
);

AOI21xp5_ASAP7_75t_L g1298 ( 
.A1(n_1165),
.A2(n_996),
.B(n_1032),
.Y(n_1298)
);

BUFx3_ASAP7_75t_L g1299 ( 
.A(n_1178),
.Y(n_1299)
);

NAND3x1_ASAP7_75t_L g1300 ( 
.A(n_1128),
.B(n_989),
.C(n_1053),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_L g1301 ( 
.A(n_1133),
.B(n_1025),
.Y(n_1301)
);

AOI21xp5_ASAP7_75t_L g1302 ( 
.A1(n_1165),
.A2(n_1213),
.B(n_1129),
.Y(n_1302)
);

OAI21x1_ASAP7_75t_L g1303 ( 
.A1(n_1152),
.A2(n_1056),
.B(n_1052),
.Y(n_1303)
);

O2A1O1Ixp33_ASAP7_75t_L g1304 ( 
.A1(n_1180),
.A2(n_981),
.B(n_1055),
.C(n_971),
.Y(n_1304)
);

OR2x2_ASAP7_75t_L g1305 ( 
.A(n_1220),
.B(n_993),
.Y(n_1305)
);

O2A1O1Ixp33_ASAP7_75t_SL g1306 ( 
.A1(n_1129),
.A2(n_1004),
.B(n_1018),
.C(n_983),
.Y(n_1306)
);

INVx2_ASAP7_75t_L g1307 ( 
.A(n_1135),
.Y(n_1307)
);

AO31x2_ASAP7_75t_L g1308 ( 
.A1(n_1280),
.A2(n_1000),
.A3(n_1034),
.B(n_1039),
.Y(n_1308)
);

OAI21x1_ASAP7_75t_L g1309 ( 
.A1(n_1179),
.A2(n_1056),
.B(n_1052),
.Y(n_1309)
);

AO32x2_ASAP7_75t_L g1310 ( 
.A1(n_1213),
.A2(n_1020),
.A3(n_966),
.B1(n_1030),
.B2(n_1021),
.Y(n_1310)
);

AOI21xp5_ASAP7_75t_L g1311 ( 
.A1(n_1150),
.A2(n_975),
.B(n_977),
.Y(n_1311)
);

AO31x2_ASAP7_75t_L g1312 ( 
.A1(n_1143),
.A2(n_1126),
.A3(n_997),
.B(n_948),
.Y(n_1312)
);

O2A1O1Ixp33_ASAP7_75t_L g1313 ( 
.A1(n_1170),
.A2(n_979),
.B(n_984),
.C(n_1033),
.Y(n_1313)
);

INVx2_ASAP7_75t_L g1314 ( 
.A(n_1162),
.Y(n_1314)
);

CKINVDCx5p33_ASAP7_75t_R g1315 ( 
.A(n_1130),
.Y(n_1315)
);

AO21x2_ASAP7_75t_L g1316 ( 
.A1(n_1179),
.A2(n_997),
.B(n_1054),
.Y(n_1316)
);

BUFx6f_ASAP7_75t_L g1317 ( 
.A(n_1166),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_L g1318 ( 
.A(n_1273),
.B(n_1038),
.Y(n_1318)
);

AOI21xp5_ASAP7_75t_L g1319 ( 
.A1(n_1136),
.A2(n_941),
.B(n_948),
.Y(n_1319)
);

AOI21x1_ASAP7_75t_L g1320 ( 
.A1(n_1270),
.A2(n_1077),
.B(n_941),
.Y(n_1320)
);

NAND2xp5_ASAP7_75t_L g1321 ( 
.A(n_1281),
.B(n_1025),
.Y(n_1321)
);

OAI21xp5_ASAP7_75t_L g1322 ( 
.A1(n_1131),
.A2(n_1077),
.B(n_987),
.Y(n_1322)
);

OAI21xp5_ASAP7_75t_L g1323 ( 
.A1(n_1154),
.A2(n_987),
.B(n_970),
.Y(n_1323)
);

NOR2xp67_ASAP7_75t_L g1324 ( 
.A(n_1233),
.B(n_1260),
.Y(n_1324)
);

OR2x6_ASAP7_75t_L g1325 ( 
.A(n_1196),
.B(n_1038),
.Y(n_1325)
);

AOI21xp5_ASAP7_75t_L g1326 ( 
.A1(n_1140),
.A2(n_970),
.B(n_1120),
.Y(n_1326)
);

BUFx6f_ASAP7_75t_L g1327 ( 
.A(n_1166),
.Y(n_1327)
);

CKINVDCx5p33_ASAP7_75t_R g1328 ( 
.A(n_1153),
.Y(n_1328)
);

NOR2x1_ASAP7_75t_SL g1329 ( 
.A(n_1156),
.B(n_1038),
.Y(n_1329)
);

OAI21xp5_ASAP7_75t_L g1330 ( 
.A1(n_1263),
.A2(n_1266),
.B(n_1138),
.Y(n_1330)
);

BUFx2_ASAP7_75t_L g1331 ( 
.A(n_1188),
.Y(n_1331)
);

BUFx6f_ASAP7_75t_L g1332 ( 
.A(n_1166),
.Y(n_1332)
);

OAI21xp5_ASAP7_75t_L g1333 ( 
.A1(n_1181),
.A2(n_1118),
.B(n_1111),
.Y(n_1333)
);

AOI21xp5_ASAP7_75t_L g1334 ( 
.A1(n_1169),
.A2(n_1118),
.B(n_1111),
.Y(n_1334)
);

AOI21xp5_ASAP7_75t_L g1335 ( 
.A1(n_1169),
.A2(n_1106),
.B(n_1098),
.Y(n_1335)
);

OAI21x1_ASAP7_75t_L g1336 ( 
.A1(n_1149),
.A2(n_1106),
.B(n_1098),
.Y(n_1336)
);

AOI21xp5_ASAP7_75t_L g1337 ( 
.A1(n_1167),
.A2(n_1096),
.B(n_989),
.Y(n_1337)
);

CKINVDCx5p33_ASAP7_75t_R g1338 ( 
.A(n_1202),
.Y(n_1338)
);

OAI21xp5_ASAP7_75t_L g1339 ( 
.A1(n_1256),
.A2(n_1096),
.B(n_578),
.Y(n_1339)
);

OAI21xp5_ASAP7_75t_L g1340 ( 
.A1(n_1256),
.A2(n_1269),
.B(n_1148),
.Y(n_1340)
);

AND2x2_ASAP7_75t_L g1341 ( 
.A(n_1186),
.B(n_1155),
.Y(n_1341)
);

NAND2xp5_ASAP7_75t_L g1342 ( 
.A(n_1146),
.B(n_1244),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_SL g1343 ( 
.A(n_1274),
.B(n_1094),
.Y(n_1343)
);

A2O1A1Ixp33_ASAP7_75t_L g1344 ( 
.A1(n_1218),
.A2(n_1094),
.B(n_48),
.C(n_50),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_L g1345 ( 
.A(n_1240),
.B(n_47),
.Y(n_1345)
);

AO31x2_ASAP7_75t_L g1346 ( 
.A1(n_1257),
.A2(n_578),
.A3(n_572),
.B(n_103),
.Y(n_1346)
);

OR2x2_ASAP7_75t_L g1347 ( 
.A(n_1145),
.B(n_48),
.Y(n_1347)
);

AOI22xp5_ASAP7_75t_L g1348 ( 
.A1(n_1184),
.A2(n_578),
.B1(n_572),
.B2(n_60),
.Y(n_1348)
);

NAND2xp5_ASAP7_75t_L g1349 ( 
.A(n_1210),
.B(n_54),
.Y(n_1349)
);

OAI21x1_ASAP7_75t_L g1350 ( 
.A1(n_1272),
.A2(n_107),
.B(n_210),
.Y(n_1350)
);

AOI21xp5_ASAP7_75t_L g1351 ( 
.A1(n_1167),
.A2(n_101),
.B(n_204),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1132),
.Y(n_1352)
);

AO31x2_ASAP7_75t_L g1353 ( 
.A1(n_1161),
.A2(n_578),
.A3(n_572),
.B(n_98),
.Y(n_1353)
);

HB1xp67_ASAP7_75t_L g1354 ( 
.A(n_1253),
.Y(n_1354)
);

OR2x2_ASAP7_75t_L g1355 ( 
.A(n_1141),
.B(n_54),
.Y(n_1355)
);

AOI21xp5_ASAP7_75t_L g1356 ( 
.A1(n_1159),
.A2(n_93),
.B(n_179),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_L g1357 ( 
.A(n_1215),
.B(n_58),
.Y(n_1357)
);

A2O1A1Ixp33_ASAP7_75t_L g1358 ( 
.A1(n_1271),
.A2(n_62),
.B(n_63),
.C(n_65),
.Y(n_1358)
);

AO31x2_ASAP7_75t_L g1359 ( 
.A1(n_1246),
.A2(n_123),
.A3(n_175),
.B(n_173),
.Y(n_1359)
);

AOI21xp5_ASAP7_75t_L g1360 ( 
.A1(n_1159),
.A2(n_115),
.B(n_160),
.Y(n_1360)
);

OR2x6_ASAP7_75t_L g1361 ( 
.A(n_1196),
.B(n_70),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1144),
.Y(n_1362)
);

AOI31xp67_ASAP7_75t_L g1363 ( 
.A1(n_1267),
.A2(n_88),
.A3(n_151),
.B(n_149),
.Y(n_1363)
);

OAI21x1_ASAP7_75t_L g1364 ( 
.A1(n_1279),
.A2(n_1261),
.B(n_1192),
.Y(n_1364)
);

AOI21xp5_ASAP7_75t_L g1365 ( 
.A1(n_1242),
.A2(n_86),
.B(n_146),
.Y(n_1365)
);

BUFx2_ASAP7_75t_R g1366 ( 
.A(n_1147),
.Y(n_1366)
);

BUFx2_ASAP7_75t_L g1367 ( 
.A(n_1208),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1173),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1185),
.Y(n_1369)
);

O2A1O1Ixp33_ASAP7_75t_SL g1370 ( 
.A1(n_1214),
.A2(n_72),
.B(n_75),
.C(n_76),
.Y(n_1370)
);

AND2x2_ASAP7_75t_L g1371 ( 
.A(n_1164),
.B(n_77),
.Y(n_1371)
);

OA22x2_ASAP7_75t_L g1372 ( 
.A1(n_1134),
.A2(n_80),
.B1(n_125),
.B2(n_140),
.Y(n_1372)
);

O2A1O1Ixp33_ASAP7_75t_SL g1373 ( 
.A1(n_1217),
.A2(n_200),
.B(n_1194),
.C(n_1175),
.Y(n_1373)
);

INVxp67_ASAP7_75t_SL g1374 ( 
.A(n_1238),
.Y(n_1374)
);

INVx2_ASAP7_75t_L g1375 ( 
.A(n_1221),
.Y(n_1375)
);

A2O1A1Ixp33_ASAP7_75t_L g1376 ( 
.A1(n_1183),
.A2(n_1241),
.B(n_1193),
.C(n_1176),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1189),
.Y(n_1377)
);

A2O1A1Ixp33_ASAP7_75t_L g1378 ( 
.A1(n_1282),
.A2(n_1219),
.B(n_1157),
.C(n_1177),
.Y(n_1378)
);

OAI21x1_ASAP7_75t_L g1379 ( 
.A1(n_1192),
.A2(n_1242),
.B(n_1223),
.Y(n_1379)
);

INVx4_ASAP7_75t_L g1380 ( 
.A(n_1209),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_L g1381 ( 
.A(n_1238),
.B(n_1208),
.Y(n_1381)
);

HB1xp67_ASAP7_75t_L g1382 ( 
.A(n_1249),
.Y(n_1382)
);

NOR2xp33_ASAP7_75t_SL g1383 ( 
.A(n_1196),
.B(n_1254),
.Y(n_1383)
);

AOI21xp5_ASAP7_75t_L g1384 ( 
.A1(n_1163),
.A2(n_1269),
.B(n_1258),
.Y(n_1384)
);

AO31x2_ASAP7_75t_L g1385 ( 
.A1(n_1224),
.A2(n_1227),
.A3(n_1229),
.B(n_1207),
.Y(n_1385)
);

NOR2xp67_ASAP7_75t_L g1386 ( 
.A(n_1260),
.B(n_1265),
.Y(n_1386)
);

INVxp67_ASAP7_75t_L g1387 ( 
.A(n_1200),
.Y(n_1387)
);

OAI21xp5_ASAP7_75t_L g1388 ( 
.A1(n_1223),
.A2(n_1158),
.B(n_1286),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_L g1389 ( 
.A(n_1174),
.B(n_1211),
.Y(n_1389)
);

AO32x2_ASAP7_75t_L g1390 ( 
.A1(n_1206),
.A2(n_1203),
.A3(n_1199),
.B1(n_1236),
.B2(n_1182),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_1174),
.B(n_1142),
.Y(n_1391)
);

OAI21x1_ASAP7_75t_L g1392 ( 
.A1(n_1207),
.A2(n_1229),
.B(n_1239),
.Y(n_1392)
);

NOR2xp33_ASAP7_75t_L g1393 ( 
.A(n_1191),
.B(n_1182),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_L g1394 ( 
.A(n_1142),
.B(n_1216),
.Y(n_1394)
);

NOR2xp67_ASAP7_75t_SL g1395 ( 
.A(n_1265),
.B(n_1268),
.Y(n_1395)
);

OAI21x1_ASAP7_75t_L g1396 ( 
.A1(n_1237),
.A2(n_1259),
.B(n_1251),
.Y(n_1396)
);

OAI21xp5_ASAP7_75t_L g1397 ( 
.A1(n_1286),
.A2(n_1230),
.B(n_1228),
.Y(n_1397)
);

INVx6_ASAP7_75t_L g1398 ( 
.A(n_1226),
.Y(n_1398)
);

AOI22xp5_ASAP7_75t_L g1399 ( 
.A1(n_1247),
.A2(n_1199),
.B1(n_1190),
.B2(n_1236),
.Y(n_1399)
);

AOI21xp5_ASAP7_75t_L g1400 ( 
.A1(n_1258),
.A2(n_1172),
.B(n_1231),
.Y(n_1400)
);

OAI21x1_ASAP7_75t_L g1401 ( 
.A1(n_1264),
.A2(n_1197),
.B(n_1201),
.Y(n_1401)
);

OAI21x1_ASAP7_75t_L g1402 ( 
.A1(n_1204),
.A2(n_1232),
.B(n_1222),
.Y(n_1402)
);

AOI21xp5_ASAP7_75t_L g1403 ( 
.A1(n_1172),
.A2(n_1205),
.B(n_1235),
.Y(n_1403)
);

AOI22xp33_ASAP7_75t_L g1404 ( 
.A1(n_1203),
.A2(n_1285),
.B1(n_1252),
.B2(n_1250),
.Y(n_1404)
);

INVxp67_ASAP7_75t_L g1405 ( 
.A(n_1226),
.Y(n_1405)
);

O2A1O1Ixp33_ASAP7_75t_SL g1406 ( 
.A1(n_1278),
.A2(n_1212),
.B(n_1206),
.C(n_1225),
.Y(n_1406)
);

AOI21x1_ASAP7_75t_L g1407 ( 
.A1(n_1235),
.A2(n_1205),
.B(n_1172),
.Y(n_1407)
);

INVx2_ASAP7_75t_SL g1408 ( 
.A(n_1255),
.Y(n_1408)
);

OAI21x1_ASAP7_75t_L g1409 ( 
.A1(n_1187),
.A2(n_1151),
.B(n_1275),
.Y(n_1409)
);

NAND2xp5_ASAP7_75t_L g1410 ( 
.A(n_1277),
.B(n_1285),
.Y(n_1410)
);

BUFx2_ASAP7_75t_L g1411 ( 
.A(n_1137),
.Y(n_1411)
);

AOI221xp5_ASAP7_75t_SL g1412 ( 
.A1(n_1206),
.A2(n_1243),
.B1(n_1276),
.B2(n_1265),
.C(n_1285),
.Y(n_1412)
);

OAI21xp5_ASAP7_75t_L g1413 ( 
.A1(n_1205),
.A2(n_1262),
.B(n_1235),
.Y(n_1413)
);

INVx2_ASAP7_75t_L g1414 ( 
.A(n_1255),
.Y(n_1414)
);

AOI21xp5_ASAP7_75t_L g1415 ( 
.A1(n_1262),
.A2(n_1171),
.B(n_1198),
.Y(n_1415)
);

AOI21xp5_ASAP7_75t_L g1416 ( 
.A1(n_1171),
.A2(n_968),
.B(n_954),
.Y(n_1416)
);

NAND2xp5_ASAP7_75t_L g1417 ( 
.A(n_1198),
.B(n_624),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1132),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1132),
.Y(n_1419)
);

AO32x2_ASAP7_75t_L g1420 ( 
.A1(n_1213),
.A2(n_1274),
.A3(n_610),
.B1(n_623),
.B2(n_962),
.Y(n_1420)
);

INVx2_ASAP7_75t_SL g1421 ( 
.A(n_1202),
.Y(n_1421)
);

AOI21xp5_ASAP7_75t_L g1422 ( 
.A1(n_1165),
.A2(n_968),
.B(n_954),
.Y(n_1422)
);

NOR2xp33_ASAP7_75t_L g1423 ( 
.A(n_1234),
.B(n_624),
.Y(n_1423)
);

OR2x2_ASAP7_75t_L g1424 ( 
.A(n_1234),
.B(n_1139),
.Y(n_1424)
);

AOI21xp5_ASAP7_75t_L g1425 ( 
.A1(n_1165),
.A2(n_968),
.B(n_954),
.Y(n_1425)
);

OAI21x1_ASAP7_75t_L g1426 ( 
.A1(n_1152),
.A2(n_1179),
.B(n_1270),
.Y(n_1426)
);

OAI21x1_ASAP7_75t_L g1427 ( 
.A1(n_1152),
.A2(n_1179),
.B(n_1270),
.Y(n_1427)
);

A2O1A1Ixp33_ASAP7_75t_L g1428 ( 
.A1(n_1245),
.A2(n_624),
.B(n_957),
.C(n_1195),
.Y(n_1428)
);

AOI22xp33_ASAP7_75t_SL g1429 ( 
.A1(n_1134),
.A2(n_715),
.B1(n_427),
.B2(n_439),
.Y(n_1429)
);

NAND3xp33_ASAP7_75t_L g1430 ( 
.A(n_1245),
.B(n_624),
.C(n_1282),
.Y(n_1430)
);

NAND2xp5_ASAP7_75t_L g1431 ( 
.A(n_1234),
.B(n_624),
.Y(n_1431)
);

BUFx6f_ASAP7_75t_L g1432 ( 
.A(n_1168),
.Y(n_1432)
);

AOI21xp5_ASAP7_75t_L g1433 ( 
.A1(n_1165),
.A2(n_968),
.B(n_954),
.Y(n_1433)
);

OAI21x1_ASAP7_75t_L g1434 ( 
.A1(n_1152),
.A2(n_1179),
.B(n_1270),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_L g1435 ( 
.A(n_1234),
.B(n_624),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1132),
.Y(n_1436)
);

AND2x2_ASAP7_75t_L g1437 ( 
.A(n_1234),
.B(n_819),
.Y(n_1437)
);

NAND2x1p5_ASAP7_75t_L g1438 ( 
.A(n_1151),
.B(n_1049),
.Y(n_1438)
);

INVx6_ASAP7_75t_L g1439 ( 
.A(n_1208),
.Y(n_1439)
);

OAI21xp5_ASAP7_75t_L g1440 ( 
.A1(n_1213),
.A2(n_1109),
.B(n_1131),
.Y(n_1440)
);

AO21x1_ASAP7_75t_L g1441 ( 
.A1(n_1245),
.A2(n_957),
.B(n_1213),
.Y(n_1441)
);

INVx1_ASAP7_75t_SL g1442 ( 
.A(n_1139),
.Y(n_1442)
);

BUFx3_ASAP7_75t_L g1443 ( 
.A(n_1168),
.Y(n_1443)
);

BUFx12f_ASAP7_75t_L g1444 ( 
.A(n_1208),
.Y(n_1444)
);

AOI221x1_ASAP7_75t_L g1445 ( 
.A1(n_1247),
.A2(n_1245),
.B1(n_1143),
.B2(n_1274),
.C(n_624),
.Y(n_1445)
);

O2A1O1Ixp33_ASAP7_75t_L g1446 ( 
.A1(n_1245),
.A2(n_624),
.B(n_623),
.C(n_957),
.Y(n_1446)
);

A2O1A1Ixp33_ASAP7_75t_L g1447 ( 
.A1(n_1245),
.A2(n_624),
.B(n_957),
.C(n_1195),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_L g1448 ( 
.A(n_1234),
.B(n_624),
.Y(n_1448)
);

OAI21x1_ASAP7_75t_L g1449 ( 
.A1(n_1152),
.A2(n_1179),
.B(n_1270),
.Y(n_1449)
);

INVx2_ASAP7_75t_SL g1450 ( 
.A(n_1202),
.Y(n_1450)
);

OAI22xp5_ASAP7_75t_L g1451 ( 
.A1(n_1245),
.A2(n_957),
.B1(n_988),
.B2(n_1072),
.Y(n_1451)
);

INVx2_ASAP7_75t_L g1452 ( 
.A(n_1135),
.Y(n_1452)
);

AO31x2_ASAP7_75t_L g1453 ( 
.A1(n_1280),
.A2(n_1008),
.A3(n_1283),
.B(n_1143),
.Y(n_1453)
);

AOI21xp5_ASAP7_75t_L g1454 ( 
.A1(n_1165),
.A2(n_968),
.B(n_954),
.Y(n_1454)
);

OAI22xp5_ASAP7_75t_L g1455 ( 
.A1(n_1245),
.A2(n_957),
.B1(n_624),
.B2(n_967),
.Y(n_1455)
);

AOI21xp5_ASAP7_75t_L g1456 ( 
.A1(n_1165),
.A2(n_968),
.B(n_954),
.Y(n_1456)
);

NOR2xp67_ASAP7_75t_SL g1457 ( 
.A(n_1284),
.B(n_668),
.Y(n_1457)
);

AOI221x1_ASAP7_75t_L g1458 ( 
.A1(n_1247),
.A2(n_1245),
.B1(n_1143),
.B2(n_1274),
.C(n_624),
.Y(n_1458)
);

AO31x2_ASAP7_75t_L g1459 ( 
.A1(n_1280),
.A2(n_1008),
.A3(n_1283),
.B(n_1143),
.Y(n_1459)
);

A2O1A1Ixp33_ASAP7_75t_L g1460 ( 
.A1(n_1245),
.A2(n_624),
.B(n_957),
.C(n_1195),
.Y(n_1460)
);

AOI22xp5_ASAP7_75t_L g1461 ( 
.A1(n_1455),
.A2(n_1451),
.B1(n_1423),
.B2(n_1430),
.Y(n_1461)
);

AOI22xp33_ASAP7_75t_L g1462 ( 
.A1(n_1451),
.A2(n_1430),
.B1(n_1429),
.B2(n_1441),
.Y(n_1462)
);

OAI21xp5_ASAP7_75t_SL g1463 ( 
.A1(n_1446),
.A2(n_1447),
.B(n_1428),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1352),
.Y(n_1464)
);

BUFx2_ASAP7_75t_SL g1465 ( 
.A(n_1288),
.Y(n_1465)
);

INVx4_ASAP7_75t_L g1466 ( 
.A(n_1338),
.Y(n_1466)
);

CKINVDCx5p33_ASAP7_75t_R g1467 ( 
.A(n_1315),
.Y(n_1467)
);

AOI22xp33_ASAP7_75t_L g1468 ( 
.A1(n_1437),
.A2(n_1393),
.B1(n_1387),
.B2(n_1293),
.Y(n_1468)
);

INVx8_ASAP7_75t_L g1469 ( 
.A(n_1444),
.Y(n_1469)
);

INVxp67_ASAP7_75t_SL g1470 ( 
.A(n_1302),
.Y(n_1470)
);

CKINVDCx11_ASAP7_75t_R g1471 ( 
.A(n_1292),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1362),
.Y(n_1472)
);

AOI22xp33_ASAP7_75t_SL g1473 ( 
.A1(n_1420),
.A2(n_1372),
.B1(n_1440),
.B2(n_1296),
.Y(n_1473)
);

BUFx2_ASAP7_75t_L g1474 ( 
.A(n_1341),
.Y(n_1474)
);

INVx2_ASAP7_75t_L g1475 ( 
.A(n_1314),
.Y(n_1475)
);

INVx4_ASAP7_75t_L g1476 ( 
.A(n_1292),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1368),
.Y(n_1477)
);

BUFx8_ASAP7_75t_L g1478 ( 
.A(n_1367),
.Y(n_1478)
);

INVx4_ASAP7_75t_L g1479 ( 
.A(n_1292),
.Y(n_1479)
);

INVx4_ASAP7_75t_SL g1480 ( 
.A(n_1361),
.Y(n_1480)
);

OAI22xp33_ASAP7_75t_SL g1481 ( 
.A1(n_1394),
.A2(n_1389),
.B1(n_1361),
.B2(n_1342),
.Y(n_1481)
);

OAI22xp5_ASAP7_75t_L g1482 ( 
.A1(n_1460),
.A2(n_1399),
.B1(n_1376),
.B2(n_1417),
.Y(n_1482)
);

CKINVDCx11_ASAP7_75t_R g1483 ( 
.A(n_1432),
.Y(n_1483)
);

BUFx4_ASAP7_75t_SL g1484 ( 
.A(n_1328),
.Y(n_1484)
);

BUFx5_ASAP7_75t_L g1485 ( 
.A(n_1369),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1377),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1418),
.Y(n_1487)
);

AOI22xp33_ASAP7_75t_L g1488 ( 
.A1(n_1420),
.A2(n_1440),
.B1(n_1399),
.B2(n_1374),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1419),
.Y(n_1489)
);

OAI22xp33_ASAP7_75t_L g1490 ( 
.A1(n_1361),
.A2(n_1445),
.B1(n_1458),
.B2(n_1420),
.Y(n_1490)
);

BUFx12f_ASAP7_75t_L g1491 ( 
.A(n_1432),
.Y(n_1491)
);

OAI22xp33_ASAP7_75t_L g1492 ( 
.A1(n_1348),
.A2(n_1355),
.B1(n_1448),
.B2(n_1431),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_L g1493 ( 
.A(n_1290),
.B(n_1442),
.Y(n_1493)
);

INVx6_ASAP7_75t_L g1494 ( 
.A(n_1380),
.Y(n_1494)
);

AOI22xp33_ASAP7_75t_L g1495 ( 
.A1(n_1435),
.A2(n_1343),
.B1(n_1452),
.B2(n_1375),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1436),
.Y(n_1496)
);

AOI22xp33_ASAP7_75t_SL g1497 ( 
.A1(n_1366),
.A2(n_1345),
.B1(n_1357),
.B2(n_1439),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_L g1498 ( 
.A(n_1290),
.B(n_1442),
.Y(n_1498)
);

AOI22xp33_ASAP7_75t_L g1499 ( 
.A1(n_1391),
.A2(n_1305),
.B1(n_1457),
.B2(n_1404),
.Y(n_1499)
);

AOI22xp5_ASAP7_75t_L g1500 ( 
.A1(n_1381),
.A2(n_1439),
.B1(n_1410),
.B2(n_1383),
.Y(n_1500)
);

INVxp67_ASAP7_75t_SL g1501 ( 
.A(n_1330),
.Y(n_1501)
);

BUFx6f_ASAP7_75t_L g1502 ( 
.A(n_1325),
.Y(n_1502)
);

AOI22xp33_ASAP7_75t_L g1503 ( 
.A1(n_1348),
.A2(n_1424),
.B1(n_1349),
.B2(n_1371),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1385),
.Y(n_1504)
);

OAI21xp33_ASAP7_75t_L g1505 ( 
.A1(n_1358),
.A2(n_1344),
.B(n_1378),
.Y(n_1505)
);

INVxp67_ASAP7_75t_L g1506 ( 
.A(n_1301),
.Y(n_1506)
);

BUFx8_ASAP7_75t_SL g1507 ( 
.A(n_1331),
.Y(n_1507)
);

INVx2_ASAP7_75t_SL g1508 ( 
.A(n_1299),
.Y(n_1508)
);

CKINVDCx11_ASAP7_75t_R g1509 ( 
.A(n_1443),
.Y(n_1509)
);

INVx2_ASAP7_75t_L g1510 ( 
.A(n_1318),
.Y(n_1510)
);

AOI22xp33_ASAP7_75t_L g1511 ( 
.A1(n_1347),
.A2(n_1321),
.B1(n_1382),
.B2(n_1291),
.Y(n_1511)
);

AOI22xp33_ASAP7_75t_SL g1512 ( 
.A1(n_1390),
.A2(n_1383),
.B1(n_1412),
.B2(n_1388),
.Y(n_1512)
);

NAND2x1p5_ASAP7_75t_L g1513 ( 
.A(n_1395),
.B(n_1288),
.Y(n_1513)
);

INVx6_ASAP7_75t_L g1514 ( 
.A(n_1380),
.Y(n_1514)
);

OAI21xp5_ASAP7_75t_L g1515 ( 
.A1(n_1294),
.A2(n_1289),
.B(n_1456),
.Y(n_1515)
);

OAI21xp33_ASAP7_75t_L g1516 ( 
.A1(n_1330),
.A2(n_1322),
.B(n_1304),
.Y(n_1516)
);

INVx1_ASAP7_75t_SL g1517 ( 
.A(n_1354),
.Y(n_1517)
);

BUFx3_ASAP7_75t_L g1518 ( 
.A(n_1421),
.Y(n_1518)
);

AOI22xp33_ASAP7_75t_L g1519 ( 
.A1(n_1291),
.A2(n_1388),
.B1(n_1298),
.B2(n_1397),
.Y(n_1519)
);

INVx3_ASAP7_75t_L g1520 ( 
.A(n_1325),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1385),
.Y(n_1521)
);

AOI22xp33_ASAP7_75t_SL g1522 ( 
.A1(n_1390),
.A2(n_1412),
.B1(n_1413),
.B2(n_1322),
.Y(n_1522)
);

AOI22xp33_ASAP7_75t_SL g1523 ( 
.A1(n_1390),
.A2(n_1413),
.B1(n_1411),
.B2(n_1397),
.Y(n_1523)
);

AOI22xp33_ASAP7_75t_L g1524 ( 
.A1(n_1450),
.A2(n_1295),
.B1(n_1415),
.B2(n_1340),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1317),
.Y(n_1525)
);

CKINVDCx20_ASAP7_75t_R g1526 ( 
.A(n_1408),
.Y(n_1526)
);

OAI22xp5_ASAP7_75t_L g1527 ( 
.A1(n_1422),
.A2(n_1433),
.B1(n_1425),
.B2(n_1454),
.Y(n_1527)
);

OAI21xp5_ASAP7_75t_SL g1528 ( 
.A1(n_1351),
.A2(n_1365),
.B(n_1438),
.Y(n_1528)
);

AOI22xp33_ASAP7_75t_L g1529 ( 
.A1(n_1340),
.A2(n_1414),
.B1(n_1402),
.B2(n_1409),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1317),
.Y(n_1530)
);

BUFx12f_ASAP7_75t_L g1531 ( 
.A(n_1327),
.Y(n_1531)
);

AOI21xp5_ASAP7_75t_L g1532 ( 
.A1(n_1416),
.A2(n_1311),
.B(n_1306),
.Y(n_1532)
);

AOI22xp33_ASAP7_75t_L g1533 ( 
.A1(n_1333),
.A2(n_1316),
.B1(n_1323),
.B2(n_1339),
.Y(n_1533)
);

OAI22xp5_ASAP7_75t_L g1534 ( 
.A1(n_1300),
.A2(n_1403),
.B1(n_1297),
.B2(n_1407),
.Y(n_1534)
);

AOI22xp33_ASAP7_75t_L g1535 ( 
.A1(n_1333),
.A2(n_1316),
.B1(n_1323),
.B2(n_1339),
.Y(n_1535)
);

AND2x2_ASAP7_75t_L g1536 ( 
.A(n_1405),
.B(n_1398),
.Y(n_1536)
);

AOI22xp33_ASAP7_75t_L g1537 ( 
.A1(n_1398),
.A2(n_1386),
.B1(n_1379),
.B2(n_1360),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1332),
.Y(n_1538)
);

INVxp67_ASAP7_75t_SL g1539 ( 
.A(n_1309),
.Y(n_1539)
);

AOI22xp33_ASAP7_75t_L g1540 ( 
.A1(n_1386),
.A2(n_1356),
.B1(n_1400),
.B2(n_1332),
.Y(n_1540)
);

AOI22xp33_ASAP7_75t_L g1541 ( 
.A1(n_1332),
.A2(n_1401),
.B1(n_1319),
.B2(n_1324),
.Y(n_1541)
);

OAI22xp33_ASAP7_75t_L g1542 ( 
.A1(n_1297),
.A2(n_1324),
.B1(n_1337),
.B2(n_1406),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_L g1543 ( 
.A(n_1329),
.B(n_1370),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1453),
.Y(n_1544)
);

AOI22xp33_ASAP7_75t_L g1545 ( 
.A1(n_1384),
.A2(n_1350),
.B1(n_1335),
.B2(n_1334),
.Y(n_1545)
);

OAI22xp33_ASAP7_75t_L g1546 ( 
.A1(n_1326),
.A2(n_1320),
.B1(n_1346),
.B2(n_1363),
.Y(n_1546)
);

NAND2xp5_ASAP7_75t_L g1547 ( 
.A(n_1459),
.B(n_1346),
.Y(n_1547)
);

OAI22xp5_ASAP7_75t_L g1548 ( 
.A1(n_1313),
.A2(n_1373),
.B1(n_1310),
.B2(n_1346),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1459),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_L g1550 ( 
.A(n_1459),
.B(n_1359),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_L g1551 ( 
.A(n_1359),
.B(n_1308),
.Y(n_1551)
);

AOI22xp33_ASAP7_75t_L g1552 ( 
.A1(n_1392),
.A2(n_1396),
.B1(n_1364),
.B2(n_1336),
.Y(n_1552)
);

BUFx2_ASAP7_75t_L g1553 ( 
.A(n_1312),
.Y(n_1553)
);

AOI22xp33_ASAP7_75t_L g1554 ( 
.A1(n_1426),
.A2(n_1449),
.B1(n_1434),
.B2(n_1427),
.Y(n_1554)
);

CKINVDCx11_ASAP7_75t_R g1555 ( 
.A(n_1310),
.Y(n_1555)
);

INVx4_ASAP7_75t_L g1556 ( 
.A(n_1310),
.Y(n_1556)
);

INVx1_ASAP7_75t_SL g1557 ( 
.A(n_1303),
.Y(n_1557)
);

INVx4_ASAP7_75t_SL g1558 ( 
.A(n_1312),
.Y(n_1558)
);

AOI22xp33_ASAP7_75t_SL g1559 ( 
.A1(n_1353),
.A2(n_1451),
.B1(n_715),
.B2(n_1072),
.Y(n_1559)
);

BUFx3_ASAP7_75t_L g1560 ( 
.A(n_1312),
.Y(n_1560)
);

AOI22xp33_ASAP7_75t_SL g1561 ( 
.A1(n_1353),
.A2(n_1451),
.B1(n_715),
.B2(n_1072),
.Y(n_1561)
);

INVx2_ASAP7_75t_L g1562 ( 
.A(n_1353),
.Y(n_1562)
);

AOI22xp33_ASAP7_75t_L g1563 ( 
.A1(n_1451),
.A2(n_1455),
.B1(n_715),
.B2(n_1072),
.Y(n_1563)
);

AND2x2_ASAP7_75t_L g1564 ( 
.A(n_1293),
.B(n_1437),
.Y(n_1564)
);

AOI22xp5_ASAP7_75t_L g1565 ( 
.A1(n_1455),
.A2(n_624),
.B1(n_1451),
.B2(n_1423),
.Y(n_1565)
);

BUFx2_ASAP7_75t_L g1566 ( 
.A(n_1341),
.Y(n_1566)
);

BUFx10_ASAP7_75t_L g1567 ( 
.A(n_1315),
.Y(n_1567)
);

OAI22xp5_ASAP7_75t_SL g1568 ( 
.A1(n_1423),
.A2(n_1153),
.B1(n_620),
.B2(n_687),
.Y(n_1568)
);

BUFx2_ASAP7_75t_L g1569 ( 
.A(n_1341),
.Y(n_1569)
);

OAI21xp33_ASAP7_75t_L g1570 ( 
.A1(n_1428),
.A2(n_624),
.B(n_1447),
.Y(n_1570)
);

OAI22xp33_ASAP7_75t_L g1571 ( 
.A1(n_1451),
.A2(n_1455),
.B1(n_957),
.B2(n_1430),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1352),
.Y(n_1572)
);

INVx6_ASAP7_75t_L g1573 ( 
.A(n_1292),
.Y(n_1573)
);

BUFx6f_ASAP7_75t_L g1574 ( 
.A(n_1325),
.Y(n_1574)
);

INVx6_ASAP7_75t_L g1575 ( 
.A(n_1292),
.Y(n_1575)
);

INVx4_ASAP7_75t_SL g1576 ( 
.A(n_1361),
.Y(n_1576)
);

CKINVDCx5p33_ASAP7_75t_R g1577 ( 
.A(n_1315),
.Y(n_1577)
);

INVx4_ASAP7_75t_L g1578 ( 
.A(n_1338),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1352),
.Y(n_1579)
);

NAND2x1p5_ASAP7_75t_L g1580 ( 
.A(n_1395),
.B(n_1049),
.Y(n_1580)
);

AOI22xp33_ASAP7_75t_SL g1581 ( 
.A1(n_1451),
.A2(n_715),
.B1(n_1072),
.B2(n_610),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1374),
.B(n_1455),
.Y(n_1582)
);

INVx2_ASAP7_75t_L g1583 ( 
.A(n_1307),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1352),
.Y(n_1584)
);

CKINVDCx20_ASAP7_75t_R g1585 ( 
.A(n_1315),
.Y(n_1585)
);

AOI22xp33_ASAP7_75t_L g1586 ( 
.A1(n_1451),
.A2(n_1455),
.B1(n_715),
.B2(n_1072),
.Y(n_1586)
);

BUFx2_ASAP7_75t_R g1587 ( 
.A(n_1338),
.Y(n_1587)
);

AOI22xp33_ASAP7_75t_L g1588 ( 
.A1(n_1451),
.A2(n_1455),
.B1(n_715),
.B2(n_1072),
.Y(n_1588)
);

INVx2_ASAP7_75t_L g1589 ( 
.A(n_1307),
.Y(n_1589)
);

CKINVDCx6p67_ASAP7_75t_R g1590 ( 
.A(n_1444),
.Y(n_1590)
);

BUFx2_ASAP7_75t_L g1591 ( 
.A(n_1341),
.Y(n_1591)
);

INVx2_ASAP7_75t_L g1592 ( 
.A(n_1307),
.Y(n_1592)
);

BUFx2_ASAP7_75t_L g1593 ( 
.A(n_1341),
.Y(n_1593)
);

BUFx8_ASAP7_75t_L g1594 ( 
.A(n_1444),
.Y(n_1594)
);

CKINVDCx20_ASAP7_75t_R g1595 ( 
.A(n_1315),
.Y(n_1595)
);

BUFx12f_ASAP7_75t_L g1596 ( 
.A(n_1315),
.Y(n_1596)
);

INVx1_ASAP7_75t_SL g1597 ( 
.A(n_1331),
.Y(n_1597)
);

CKINVDCx11_ASAP7_75t_R g1598 ( 
.A(n_1444),
.Y(n_1598)
);

HB1xp67_ASAP7_75t_L g1599 ( 
.A(n_1453),
.Y(n_1599)
);

INVx5_ASAP7_75t_L g1600 ( 
.A(n_1361),
.Y(n_1600)
);

AOI22xp33_ASAP7_75t_L g1601 ( 
.A1(n_1451),
.A2(n_1455),
.B1(n_715),
.B2(n_1072),
.Y(n_1601)
);

INVx6_ASAP7_75t_L g1602 ( 
.A(n_1292),
.Y(n_1602)
);

BUFx3_ASAP7_75t_L g1603 ( 
.A(n_1338),
.Y(n_1603)
);

CKINVDCx11_ASAP7_75t_R g1604 ( 
.A(n_1444),
.Y(n_1604)
);

INVx4_ASAP7_75t_L g1605 ( 
.A(n_1338),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1352),
.Y(n_1606)
);

CKINVDCx5p33_ASAP7_75t_R g1607 ( 
.A(n_1315),
.Y(n_1607)
);

AOI22xp33_ASAP7_75t_L g1608 ( 
.A1(n_1451),
.A2(n_1455),
.B1(n_715),
.B2(n_1072),
.Y(n_1608)
);

CKINVDCx20_ASAP7_75t_R g1609 ( 
.A(n_1315),
.Y(n_1609)
);

AOI22xp33_ASAP7_75t_L g1610 ( 
.A1(n_1429),
.A2(n_715),
.B1(n_1451),
.B2(n_846),
.Y(n_1610)
);

CKINVDCx20_ASAP7_75t_R g1611 ( 
.A(n_1315),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1352),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1352),
.Y(n_1613)
);

AND2x2_ASAP7_75t_L g1614 ( 
.A(n_1522),
.B(n_1501),
.Y(n_1614)
);

BUFx3_ASAP7_75t_L g1615 ( 
.A(n_1600),
.Y(n_1615)
);

OR2x2_ASAP7_75t_L g1616 ( 
.A(n_1582),
.B(n_1556),
.Y(n_1616)
);

BUFx2_ASAP7_75t_L g1617 ( 
.A(n_1501),
.Y(n_1617)
);

INVx3_ASAP7_75t_L g1618 ( 
.A(n_1557),
.Y(n_1618)
);

INVx2_ASAP7_75t_SL g1619 ( 
.A(n_1485),
.Y(n_1619)
);

HB1xp67_ASAP7_75t_L g1620 ( 
.A(n_1493),
.Y(n_1620)
);

BUFx3_ASAP7_75t_L g1621 ( 
.A(n_1600),
.Y(n_1621)
);

INVx1_ASAP7_75t_SL g1622 ( 
.A(n_1526),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1504),
.Y(n_1623)
);

INVx1_ASAP7_75t_SL g1624 ( 
.A(n_1597),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1521),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1544),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1549),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1485),
.Y(n_1628)
);

BUFx2_ASAP7_75t_L g1629 ( 
.A(n_1485),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1522),
.B(n_1556),
.Y(n_1630)
);

INVx2_ASAP7_75t_SL g1631 ( 
.A(n_1485),
.Y(n_1631)
);

OAI21x1_ASAP7_75t_L g1632 ( 
.A1(n_1532),
.A2(n_1527),
.B(n_1554),
.Y(n_1632)
);

OAI21x1_ASAP7_75t_L g1633 ( 
.A1(n_1545),
.A2(n_1515),
.B(n_1552),
.Y(n_1633)
);

BUFx6f_ASAP7_75t_L g1634 ( 
.A(n_1600),
.Y(n_1634)
);

AO21x2_ASAP7_75t_L g1635 ( 
.A1(n_1550),
.A2(n_1547),
.B(n_1546),
.Y(n_1635)
);

BUFx2_ASAP7_75t_L g1636 ( 
.A(n_1470),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1599),
.Y(n_1637)
);

INVx5_ASAP7_75t_L g1638 ( 
.A(n_1600),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1506),
.B(n_1498),
.Y(n_1639)
);

AND2x2_ASAP7_75t_L g1640 ( 
.A(n_1523),
.B(n_1555),
.Y(n_1640)
);

NOR2x1_ASAP7_75t_L g1641 ( 
.A(n_1534),
.B(n_1528),
.Y(n_1641)
);

AND2x2_ASAP7_75t_L g1642 ( 
.A(n_1523),
.B(n_1464),
.Y(n_1642)
);

AND2x2_ASAP7_75t_L g1643 ( 
.A(n_1472),
.B(n_1477),
.Y(n_1643)
);

AND2x2_ASAP7_75t_L g1644 ( 
.A(n_1486),
.B(n_1487),
.Y(n_1644)
);

OR2x2_ASAP7_75t_L g1645 ( 
.A(n_1488),
.B(n_1506),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1599),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1470),
.Y(n_1647)
);

BUFx4f_ASAP7_75t_SL g1648 ( 
.A(n_1585),
.Y(n_1648)
);

OAI21x1_ASAP7_75t_L g1649 ( 
.A1(n_1545),
.A2(n_1562),
.B(n_1541),
.Y(n_1649)
);

AO21x2_ASAP7_75t_L g1650 ( 
.A1(n_1546),
.A2(n_1551),
.B(n_1548),
.Y(n_1650)
);

CKINVDCx5p33_ASAP7_75t_R g1651 ( 
.A(n_1598),
.Y(n_1651)
);

INVx4_ASAP7_75t_L g1652 ( 
.A(n_1480),
.Y(n_1652)
);

INVx8_ASAP7_75t_L g1653 ( 
.A(n_1531),
.Y(n_1653)
);

INVx3_ASAP7_75t_L g1654 ( 
.A(n_1560),
.Y(n_1654)
);

INVxp33_ASAP7_75t_L g1655 ( 
.A(n_1568),
.Y(n_1655)
);

INVx1_ASAP7_75t_SL g1656 ( 
.A(n_1474),
.Y(n_1656)
);

HB1xp67_ASAP7_75t_L g1657 ( 
.A(n_1489),
.Y(n_1657)
);

BUFx2_ASAP7_75t_L g1658 ( 
.A(n_1539),
.Y(n_1658)
);

CKINVDCx6p67_ASAP7_75t_R g1659 ( 
.A(n_1469),
.Y(n_1659)
);

INVxp67_ASAP7_75t_L g1660 ( 
.A(n_1566),
.Y(n_1660)
);

INVx2_ASAP7_75t_SL g1661 ( 
.A(n_1494),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1613),
.Y(n_1662)
);

OAI21x1_ASAP7_75t_L g1663 ( 
.A1(n_1541),
.A2(n_1529),
.B(n_1539),
.Y(n_1663)
);

AND2x2_ASAP7_75t_L g1664 ( 
.A(n_1496),
.B(n_1572),
.Y(n_1664)
);

INVx1_ASAP7_75t_SL g1665 ( 
.A(n_1569),
.Y(n_1665)
);

OR2x2_ASAP7_75t_L g1666 ( 
.A(n_1488),
.B(n_1553),
.Y(n_1666)
);

OAI21x1_ASAP7_75t_L g1667 ( 
.A1(n_1533),
.A2(n_1535),
.B(n_1519),
.Y(n_1667)
);

OAI21x1_ASAP7_75t_L g1668 ( 
.A1(n_1533),
.A2(n_1535),
.B(n_1519),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1612),
.Y(n_1669)
);

INVxp67_ASAP7_75t_L g1670 ( 
.A(n_1591),
.Y(n_1670)
);

AND2x2_ASAP7_75t_L g1671 ( 
.A(n_1579),
.B(n_1584),
.Y(n_1671)
);

OAI21xp33_ASAP7_75t_SL g1672 ( 
.A1(n_1565),
.A2(n_1461),
.B(n_1462),
.Y(n_1672)
);

OA21x2_ASAP7_75t_L g1673 ( 
.A1(n_1516),
.A2(n_1463),
.B(n_1570),
.Y(n_1673)
);

INVx2_ASAP7_75t_L g1674 ( 
.A(n_1558),
.Y(n_1674)
);

HB1xp67_ASAP7_75t_L g1675 ( 
.A(n_1606),
.Y(n_1675)
);

INVx2_ASAP7_75t_L g1676 ( 
.A(n_1558),
.Y(n_1676)
);

BUFx2_ASAP7_75t_L g1677 ( 
.A(n_1558),
.Y(n_1677)
);

AOI21xp33_ASAP7_75t_L g1678 ( 
.A1(n_1505),
.A2(n_1490),
.B(n_1581),
.Y(n_1678)
);

AND2x2_ASAP7_75t_L g1679 ( 
.A(n_1512),
.B(n_1473),
.Y(n_1679)
);

AND2x4_ASAP7_75t_L g1680 ( 
.A(n_1480),
.B(n_1576),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1510),
.Y(n_1681)
);

NAND2xp5_ASAP7_75t_L g1682 ( 
.A(n_1473),
.B(n_1571),
.Y(n_1682)
);

CKINVDCx20_ASAP7_75t_R g1683 ( 
.A(n_1595),
.Y(n_1683)
);

AND2x2_ASAP7_75t_L g1684 ( 
.A(n_1512),
.B(n_1593),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1475),
.Y(n_1685)
);

AOI21x1_ASAP7_75t_L g1686 ( 
.A1(n_1543),
.A2(n_1482),
.B(n_1538),
.Y(n_1686)
);

OAI21x1_ASAP7_75t_L g1687 ( 
.A1(n_1537),
.A2(n_1540),
.B(n_1495),
.Y(n_1687)
);

INVx3_ASAP7_75t_L g1688 ( 
.A(n_1494),
.Y(n_1688)
);

OR2x2_ASAP7_75t_L g1689 ( 
.A(n_1468),
.B(n_1511),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1583),
.Y(n_1690)
);

INVx1_ASAP7_75t_SL g1691 ( 
.A(n_1465),
.Y(n_1691)
);

AND2x2_ASAP7_75t_L g1692 ( 
.A(n_1564),
.B(n_1462),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1589),
.Y(n_1693)
);

BUFx3_ASAP7_75t_L g1694 ( 
.A(n_1494),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1592),
.Y(n_1695)
);

HB1xp67_ASAP7_75t_L g1696 ( 
.A(n_1525),
.Y(n_1696)
);

BUFx2_ASAP7_75t_L g1697 ( 
.A(n_1480),
.Y(n_1697)
);

INVx2_ASAP7_75t_SL g1698 ( 
.A(n_1514),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1542),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1542),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1571),
.Y(n_1701)
);

OAI21x1_ASAP7_75t_L g1702 ( 
.A1(n_1537),
.A2(n_1540),
.B(n_1520),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1490),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1530),
.Y(n_1704)
);

INVx2_ASAP7_75t_L g1705 ( 
.A(n_1576),
.Y(n_1705)
);

HB1xp67_ASAP7_75t_L g1706 ( 
.A(n_1536),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1576),
.Y(n_1707)
);

AND2x2_ASAP7_75t_L g1708 ( 
.A(n_1559),
.B(n_1561),
.Y(n_1708)
);

NOR2xp33_ASAP7_75t_R g1709 ( 
.A(n_1609),
.B(n_1611),
.Y(n_1709)
);

OR2x6_ASAP7_75t_L g1710 ( 
.A(n_1580),
.B(n_1502),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1520),
.Y(n_1711)
);

AND2x2_ASAP7_75t_L g1712 ( 
.A(n_1559),
.B(n_1561),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1481),
.Y(n_1713)
);

OAI21x1_ASAP7_75t_L g1714 ( 
.A1(n_1524),
.A2(n_1513),
.B(n_1499),
.Y(n_1714)
);

OA21x2_ASAP7_75t_L g1715 ( 
.A1(n_1563),
.A2(n_1601),
.B(n_1608),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1502),
.Y(n_1716)
);

BUFx3_ASAP7_75t_L g1717 ( 
.A(n_1514),
.Y(n_1717)
);

AOI221xp5_ASAP7_75t_L g1718 ( 
.A1(n_1581),
.A2(n_1586),
.B1(n_1608),
.B2(n_1601),
.C(n_1588),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1574),
.Y(n_1719)
);

OAI21x1_ASAP7_75t_L g1720 ( 
.A1(n_1513),
.A2(n_1580),
.B(n_1500),
.Y(n_1720)
);

AOI22xp33_ASAP7_75t_L g1721 ( 
.A1(n_1563),
.A2(n_1588),
.B1(n_1586),
.B2(n_1610),
.Y(n_1721)
);

INVx3_ASAP7_75t_L g1722 ( 
.A(n_1514),
.Y(n_1722)
);

OAI22xp5_ASAP7_75t_SL g1723 ( 
.A1(n_1497),
.A2(n_1503),
.B1(n_1517),
.B2(n_1511),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1492),
.Y(n_1724)
);

BUFx2_ASAP7_75t_L g1725 ( 
.A(n_1518),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1492),
.Y(n_1726)
);

AND2x2_ASAP7_75t_L g1727 ( 
.A(n_1503),
.B(n_1497),
.Y(n_1727)
);

INVx3_ASAP7_75t_L g1728 ( 
.A(n_1476),
.Y(n_1728)
);

INVx3_ASAP7_75t_L g1729 ( 
.A(n_1476),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1573),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1575),
.Y(n_1731)
);

BUFx3_ASAP7_75t_L g1732 ( 
.A(n_1575),
.Y(n_1732)
);

AOI22xp33_ASAP7_75t_L g1733 ( 
.A1(n_1508),
.A2(n_1478),
.B1(n_1471),
.B2(n_1483),
.Y(n_1733)
);

AOI22xp5_ASAP7_75t_L g1734 ( 
.A1(n_1718),
.A2(n_1602),
.B1(n_1590),
.B2(n_1478),
.Y(n_1734)
);

NOR2xp33_ASAP7_75t_L g1735 ( 
.A(n_1648),
.B(n_1466),
.Y(n_1735)
);

OAI21xp5_ASAP7_75t_L g1736 ( 
.A1(n_1672),
.A2(n_1479),
.B(n_1605),
.Y(n_1736)
);

AND2x2_ASAP7_75t_L g1737 ( 
.A(n_1706),
.B(n_1466),
.Y(n_1737)
);

NAND4xp25_ASAP7_75t_L g1738 ( 
.A(n_1678),
.B(n_1682),
.C(n_1701),
.D(n_1721),
.Y(n_1738)
);

OR2x2_ASAP7_75t_L g1739 ( 
.A(n_1620),
.B(n_1578),
.Y(n_1739)
);

INVx3_ASAP7_75t_L g1740 ( 
.A(n_1694),
.Y(n_1740)
);

OAI22xp5_ASAP7_75t_L g1741 ( 
.A1(n_1701),
.A2(n_1602),
.B1(n_1578),
.B2(n_1605),
.Y(n_1741)
);

O2A1O1Ixp33_ASAP7_75t_SL g1742 ( 
.A1(n_1691),
.A2(n_1484),
.B(n_1587),
.C(n_1507),
.Y(n_1742)
);

AND2x2_ASAP7_75t_L g1743 ( 
.A(n_1630),
.B(n_1603),
.Y(n_1743)
);

AOI221xp5_ASAP7_75t_L g1744 ( 
.A1(n_1672),
.A2(n_1469),
.B1(n_1467),
.B2(n_1607),
.C(n_1577),
.Y(n_1744)
);

AND2x2_ASAP7_75t_L g1745 ( 
.A(n_1630),
.B(n_1567),
.Y(n_1745)
);

A2O1A1Ixp33_ASAP7_75t_L g1746 ( 
.A1(n_1727),
.A2(n_1604),
.B(n_1594),
.C(n_1602),
.Y(n_1746)
);

AND2x4_ASAP7_75t_L g1747 ( 
.A(n_1680),
.B(n_1484),
.Y(n_1747)
);

OA21x2_ASAP7_75t_L g1748 ( 
.A1(n_1632),
.A2(n_1491),
.B(n_1567),
.Y(n_1748)
);

NOR2xp33_ASAP7_75t_R g1749 ( 
.A(n_1683),
.B(n_1594),
.Y(n_1749)
);

AND2x2_ASAP7_75t_L g1750 ( 
.A(n_1656),
.B(n_1509),
.Y(n_1750)
);

OR2x2_ASAP7_75t_L g1751 ( 
.A(n_1616),
.B(n_1596),
.Y(n_1751)
);

AND2x2_ASAP7_75t_L g1752 ( 
.A(n_1665),
.B(n_1660),
.Y(n_1752)
);

NOR2x1_ASAP7_75t_R g1753 ( 
.A(n_1651),
.B(n_1652),
.Y(n_1753)
);

AND2x2_ASAP7_75t_L g1754 ( 
.A(n_1670),
.B(n_1614),
.Y(n_1754)
);

AND2x4_ASAP7_75t_L g1755 ( 
.A(n_1680),
.B(n_1697),
.Y(n_1755)
);

A2O1A1Ixp33_ASAP7_75t_L g1756 ( 
.A1(n_1727),
.A2(n_1712),
.B(n_1708),
.C(n_1679),
.Y(n_1756)
);

AND2x4_ASAP7_75t_L g1757 ( 
.A(n_1680),
.B(n_1697),
.Y(n_1757)
);

AOI21xp5_ASAP7_75t_L g1758 ( 
.A1(n_1641),
.A2(n_1673),
.B(n_1636),
.Y(n_1758)
);

BUFx2_ASAP7_75t_L g1759 ( 
.A(n_1694),
.Y(n_1759)
);

OR2x2_ASAP7_75t_L g1760 ( 
.A(n_1657),
.B(n_1675),
.Y(n_1760)
);

INVx6_ASAP7_75t_L g1761 ( 
.A(n_1653),
.Y(n_1761)
);

AND2x2_ASAP7_75t_L g1762 ( 
.A(n_1614),
.B(n_1725),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1662),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1662),
.Y(n_1764)
);

AO32x2_ASAP7_75t_L g1765 ( 
.A1(n_1723),
.A2(n_1619),
.A3(n_1631),
.B1(n_1661),
.B2(n_1698),
.Y(n_1765)
);

AOI22xp5_ASAP7_75t_L g1766 ( 
.A1(n_1723),
.A2(n_1715),
.B1(n_1679),
.B2(n_1708),
.Y(n_1766)
);

AND2x2_ASAP7_75t_L g1767 ( 
.A(n_1643),
.B(n_1644),
.Y(n_1767)
);

AND2x4_ASAP7_75t_L g1768 ( 
.A(n_1615),
.B(n_1621),
.Y(n_1768)
);

OAI22xp5_ASAP7_75t_L g1769 ( 
.A1(n_1673),
.A2(n_1715),
.B1(n_1726),
.B2(n_1724),
.Y(n_1769)
);

AND2x2_ASAP7_75t_L g1770 ( 
.A(n_1644),
.B(n_1664),
.Y(n_1770)
);

AO32x2_ASAP7_75t_L g1771 ( 
.A1(n_1619),
.A2(n_1631),
.A3(n_1698),
.B1(n_1661),
.B2(n_1652),
.Y(n_1771)
);

OAI21x1_ASAP7_75t_L g1772 ( 
.A1(n_1632),
.A2(n_1649),
.B(n_1633),
.Y(n_1772)
);

AND2x2_ASAP7_75t_L g1773 ( 
.A(n_1664),
.B(n_1671),
.Y(n_1773)
);

NAND2xp5_ASAP7_75t_L g1774 ( 
.A(n_1639),
.B(n_1724),
.Y(n_1774)
);

NOR2xp33_ASAP7_75t_L g1775 ( 
.A(n_1624),
.B(n_1622),
.Y(n_1775)
);

CKINVDCx8_ASAP7_75t_R g1776 ( 
.A(n_1653),
.Y(n_1776)
);

CKINVDCx5p33_ASAP7_75t_R g1777 ( 
.A(n_1709),
.Y(n_1777)
);

O2A1O1Ixp33_ASAP7_75t_L g1778 ( 
.A1(n_1726),
.A2(n_1673),
.B(n_1655),
.C(n_1703),
.Y(n_1778)
);

O2A1O1Ixp33_ASAP7_75t_L g1779 ( 
.A1(n_1673),
.A2(n_1703),
.B(n_1641),
.C(n_1699),
.Y(n_1779)
);

NAND2xp5_ASAP7_75t_L g1780 ( 
.A(n_1671),
.B(n_1669),
.Y(n_1780)
);

AOI22xp5_ASAP7_75t_L g1781 ( 
.A1(n_1715),
.A2(n_1712),
.B1(n_1640),
.B2(n_1692),
.Y(n_1781)
);

A2O1A1Ixp33_ASAP7_75t_L g1782 ( 
.A1(n_1714),
.A2(n_1687),
.B(n_1689),
.C(n_1642),
.Y(n_1782)
);

AND2x2_ASAP7_75t_L g1783 ( 
.A(n_1684),
.B(n_1696),
.Y(n_1783)
);

BUFx4f_ASAP7_75t_L g1784 ( 
.A(n_1659),
.Y(n_1784)
);

AOI22xp5_ASAP7_75t_L g1785 ( 
.A1(n_1715),
.A2(n_1692),
.B1(n_1689),
.B2(n_1642),
.Y(n_1785)
);

OAI22xp5_ASAP7_75t_L g1786 ( 
.A1(n_1699),
.A2(n_1700),
.B1(n_1636),
.B2(n_1645),
.Y(n_1786)
);

OA21x2_ASAP7_75t_L g1787 ( 
.A1(n_1633),
.A2(n_1687),
.B(n_1649),
.Y(n_1787)
);

HB1xp67_ASAP7_75t_L g1788 ( 
.A(n_1704),
.Y(n_1788)
);

AOI21xp5_ASAP7_75t_L g1789 ( 
.A1(n_1647),
.A2(n_1629),
.B(n_1650),
.Y(n_1789)
);

OR2x6_ASAP7_75t_L g1790 ( 
.A(n_1634),
.B(n_1652),
.Y(n_1790)
);

INVx3_ASAP7_75t_L g1791 ( 
.A(n_1717),
.Y(n_1791)
);

A2O1A1Ixp33_ASAP7_75t_L g1792 ( 
.A1(n_1714),
.A2(n_1668),
.B(n_1667),
.C(n_1720),
.Y(n_1792)
);

OAI22xp5_ASAP7_75t_L g1793 ( 
.A1(n_1700),
.A2(n_1645),
.B1(n_1666),
.B2(n_1617),
.Y(n_1793)
);

OAI21xp5_ASAP7_75t_L g1794 ( 
.A1(n_1667),
.A2(n_1668),
.B(n_1686),
.Y(n_1794)
);

OR2x6_ASAP7_75t_L g1795 ( 
.A(n_1634),
.B(n_1652),
.Y(n_1795)
);

AOI21xp5_ASAP7_75t_L g1796 ( 
.A1(n_1647),
.A2(n_1629),
.B(n_1650),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1681),
.Y(n_1797)
);

AND2x2_ASAP7_75t_L g1798 ( 
.A(n_1730),
.B(n_1731),
.Y(n_1798)
);

INVx4_ASAP7_75t_L g1799 ( 
.A(n_1688),
.Y(n_1799)
);

A2O1A1Ixp33_ASAP7_75t_L g1800 ( 
.A1(n_1720),
.A2(n_1713),
.B(n_1702),
.C(n_1617),
.Y(n_1800)
);

AND2x4_ASAP7_75t_L g1801 ( 
.A(n_1638),
.B(n_1677),
.Y(n_1801)
);

NAND2xp5_ASAP7_75t_L g1802 ( 
.A(n_1688),
.B(n_1722),
.Y(n_1802)
);

NAND2xp5_ASAP7_75t_L g1803 ( 
.A(n_1688),
.B(n_1722),
.Y(n_1803)
);

AND2x2_ASAP7_75t_L g1804 ( 
.A(n_1732),
.B(n_1711),
.Y(n_1804)
);

AND2x2_ASAP7_75t_L g1805 ( 
.A(n_1732),
.B(n_1711),
.Y(n_1805)
);

A2O1A1Ixp33_ASAP7_75t_L g1806 ( 
.A1(n_1713),
.A2(n_1702),
.B(n_1663),
.C(n_1707),
.Y(n_1806)
);

NAND2xp5_ASAP7_75t_L g1807 ( 
.A(n_1637),
.B(n_1646),
.Y(n_1807)
);

INVx2_ASAP7_75t_L g1808 ( 
.A(n_1763),
.Y(n_1808)
);

INVx2_ASAP7_75t_L g1809 ( 
.A(n_1764),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1807),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1807),
.Y(n_1811)
);

BUFx3_ASAP7_75t_L g1812 ( 
.A(n_1747),
.Y(n_1812)
);

BUFx2_ASAP7_75t_L g1813 ( 
.A(n_1771),
.Y(n_1813)
);

AND2x2_ASAP7_75t_L g1814 ( 
.A(n_1767),
.B(n_1650),
.Y(n_1814)
);

INVxp67_ASAP7_75t_SL g1815 ( 
.A(n_1779),
.Y(n_1815)
);

HB1xp67_ASAP7_75t_L g1816 ( 
.A(n_1788),
.Y(n_1816)
);

INVx2_ASAP7_75t_L g1817 ( 
.A(n_1787),
.Y(n_1817)
);

BUFx3_ASAP7_75t_L g1818 ( 
.A(n_1747),
.Y(n_1818)
);

AND2x2_ASAP7_75t_L g1819 ( 
.A(n_1770),
.B(n_1635),
.Y(n_1819)
);

AND2x2_ASAP7_75t_L g1820 ( 
.A(n_1773),
.B(n_1635),
.Y(n_1820)
);

OR2x2_ASAP7_75t_L g1821 ( 
.A(n_1760),
.B(n_1635),
.Y(n_1821)
);

BUFx8_ASAP7_75t_SL g1822 ( 
.A(n_1777),
.Y(n_1822)
);

BUFx2_ASAP7_75t_L g1823 ( 
.A(n_1771),
.Y(n_1823)
);

NOR2xp33_ASAP7_75t_L g1824 ( 
.A(n_1739),
.B(n_1686),
.Y(n_1824)
);

NAND2xp5_ASAP7_75t_L g1825 ( 
.A(n_1758),
.B(n_1646),
.Y(n_1825)
);

INVx3_ASAP7_75t_L g1826 ( 
.A(n_1772),
.Y(n_1826)
);

AOI22xp33_ASAP7_75t_L g1827 ( 
.A1(n_1738),
.A2(n_1626),
.B1(n_1627),
.B2(n_1693),
.Y(n_1827)
);

INVxp67_ASAP7_75t_SL g1828 ( 
.A(n_1789),
.Y(n_1828)
);

AND2x2_ASAP7_75t_L g1829 ( 
.A(n_1762),
.B(n_1658),
.Y(n_1829)
);

OR2x2_ASAP7_75t_L g1830 ( 
.A(n_1793),
.B(n_1658),
.Y(n_1830)
);

INVx2_ASAP7_75t_L g1831 ( 
.A(n_1787),
.Y(n_1831)
);

NAND2xp5_ASAP7_75t_L g1832 ( 
.A(n_1786),
.B(n_1769),
.Y(n_1832)
);

AND2x2_ASAP7_75t_L g1833 ( 
.A(n_1754),
.B(n_1663),
.Y(n_1833)
);

INVx2_ASAP7_75t_L g1834 ( 
.A(n_1771),
.Y(n_1834)
);

NAND2xp5_ASAP7_75t_L g1835 ( 
.A(n_1769),
.B(n_1625),
.Y(n_1835)
);

BUFx3_ASAP7_75t_L g1836 ( 
.A(n_1748),
.Y(n_1836)
);

BUFx6f_ASAP7_75t_L g1837 ( 
.A(n_1748),
.Y(n_1837)
);

BUFx2_ASAP7_75t_L g1838 ( 
.A(n_1759),
.Y(n_1838)
);

INVx2_ASAP7_75t_L g1839 ( 
.A(n_1797),
.Y(n_1839)
);

AOI22xp33_ASAP7_75t_L g1840 ( 
.A1(n_1738),
.A2(n_1627),
.B1(n_1626),
.B2(n_1695),
.Y(n_1840)
);

AND2x2_ASAP7_75t_L g1841 ( 
.A(n_1783),
.B(n_1628),
.Y(n_1841)
);

AND2x2_ASAP7_75t_L g1842 ( 
.A(n_1780),
.B(n_1628),
.Y(n_1842)
);

INVxp67_ASAP7_75t_SL g1843 ( 
.A(n_1796),
.Y(n_1843)
);

INVxp67_ASAP7_75t_SL g1844 ( 
.A(n_1778),
.Y(n_1844)
);

OR2x2_ASAP7_75t_L g1845 ( 
.A(n_1774),
.B(n_1618),
.Y(n_1845)
);

NAND2xp5_ASAP7_75t_L g1846 ( 
.A(n_1785),
.B(n_1625),
.Y(n_1846)
);

NAND2xp5_ASAP7_75t_L g1847 ( 
.A(n_1785),
.B(n_1623),
.Y(n_1847)
);

NAND2xp5_ASAP7_75t_L g1848 ( 
.A(n_1781),
.B(n_1623),
.Y(n_1848)
);

INVx2_ASAP7_75t_L g1849 ( 
.A(n_1765),
.Y(n_1849)
);

AOI22xp33_ASAP7_75t_L g1850 ( 
.A1(n_1766),
.A2(n_1695),
.B1(n_1685),
.B2(n_1690),
.Y(n_1850)
);

NAND2xp5_ASAP7_75t_L g1851 ( 
.A(n_1781),
.B(n_1618),
.Y(n_1851)
);

AND2x2_ASAP7_75t_L g1852 ( 
.A(n_1813),
.B(n_1743),
.Y(n_1852)
);

OAI33xp33_ASAP7_75t_L g1853 ( 
.A1(n_1832),
.A2(n_1741),
.A3(n_1751),
.B1(n_1802),
.B2(n_1803),
.B3(n_1756),
.Y(n_1853)
);

NAND3xp33_ASAP7_75t_L g1854 ( 
.A(n_1815),
.B(n_1744),
.C(n_1766),
.Y(n_1854)
);

OR2x2_ASAP7_75t_L g1855 ( 
.A(n_1832),
.B(n_1782),
.Y(n_1855)
);

AND2x2_ASAP7_75t_L g1856 ( 
.A(n_1813),
.B(n_1745),
.Y(n_1856)
);

NOR2xp67_ASAP7_75t_L g1857 ( 
.A(n_1834),
.B(n_1794),
.Y(n_1857)
);

AND2x2_ASAP7_75t_L g1858 ( 
.A(n_1813),
.B(n_1752),
.Y(n_1858)
);

AOI22xp33_ASAP7_75t_SL g1859 ( 
.A1(n_1815),
.A2(n_1794),
.B1(n_1736),
.B2(n_1765),
.Y(n_1859)
);

AND2x2_ASAP7_75t_L g1860 ( 
.A(n_1823),
.B(n_1737),
.Y(n_1860)
);

AND2x2_ASAP7_75t_L g1861 ( 
.A(n_1823),
.B(n_1804),
.Y(n_1861)
);

INVx2_ASAP7_75t_L g1862 ( 
.A(n_1817),
.Y(n_1862)
);

AOI211xp5_ASAP7_75t_SL g1863 ( 
.A1(n_1844),
.A2(n_1742),
.B(n_1741),
.C(n_1746),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1839),
.Y(n_1864)
);

NAND2xp5_ASAP7_75t_L g1865 ( 
.A(n_1814),
.B(n_1800),
.Y(n_1865)
);

INVx2_ASAP7_75t_L g1866 ( 
.A(n_1817),
.Y(n_1866)
);

NAND2xp5_ASAP7_75t_L g1867 ( 
.A(n_1814),
.B(n_1798),
.Y(n_1867)
);

INVxp67_ASAP7_75t_L g1868 ( 
.A(n_1824),
.Y(n_1868)
);

INVx2_ASAP7_75t_L g1869 ( 
.A(n_1817),
.Y(n_1869)
);

HB1xp67_ASAP7_75t_L g1870 ( 
.A(n_1816),
.Y(n_1870)
);

AND2x2_ASAP7_75t_L g1871 ( 
.A(n_1823),
.B(n_1805),
.Y(n_1871)
);

NOR2x1_ASAP7_75t_L g1872 ( 
.A(n_1812),
.B(n_1740),
.Y(n_1872)
);

INVx3_ASAP7_75t_L g1873 ( 
.A(n_1826),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1808),
.Y(n_1874)
);

AND2x2_ASAP7_75t_L g1875 ( 
.A(n_1829),
.B(n_1791),
.Y(n_1875)
);

AND2x2_ASAP7_75t_L g1876 ( 
.A(n_1829),
.B(n_1791),
.Y(n_1876)
);

NOR2xp33_ASAP7_75t_L g1877 ( 
.A(n_1822),
.B(n_1735),
.Y(n_1877)
);

AOI221xp5_ASAP7_75t_L g1878 ( 
.A1(n_1844),
.A2(n_1792),
.B1(n_1806),
.B2(n_1734),
.C(n_1736),
.Y(n_1878)
);

INVx1_ASAP7_75t_L g1879 ( 
.A(n_1808),
.Y(n_1879)
);

INVx5_ASAP7_75t_L g1880 ( 
.A(n_1837),
.Y(n_1880)
);

OAI31xp33_ASAP7_75t_L g1881 ( 
.A1(n_1827),
.A2(n_1765),
.A3(n_1750),
.B(n_1734),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1808),
.Y(n_1882)
);

BUFx2_ASAP7_75t_L g1883 ( 
.A(n_1812),
.Y(n_1883)
);

OR2x6_ASAP7_75t_L g1884 ( 
.A(n_1849),
.B(n_1790),
.Y(n_1884)
);

INVx2_ASAP7_75t_L g1885 ( 
.A(n_1817),
.Y(n_1885)
);

INVx2_ASAP7_75t_L g1886 ( 
.A(n_1831),
.Y(n_1886)
);

INVx4_ASAP7_75t_L g1887 ( 
.A(n_1822),
.Y(n_1887)
);

AOI22xp33_ASAP7_75t_SL g1888 ( 
.A1(n_1849),
.A2(n_1707),
.B1(n_1705),
.B2(n_1638),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1809),
.Y(n_1889)
);

AOI22xp5_ASAP7_75t_L g1890 ( 
.A1(n_1827),
.A2(n_1710),
.B1(n_1775),
.B2(n_1705),
.Y(n_1890)
);

INVx1_ASAP7_75t_SL g1891 ( 
.A(n_1838),
.Y(n_1891)
);

OAI31xp33_ASAP7_75t_L g1892 ( 
.A1(n_1840),
.A2(n_1733),
.A3(n_1757),
.B(n_1755),
.Y(n_1892)
);

OAI22xp5_ASAP7_75t_L g1893 ( 
.A1(n_1840),
.A2(n_1776),
.B1(n_1761),
.B2(n_1784),
.Y(n_1893)
);

INVx2_ASAP7_75t_L g1894 ( 
.A(n_1831),
.Y(n_1894)
);

BUFx2_ASAP7_75t_L g1895 ( 
.A(n_1812),
.Y(n_1895)
);

BUFx2_ASAP7_75t_L g1896 ( 
.A(n_1812),
.Y(n_1896)
);

INVx2_ASAP7_75t_L g1897 ( 
.A(n_1831),
.Y(n_1897)
);

AOI22xp33_ASAP7_75t_L g1898 ( 
.A1(n_1850),
.A2(n_1674),
.B1(n_1676),
.B2(n_1654),
.Y(n_1898)
);

AND2x2_ASAP7_75t_L g1899 ( 
.A(n_1819),
.B(n_1820),
.Y(n_1899)
);

INVx2_ASAP7_75t_L g1900 ( 
.A(n_1831),
.Y(n_1900)
);

NAND3xp33_ASAP7_75t_L g1901 ( 
.A(n_1828),
.B(n_1799),
.C(n_1729),
.Y(n_1901)
);

NAND2x1_ASAP7_75t_L g1902 ( 
.A(n_1834),
.B(n_1801),
.Y(n_1902)
);

INVx2_ASAP7_75t_L g1903 ( 
.A(n_1834),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1809),
.Y(n_1904)
);

INVx1_ASAP7_75t_SL g1905 ( 
.A(n_1838),
.Y(n_1905)
);

OAI321xp33_ASAP7_75t_L g1906 ( 
.A1(n_1828),
.A2(n_1710),
.A3(n_1795),
.B1(n_1790),
.B2(n_1719),
.C(n_1716),
.Y(n_1906)
);

AND2x2_ASAP7_75t_L g1907 ( 
.A(n_1820),
.B(n_1768),
.Y(n_1907)
);

AND2x2_ASAP7_75t_L g1908 ( 
.A(n_1833),
.B(n_1768),
.Y(n_1908)
);

AND2x2_ASAP7_75t_L g1909 ( 
.A(n_1883),
.B(n_1838),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1903),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1903),
.Y(n_1911)
);

AND2x2_ASAP7_75t_L g1912 ( 
.A(n_1883),
.B(n_1818),
.Y(n_1912)
);

AND2x4_ASAP7_75t_L g1913 ( 
.A(n_1880),
.B(n_1836),
.Y(n_1913)
);

AND2x2_ASAP7_75t_L g1914 ( 
.A(n_1895),
.B(n_1818),
.Y(n_1914)
);

INVx2_ASAP7_75t_L g1915 ( 
.A(n_1862),
.Y(n_1915)
);

INVx1_ASAP7_75t_L g1916 ( 
.A(n_1903),
.Y(n_1916)
);

NAND2xp5_ASAP7_75t_L g1917 ( 
.A(n_1868),
.B(n_1810),
.Y(n_1917)
);

AOI221xp5_ASAP7_75t_L g1918 ( 
.A1(n_1854),
.A2(n_1849),
.B1(n_1843),
.B2(n_1848),
.C(n_1835),
.Y(n_1918)
);

INVx1_ASAP7_75t_L g1919 ( 
.A(n_1874),
.Y(n_1919)
);

INVx1_ASAP7_75t_L g1920 ( 
.A(n_1874),
.Y(n_1920)
);

AND2x2_ASAP7_75t_L g1921 ( 
.A(n_1895),
.B(n_1818),
.Y(n_1921)
);

BUFx3_ASAP7_75t_L g1922 ( 
.A(n_1887),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1879),
.Y(n_1923)
);

AND2x2_ASAP7_75t_L g1924 ( 
.A(n_1896),
.B(n_1833),
.Y(n_1924)
);

NOR2xp33_ASAP7_75t_L g1925 ( 
.A(n_1887),
.B(n_1659),
.Y(n_1925)
);

INVx1_ASAP7_75t_L g1926 ( 
.A(n_1879),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_1882),
.Y(n_1927)
);

INVx1_ASAP7_75t_L g1928 ( 
.A(n_1882),
.Y(n_1928)
);

AND2x2_ASAP7_75t_L g1929 ( 
.A(n_1896),
.B(n_1833),
.Y(n_1929)
);

NAND2x1p5_ASAP7_75t_L g1930 ( 
.A(n_1872),
.B(n_1836),
.Y(n_1930)
);

AND2x2_ASAP7_75t_L g1931 ( 
.A(n_1852),
.B(n_1842),
.Y(n_1931)
);

INVx1_ASAP7_75t_SL g1932 ( 
.A(n_1891),
.Y(n_1932)
);

NAND2xp5_ASAP7_75t_L g1933 ( 
.A(n_1855),
.B(n_1810),
.Y(n_1933)
);

INVx1_ASAP7_75t_L g1934 ( 
.A(n_1889),
.Y(n_1934)
);

NAND2xp5_ASAP7_75t_L g1935 ( 
.A(n_1855),
.B(n_1811),
.Y(n_1935)
);

AND2x4_ASAP7_75t_L g1936 ( 
.A(n_1880),
.B(n_1836),
.Y(n_1936)
);

AND2x2_ASAP7_75t_L g1937 ( 
.A(n_1852),
.B(n_1842),
.Y(n_1937)
);

INVx1_ASAP7_75t_SL g1938 ( 
.A(n_1891),
.Y(n_1938)
);

INVx1_ASAP7_75t_SL g1939 ( 
.A(n_1905),
.Y(n_1939)
);

OR2x2_ASAP7_75t_L g1940 ( 
.A(n_1870),
.B(n_1821),
.Y(n_1940)
);

OR2x2_ASAP7_75t_L g1941 ( 
.A(n_1867),
.B(n_1821),
.Y(n_1941)
);

AND2x2_ASAP7_75t_L g1942 ( 
.A(n_1856),
.B(n_1899),
.Y(n_1942)
);

INVx1_ASAP7_75t_L g1943 ( 
.A(n_1889),
.Y(n_1943)
);

AND2x4_ASAP7_75t_L g1944 ( 
.A(n_1880),
.B(n_1836),
.Y(n_1944)
);

AND2x2_ASAP7_75t_L g1945 ( 
.A(n_1908),
.B(n_1818),
.Y(n_1945)
);

INVx1_ASAP7_75t_L g1946 ( 
.A(n_1904),
.Y(n_1946)
);

INVx1_ASAP7_75t_SL g1947 ( 
.A(n_1905),
.Y(n_1947)
);

INVx1_ASAP7_75t_L g1948 ( 
.A(n_1904),
.Y(n_1948)
);

INVx3_ASAP7_75t_L g1949 ( 
.A(n_1880),
.Y(n_1949)
);

AND2x4_ASAP7_75t_SL g1950 ( 
.A(n_1907),
.B(n_1908),
.Y(n_1950)
);

AND2x2_ASAP7_75t_L g1951 ( 
.A(n_1856),
.B(n_1841),
.Y(n_1951)
);

AND2x4_ASAP7_75t_L g1952 ( 
.A(n_1880),
.B(n_1843),
.Y(n_1952)
);

INVx2_ASAP7_75t_L g1953 ( 
.A(n_1862),
.Y(n_1953)
);

AND2x2_ASAP7_75t_L g1954 ( 
.A(n_1899),
.B(n_1842),
.Y(n_1954)
);

HB1xp67_ASAP7_75t_L g1955 ( 
.A(n_1864),
.Y(n_1955)
);

INVx1_ASAP7_75t_L g1956 ( 
.A(n_1864),
.Y(n_1956)
);

NOR2xp67_ASAP7_75t_L g1957 ( 
.A(n_1949),
.B(n_1887),
.Y(n_1957)
);

AOI22xp33_ASAP7_75t_L g1958 ( 
.A1(n_1918),
.A2(n_1854),
.B1(n_1881),
.B2(n_1853),
.Y(n_1958)
);

AND2x4_ASAP7_75t_L g1959 ( 
.A(n_1950),
.B(n_1880),
.Y(n_1959)
);

HB1xp67_ASAP7_75t_L g1960 ( 
.A(n_1917),
.Y(n_1960)
);

AND2x4_ASAP7_75t_L g1961 ( 
.A(n_1950),
.B(n_1872),
.Y(n_1961)
);

OR2x6_ASAP7_75t_L g1962 ( 
.A(n_1913),
.B(n_1837),
.Y(n_1962)
);

INVx2_ASAP7_75t_SL g1963 ( 
.A(n_1922),
.Y(n_1963)
);

INVx2_ASAP7_75t_L g1964 ( 
.A(n_1915),
.Y(n_1964)
);

INVx1_ASAP7_75t_L g1965 ( 
.A(n_1933),
.Y(n_1965)
);

INVx1_ASAP7_75t_SL g1966 ( 
.A(n_1922),
.Y(n_1966)
);

NAND2xp5_ASAP7_75t_L g1967 ( 
.A(n_1933),
.B(n_1858),
.Y(n_1967)
);

INVx1_ASAP7_75t_L g1968 ( 
.A(n_1935),
.Y(n_1968)
);

OAI33xp33_ASAP7_75t_L g1969 ( 
.A1(n_1935),
.A2(n_1865),
.A3(n_1835),
.B1(n_1821),
.B2(n_1825),
.B3(n_1848),
.Y(n_1969)
);

NAND2xp67_ASAP7_75t_L g1970 ( 
.A(n_1915),
.B(n_1858),
.Y(n_1970)
);

OR2x6_ASAP7_75t_L g1971 ( 
.A(n_1913),
.B(n_1837),
.Y(n_1971)
);

OR2x2_ASAP7_75t_L g1972 ( 
.A(n_1917),
.B(n_1867),
.Y(n_1972)
);

OR2x2_ASAP7_75t_L g1973 ( 
.A(n_1941),
.B(n_1845),
.Y(n_1973)
);

AND2x2_ASAP7_75t_L g1974 ( 
.A(n_1950),
.B(n_1860),
.Y(n_1974)
);

INVx2_ASAP7_75t_L g1975 ( 
.A(n_1915),
.Y(n_1975)
);

HB1xp67_ASAP7_75t_L g1976 ( 
.A(n_1932),
.Y(n_1976)
);

INVx1_ASAP7_75t_L g1977 ( 
.A(n_1919),
.Y(n_1977)
);

AND2x2_ASAP7_75t_L g1978 ( 
.A(n_1942),
.B(n_1860),
.Y(n_1978)
);

INVx1_ASAP7_75t_L g1979 ( 
.A(n_1919),
.Y(n_1979)
);

OR2x2_ASAP7_75t_L g1980 ( 
.A(n_1941),
.B(n_1845),
.Y(n_1980)
);

NOR2x1_ASAP7_75t_L g1981 ( 
.A(n_1922),
.B(n_1887),
.Y(n_1981)
);

INVx2_ASAP7_75t_L g1982 ( 
.A(n_1953),
.Y(n_1982)
);

INVx1_ASAP7_75t_L g1983 ( 
.A(n_1920),
.Y(n_1983)
);

OR2x2_ASAP7_75t_L g1984 ( 
.A(n_1940),
.B(n_1816),
.Y(n_1984)
);

HB1xp67_ASAP7_75t_L g1985 ( 
.A(n_1932),
.Y(n_1985)
);

INVx1_ASAP7_75t_L g1986 ( 
.A(n_1920),
.Y(n_1986)
);

AND2x2_ASAP7_75t_L g1987 ( 
.A(n_1942),
.B(n_1861),
.Y(n_1987)
);

AND2x4_ASAP7_75t_L g1988 ( 
.A(n_1942),
.B(n_1901),
.Y(n_1988)
);

NOR2xp33_ASAP7_75t_SL g1989 ( 
.A(n_1925),
.B(n_1753),
.Y(n_1989)
);

AOI21xp33_ASAP7_75t_L g1990 ( 
.A1(n_1918),
.A2(n_1881),
.B(n_1878),
.Y(n_1990)
);

A2O1A1Ixp33_ASAP7_75t_L g1991 ( 
.A1(n_1952),
.A2(n_1863),
.B(n_1892),
.C(n_1859),
.Y(n_1991)
);

INVx2_ASAP7_75t_L g1992 ( 
.A(n_1953),
.Y(n_1992)
);

INVx1_ASAP7_75t_L g1993 ( 
.A(n_1923),
.Y(n_1993)
);

INVx1_ASAP7_75t_L g1994 ( 
.A(n_1923),
.Y(n_1994)
);

O2A1O1Ixp33_ASAP7_75t_SL g1995 ( 
.A1(n_1938),
.A2(n_1863),
.B(n_1877),
.C(n_1902),
.Y(n_1995)
);

HB1xp67_ASAP7_75t_L g1996 ( 
.A(n_1938),
.Y(n_1996)
);

INVx1_ASAP7_75t_L g1997 ( 
.A(n_1926),
.Y(n_1997)
);

INVx1_ASAP7_75t_L g1998 ( 
.A(n_1926),
.Y(n_1998)
);

NAND2xp5_ASAP7_75t_L g1999 ( 
.A(n_1939),
.B(n_1857),
.Y(n_1999)
);

OR2x2_ASAP7_75t_L g2000 ( 
.A(n_1940),
.B(n_1865),
.Y(n_2000)
);

INVx2_ASAP7_75t_L g2001 ( 
.A(n_1953),
.Y(n_2001)
);

INVx1_ASAP7_75t_L g2002 ( 
.A(n_1927),
.Y(n_2002)
);

AOI22xp5_ASAP7_75t_L g2003 ( 
.A1(n_1924),
.A2(n_1890),
.B1(n_1857),
.B2(n_1847),
.Y(n_2003)
);

OR2x2_ASAP7_75t_L g2004 ( 
.A(n_1972),
.B(n_1939),
.Y(n_2004)
);

NOR2xp33_ASAP7_75t_L g2005 ( 
.A(n_1966),
.B(n_1947),
.Y(n_2005)
);

NAND2xp5_ASAP7_75t_L g2006 ( 
.A(n_1958),
.B(n_1931),
.Y(n_2006)
);

INVx1_ASAP7_75t_L g2007 ( 
.A(n_1977),
.Y(n_2007)
);

AND2x2_ASAP7_75t_L g2008 ( 
.A(n_1974),
.B(n_1912),
.Y(n_2008)
);

OR2x2_ASAP7_75t_L g2009 ( 
.A(n_1972),
.B(n_1947),
.Y(n_2009)
);

AND2x4_ASAP7_75t_L g2010 ( 
.A(n_1957),
.B(n_1913),
.Y(n_2010)
);

OR2x2_ASAP7_75t_L g2011 ( 
.A(n_2000),
.B(n_1927),
.Y(n_2011)
);

AND4x1_ASAP7_75t_L g2012 ( 
.A(n_1991),
.B(n_1958),
.C(n_1981),
.D(n_1989),
.Y(n_2012)
);

AND2x2_ASAP7_75t_L g2013 ( 
.A(n_1974),
.B(n_1912),
.Y(n_2013)
);

NAND2x1p5_ASAP7_75t_L g2014 ( 
.A(n_1963),
.B(n_1784),
.Y(n_2014)
);

NAND2xp5_ASAP7_75t_L g2015 ( 
.A(n_1976),
.B(n_1931),
.Y(n_2015)
);

OAI31xp33_ASAP7_75t_L g2016 ( 
.A1(n_1990),
.A2(n_1892),
.A3(n_1824),
.B(n_1893),
.Y(n_2016)
);

INVx2_ASAP7_75t_L g2017 ( 
.A(n_1964),
.Y(n_2017)
);

INVx3_ASAP7_75t_L g2018 ( 
.A(n_1959),
.Y(n_2018)
);

OR2x2_ASAP7_75t_L g2019 ( 
.A(n_2000),
.B(n_1965),
.Y(n_2019)
);

AND2x2_ASAP7_75t_L g2020 ( 
.A(n_1978),
.B(n_1914),
.Y(n_2020)
);

INVx1_ASAP7_75t_L g2021 ( 
.A(n_1979),
.Y(n_2021)
);

INVx1_ASAP7_75t_L g2022 ( 
.A(n_1983),
.Y(n_2022)
);

OAI31xp33_ASAP7_75t_L g2023 ( 
.A1(n_1991),
.A2(n_1893),
.A3(n_1851),
.B(n_1846),
.Y(n_2023)
);

INVx2_ASAP7_75t_L g2024 ( 
.A(n_1964),
.Y(n_2024)
);

INVx2_ASAP7_75t_L g2025 ( 
.A(n_1975),
.Y(n_2025)
);

INVxp67_ASAP7_75t_SL g2026 ( 
.A(n_1985),
.Y(n_2026)
);

NAND2xp5_ASAP7_75t_L g2027 ( 
.A(n_1996),
.B(n_1931),
.Y(n_2027)
);

INVx1_ASAP7_75t_SL g2028 ( 
.A(n_1963),
.Y(n_2028)
);

INVx1_ASAP7_75t_L g2029 ( 
.A(n_1986),
.Y(n_2029)
);

INVx1_ASAP7_75t_L g2030 ( 
.A(n_1993),
.Y(n_2030)
);

INVx1_ASAP7_75t_L g2031 ( 
.A(n_1994),
.Y(n_2031)
);

NAND4xp75_ASAP7_75t_L g2032 ( 
.A(n_2003),
.B(n_1890),
.C(n_1851),
.D(n_1846),
.Y(n_2032)
);

AND2x2_ASAP7_75t_L g2033 ( 
.A(n_1978),
.B(n_1914),
.Y(n_2033)
);

NAND2xp5_ASAP7_75t_L g2034 ( 
.A(n_1960),
.B(n_1937),
.Y(n_2034)
);

AND2x2_ASAP7_75t_L g2035 ( 
.A(n_1987),
.B(n_1921),
.Y(n_2035)
);

OR2x2_ASAP7_75t_L g2036 ( 
.A(n_1968),
.B(n_1928),
.Y(n_2036)
);

INVxp67_ASAP7_75t_L g2037 ( 
.A(n_1999),
.Y(n_2037)
);

AND2x2_ASAP7_75t_L g2038 ( 
.A(n_1987),
.B(n_1921),
.Y(n_2038)
);

INVx1_ASAP7_75t_L g2039 ( 
.A(n_1997),
.Y(n_2039)
);

AND2x2_ASAP7_75t_L g2040 ( 
.A(n_1959),
.B(n_1924),
.Y(n_2040)
);

NAND2xp5_ASAP7_75t_SL g2041 ( 
.A(n_1959),
.B(n_1913),
.Y(n_2041)
);

NAND4xp25_ASAP7_75t_L g2042 ( 
.A(n_1995),
.B(n_1988),
.C(n_1901),
.D(n_1961),
.Y(n_2042)
);

NAND2xp5_ASAP7_75t_L g2043 ( 
.A(n_2026),
.B(n_1967),
.Y(n_2043)
);

AOI221xp5_ASAP7_75t_L g2044 ( 
.A1(n_2006),
.A2(n_1969),
.B1(n_1995),
.B2(n_1982),
.C(n_2001),
.Y(n_2044)
);

NOR4xp25_ASAP7_75t_L g2045 ( 
.A(n_2028),
.B(n_1998),
.C(n_2002),
.D(n_2001),
.Y(n_2045)
);

AOI31xp33_ASAP7_75t_SL g2046 ( 
.A1(n_2037),
.A2(n_1984),
.A3(n_1980),
.B(n_1973),
.Y(n_2046)
);

AOI22xp5_ASAP7_75t_L g2047 ( 
.A1(n_2032),
.A2(n_2042),
.B1(n_2005),
.B2(n_2012),
.Y(n_2047)
);

INVx1_ASAP7_75t_L g2048 ( 
.A(n_2007),
.Y(n_2048)
);

O2A1O1Ixp33_ASAP7_75t_SL g2049 ( 
.A1(n_2012),
.A2(n_1970),
.B(n_1749),
.C(n_1984),
.Y(n_2049)
);

OAI22xp5_ASAP7_75t_L g2050 ( 
.A1(n_2032),
.A2(n_2015),
.B1(n_2027),
.B2(n_1988),
.Y(n_2050)
);

OAI221xp5_ASAP7_75t_L g2051 ( 
.A1(n_2023),
.A2(n_1930),
.B1(n_1971),
.B2(n_1962),
.C(n_1847),
.Y(n_2051)
);

OR2x2_ASAP7_75t_L g2052 ( 
.A(n_2004),
.B(n_1954),
.Y(n_2052)
);

INVx1_ASAP7_75t_L g2053 ( 
.A(n_2007),
.Y(n_2053)
);

INVx1_ASAP7_75t_SL g2054 ( 
.A(n_2004),
.Y(n_2054)
);

NOR3xp33_ASAP7_75t_L g2055 ( 
.A(n_2009),
.B(n_1982),
.C(n_1975),
.Y(n_2055)
);

AOI22xp5_ASAP7_75t_L g2056 ( 
.A1(n_2017),
.A2(n_1884),
.B1(n_1988),
.B2(n_1916),
.Y(n_2056)
);

NAND2x1p5_ASAP7_75t_L g2057 ( 
.A(n_2018),
.B(n_1961),
.Y(n_2057)
);

INVx1_ASAP7_75t_L g2058 ( 
.A(n_2021),
.Y(n_2058)
);

INVx2_ASAP7_75t_L g2059 ( 
.A(n_2020),
.Y(n_2059)
);

OAI32xp33_ASAP7_75t_L g2060 ( 
.A1(n_2009),
.A2(n_1930),
.A3(n_1949),
.B1(n_1830),
.B2(n_1873),
.Y(n_2060)
);

INVx2_ASAP7_75t_L g2061 ( 
.A(n_2020),
.Y(n_2061)
);

HB1xp67_ASAP7_75t_L g2062 ( 
.A(n_2021),
.Y(n_2062)
);

INVx2_ASAP7_75t_L g2063 ( 
.A(n_2033),
.Y(n_2063)
);

AOI222xp33_ASAP7_75t_L g2064 ( 
.A1(n_2023),
.A2(n_1916),
.B1(n_1910),
.B2(n_1911),
.C1(n_1850),
.C2(n_1825),
.Y(n_2064)
);

NAND2xp5_ASAP7_75t_L g2065 ( 
.A(n_2019),
.B(n_1937),
.Y(n_2065)
);

NAND2xp5_ASAP7_75t_L g2066 ( 
.A(n_2019),
.B(n_1937),
.Y(n_2066)
);

INVx1_ASAP7_75t_L g2067 ( 
.A(n_2022),
.Y(n_2067)
);

O2A1O1Ixp33_ASAP7_75t_L g2068 ( 
.A1(n_2016),
.A2(n_1971),
.B(n_1962),
.C(n_1930),
.Y(n_2068)
);

AOI22xp33_ASAP7_75t_L g2069 ( 
.A1(n_2016),
.A2(n_2024),
.B1(n_2025),
.B2(n_2017),
.Y(n_2069)
);

OR2x2_ASAP7_75t_L g2070 ( 
.A(n_2034),
.B(n_1954),
.Y(n_2070)
);

OAI22xp5_ASAP7_75t_L g2071 ( 
.A1(n_2018),
.A2(n_1961),
.B1(n_1930),
.B2(n_1924),
.Y(n_2071)
);

NAND2xp5_ASAP7_75t_SL g2072 ( 
.A(n_2047),
.B(n_2018),
.Y(n_2072)
);

INVx1_ASAP7_75t_L g2073 ( 
.A(n_2062),
.Y(n_2073)
);

INVx1_ASAP7_75t_SL g2074 ( 
.A(n_2054),
.Y(n_2074)
);

INVx2_ASAP7_75t_L g2075 ( 
.A(n_2059),
.Y(n_2075)
);

INVx1_ASAP7_75t_L g2076 ( 
.A(n_2062),
.Y(n_2076)
);

AOI221xp5_ASAP7_75t_L g2077 ( 
.A1(n_2044),
.A2(n_2029),
.B1(n_2030),
.B2(n_2039),
.C(n_2022),
.Y(n_2077)
);

OR2x2_ASAP7_75t_L g2078 ( 
.A(n_2045),
.B(n_2011),
.Y(n_2078)
);

INVx2_ASAP7_75t_L g2079 ( 
.A(n_2059),
.Y(n_2079)
);

INVx1_ASAP7_75t_L g2080 ( 
.A(n_2048),
.Y(n_2080)
);

INVx1_ASAP7_75t_L g2081 ( 
.A(n_2053),
.Y(n_2081)
);

NAND2xp33_ASAP7_75t_SL g2082 ( 
.A(n_2050),
.B(n_2018),
.Y(n_2082)
);

INVx1_ASAP7_75t_SL g2083 ( 
.A(n_2043),
.Y(n_2083)
);

INVx2_ASAP7_75t_L g2084 ( 
.A(n_2061),
.Y(n_2084)
);

INVx1_ASAP7_75t_L g2085 ( 
.A(n_2058),
.Y(n_2085)
);

NOR4xp25_ASAP7_75t_L g2086 ( 
.A(n_2069),
.B(n_2029),
.C(n_2030),
.D(n_2039),
.Y(n_2086)
);

INVx1_ASAP7_75t_L g2087 ( 
.A(n_2067),
.Y(n_2087)
);

OAI221xp5_ASAP7_75t_L g2088 ( 
.A1(n_2069),
.A2(n_2014),
.B1(n_1971),
.B2(n_1962),
.C(n_2011),
.Y(n_2088)
);

INVx1_ASAP7_75t_L g2089 ( 
.A(n_2055),
.Y(n_2089)
);

INVxp67_ASAP7_75t_SL g2090 ( 
.A(n_2057),
.Y(n_2090)
);

INVx1_ASAP7_75t_L g2091 ( 
.A(n_2052),
.Y(n_2091)
);

OAI31xp33_ASAP7_75t_L g2092 ( 
.A1(n_2051),
.A2(n_2014),
.A3(n_2024),
.B(n_2025),
.Y(n_2092)
);

AOI22xp5_ASAP7_75t_L g2093 ( 
.A1(n_2064),
.A2(n_2008),
.B1(n_2013),
.B2(n_2040),
.Y(n_2093)
);

NAND2xp5_ASAP7_75t_L g2094 ( 
.A(n_2063),
.B(n_2033),
.Y(n_2094)
);

NAND2xp5_ASAP7_75t_L g2095 ( 
.A(n_2074),
.B(n_2055),
.Y(n_2095)
);

OAI21xp5_ASAP7_75t_SL g2096 ( 
.A1(n_2077),
.A2(n_2068),
.B(n_2057),
.Y(n_2096)
);

INVxp67_ASAP7_75t_L g2097 ( 
.A(n_2082),
.Y(n_2097)
);

OAI21xp5_ASAP7_75t_SL g2098 ( 
.A1(n_2078),
.A2(n_2014),
.B(n_2046),
.Y(n_2098)
);

OAI22xp5_ASAP7_75t_L g2099 ( 
.A1(n_2078),
.A2(n_2056),
.B1(n_2066),
.B2(n_2065),
.Y(n_2099)
);

OAI32xp33_ASAP7_75t_L g2100 ( 
.A1(n_2082),
.A2(n_2049),
.A3(n_2071),
.B1(n_2070),
.B2(n_2041),
.Y(n_2100)
);

NAND2xp5_ASAP7_75t_L g2101 ( 
.A(n_2083),
.B(n_2035),
.Y(n_2101)
);

AOI22xp33_ASAP7_75t_L g2102 ( 
.A1(n_2089),
.A2(n_2072),
.B1(n_2092),
.B2(n_2088),
.Y(n_2102)
);

INVx1_ASAP7_75t_L g2103 ( 
.A(n_2075),
.Y(n_2103)
);

O2A1O1Ixp33_ASAP7_75t_L g2104 ( 
.A1(n_2086),
.A2(n_2049),
.B(n_2060),
.C(n_2031),
.Y(n_2104)
);

AOI22xp33_ASAP7_75t_L g2105 ( 
.A1(n_2089),
.A2(n_1992),
.B1(n_1837),
.B2(n_2040),
.Y(n_2105)
);

AND2x2_ASAP7_75t_L g2106 ( 
.A(n_2090),
.B(n_2008),
.Y(n_2106)
);

INVxp67_ASAP7_75t_L g2107 ( 
.A(n_2072),
.Y(n_2107)
);

INVx2_ASAP7_75t_L g2108 ( 
.A(n_2075),
.Y(n_2108)
);

AOI221xp5_ASAP7_75t_L g2109 ( 
.A1(n_2076),
.A2(n_2031),
.B1(n_1992),
.B2(n_2036),
.C(n_1866),
.Y(n_2109)
);

AND2x2_ASAP7_75t_L g2110 ( 
.A(n_2106),
.B(n_2091),
.Y(n_2110)
);

NOR4xp75_ASAP7_75t_L g2111 ( 
.A(n_2095),
.B(n_2094),
.C(n_2013),
.D(n_2035),
.Y(n_2111)
);

INVx1_ASAP7_75t_L g2112 ( 
.A(n_2101),
.Y(n_2112)
);

NOR2xp33_ASAP7_75t_L g2113 ( 
.A(n_2107),
.B(n_2079),
.Y(n_2113)
);

NOR4xp25_ASAP7_75t_L g2114 ( 
.A(n_2097),
.B(n_2076),
.C(n_2073),
.D(n_2085),
.Y(n_2114)
);

INVx2_ASAP7_75t_L g2115 ( 
.A(n_2108),
.Y(n_2115)
);

AOI221xp5_ASAP7_75t_L g2116 ( 
.A1(n_2099),
.A2(n_2098),
.B1(n_2104),
.B2(n_2102),
.C(n_2096),
.Y(n_2116)
);

NOR3xp33_ASAP7_75t_SL g2117 ( 
.A(n_2100),
.B(n_2081),
.C(n_2080),
.Y(n_2117)
);

NAND3xp33_ASAP7_75t_L g2118 ( 
.A(n_2103),
.B(n_2087),
.C(n_2079),
.Y(n_2118)
);

NOR2xp33_ASAP7_75t_L g2119 ( 
.A(n_2099),
.B(n_2084),
.Y(n_2119)
);

NOR2x1_ASAP7_75t_L g2120 ( 
.A(n_2109),
.B(n_2084),
.Y(n_2120)
);

XNOR2x1_ASAP7_75t_L g2121 ( 
.A(n_2105),
.B(n_2093),
.Y(n_2121)
);

NAND3xp33_ASAP7_75t_L g2122 ( 
.A(n_2107),
.B(n_2036),
.C(n_2038),
.Y(n_2122)
);

O2A1O1Ixp33_ASAP7_75t_L g2123 ( 
.A1(n_2107),
.A2(n_1971),
.B(n_1962),
.C(n_1952),
.Y(n_2123)
);

NOR2xp33_ASAP7_75t_L g2124 ( 
.A(n_2107),
.B(n_2010),
.Y(n_2124)
);

AOI321xp33_ASAP7_75t_L g2125 ( 
.A1(n_2099),
.A2(n_2010),
.A3(n_2038),
.B1(n_1906),
.B2(n_1936),
.C(n_1944),
.Y(n_2125)
);

AOI221xp5_ASAP7_75t_L g2126 ( 
.A1(n_2119),
.A2(n_2010),
.B1(n_1952),
.B2(n_1885),
.C(n_1886),
.Y(n_2126)
);

AOI21xp5_ASAP7_75t_L g2127 ( 
.A1(n_2116),
.A2(n_2010),
.B(n_1944),
.Y(n_2127)
);

NAND4xp25_ASAP7_75t_L g2128 ( 
.A(n_2124),
.B(n_1952),
.C(n_1949),
.D(n_1944),
.Y(n_2128)
);

O2A1O1Ixp33_ASAP7_75t_L g2129 ( 
.A1(n_2117),
.A2(n_1936),
.B(n_1944),
.C(n_1949),
.Y(n_2129)
);

AOI221xp5_ASAP7_75t_L g2130 ( 
.A1(n_2114),
.A2(n_1886),
.B1(n_1885),
.B2(n_1869),
.C(n_1894),
.Y(n_2130)
);

OAI221xp5_ASAP7_75t_L g2131 ( 
.A1(n_2125),
.A2(n_1902),
.B1(n_1897),
.B2(n_1862),
.C(n_1885),
.Y(n_2131)
);

AOI21xp5_ASAP7_75t_L g2132 ( 
.A1(n_2120),
.A2(n_1936),
.B(n_1955),
.Y(n_2132)
);

INVx1_ASAP7_75t_L g2133 ( 
.A(n_2110),
.Y(n_2133)
);

AOI211xp5_ASAP7_75t_L g2134 ( 
.A1(n_2113),
.A2(n_1936),
.B(n_1753),
.C(n_1929),
.Y(n_2134)
);

AOI221xp5_ASAP7_75t_L g2135 ( 
.A1(n_2118),
.A2(n_1869),
.B1(n_1886),
.B2(n_1894),
.C(n_1897),
.Y(n_2135)
);

OAI22xp33_ASAP7_75t_L g2136 ( 
.A1(n_2131),
.A2(n_2118),
.B1(n_2115),
.B2(n_2112),
.Y(n_2136)
);

AOI21xp5_ASAP7_75t_L g2137 ( 
.A1(n_2129),
.A2(n_2121),
.B(n_2122),
.Y(n_2137)
);

AOI211xp5_ASAP7_75t_L g2138 ( 
.A1(n_2127),
.A2(n_2123),
.B(n_2111),
.C(n_1929),
.Y(n_2138)
);

AO22x2_ASAP7_75t_L g2139 ( 
.A1(n_2133),
.A2(n_2132),
.B1(n_2128),
.B2(n_2134),
.Y(n_2139)
);

OAI221xp5_ASAP7_75t_L g2140 ( 
.A1(n_2126),
.A2(n_1866),
.B1(n_1869),
.B2(n_1894),
.C(n_1897),
.Y(n_2140)
);

NAND5xp2_ASAP7_75t_L g2141 ( 
.A(n_2130),
.B(n_1929),
.C(n_1909),
.D(n_1906),
.E(n_1945),
.Y(n_2141)
);

AOI22xp5_ASAP7_75t_L g2142 ( 
.A1(n_2135),
.A2(n_1900),
.B1(n_1866),
.B2(n_1910),
.Y(n_2142)
);

AOI321xp33_ASAP7_75t_L g2143 ( 
.A1(n_2129),
.A2(n_1911),
.A3(n_1898),
.B1(n_1900),
.B2(n_1826),
.C(n_1861),
.Y(n_2143)
);

NAND3xp33_ASAP7_75t_L g2144 ( 
.A(n_2133),
.B(n_1909),
.C(n_1873),
.Y(n_2144)
);

INVx1_ASAP7_75t_L g2145 ( 
.A(n_2136),
.Y(n_2145)
);

NAND2xp5_ASAP7_75t_L g2146 ( 
.A(n_2137),
.B(n_1955),
.Y(n_2146)
);

INVx1_ASAP7_75t_L g2147 ( 
.A(n_2139),
.Y(n_2147)
);

NAND4xp75_ASAP7_75t_L g2148 ( 
.A(n_2138),
.B(n_1954),
.C(n_1951),
.D(n_1945),
.Y(n_2148)
);

NOR2xp67_ASAP7_75t_L g2149 ( 
.A(n_2144),
.B(n_1873),
.Y(n_2149)
);

NOR2x1_ASAP7_75t_L g2150 ( 
.A(n_2141),
.B(n_2140),
.Y(n_2150)
);

AOI221xp5_ASAP7_75t_L g2151 ( 
.A1(n_2147),
.A2(n_2143),
.B1(n_2142),
.B2(n_1900),
.C(n_1948),
.Y(n_2151)
);

NOR4xp75_ASAP7_75t_L g2152 ( 
.A(n_2146),
.B(n_1873),
.C(n_1871),
.D(n_1951),
.Y(n_2152)
);

OR2x2_ASAP7_75t_L g2153 ( 
.A(n_2145),
.B(n_1956),
.Y(n_2153)
);

NOR3xp33_ASAP7_75t_L g2154 ( 
.A(n_2150),
.B(n_1826),
.C(n_1888),
.Y(n_2154)
);

INVx1_ASAP7_75t_L g2155 ( 
.A(n_2153),
.Y(n_2155)
);

AOI22xp5_ASAP7_75t_L g2156 ( 
.A1(n_2154),
.A2(n_2148),
.B1(n_2149),
.B2(n_1956),
.Y(n_2156)
);

INVx1_ASAP7_75t_L g2157 ( 
.A(n_2155),
.Y(n_2157)
);

AOI221xp5_ASAP7_75t_L g2158 ( 
.A1(n_2157),
.A2(n_2151),
.B1(n_2156),
.B2(n_2152),
.C(n_1948),
.Y(n_2158)
);

OAI22xp5_ASAP7_75t_L g2159 ( 
.A1(n_2157),
.A2(n_1946),
.B1(n_1943),
.B2(n_1934),
.Y(n_2159)
);

OR2x2_ASAP7_75t_L g2160 ( 
.A(n_2159),
.B(n_1928),
.Y(n_2160)
);

XNOR2x1_ASAP7_75t_L g2161 ( 
.A(n_2158),
.B(n_1837),
.Y(n_2161)
);

INVx2_ASAP7_75t_L g2162 ( 
.A(n_2160),
.Y(n_2162)
);

AOI21xp5_ASAP7_75t_L g2163 ( 
.A1(n_2161),
.A2(n_1653),
.B(n_1943),
.Y(n_2163)
);

AOI221xp5_ASAP7_75t_L g2164 ( 
.A1(n_2162),
.A2(n_1946),
.B1(n_1934),
.B2(n_1837),
.C(n_1826),
.Y(n_2164)
);

OAI21xp5_ASAP7_75t_L g2165 ( 
.A1(n_2164),
.A2(n_2163),
.B(n_1871),
.Y(n_2165)
);

INVx1_ASAP7_75t_L g2166 ( 
.A(n_2165),
.Y(n_2166)
);

OAI221xp5_ASAP7_75t_R g2167 ( 
.A1(n_2166),
.A2(n_1653),
.B1(n_1761),
.B2(n_1875),
.C(n_1876),
.Y(n_2167)
);

AOI211xp5_ASAP7_75t_L g2168 ( 
.A1(n_2167),
.A2(n_1837),
.B(n_1653),
.C(n_1728),
.Y(n_2168)
);


endmodule