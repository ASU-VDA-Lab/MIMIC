module fake_jpeg_24097_n_164 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_164);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_164;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx2_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

INVx8_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_9),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_12),
.Y(n_17)
);

INVx6_ASAP7_75t_SL g18 ( 
.A(n_10),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx16f_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx16f_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx16f_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_13),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_9),
.Y(n_30)
);

INVx13_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_31),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_19),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

AOI21xp5_ASAP7_75t_L g33 ( 
.A1(n_14),
.A2(n_0),
.B(n_1),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_33),
.B(n_29),
.C(n_25),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

BUFx2_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_16),
.B(n_0),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_35),
.B(n_36),
.Y(n_48)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

NAND3xp33_ASAP7_75t_L g37 ( 
.A(n_29),
.B(n_10),
.C(n_8),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_42),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

BUFx2_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_16),
.B(n_0),
.Y(n_39)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

HAxp5_ASAP7_75t_SL g53 ( 
.A(n_40),
.B(n_41),
.CON(n_53),
.SN(n_53)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_25),
.B(n_1),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

BUFx10_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

CKINVDCx14_ASAP7_75t_R g72 ( 
.A(n_45),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_42),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_46),
.B(n_50),
.Y(n_90)
);

INVx13_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_51),
.Y(n_79)
);

OR2x2_ASAP7_75t_L g54 ( 
.A(n_31),
.B(n_30),
.Y(n_54)
);

NAND3xp33_ASAP7_75t_L g83 ( 
.A(n_54),
.B(n_58),
.C(n_47),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_SL g76 ( 
.A1(n_55),
.A2(n_62),
.B(n_17),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_33),
.A2(n_14),
.B1(n_20),
.B2(n_15),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_56),
.A2(n_57),
.B1(n_59),
.B2(n_64),
.Y(n_74)
);

OAI32xp33_ASAP7_75t_L g57 ( 
.A1(n_38),
.A2(n_23),
.A3(n_18),
.B1(n_20),
.B2(n_24),
.Y(n_57)
);

AND2x6_ASAP7_75t_L g58 ( 
.A(n_41),
.B(n_2),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_40),
.A2(n_15),
.B1(n_21),
.B2(n_32),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_44),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_61),
.B(n_3),
.Y(n_78)
);

O2A1O1Ixp33_ASAP7_75t_SL g62 ( 
.A1(n_43),
.A2(n_24),
.B(n_23),
.C(n_26),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_36),
.A2(n_21),
.B1(n_28),
.B2(n_30),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g91 ( 
.A(n_65),
.Y(n_91)
);

OA22x2_ASAP7_75t_L g69 ( 
.A1(n_31),
.A2(n_23),
.B1(n_28),
.B2(n_17),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_69),
.A2(n_18),
.B1(n_27),
.B2(n_22),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_53),
.B(n_2),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_70),
.B(n_4),
.C(n_7),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_54),
.B(n_27),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_71),
.B(n_75),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_65),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_73),
.B(n_76),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_48),
.B(n_27),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_69),
.B(n_27),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_77),
.B(n_82),
.Y(n_95)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_78),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_80),
.B(n_52),
.Y(n_111)
);

NOR2x1_ASAP7_75t_L g81 ( 
.A(n_47),
.B(n_18),
.Y(n_81)
);

OR2x2_ASAP7_75t_L g98 ( 
.A(n_81),
.B(n_63),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_69),
.B(n_22),
.Y(n_82)
);

NOR3xp33_ASAP7_75t_L g100 ( 
.A(n_83),
.B(n_6),
.C(n_7),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_62),
.B(n_22),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_84),
.B(n_70),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_53),
.A2(n_22),
.B(n_26),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_85),
.A2(n_87),
.B(n_26),
.Y(n_103)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_49),
.Y(n_86)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_86),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_58),
.A2(n_26),
.B(n_5),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_68),
.B(n_4),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_88),
.B(n_92),
.Y(n_107)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_50),
.Y(n_89)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_89),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_59),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_91),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_93),
.B(n_100),
.Y(n_117)
);

AND2x6_ASAP7_75t_L g96 ( 
.A(n_81),
.B(n_6),
.Y(n_96)
);

BUFx12_ASAP7_75t_L g126 ( 
.A(n_96),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_98),
.B(n_106),
.Y(n_123)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_90),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_102),
.B(n_111),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_103),
.A2(n_108),
.B(n_73),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_85),
.B(n_45),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_104),
.B(n_77),
.C(n_76),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_71),
.B(n_45),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_109),
.B(n_70),
.Y(n_114)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_91),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_110),
.B(n_66),
.Y(n_124)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_109),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_113),
.B(n_114),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_97),
.A2(n_87),
.B1(n_84),
.B2(n_82),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_115),
.A2(n_95),
.B1(n_103),
.B2(n_101),
.Y(n_127)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_94),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_116),
.B(n_118),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_94),
.B(n_108),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_119),
.B(n_74),
.C(n_106),
.Y(n_130)
);

OA21x2_ASAP7_75t_SL g120 ( 
.A1(n_104),
.A2(n_75),
.B(n_80),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_120),
.A2(n_122),
.B(n_98),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_107),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_121),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_124),
.A2(n_125),
.B(n_92),
.Y(n_135)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_111),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_127),
.A2(n_120),
.B1(n_118),
.B2(n_114),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_125),
.B(n_112),
.C(n_113),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_128),
.B(n_129),
.C(n_130),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_119),
.B(n_95),
.C(n_102),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_131),
.B(n_133),
.C(n_123),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_122),
.B(n_74),
.C(n_101),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_135),
.B(n_137),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_115),
.A2(n_96),
.B(n_89),
.Y(n_137)
);

HB1xp67_ASAP7_75t_L g139 ( 
.A(n_132),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_139),
.A2(n_99),
.B1(n_105),
.B2(n_86),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_132),
.B(n_116),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_140),
.A2(n_141),
.B(n_144),
.Y(n_147)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_136),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_143),
.B(n_145),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_134),
.B(n_121),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_128),
.B(n_117),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_146),
.B(n_123),
.Y(n_151)
);

NAND3xp33_ASAP7_75t_L g149 ( 
.A(n_138),
.B(n_126),
.C(n_129),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_149),
.A2(n_150),
.B(n_126),
.Y(n_156)
);

XOR2x1_ASAP7_75t_SL g150 ( 
.A(n_146),
.B(n_126),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_151),
.B(n_148),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_152),
.A2(n_79),
.B1(n_72),
.B2(n_67),
.Y(n_157)
);

AO21x1_ASAP7_75t_L g158 ( 
.A1(n_153),
.A2(n_154),
.B(n_156),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_147),
.B(n_142),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_149),
.A2(n_126),
.B1(n_142),
.B2(n_66),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_155),
.B(n_157),
.Y(n_160)
);

NOR2xp67_ASAP7_75t_SL g159 ( 
.A(n_155),
.B(n_60),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_159),
.A2(n_60),
.B(n_52),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_160),
.B(n_49),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_161),
.B(n_162),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_163),
.B(n_158),
.Y(n_164)
);


endmodule