module fake_jpeg_28071_n_264 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_264);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_264;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_14;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_11;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

BUFx5_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

CKINVDCx16_ASAP7_75t_R g15 ( 
.A(n_4),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx2_ASAP7_75t_SL g20 ( 
.A(n_6),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_18),
.Y(n_24)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_21),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_25),
.B(n_34),
.Y(n_38)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

INVx2_ASAP7_75t_SL g43 ( 
.A(n_28),
.Y(n_43)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_30),
.B(n_33),
.Y(n_41)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

INVxp67_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

OAI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_31),
.A2(n_20),
.B1(n_21),
.B2(n_22),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_36),
.A2(n_32),
.B1(n_34),
.B2(n_29),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_39),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_45),
.B(n_48),
.Y(n_62)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_47),
.Y(n_78)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_49),
.Y(n_61)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_50),
.B(n_59),
.Y(n_74)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_51),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

BUFx12_ASAP7_75t_L g77 ( 
.A(n_52),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_39),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_53),
.Y(n_67)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_54),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_38),
.A2(n_34),
.B1(n_32),
.B2(n_31),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_55),
.A2(n_40),
.B1(n_35),
.B2(n_44),
.Y(n_72)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_56),
.Y(n_75)
);

HB1xp67_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_57),
.Y(n_76)
);

INVx3_ASAP7_75t_SL g58 ( 
.A(n_37),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_58),
.B(n_60),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

O2A1O1Ixp33_ASAP7_75t_SL g65 ( 
.A1(n_50),
.A2(n_60),
.B(n_41),
.C(n_36),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_65),
.A2(n_26),
.B1(n_28),
.B2(n_24),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g68 ( 
.A1(n_45),
.A2(n_38),
.B(n_41),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_68),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_48),
.A2(n_30),
.B1(n_29),
.B2(n_40),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_70),
.A2(n_72),
.B1(n_73),
.B2(n_41),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_L g71 ( 
.A1(n_51),
.A2(n_41),
.B(n_25),
.Y(n_71)
);

CKINVDCx14_ASAP7_75t_R g90 ( 
.A(n_71),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_46),
.A2(n_40),
.B1(n_41),
.B2(n_27),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_74),
.B(n_52),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_79),
.B(n_80),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_67),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_81),
.A2(n_86),
.B1(n_92),
.B2(n_66),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_74),
.B(n_53),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_82),
.B(n_83),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_71),
.B(n_56),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_62),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_84),
.B(n_88),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_65),
.A2(n_49),
.B1(n_58),
.B2(n_20),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_85),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_63),
.A2(n_58),
.B1(n_54),
.B2(n_47),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_67),
.B(n_59),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_65),
.A2(n_24),
.B1(n_28),
.B2(n_27),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_89),
.A2(n_91),
.B1(n_37),
.B2(n_43),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_63),
.A2(n_37),
.B1(n_43),
.B2(n_33),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_73),
.B(n_33),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_93),
.A2(n_65),
.B(n_66),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_76),
.B(n_59),
.Y(n_94)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_94),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_68),
.B(n_14),
.Y(n_95)
);

OAI32xp33_ASAP7_75t_L g109 ( 
.A1(n_95),
.A2(n_12),
.A3(n_75),
.B1(n_69),
.B2(n_14),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_80),
.B(n_61),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_96),
.B(n_100),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_90),
.B(n_62),
.C(n_61),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_97),
.B(n_116),
.C(n_103),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_83),
.B(n_72),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_99),
.A2(n_102),
.B(n_103),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_88),
.B(n_76),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_85),
.B(n_82),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_85),
.B(n_70),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_105),
.A2(n_114),
.B(n_118),
.Y(n_135)
);

NOR2x1p5_ASAP7_75t_L g106 ( 
.A(n_91),
.B(n_90),
.Y(n_106)
);

OR2x2_ASAP7_75t_L g131 ( 
.A(n_106),
.B(n_112),
.Y(n_131)
);

NAND3xp33_ASAP7_75t_L g107 ( 
.A(n_95),
.B(n_6),
.C(n_10),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_107),
.B(n_111),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_108),
.A2(n_113),
.B1(n_93),
.B2(n_91),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_109),
.B(n_118),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_110),
.A2(n_81),
.B1(n_86),
.B2(n_92),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_94),
.Y(n_111)
);

OR2x2_ASAP7_75t_L g112 ( 
.A(n_89),
.B(n_17),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_81),
.A2(n_64),
.B1(n_75),
.B2(n_69),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_87),
.A2(n_12),
.B(n_15),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_84),
.B(n_77),
.C(n_78),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_79),
.A2(n_15),
.B(n_13),
.Y(n_118)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_101),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_120),
.B(n_121),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_122),
.A2(n_127),
.B1(n_77),
.B2(n_20),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_123),
.B(n_129),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_116),
.B(n_86),
.Y(n_125)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_125),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_126),
.A2(n_43),
.B1(n_33),
.B2(n_77),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_102),
.A2(n_92),
.B1(n_93),
.B2(n_64),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_117),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_128),
.B(n_133),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_97),
.B(n_93),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_98),
.B(n_103),
.C(n_106),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_130),
.B(n_123),
.C(n_129),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_110),
.A2(n_104),
.B1(n_106),
.B2(n_98),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_132),
.A2(n_143),
.B1(n_140),
.B2(n_134),
.Y(n_151)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_113),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_108),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_134),
.B(n_138),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_111),
.B(n_78),
.Y(n_136)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_136),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_115),
.B(n_64),
.Y(n_137)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_137),
.Y(n_158)
);

INVx1_ASAP7_75t_SL g138 ( 
.A(n_99),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_99),
.B(n_105),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_139),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_105),
.B(n_78),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_140),
.Y(n_168)
);

MAJx2_ASAP7_75t_L g141 ( 
.A(n_104),
.B(n_109),
.C(n_114),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_SL g161 ( 
.A(n_141),
.B(n_13),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_112),
.B(n_17),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_142),
.B(n_77),
.Y(n_164)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_96),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_96),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_144),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_96),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_146),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_149),
.A2(n_145),
.B1(n_19),
.B2(n_11),
.Y(n_183)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_151),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_152),
.B(n_161),
.Y(n_175)
);

NOR2xp67_ASAP7_75t_L g153 ( 
.A(n_121),
.B(n_22),
.Y(n_153)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_153),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_130),
.B(n_119),
.C(n_133),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_157),
.B(n_159),
.C(n_135),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_119),
.B(n_126),
.C(n_127),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_160),
.A2(n_23),
.B1(n_19),
.B2(n_7),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_164),
.B(n_142),
.Y(n_182)
);

OA21x2_ASAP7_75t_L g165 ( 
.A1(n_139),
.A2(n_77),
.B(n_23),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_165),
.A2(n_131),
.B(n_138),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_124),
.B(n_17),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_166),
.B(n_169),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_136),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_167),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_135),
.B(n_23),
.Y(n_169)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_155),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_173),
.B(n_174),
.Y(n_196)
);

BUFx12_ASAP7_75t_L g174 ( 
.A(n_162),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_177),
.B(n_188),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_154),
.B(n_144),
.Y(n_179)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_179),
.Y(n_194)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_180),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_163),
.A2(n_131),
.B(n_141),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_181),
.A2(n_184),
.B(n_185),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_SL g201 ( 
.A(n_182),
.B(n_178),
.Y(n_201)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_183),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_163),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_155),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g193 ( 
.A(n_186),
.B(n_189),
.Y(n_193)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_149),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_187),
.B(n_159),
.C(n_147),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_152),
.B(n_19),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_154),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_188),
.B(n_150),
.C(n_157),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_190),
.B(n_197),
.C(n_198),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_191),
.A2(n_156),
.B1(n_183),
.B2(n_160),
.Y(n_218)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_174),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_192),
.B(n_195),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_177),
.B(n_158),
.C(n_148),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_175),
.B(n_150),
.C(n_147),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_175),
.B(n_166),
.C(n_161),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_174),
.B(n_164),
.C(n_170),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_200),
.B(n_205),
.C(n_179),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_201),
.B(n_206),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_171),
.B(n_178),
.C(n_181),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_182),
.B(n_169),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_202),
.A2(n_193),
.B1(n_184),
.B2(n_203),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_208),
.A2(n_213),
.B1(n_165),
.B2(n_201),
.Y(n_222)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_193),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_209),
.B(n_215),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_199),
.B(n_190),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_210),
.B(n_212),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_194),
.A2(n_176),
.B1(n_172),
.B2(n_186),
.Y(n_213)
);

XOR2x2_ASAP7_75t_SL g214 ( 
.A(n_204),
.B(n_180),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_214),
.B(n_216),
.Y(n_231)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_196),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_192),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_199),
.B(n_170),
.C(n_168),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_217),
.B(n_165),
.C(n_5),
.Y(n_223)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_218),
.Y(n_225)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_206),
.Y(n_220)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_220),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_207),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_221),
.Y(n_234)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_222),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_223),
.B(n_227),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_214),
.A2(n_5),
.B1(n_9),
.B2(n_8),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_224),
.A2(n_10),
.B1(n_4),
.B2(n_3),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_208),
.A2(n_5),
.B(n_9),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_210),
.B(n_0),
.C(n_1),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_228),
.B(n_211),
.C(n_219),
.Y(n_238)
);

AND2x2_ASAP7_75t_L g232 ( 
.A(n_231),
.B(n_217),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_232),
.B(n_237),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_229),
.B(n_219),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_235),
.B(n_223),
.C(n_226),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_228),
.B(n_212),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_236),
.B(n_226),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_229),
.B(n_211),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_238),
.B(n_235),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_240),
.B(n_227),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_242),
.B(n_245),
.Y(n_253)
);

AND2x6_ASAP7_75t_L g243 ( 
.A(n_234),
.B(n_232),
.Y(n_243)
);

NOR2xp67_ASAP7_75t_L g249 ( 
.A(n_243),
.B(n_239),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_244),
.B(n_246),
.C(n_248),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_238),
.B(n_230),
.C(n_225),
.Y(n_245)
);

XNOR2x2_ASAP7_75t_SL g247 ( 
.A(n_233),
.B(n_4),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_247),
.A2(n_241),
.B1(n_7),
.B2(n_3),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_249),
.A2(n_251),
.B(n_8),
.Y(n_256)
);

NOR2xp67_ASAP7_75t_L g251 ( 
.A(n_241),
.B(n_7),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_252),
.B(n_3),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_253),
.B(n_3),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_254),
.A2(n_255),
.B(n_8),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_256),
.B(n_250),
.C(n_8),
.Y(n_258)
);

OAI31xp33_ASAP7_75t_SL g259 ( 
.A1(n_257),
.A2(n_258),
.A3(n_9),
.B(n_10),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_259),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_260),
.B(n_250),
.Y(n_261)
);

A2O1A1Ixp33_ASAP7_75t_L g262 ( 
.A1(n_261),
.A2(n_10),
.B(n_1),
.C(n_2),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_262),
.B(n_0),
.Y(n_263)
);

AO21x1_ASAP7_75t_L g264 ( 
.A1(n_263),
.A2(n_0),
.B(n_1),
.Y(n_264)
);


endmodule