module fake_jpeg_13777_n_527 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_527);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_527;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_15),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_13),
.B(n_6),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx24_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

INVx2_ASAP7_75t_SL g32 ( 
.A(n_7),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

INVx2_ASAP7_75t_SL g36 ( 
.A(n_8),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_8),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_4),
.B(n_14),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_5),
.Y(n_43)
);

BUFx16f_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_10),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_1),
.Y(n_46)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_5),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_10),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_13),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_9),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_9),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_16),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_52),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_42),
.B(n_14),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_53),
.B(n_68),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_16),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_54),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_16),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_55),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_18),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_56),
.Y(n_134)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_17),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g149 ( 
.A(n_57),
.Y(n_149)
);

INVx2_ASAP7_75t_SL g58 ( 
.A(n_31),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g148 ( 
.A(n_58),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_18),
.Y(n_59)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_59),
.Y(n_119)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_30),
.Y(n_60)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_60),
.Y(n_105)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_61),
.Y(n_106)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_30),
.Y(n_62)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_62),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_18),
.Y(n_63)
);

INVx8_ASAP7_75t_L g133 ( 
.A(n_63),
.Y(n_133)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_24),
.Y(n_64)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_64),
.Y(n_121)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_65),
.Y(n_116)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_22),
.Y(n_66)
);

INVx3_ASAP7_75t_SL g139 ( 
.A(n_66),
.Y(n_139)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_17),
.Y(n_67)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_67),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_42),
.B(n_14),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_22),
.Y(n_69)
);

INVx8_ASAP7_75t_L g140 ( 
.A(n_69),
.Y(n_140)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_22),
.Y(n_70)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_70),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_23),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g156 ( 
.A(n_71),
.Y(n_156)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_31),
.Y(n_72)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_72),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_23),
.Y(n_73)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_73),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_25),
.B(n_0),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_74),
.B(n_76),
.Y(n_142)
);

BUFx10_ASAP7_75t_L g75 ( 
.A(n_31),
.Y(n_75)
);

INVx4_ASAP7_75t_SL g132 ( 
.A(n_75),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_25),
.B(n_0),
.Y(n_76)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_20),
.Y(n_77)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_77),
.Y(n_147)
);

INVx11_ASAP7_75t_L g78 ( 
.A(n_31),
.Y(n_78)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_78),
.Y(n_129)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_51),
.Y(n_79)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_79),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_19),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_80),
.B(n_87),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_19),
.B(n_0),
.Y(n_81)
);

OR2x2_ASAP7_75t_L g103 ( 
.A(n_81),
.B(n_28),
.Y(n_103)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_51),
.Y(n_82)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_82),
.Y(n_137)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_44),
.Y(n_83)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_83),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_26),
.B(n_0),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_84),
.B(n_101),
.Y(n_111)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_35),
.Y(n_85)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_85),
.Y(n_138)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_35),
.Y(n_86)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_86),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_21),
.B(n_12),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_23),
.Y(n_88)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_88),
.Y(n_145)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_20),
.Y(n_89)
);

BUFx4f_ASAP7_75t_L g115 ( 
.A(n_89),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_21),
.B(n_50),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_90),
.B(n_95),
.Y(n_114)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_44),
.Y(n_91)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_91),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_34),
.Y(n_92)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_92),
.Y(n_150)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_44),
.Y(n_93)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_93),
.Y(n_152)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_35),
.Y(n_94)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_94),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_24),
.B(n_1),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_24),
.Y(n_96)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_96),
.Y(n_124)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_47),
.Y(n_97)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_97),
.Y(n_154)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_41),
.Y(n_98)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_98),
.Y(n_155)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_26),
.Y(n_99)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_99),
.Y(n_161)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_41),
.Y(n_100)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_100),
.Y(n_128)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_47),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_32),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_102),
.A2(n_36),
.B1(n_32),
.B2(n_38),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_103),
.B(n_104),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_72),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_66),
.A2(n_36),
.B1(n_32),
.B2(n_47),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_107),
.A2(n_144),
.B1(n_102),
.B2(n_89),
.Y(n_172)
);

OR2x2_ASAP7_75t_L g108 ( 
.A(n_75),
.B(n_26),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_108),
.B(n_151),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_83),
.B(n_91),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_117),
.B(n_141),
.Y(n_182)
);

BUFx12_ASAP7_75t_L g123 ( 
.A(n_75),
.Y(n_123)
);

INVx6_ASAP7_75t_SL g200 ( 
.A(n_123),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_93),
.B(n_50),
.Y(n_127)
);

OR2x2_ASAP7_75t_L g186 ( 
.A(n_127),
.B(n_130),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_97),
.B(n_43),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_131),
.A2(n_157),
.B1(n_48),
.B2(n_39),
.Y(n_163)
);

INVx4_ASAP7_75t_SL g141 ( 
.A(n_78),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_58),
.A2(n_36),
.B1(n_34),
.B2(n_41),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_98),
.Y(n_151)
);

OAI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_52),
.A2(n_49),
.B1(n_40),
.B2(n_39),
.Y(n_157)
);

INVx4_ASAP7_75t_SL g158 ( 
.A(n_92),
.Y(n_158)
);

INVx4_ASAP7_75t_L g183 ( 
.A(n_158),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_100),
.B(n_48),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_159),
.B(n_48),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_70),
.B(n_43),
.Y(n_160)
);

OR2x2_ASAP7_75t_L g190 ( 
.A(n_160),
.B(n_49),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_163),
.A2(n_184),
.B1(n_144),
.B2(n_126),
.Y(n_216)
);

HB1xp67_ASAP7_75t_L g164 ( 
.A(n_128),
.Y(n_164)
);

INVx1_ASAP7_75t_SL g247 ( 
.A(n_164),
.Y(n_247)
);

BUFx3_ASAP7_75t_L g165 ( 
.A(n_149),
.Y(n_165)
);

BUFx3_ASAP7_75t_L g243 ( 
.A(n_165),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_114),
.B(n_37),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_166),
.B(n_170),
.Y(n_218)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_115),
.Y(n_167)
);

INVx4_ASAP7_75t_L g233 ( 
.A(n_167),
.Y(n_233)
);

INVx2_ASAP7_75t_SL g168 ( 
.A(n_117),
.Y(n_168)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_168),
.Y(n_220)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_105),
.Y(n_169)
);

INVx2_ASAP7_75t_SL g249 ( 
.A(n_169),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_111),
.B(n_37),
.Y(n_170)
);

INVx1_ASAP7_75t_SL g171 ( 
.A(n_148),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_171),
.B(n_180),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_172),
.A2(n_189),
.B1(n_192),
.B2(n_122),
.Y(n_239)
);

INVx11_ASAP7_75t_L g173 ( 
.A(n_141),
.Y(n_173)
);

INVx8_ASAP7_75t_L g227 ( 
.A(n_173),
.Y(n_227)
);

BUFx3_ASAP7_75t_L g174 ( 
.A(n_149),
.Y(n_174)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_174),
.Y(n_229)
);

INVx6_ASAP7_75t_L g176 ( 
.A(n_118),
.Y(n_176)
);

INVx8_ASAP7_75t_L g234 ( 
.A(n_176),
.Y(n_234)
);

INVx8_ASAP7_75t_L g177 ( 
.A(n_118),
.Y(n_177)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_177),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_159),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_178),
.B(n_190),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_147),
.A2(n_34),
.B1(n_77),
.B2(n_67),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_181),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_L g184 ( 
.A1(n_111),
.A2(n_88),
.B1(n_73),
.B2(n_71),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_110),
.A2(n_40),
.B1(n_28),
.B2(n_33),
.Y(n_185)
);

CKINVDCx16_ASAP7_75t_R g240 ( 
.A(n_185),
.Y(n_240)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_112),
.Y(n_187)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_187),
.Y(n_221)
);

INVx5_ASAP7_75t_L g188 ( 
.A(n_133),
.Y(n_188)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_188),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_142),
.A2(n_69),
.B1(n_63),
.B2(n_59),
.Y(n_189)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_135),
.Y(n_191)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_191),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_142),
.A2(n_56),
.B1(n_55),
.B2(n_54),
.Y(n_192)
);

INVx6_ASAP7_75t_L g193 ( 
.A(n_120),
.Y(n_193)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_193),
.Y(n_245)
);

INVx5_ASAP7_75t_L g194 ( 
.A(n_133),
.Y(n_194)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_194),
.Y(n_246)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_155),
.Y(n_195)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_195),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_103),
.B(n_49),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_196),
.B(n_212),
.Y(n_244)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_139),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g231 ( 
.A(n_197),
.B(n_199),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_113),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_198),
.B(n_206),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_121),
.B(n_38),
.C(n_33),
.Y(n_199)
);

INVx8_ASAP7_75t_L g201 ( 
.A(n_120),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_201),
.B(n_205),
.Y(n_241)
);

OA22x2_ASAP7_75t_L g202 ( 
.A1(n_107),
.A2(n_29),
.B1(n_46),
.B2(n_45),
.Y(n_202)
);

OAI32xp33_ASAP7_75t_L g251 ( 
.A1(n_202),
.A2(n_129),
.A3(n_140),
.B1(n_134),
.B2(n_125),
.Y(n_251)
);

HAxp5_ASAP7_75t_SL g203 ( 
.A(n_108),
.B(n_48),
.CON(n_203),
.SN(n_203)
);

CKINVDCx14_ASAP7_75t_R g235 ( 
.A(n_203),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_139),
.A2(n_29),
.B1(n_48),
.B2(n_45),
.Y(n_204)
);

CKINVDCx16_ASAP7_75t_R g248 ( 
.A(n_204),
.Y(n_248)
);

INVx4_ASAP7_75t_L g205 ( 
.A(n_158),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_124),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_145),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_207),
.B(n_210),
.Y(n_225)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_138),
.Y(n_208)
);

OR2x2_ASAP7_75t_L g215 ( 
.A(n_208),
.B(n_211),
.Y(n_215)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_115),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_209),
.Y(n_214)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_146),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_143),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_149),
.A2(n_46),
.B1(n_27),
.B2(n_4),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_150),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_213),
.B(n_137),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_216),
.A2(n_238),
.B1(n_168),
.B2(n_182),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_173),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_223),
.B(n_242),
.Y(n_256)
);

A2O1A1Ixp33_ASAP7_75t_L g228 ( 
.A1(n_186),
.A2(n_109),
.B(n_157),
.C(n_132),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_228),
.B(n_230),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_186),
.B(n_153),
.Y(n_230)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_236),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_170),
.B(n_109),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_237),
.B(n_251),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_163),
.A2(n_136),
.B1(n_116),
.B2(n_119),
.Y(n_238)
);

OAI22xp33_ASAP7_75t_SL g271 ( 
.A1(n_239),
.A2(n_202),
.B1(n_199),
.B2(n_134),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_200),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_200),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_252),
.B(n_171),
.Y(n_264)
);

INVx2_ASAP7_75t_SL g254 ( 
.A(n_245),
.Y(n_254)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_254),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_255),
.A2(n_208),
.B1(n_161),
.B2(n_197),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_244),
.A2(n_168),
.B(n_182),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_257),
.A2(n_275),
.B(n_205),
.Y(n_311)
);

AND2x6_ASAP7_75t_L g258 ( 
.A(n_228),
.B(n_203),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_258),
.B(n_260),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_218),
.B(n_166),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_259),
.B(n_288),
.Y(n_312)
);

AND2x6_ASAP7_75t_L g260 ( 
.A(n_235),
.B(n_190),
.Y(n_260)
);

NAND2x1_ASAP7_75t_SL g261 ( 
.A(n_220),
.B(n_182),
.Y(n_261)
);

INVx1_ASAP7_75t_SL g315 ( 
.A(n_261),
.Y(n_315)
);

INVx3_ASAP7_75t_L g262 ( 
.A(n_232),
.Y(n_262)
);

INVx1_ASAP7_75t_SL g320 ( 
.A(n_262),
.Y(n_320)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_234),
.Y(n_263)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_263),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_264),
.B(n_266),
.Y(n_297)
);

INVx3_ASAP7_75t_L g265 ( 
.A(n_232),
.Y(n_265)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_265),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_219),
.B(n_175),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_225),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_267),
.B(n_268),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_237),
.B(n_187),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_271),
.A2(n_216),
.B1(n_231),
.B2(n_238),
.Y(n_296)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_221),
.Y(n_272)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_272),
.Y(n_305)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_221),
.Y(n_273)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_273),
.Y(n_323)
);

INVx13_ASAP7_75t_L g274 ( 
.A(n_242),
.Y(n_274)
);

CKINVDCx14_ASAP7_75t_R g304 ( 
.A(n_274),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_244),
.A2(n_179),
.B(n_183),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_250),
.Y(n_276)
);

AND2x2_ASAP7_75t_L g322 ( 
.A(n_276),
.B(n_280),
.Y(n_322)
);

CKINVDCx16_ASAP7_75t_R g277 ( 
.A(n_241),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_277),
.B(n_281),
.Y(n_313)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_250),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_278),
.B(n_283),
.Y(n_300)
);

AND2x2_ASAP7_75t_L g280 ( 
.A(n_220),
.B(n_202),
.Y(n_280)
);

CKINVDCx16_ASAP7_75t_R g281 ( 
.A(n_241),
.Y(n_281)
);

INVx13_ASAP7_75t_L g282 ( 
.A(n_252),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g307 ( 
.A(n_282),
.Y(n_307)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_249),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_249),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_284),
.B(n_285),
.Y(n_314)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_249),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_SL g286 ( 
.A1(n_222),
.A2(n_215),
.B(n_230),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_286),
.A2(n_247),
.B(n_202),
.Y(n_319)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_215),
.Y(n_287)
);

AOI22xp33_ASAP7_75t_SL g301 ( 
.A1(n_287),
.A2(n_289),
.B1(n_227),
.B2(n_183),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_218),
.B(n_211),
.Y(n_288)
);

INVx3_ASAP7_75t_SL g289 ( 
.A(n_227),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_279),
.A2(n_239),
.B1(n_217),
.B2(n_248),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_291),
.A2(n_295),
.B1(n_310),
.B2(n_321),
.Y(n_356)
);

OAI21xp5_ASAP7_75t_L g294 ( 
.A1(n_269),
.A2(n_222),
.B(n_215),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_L g333 ( 
.A1(n_294),
.A2(n_303),
.B(n_261),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_279),
.A2(n_217),
.B1(n_248),
.B2(n_240),
.Y(n_295)
);

AO21x1_ASAP7_75t_L g345 ( 
.A1(n_296),
.A2(n_285),
.B(n_284),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_280),
.A2(n_240),
.B1(n_251),
.B2(n_231),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_298),
.B(n_306),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_280),
.A2(n_226),
.B1(n_231),
.B2(n_246),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_SL g344 ( 
.A1(n_299),
.A2(n_311),
.B(n_317),
.Y(n_344)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_301),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_L g303 ( 
.A1(n_269),
.A2(n_226),
.B(n_223),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_287),
.A2(n_226),
.B1(n_245),
.B2(n_246),
.Y(n_306)
);

CKINVDCx16_ASAP7_75t_R g309 ( 
.A(n_256),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_309),
.B(n_272),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_288),
.B(n_247),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_316),
.B(n_259),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_270),
.A2(n_253),
.B1(n_229),
.B2(n_214),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_270),
.A2(n_234),
.B1(n_253),
.B2(n_214),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_318),
.B(n_324),
.Y(n_338)
);

A2O1A1Ixp33_ASAP7_75t_L g340 ( 
.A1(n_319),
.A2(n_260),
.B(n_282),
.C(n_274),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_L g321 ( 
.A1(n_255),
.A2(n_193),
.B1(n_176),
.B2(n_201),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_286),
.A2(n_119),
.B1(n_125),
.B2(n_140),
.Y(n_324)
);

CKINVDCx14_ASAP7_75t_R g325 ( 
.A(n_308),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_325),
.Y(n_386)
);

INVxp33_ASAP7_75t_L g326 ( 
.A(n_297),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_326),
.B(n_346),
.Y(n_360)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_300),
.Y(n_328)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_328),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_314),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_329),
.B(n_350),
.Y(n_369)
);

AOI21xp5_ASAP7_75t_L g330 ( 
.A1(n_315),
.A2(n_257),
.B(n_275),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_SL g362 ( 
.A1(n_330),
.A2(n_340),
.B(n_311),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_331),
.B(n_335),
.C(n_355),
.Y(n_366)
);

INVx8_ASAP7_75t_L g332 ( 
.A(n_304),
.Y(n_332)
);

INVxp67_ASAP7_75t_L g368 ( 
.A(n_332),
.Y(n_368)
);

XNOR2x2_ASAP7_75t_SL g378 ( 
.A(n_333),
.B(n_323),
.Y(n_378)
);

AND2x2_ASAP7_75t_L g334 ( 
.A(n_315),
.B(n_278),
.Y(n_334)
);

INVxp67_ASAP7_75t_L g373 ( 
.A(n_334),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_312),
.B(n_258),
.Y(n_335)
);

AOI22xp33_ASAP7_75t_SL g337 ( 
.A1(n_295),
.A2(n_289),
.B1(n_262),
.B2(n_265),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_L g370 ( 
.A1(n_337),
.A2(n_324),
.B(n_319),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_313),
.B(n_243),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_339),
.B(n_342),
.Y(n_381)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_305),
.Y(n_341)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_341),
.Y(n_375)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_300),
.Y(n_343)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_343),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_345),
.A2(n_298),
.B1(n_299),
.B2(n_296),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_SL g346 ( 
.A(n_292),
.B(n_276),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_312),
.B(n_243),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_347),
.B(n_349),
.Y(n_367)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_314),
.Y(n_348)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_348),
.Y(n_385)
);

INVx4_ASAP7_75t_L g349 ( 
.A(n_290),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_305),
.Y(n_350)
);

INVx13_ASAP7_75t_L g351 ( 
.A(n_307),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_351),
.Y(n_363)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_323),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_352),
.B(n_353),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_307),
.B(n_322),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_322),
.B(n_254),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_354),
.B(n_357),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_294),
.B(n_283),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_322),
.B(n_254),
.Y(n_357)
);

CKINVDCx16_ASAP7_75t_R g358 ( 
.A(n_317),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_358),
.B(n_306),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_336),
.A2(n_291),
.B1(n_303),
.B2(n_321),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_L g396 ( 
.A1(n_359),
.A2(n_370),
.B1(n_376),
.B2(n_379),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g392 ( 
.A1(n_361),
.A2(n_391),
.B1(n_334),
.B2(n_338),
.Y(n_392)
);

AOI21x1_ASAP7_75t_SL g394 ( 
.A1(n_362),
.A2(n_384),
.B(n_344),
.Y(n_394)
);

XOR2x1_ASAP7_75t_L g364 ( 
.A(n_355),
.B(n_316),
.Y(n_364)
);

XNOR2x1_ASAP7_75t_L g409 ( 
.A(n_364),
.B(n_378),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_354),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_372),
.B(n_377),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_335),
.B(n_331),
.C(n_330),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_374),
.B(n_380),
.C(n_356),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_357),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_336),
.A2(n_348),
.B1(n_329),
.B2(n_343),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_333),
.B(n_318),
.C(n_290),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_353),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_382),
.B(n_340),
.Y(n_399)
);

OAI21xp5_ASAP7_75t_L g384 ( 
.A1(n_344),
.A2(n_302),
.B(n_320),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_328),
.B(n_302),
.Y(n_388)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_388),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_332),
.B(n_233),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_SL g420 ( 
.A(n_389),
.B(n_390),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_352),
.B(n_233),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_SL g391 ( 
.A1(n_345),
.A2(n_293),
.B1(n_320),
.B2(n_263),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_SL g427 ( 
.A1(n_392),
.A2(n_370),
.B1(n_385),
.B2(n_365),
.Y(n_427)
);

XOR2xp5_ASAP7_75t_L g440 ( 
.A(n_394),
.B(n_400),
.Y(n_440)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_369),
.Y(n_395)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_395),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_366),
.B(n_334),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g422 ( 
.A(n_397),
.B(n_404),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_399),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g400 ( 
.A(n_366),
.B(n_356),
.Y(n_400)
);

OAI21xp5_ASAP7_75t_L g401 ( 
.A1(n_362),
.A2(n_327),
.B(n_338),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_401),
.B(n_411),
.Y(n_437)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_369),
.Y(n_402)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_402),
.Y(n_428)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_371),
.Y(n_403)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_403),
.Y(n_436)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_371),
.Y(n_405)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_405),
.Y(n_438)
);

CKINVDCx16_ASAP7_75t_R g406 ( 
.A(n_386),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_SL g432 ( 
.A(n_406),
.B(n_412),
.Y(n_432)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_386),
.Y(n_407)
);

HB1xp67_ASAP7_75t_L g429 ( 
.A(n_407),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_364),
.B(n_350),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_L g424 ( 
.A(n_408),
.B(n_416),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_374),
.B(n_341),
.C(n_327),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_410),
.B(n_414),
.C(n_384),
.Y(n_426)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_360),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_387),
.Y(n_412)
);

XOR2xp5_ASAP7_75t_L g413 ( 
.A(n_379),
.B(n_361),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_L g421 ( 
.A(n_413),
.B(n_417),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_380),
.B(n_385),
.C(n_378),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_L g415 ( 
.A1(n_359),
.A2(n_349),
.B1(n_293),
.B2(n_351),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_415),
.A2(n_391),
.B1(n_363),
.B2(n_368),
.Y(n_423)
);

OAI21xp5_ASAP7_75t_L g416 ( 
.A1(n_373),
.A2(n_229),
.B(n_165),
.Y(n_416)
);

XOR2xp5_ASAP7_75t_L g417 ( 
.A(n_387),
.B(n_224),
.Y(n_417)
);

XOR2xp5_ASAP7_75t_L g418 ( 
.A(n_388),
.B(n_224),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_SL g444 ( 
.A(n_418),
.B(n_419),
.Y(n_444)
);

XOR2xp5_ASAP7_75t_L g419 ( 
.A(n_367),
.B(n_195),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_L g460 ( 
.A1(n_423),
.A2(n_443),
.B1(n_227),
.B2(n_194),
.Y(n_460)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_426),
.B(n_435),
.Y(n_461)
);

AOI22xp5_ASAP7_75t_L g464 ( 
.A1(n_427),
.A2(n_188),
.B1(n_177),
.B2(n_209),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_400),
.B(n_373),
.C(n_382),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_430),
.B(n_439),
.Y(n_449)
);

INVx1_ASAP7_75t_SL g433 ( 
.A(n_407),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_433),
.B(n_363),
.Y(n_445)
);

FAx1_ASAP7_75t_SL g434 ( 
.A(n_414),
.B(n_377),
.CI(n_372),
.CON(n_434),
.SN(n_434)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_434),
.B(n_442),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_L g435 ( 
.A(n_397),
.B(n_383),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_398),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_404),
.B(n_410),
.C(n_408),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_441),
.B(n_413),
.C(n_394),
.Y(n_447)
);

BUFx24_ASAP7_75t_SL g442 ( 
.A(n_420),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_396),
.A2(n_383),
.B1(n_365),
.B2(n_368),
.Y(n_443)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_445),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_SL g479 ( 
.A(n_447),
.B(n_457),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_422),
.B(n_418),
.C(n_417),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_448),
.B(n_450),
.Y(n_471)
);

NAND3xp33_ASAP7_75t_L g450 ( 
.A(n_437),
.B(n_381),
.C(n_432),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_SL g451 ( 
.A1(n_431),
.A2(n_392),
.B1(n_393),
.B2(n_401),
.Y(n_451)
);

AOI22xp5_ASAP7_75t_L g467 ( 
.A1(n_451),
.A2(n_460),
.B1(n_438),
.B2(n_436),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_434),
.B(n_419),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_SL g468 ( 
.A(n_452),
.B(n_454),
.Y(n_468)
);

HB1xp67_ASAP7_75t_L g453 ( 
.A(n_429),
.Y(n_453)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_453),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_435),
.B(n_375),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_433),
.B(n_375),
.Y(n_455)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_455),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_430),
.B(n_234),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_SL g470 ( 
.A(n_456),
.B(n_462),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_422),
.B(n_409),
.C(n_416),
.Y(n_457)
);

OAI21xp5_ASAP7_75t_SL g458 ( 
.A1(n_426),
.A2(n_409),
.B(n_174),
.Y(n_458)
);

AOI21xp5_ASAP7_75t_L g482 ( 
.A1(n_458),
.A2(n_459),
.B(n_445),
.Y(n_482)
);

INVx13_ASAP7_75t_L g459 ( 
.A(n_425),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_421),
.B(n_191),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_441),
.B(n_213),
.C(n_207),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_463),
.B(n_424),
.C(n_444),
.Y(n_469)
);

XNOR2x1_ASAP7_75t_L g475 ( 
.A(n_464),
.B(n_455),
.Y(n_475)
);

AOI21xp33_ASAP7_75t_SL g466 ( 
.A1(n_446),
.A2(n_440),
.B(n_428),
.Y(n_466)
);

XNOR2xp5_ASAP7_75t_L g496 ( 
.A(n_466),
.B(n_469),
.Y(n_496)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_467),
.Y(n_490)
);

AND2x2_ASAP7_75t_L g472 ( 
.A(n_449),
.B(n_440),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_472),
.B(n_474),
.Y(n_483)
);

AOI22xp5_ASAP7_75t_L g473 ( 
.A1(n_451),
.A2(n_424),
.B1(n_444),
.B2(n_156),
.Y(n_473)
);

HB1xp67_ASAP7_75t_L g486 ( 
.A(n_473),
.Y(n_486)
);

OAI21xp5_ASAP7_75t_L g474 ( 
.A1(n_457),
.A2(n_167),
.B(n_162),
.Y(n_474)
);

OR2x2_ASAP7_75t_L g497 ( 
.A(n_475),
.B(n_27),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_461),
.B(n_447),
.C(n_448),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_476),
.B(n_482),
.Y(n_484)
);

XOR2xp5_ASAP7_75t_L g477 ( 
.A(n_461),
.B(n_106),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_477),
.B(n_478),
.C(n_459),
.Y(n_487)
);

XOR2xp5_ASAP7_75t_L g478 ( 
.A(n_458),
.B(n_463),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_SL g485 ( 
.A(n_471),
.B(n_464),
.Y(n_485)
);

CKINVDCx20_ASAP7_75t_R g505 ( 
.A(n_485),
.Y(n_505)
);

XOR2xp5_ASAP7_75t_L g498 ( 
.A(n_487),
.B(n_477),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_SL g488 ( 
.A(n_476),
.B(n_152),
.Y(n_488)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_488),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_SL g489 ( 
.A(n_468),
.B(n_154),
.Y(n_489)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_489),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_SL g491 ( 
.A(n_479),
.B(n_2),
.Y(n_491)
);

AOI21xp5_ASAP7_75t_L g499 ( 
.A1(n_491),
.A2(n_493),
.B(n_494),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_480),
.B(n_2),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_492),
.B(n_495),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_478),
.B(n_123),
.C(n_132),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_SL g494 ( 
.A(n_472),
.B(n_470),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_465),
.B(n_3),
.Y(n_495)
);

INVxp67_ASAP7_75t_L g502 ( 
.A(n_497),
.Y(n_502)
);

AND2x2_ASAP7_75t_L g513 ( 
.A(n_498),
.B(n_11),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_496),
.B(n_467),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_501),
.B(n_503),
.Y(n_515)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_490),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_484),
.B(n_475),
.C(n_481),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_507),
.B(n_508),
.Y(n_516)
);

OAI22xp5_ASAP7_75t_L g508 ( 
.A1(n_486),
.A2(n_473),
.B1(n_474),
.B2(n_469),
.Y(n_508)
);

AND2x2_ASAP7_75t_L g509 ( 
.A(n_486),
.B(n_3),
.Y(n_509)
);

AOI21xp5_ASAP7_75t_L g514 ( 
.A1(n_509),
.A2(n_11),
.B(n_500),
.Y(n_514)
);

INVxp67_ASAP7_75t_L g510 ( 
.A(n_509),
.Y(n_510)
);

OAI21xp5_ASAP7_75t_L g517 ( 
.A1(n_510),
.A2(n_512),
.B(n_504),
.Y(n_517)
);

AOI322xp5_ASAP7_75t_L g511 ( 
.A1(n_505),
.A2(n_483),
.A3(n_497),
.B1(n_493),
.B2(n_7),
.C1(n_12),
.C2(n_11),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_511),
.B(n_513),
.Y(n_518)
);

OAI21xp5_ASAP7_75t_SL g512 ( 
.A1(n_499),
.A2(n_11),
.B(n_12),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_514),
.B(n_506),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_517),
.B(n_519),
.Y(n_522)
);

CKINVDCx20_ASAP7_75t_R g519 ( 
.A(n_515),
.Y(n_519)
);

XNOR2xp5_ASAP7_75t_L g521 ( 
.A(n_520),
.B(n_498),
.Y(n_521)
);

INVxp67_ASAP7_75t_L g523 ( 
.A(n_521),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_523),
.B(n_522),
.Y(n_524)
);

AOI21xp5_ASAP7_75t_L g525 ( 
.A1(n_524),
.A2(n_516),
.B(n_518),
.Y(n_525)
);

XOR2xp5_ASAP7_75t_L g526 ( 
.A(n_525),
.B(n_502),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_SL g527 ( 
.A(n_526),
.B(n_502),
.Y(n_527)
);


endmodule