module fake_ariane_2534_n_856 (n_83, n_8, n_56, n_60, n_170, n_160, n_64, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_856);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_160;
input n_64;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_856;

wire n_295;
wire n_356;
wire n_556;
wire n_190;
wire n_698;
wire n_695;
wire n_180;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_581;
wire n_294;
wire n_646;
wire n_197;
wire n_640;
wire n_463;
wire n_830;
wire n_691;
wire n_404;
wire n_678;
wire n_651;
wire n_347;
wire n_423;
wire n_183;
wire n_469;
wire n_479;
wire n_726;
wire n_603;
wire n_373;
wire n_299;
wire n_836;
wire n_541;
wire n_499;
wire n_789;
wire n_788;
wire n_850;
wire n_771;
wire n_564;
wire n_610;
wire n_205;
wire n_752;
wire n_341;
wire n_421;
wire n_245;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_760;
wire n_690;
wire n_416;
wire n_283;
wire n_525;
wire n_187;
wire n_806;
wire n_367;
wire n_713;
wire n_649;
wire n_598;
wire n_345;
wire n_374;
wire n_318;
wire n_817;
wire n_244;
wire n_643;
wire n_679;
wire n_226;
wire n_781;
wire n_220;
wire n_261;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_189;
wire n_717;
wire n_819;
wire n_286;
wire n_586;
wire n_443;
wire n_686;
wire n_605;
wire n_776;
wire n_528;
wire n_584;
wire n_424;
wire n_387;
wire n_406;
wire n_826;
wire n_524;
wire n_634;
wire n_391;
wire n_349;
wire n_756;
wire n_466;
wire n_346;
wire n_214;
wire n_764;
wire n_348;
wire n_552;
wire n_462;
wire n_607;
wire n_670;
wire n_410;
wire n_379;
wire n_445;
wire n_515;
wire n_807;
wire n_765;
wire n_264;
wire n_737;
wire n_198;
wire n_232;
wire n_441;
wire n_568;
wire n_385;
wire n_637;
wire n_327;
wire n_766;
wire n_372;
wire n_377;
wire n_396;
wire n_802;
wire n_631;
wire n_399;
wire n_554;
wire n_520;
wire n_714;
wire n_279;
wire n_702;
wire n_207;
wire n_790;
wire n_363;
wire n_720;
wire n_354;
wire n_813;
wire n_725;
wire n_419;
wire n_230;
wire n_270;
wire n_194;
wire n_633;
wire n_338;
wire n_285;
wire n_473;
wire n_186;
wire n_801;
wire n_202;
wire n_193;
wire n_761;
wire n_733;
wire n_818;
wire n_500;
wire n_665;
wire n_336;
wire n_731;
wire n_754;
wire n_779;
wire n_315;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_829;
wire n_668;
wire n_339;
wire n_738;
wire n_758;
wire n_833;
wire n_672;
wire n_487;
wire n_740;
wire n_422;
wire n_648;
wire n_784;
wire n_269;
wire n_597;
wire n_816;
wire n_855;
wire n_259;
wire n_835;
wire n_808;
wire n_553;
wire n_446;
wire n_753;
wire n_566;
wire n_814;
wire n_578;
wire n_701;
wire n_625;
wire n_405;
wire n_557;
wire n_242;
wire n_645;
wire n_309;
wire n_320;
wire n_331;
wire n_559;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_822;
wire n_344;
wire n_381;
wire n_795;
wire n_426;
wire n_481;
wire n_600;
wire n_433;
wire n_721;
wire n_840;
wire n_398;
wire n_210;
wire n_200;
wire n_529;
wire n_502;
wire n_253;
wire n_561;
wire n_770;
wire n_218;
wire n_821;
wire n_839;
wire n_271;
wire n_507;
wire n_486;
wire n_465;
wire n_759;
wire n_247;
wire n_569;
wire n_567;
wire n_825;
wire n_732;
wire n_240;
wire n_369;
wire n_224;
wire n_787;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_222;
wire n_478;
wire n_703;
wire n_748;
wire n_786;
wire n_510;
wire n_831;
wire n_256;
wire n_326;
wire n_681;
wire n_778;
wire n_227;
wire n_188;
wire n_323;
wire n_550;
wire n_635;
wire n_707;
wire n_330;
wire n_400;
wire n_689;
wire n_694;
wire n_282;
wire n_328;
wire n_368;
wire n_590;
wire n_699;
wire n_727;
wire n_277;
wire n_248;
wire n_301;
wire n_467;
wire n_432;
wire n_545;
wire n_536;
wire n_644;
wire n_293;
wire n_823;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_693;
wire n_303;
wire n_671;
wire n_442;
wire n_777;
wire n_206;
wire n_352;
wire n_538;
wire n_576;
wire n_843;
wire n_511;
wire n_611;
wire n_238;
wire n_365;
wire n_429;
wire n_455;
wire n_654;
wire n_588;
wire n_638;
wire n_334;
wire n_192;
wire n_729;
wire n_661;
wire n_488;
wire n_775;
wire n_667;
wire n_300;
wire n_533;
wire n_505;
wire n_846;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_512;
wire n_715;
wire n_579;
wire n_844;
wire n_459;
wire n_685;
wire n_221;
wire n_321;
wire n_361;
wire n_458;
wire n_383;
wire n_623;
wire n_838;
wire n_237;
wire n_780;
wire n_711;
wire n_453;
wire n_734;
wire n_491;
wire n_810;
wire n_181;
wire n_723;
wire n_616;
wire n_658;
wire n_617;
wire n_630;
wire n_705;
wire n_570;
wire n_260;
wire n_362;
wire n_543;
wire n_310;
wire n_709;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_281;
wire n_628;
wire n_809;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_743;
wire n_225;
wire n_235;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_297;
wire n_662;
wire n_641;
wire n_503;
wire n_700;
wire n_290;
wire n_527;
wire n_741;
wire n_772;
wire n_747;
wire n_847;
wire n_371;
wire n_845;
wire n_199;
wire n_639;
wire n_217;
wire n_452;
wire n_673;
wire n_676;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_201;
wire n_572;
wire n_343;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_582;
wire n_284;
wire n_448;
wire n_593;
wire n_755;
wire n_710;
wire n_249;
wire n_534;
wire n_212;
wire n_355;
wire n_444;
wire n_609;
wire n_278;
wire n_851;
wire n_255;
wire n_560;
wire n_450;
wire n_257;
wire n_842;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_409;
wire n_519;
wire n_384;
wire n_468;
wire n_853;
wire n_526;
wire n_716;
wire n_742;
wire n_182;
wire n_696;
wire n_674;
wire n_482;
wire n_316;
wire n_196;
wire n_798;
wire n_769;
wire n_820;
wire n_577;
wire n_407;
wire n_774;
wire n_254;
wire n_596;
wire n_476;
wire n_460;
wire n_219;
wire n_832;
wire n_535;
wire n_231;
wire n_366;
wire n_744;
wire n_762;
wire n_656;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_848;
wire n_804;
wire n_280;
wire n_215;
wire n_252;
wire n_629;
wire n_664;
wire n_454;
wire n_298;
wire n_532;
wire n_415;
wire n_794;
wire n_763;
wire n_655;
wire n_544;
wire n_540;
wire n_216;
wire n_692;
wire n_599;
wire n_768;
wire n_514;
wire n_418;
wire n_537;
wire n_223;
wire n_403;
wire n_750;
wire n_834;
wire n_389;
wire n_800;
wire n_657;
wire n_513;
wire n_837;
wire n_288;
wire n_179;
wire n_812;
wire n_395;
wire n_621;
wire n_195;
wire n_606;
wire n_213;
wire n_304;
wire n_659;
wire n_509;
wire n_583;
wire n_724;
wire n_306;
wire n_666;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_203;
wire n_378;
wire n_436;
wire n_757;
wire n_375;
wire n_324;
wire n_585;
wire n_669;
wire n_785;
wire n_827;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_622;
wire n_697;
wire n_472;
wire n_296;
wire n_265;
wire n_746;
wire n_208;
wire n_456;
wire n_292;
wire n_793;
wire n_852;
wire n_275;
wire n_704;
wire n_204;
wire n_751;
wire n_615;
wire n_521;
wire n_496;
wire n_739;
wire n_342;
wire n_246;
wire n_517;
wire n_530;
wire n_792;
wire n_824;
wire n_428;
wire n_358;
wire n_580;
wire n_608;
wire n_494;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_563;
wire n_229;
wire n_394;
wire n_250;
wire n_773;
wire n_317;
wire n_243;
wire n_803;
wire n_329;
wire n_718;
wire n_185;
wire n_340;
wire n_749;
wire n_289;
wire n_548;
wire n_542;
wire n_815;
wire n_523;
wire n_268;
wire n_266;
wire n_470;
wire n_457;
wire n_632;
wire n_184;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_782;
wire n_425;
wire n_431;
wire n_811;
wire n_508;
wire n_624;
wire n_791;
wire n_618;
wire n_411;
wire n_484;
wire n_712;
wire n_849;
wire n_353;
wire n_736;
wire n_767;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_191;
wire n_382;
wire n_797;
wire n_489;
wire n_480;
wire n_211;
wire n_642;
wire n_408;
wire n_828;
wire n_595;
wire n_322;
wire n_251;
wire n_506;
wire n_602;
wire n_799;
wire n_558;
wire n_592;
wire n_397;
wire n_841;
wire n_854;
wire n_471;
wire n_351;
wire n_393;
wire n_474;
wire n_653;
wire n_359;
wire n_573;
wire n_796;
wire n_805;
wire n_531;
wire n_783;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_27),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_35),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_137),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_75),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_92),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_15),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_67),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_164),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_49),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_26),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_62),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_134),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_22),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_144),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_117),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_89),
.Y(n_194)
);

BUFx2_ASAP7_75t_L g195 ( 
.A(n_178),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_142),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_11),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_118),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_119),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_29),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_145),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_162),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_108),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_21),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_37),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_158),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_25),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_166),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_84),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_48),
.Y(n_210)
);

INVx1_ASAP7_75t_SL g211 ( 
.A(n_135),
.Y(n_211)
);

BUFx8_ASAP7_75t_SL g212 ( 
.A(n_167),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_46),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_129),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_5),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_23),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_72),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_57),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_11),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_77),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_147),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_16),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_82),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_136),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_171),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_138),
.Y(n_226)
);

INVx1_ASAP7_75t_SL g227 ( 
.A(n_30),
.Y(n_227)
);

CKINVDCx14_ASAP7_75t_R g228 ( 
.A(n_116),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_23),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_96),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_105),
.Y(n_231)
);

HB1xp67_ASAP7_75t_L g232 ( 
.A(n_9),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_54),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_28),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_100),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_170),
.Y(n_236)
);

INVx1_ASAP7_75t_SL g237 ( 
.A(n_173),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_163),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_83),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_168),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_114),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_33),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_81),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_120),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_90),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_165),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_169),
.Y(n_247)
);

INVxp67_ASAP7_75t_SL g248 ( 
.A(n_14),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_140),
.Y(n_249)
);

BUFx10_ASAP7_75t_L g250 ( 
.A(n_76),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_204),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g252 ( 
.A(n_204),
.Y(n_252)
);

AND2x4_ASAP7_75t_L g253 ( 
.A(n_184),
.B(n_0),
.Y(n_253)
);

BUFx12f_ASAP7_75t_L g254 ( 
.A(n_250),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_195),
.B(n_0),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_204),
.Y(n_256)
);

INVx4_ASAP7_75t_L g257 ( 
.A(n_250),
.Y(n_257)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_204),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_180),
.B(n_1),
.Y(n_259)
);

INVx5_ASAP7_75t_L g260 ( 
.A(n_250),
.Y(n_260)
);

BUFx12f_ASAP7_75t_L g261 ( 
.A(n_182),
.Y(n_261)
);

AND2x2_ASAP7_75t_L g262 ( 
.A(n_232),
.B(n_1),
.Y(n_262)
);

AND2x4_ASAP7_75t_L g263 ( 
.A(n_184),
.B(n_2),
.Y(n_263)
);

INVx6_ASAP7_75t_L g264 ( 
.A(n_204),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_220),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_185),
.B(n_2),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_219),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_186),
.B(n_3),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_220),
.B(n_3),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_187),
.Y(n_270)
);

INVx5_ASAP7_75t_L g271 ( 
.A(n_230),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_189),
.B(n_4),
.Y(n_272)
);

AND2x4_ASAP7_75t_L g273 ( 
.A(n_219),
.B(n_4),
.Y(n_273)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_230),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_212),
.B(n_34),
.Y(n_275)
);

INVx2_ASAP7_75t_SL g276 ( 
.A(n_215),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_249),
.B(n_5),
.Y(n_277)
);

BUFx6f_ASAP7_75t_L g278 ( 
.A(n_192),
.Y(n_278)
);

INVx5_ASAP7_75t_L g279 ( 
.A(n_228),
.Y(n_279)
);

INVxp33_ASAP7_75t_SL g280 ( 
.A(n_188),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_196),
.B(n_6),
.Y(n_281)
);

AND2x2_ASAP7_75t_L g282 ( 
.A(n_216),
.B(n_188),
.Y(n_282)
);

BUFx3_ASAP7_75t_L g283 ( 
.A(n_206),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_209),
.B(n_6),
.Y(n_284)
);

INVx5_ASAP7_75t_L g285 ( 
.A(n_181),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_233),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_236),
.B(n_7),
.Y(n_287)
);

AND2x4_ASAP7_75t_L g288 ( 
.A(n_238),
.B(n_239),
.Y(n_288)
);

BUFx2_ASAP7_75t_L g289 ( 
.A(n_179),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_241),
.Y(n_290)
);

AND2x4_ASAP7_75t_L g291 ( 
.A(n_242),
.B(n_243),
.Y(n_291)
);

INVx4_ASAP7_75t_L g292 ( 
.A(n_182),
.Y(n_292)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_190),
.Y(n_293)
);

INVx4_ASAP7_75t_L g294 ( 
.A(n_183),
.Y(n_294)
);

BUFx6f_ASAP7_75t_L g295 ( 
.A(n_193),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_183),
.B(n_7),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_235),
.B(n_8),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_235),
.B(n_240),
.Y(n_298)
);

NAND3x1_ASAP7_75t_L g299 ( 
.A(n_262),
.B(n_207),
.C(n_221),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_257),
.B(n_211),
.Y(n_300)
);

OR2x2_ASAP7_75t_L g301 ( 
.A(n_289),
.B(n_227),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_292),
.B(n_237),
.Y(n_302)
);

OAI22x1_ASAP7_75t_L g303 ( 
.A1(n_257),
.A2(n_248),
.B1(n_207),
.B2(n_191),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_264),
.Y(n_304)
);

OAI22xp33_ASAP7_75t_SL g305 ( 
.A1(n_275),
.A2(n_197),
.B1(n_229),
.B2(n_200),
.Y(n_305)
);

OAI22xp33_ASAP7_75t_L g306 ( 
.A1(n_257),
.A2(n_221),
.B1(n_234),
.B2(n_222),
.Y(n_306)
);

OAI22xp33_ASAP7_75t_L g307 ( 
.A1(n_254),
.A2(n_240),
.B1(n_246),
.B2(n_245),
.Y(n_307)
);

AND2x4_ASAP7_75t_L g308 ( 
.A(n_260),
.B(n_244),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_280),
.B(n_289),
.Y(n_309)
);

AO22x2_ASAP7_75t_L g310 ( 
.A1(n_288),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_280),
.A2(n_244),
.B1(n_246),
.B2(n_245),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_292),
.B(n_194),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_278),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_278),
.Y(n_314)
);

OAI22xp33_ASAP7_75t_SL g315 ( 
.A1(n_255),
.A2(n_247),
.B1(n_231),
.B2(n_226),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_264),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_264),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_262),
.A2(n_261),
.B1(n_282),
.B2(n_254),
.Y(n_318)
);

OAI22xp33_ASAP7_75t_SL g319 ( 
.A1(n_287),
.A2(n_225),
.B1(n_224),
.B2(n_223),
.Y(n_319)
);

AND2x2_ASAP7_75t_L g320 ( 
.A(n_260),
.B(n_198),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_261),
.A2(n_218),
.B1(n_217),
.B2(n_214),
.Y(n_321)
);

AND2x2_ASAP7_75t_SL g322 ( 
.A(n_253),
.B(n_199),
.Y(n_322)
);

OR2x6_ASAP7_75t_L g323 ( 
.A(n_282),
.B(n_10),
.Y(n_323)
);

HB1xp67_ASAP7_75t_L g324 ( 
.A(n_298),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_293),
.Y(n_325)
);

AND2x2_ASAP7_75t_L g326 ( 
.A(n_260),
.B(n_201),
.Y(n_326)
);

OAI22xp33_ASAP7_75t_SL g327 ( 
.A1(n_269),
.A2(n_213),
.B1(n_210),
.B2(n_208),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_264),
.Y(n_328)
);

OAI22xp33_ASAP7_75t_L g329 ( 
.A1(n_276),
.A2(n_205),
.B1(n_203),
.B2(n_202),
.Y(n_329)
);

AND2x2_ASAP7_75t_L g330 ( 
.A(n_260),
.B(n_12),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_253),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_272),
.A2(n_13),
.B1(n_15),
.B2(n_16),
.Y(n_332)
);

AND2x2_ASAP7_75t_L g333 ( 
.A(n_260),
.B(n_17),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_277),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_288),
.B(n_36),
.Y(n_335)
);

OAI22xp33_ASAP7_75t_L g336 ( 
.A1(n_276),
.A2(n_18),
.B1(n_19),
.B2(n_20),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_281),
.A2(n_20),
.B1(n_21),
.B2(n_22),
.Y(n_337)
);

OAI22xp33_ASAP7_75t_L g338 ( 
.A1(n_253),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_338)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_251),
.Y(n_339)
);

AND2x2_ASAP7_75t_L g340 ( 
.A(n_260),
.B(n_24),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_251),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_256),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_263),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_278),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_288),
.A2(n_30),
.B1(n_31),
.B2(n_32),
.Y(n_345)
);

OAI22xp33_ASAP7_75t_L g346 ( 
.A1(n_259),
.A2(n_31),
.B1(n_32),
.B2(n_38),
.Y(n_346)
);

AND2x2_ASAP7_75t_L g347 ( 
.A(n_292),
.B(n_39),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_256),
.Y(n_348)
);

OAI22xp33_ASAP7_75t_L g349 ( 
.A1(n_266),
.A2(n_40),
.B1(n_41),
.B2(n_42),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_294),
.B(n_43),
.Y(n_350)
);

INVx3_ASAP7_75t_L g351 ( 
.A(n_278),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_324),
.B(n_294),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_339),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_351),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_351),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_SL g356 ( 
.A(n_322),
.B(n_296),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_341),
.Y(n_357)
);

INVxp33_ASAP7_75t_L g358 ( 
.A(n_309),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_313),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_314),
.Y(n_360)
);

INVx2_ASAP7_75t_SL g361 ( 
.A(n_301),
.Y(n_361)
);

INVxp67_ASAP7_75t_SL g362 ( 
.A(n_344),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_342),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_348),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_304),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_316),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_317),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_328),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_335),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_335),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_324),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_300),
.B(n_294),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_330),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_333),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_302),
.B(n_293),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_340),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_302),
.B(n_293),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_325),
.Y(n_378)
);

XOR2xp5_ASAP7_75t_L g379 ( 
.A(n_306),
.B(n_297),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_312),
.B(n_293),
.Y(n_380)
);

AND2x4_ASAP7_75t_L g381 ( 
.A(n_323),
.B(n_263),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_SL g382 ( 
.A(n_322),
.B(n_263),
.Y(n_382)
);

NOR2xp67_ASAP7_75t_L g383 ( 
.A(n_321),
.B(n_279),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_311),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_308),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_308),
.Y(n_386)
);

AND2x2_ASAP7_75t_L g387 ( 
.A(n_323),
.B(n_283),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_347),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_320),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_326),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_323),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_345),
.Y(n_392)
);

BUFx3_ASAP7_75t_L g393 ( 
.A(n_350),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_310),
.Y(n_394)
);

XOR2x2_ASAP7_75t_L g395 ( 
.A(n_299),
.B(n_288),
.Y(n_395)
);

XOR2x2_ASAP7_75t_L g396 ( 
.A(n_318),
.B(n_291),
.Y(n_396)
);

XNOR2x2_ASAP7_75t_L g397 ( 
.A(n_310),
.B(n_268),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_329),
.B(n_293),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_329),
.B(n_295),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_310),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_332),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_334),
.Y(n_402)
);

AND2x2_ASAP7_75t_L g403 ( 
.A(n_303),
.B(n_283),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_337),
.Y(n_404)
);

OR2x2_ASAP7_75t_L g405 ( 
.A(n_306),
.B(n_291),
.Y(n_405)
);

BUFx12f_ASAP7_75t_L g406 ( 
.A(n_307),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_350),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_336),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_336),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_327),
.Y(n_410)
);

NAND2x1p5_ASAP7_75t_L g411 ( 
.A(n_305),
.B(n_263),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_338),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_343),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_315),
.B(n_295),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_338),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_319),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_331),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_346),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_346),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_SL g420 ( 
.A(n_349),
.B(n_291),
.Y(n_420)
);

NOR2xp67_ASAP7_75t_L g421 ( 
.A(n_407),
.B(n_271),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_353),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_369),
.B(n_291),
.Y(n_423)
);

INVx3_ASAP7_75t_L g424 ( 
.A(n_353),
.Y(n_424)
);

INVxp67_ASAP7_75t_L g425 ( 
.A(n_361),
.Y(n_425)
);

INVx1_ASAP7_75t_SL g426 ( 
.A(n_387),
.Y(n_426)
);

AND2x2_ASAP7_75t_L g427 ( 
.A(n_381),
.B(n_382),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_370),
.B(n_307),
.Y(n_428)
);

AND2x4_ASAP7_75t_L g429 ( 
.A(n_381),
.B(n_273),
.Y(n_429)
);

AND2x2_ASAP7_75t_L g430 ( 
.A(n_381),
.B(n_273),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_357),
.Y(n_431)
);

AND2x2_ASAP7_75t_L g432 ( 
.A(n_371),
.B(n_273),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_356),
.B(n_295),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_372),
.B(n_398),
.Y(n_434)
);

AND2x4_ASAP7_75t_L g435 ( 
.A(n_394),
.B(n_400),
.Y(n_435)
);

AND2x2_ASAP7_75t_L g436 ( 
.A(n_408),
.B(n_273),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_357),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_372),
.B(n_270),
.Y(n_438)
);

AND2x2_ASAP7_75t_L g439 ( 
.A(n_352),
.B(n_270),
.Y(n_439)
);

AND2x2_ASAP7_75t_L g440 ( 
.A(n_352),
.B(n_286),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_398),
.B(n_286),
.Y(n_441)
);

OR2x2_ASAP7_75t_L g442 ( 
.A(n_405),
.B(n_290),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_399),
.B(n_290),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_399),
.B(n_278),
.Y(n_444)
);

BUFx3_ASAP7_75t_L g445 ( 
.A(n_385),
.Y(n_445)
);

AND2x2_ASAP7_75t_L g446 ( 
.A(n_418),
.B(n_267),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_389),
.B(n_265),
.Y(n_447)
);

HB1xp67_ASAP7_75t_L g448 ( 
.A(n_412),
.Y(n_448)
);

INVxp67_ASAP7_75t_L g449 ( 
.A(n_390),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_373),
.B(n_265),
.Y(n_450)
);

AND2x2_ASAP7_75t_L g451 ( 
.A(n_419),
.B(n_267),
.Y(n_451)
);

HB1xp67_ASAP7_75t_L g452 ( 
.A(n_415),
.Y(n_452)
);

AND2x2_ASAP7_75t_L g453 ( 
.A(n_409),
.B(n_265),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_359),
.Y(n_454)
);

AND2x2_ASAP7_75t_L g455 ( 
.A(n_401),
.B(n_265),
.Y(n_455)
);

AND2x2_ASAP7_75t_L g456 ( 
.A(n_402),
.B(n_404),
.Y(n_456)
);

AND2x2_ASAP7_75t_L g457 ( 
.A(n_403),
.B(n_265),
.Y(n_457)
);

AND2x2_ASAP7_75t_L g458 ( 
.A(n_392),
.B(n_274),
.Y(n_458)
);

AND2x2_ASAP7_75t_L g459 ( 
.A(n_386),
.B(n_274),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_374),
.B(n_274),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_376),
.B(n_274),
.Y(n_461)
);

BUFx3_ASAP7_75t_L g462 ( 
.A(n_354),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_360),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_363),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_364),
.Y(n_465)
);

AND2x2_ASAP7_75t_L g466 ( 
.A(n_413),
.B(n_274),
.Y(n_466)
);

AND2x2_ASAP7_75t_L g467 ( 
.A(n_413),
.B(n_284),
.Y(n_467)
);

AND2x2_ASAP7_75t_L g468 ( 
.A(n_411),
.B(n_258),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_355),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_362),
.Y(n_470)
);

AND2x2_ASAP7_75t_L g471 ( 
.A(n_411),
.B(n_258),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_388),
.B(n_375),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_365),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_366),
.Y(n_474)
);

BUFx3_ASAP7_75t_L g475 ( 
.A(n_367),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_368),
.Y(n_476)
);

INVx3_ASAP7_75t_L g477 ( 
.A(n_388),
.Y(n_477)
);

HB1xp67_ASAP7_75t_L g478 ( 
.A(n_391),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_420),
.Y(n_479)
);

AND2x4_ASAP7_75t_L g480 ( 
.A(n_410),
.B(n_295),
.Y(n_480)
);

AND2x2_ASAP7_75t_L g481 ( 
.A(n_395),
.B(n_295),
.Y(n_481)
);

AND2x4_ASAP7_75t_L g482 ( 
.A(n_416),
.B(n_417),
.Y(n_482)
);

AND2x2_ASAP7_75t_L g483 ( 
.A(n_395),
.B(n_252),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_420),
.Y(n_484)
);

NOR2x1p5_ASAP7_75t_L g485 ( 
.A(n_406),
.B(n_349),
.Y(n_485)
);

INVx2_ASAP7_75t_SL g486 ( 
.A(n_393),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_375),
.B(n_271),
.Y(n_487)
);

HB1xp67_ASAP7_75t_L g488 ( 
.A(n_397),
.Y(n_488)
);

AND2x2_ASAP7_75t_L g489 ( 
.A(n_379),
.B(n_252),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_414),
.Y(n_490)
);

AND2x2_ASAP7_75t_L g491 ( 
.A(n_456),
.B(n_384),
.Y(n_491)
);

INVx1_ASAP7_75t_SL g492 ( 
.A(n_489),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_459),
.Y(n_493)
);

CKINVDCx8_ASAP7_75t_R g494 ( 
.A(n_482),
.Y(n_494)
);

AND2x4_ASAP7_75t_L g495 ( 
.A(n_427),
.B(n_482),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_459),
.Y(n_496)
);

HB1xp67_ASAP7_75t_L g497 ( 
.A(n_429),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_450),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_450),
.Y(n_499)
);

OR2x6_ASAP7_75t_L g500 ( 
.A(n_427),
.B(n_406),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_434),
.B(n_378),
.Y(n_501)
);

NAND2x1p5_ASAP7_75t_L g502 ( 
.A(n_435),
.B(n_383),
.Y(n_502)
);

BUFx10_ASAP7_75t_L g503 ( 
.A(n_429),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_422),
.Y(n_504)
);

INVxp67_ASAP7_75t_SL g505 ( 
.A(n_434),
.Y(n_505)
);

INVx5_ASAP7_75t_L g506 ( 
.A(n_435),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_422),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_431),
.Y(n_508)
);

BUFx6f_ASAP7_75t_L g509 ( 
.A(n_462),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_426),
.B(n_428),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_SL g511 ( 
.A(n_425),
.B(n_358),
.Y(n_511)
);

OR2x6_ASAP7_75t_L g512 ( 
.A(n_482),
.B(n_414),
.Y(n_512)
);

AND2x4_ASAP7_75t_L g513 ( 
.A(n_482),
.B(n_384),
.Y(n_513)
);

BUFx4f_ASAP7_75t_L g514 ( 
.A(n_435),
.Y(n_514)
);

BUFx2_ASAP7_75t_L g515 ( 
.A(n_425),
.Y(n_515)
);

AND2x2_ASAP7_75t_L g516 ( 
.A(n_456),
.B(n_396),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_439),
.B(n_377),
.Y(n_517)
);

OR2x2_ASAP7_75t_L g518 ( 
.A(n_489),
.B(n_358),
.Y(n_518)
);

AND2x2_ASAP7_75t_L g519 ( 
.A(n_456),
.B(n_396),
.Y(n_519)
);

NAND2x1p5_ASAP7_75t_L g520 ( 
.A(n_435),
.B(n_377),
.Y(n_520)
);

HB1xp67_ASAP7_75t_L g521 ( 
.A(n_429),
.Y(n_521)
);

NAND2x1p5_ASAP7_75t_L g522 ( 
.A(n_445),
.B(n_393),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_439),
.B(n_380),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_460),
.Y(n_524)
);

AND2x4_ASAP7_75t_L g525 ( 
.A(n_429),
.B(n_380),
.Y(n_525)
);

INVx4_ASAP7_75t_L g526 ( 
.A(n_445),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_460),
.Y(n_527)
);

HB1xp67_ASAP7_75t_L g528 ( 
.A(n_430),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_440),
.B(n_279),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_461),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_440),
.B(n_279),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_467),
.B(n_279),
.Y(n_532)
);

CKINVDCx20_ASAP7_75t_R g533 ( 
.A(n_426),
.Y(n_533)
);

AND2x2_ASAP7_75t_L g534 ( 
.A(n_467),
.B(n_279),
.Y(n_534)
);

AND2x4_ASAP7_75t_L g535 ( 
.A(n_430),
.B(n_44),
.Y(n_535)
);

AND2x2_ASAP7_75t_L g536 ( 
.A(n_481),
.B(n_442),
.Y(n_536)
);

NAND2x1p5_ASAP7_75t_L g537 ( 
.A(n_445),
.B(n_271),
.Y(n_537)
);

NAND2x1p5_ASAP7_75t_L g538 ( 
.A(n_477),
.B(n_271),
.Y(n_538)
);

BUFx4f_ASAP7_75t_L g539 ( 
.A(n_480),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_428),
.B(n_279),
.Y(n_540)
);

BUFx8_ASAP7_75t_L g541 ( 
.A(n_481),
.Y(n_541)
);

AND2x2_ASAP7_75t_L g542 ( 
.A(n_442),
.B(n_271),
.Y(n_542)
);

AND2x2_ASAP7_75t_L g543 ( 
.A(n_448),
.B(n_271),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_466),
.B(n_285),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_431),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_461),
.Y(n_546)
);

BUFx3_ASAP7_75t_L g547 ( 
.A(n_468),
.Y(n_547)
);

OR2x6_ASAP7_75t_L g548 ( 
.A(n_488),
.B(n_252),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_437),
.Y(n_549)
);

AND2x4_ASAP7_75t_L g550 ( 
.A(n_480),
.B(n_45),
.Y(n_550)
);

INVx4_ASAP7_75t_L g551 ( 
.A(n_506),
.Y(n_551)
);

BUFx2_ASAP7_75t_SL g552 ( 
.A(n_506),
.Y(n_552)
);

BUFx3_ASAP7_75t_L g553 ( 
.A(n_514),
.Y(n_553)
);

AND2x4_ASAP7_75t_L g554 ( 
.A(n_495),
.B(n_468),
.Y(n_554)
);

INVx3_ASAP7_75t_L g555 ( 
.A(n_514),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_504),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_504),
.Y(n_557)
);

INVx2_ASAP7_75t_SL g558 ( 
.A(n_506),
.Y(n_558)
);

INVx3_ASAP7_75t_L g559 ( 
.A(n_506),
.Y(n_559)
);

INVx1_ASAP7_75t_SL g560 ( 
.A(n_533),
.Y(n_560)
);

BUFx3_ASAP7_75t_L g561 ( 
.A(n_533),
.Y(n_561)
);

NAND2x1p5_ASAP7_75t_L g562 ( 
.A(n_539),
.B(n_479),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_507),
.Y(n_563)
);

INVx5_ASAP7_75t_L g564 ( 
.A(n_503),
.Y(n_564)
);

AND2x2_ASAP7_75t_L g565 ( 
.A(n_495),
.B(n_466),
.Y(n_565)
);

BUFx2_ASAP7_75t_L g566 ( 
.A(n_497),
.Y(n_566)
);

AND2x2_ASAP7_75t_L g567 ( 
.A(n_495),
.B(n_490),
.Y(n_567)
);

BUFx2_ASAP7_75t_SL g568 ( 
.A(n_494),
.Y(n_568)
);

BUFx8_ASAP7_75t_L g569 ( 
.A(n_515),
.Y(n_569)
);

BUFx12f_ASAP7_75t_L g570 ( 
.A(n_513),
.Y(n_570)
);

BUFx12f_ASAP7_75t_L g571 ( 
.A(n_513),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_510),
.B(n_505),
.Y(n_572)
);

AND2x4_ASAP7_75t_L g573 ( 
.A(n_547),
.B(n_513),
.Y(n_573)
);

BUFx2_ASAP7_75t_SL g574 ( 
.A(n_494),
.Y(n_574)
);

INVx1_ASAP7_75t_SL g575 ( 
.A(n_518),
.Y(n_575)
);

INVx4_ASAP7_75t_L g576 ( 
.A(n_539),
.Y(n_576)
);

INVx6_ASAP7_75t_L g577 ( 
.A(n_503),
.Y(n_577)
);

INVx3_ASAP7_75t_SL g578 ( 
.A(n_503),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_510),
.B(n_448),
.Y(n_579)
);

CKINVDCx16_ASAP7_75t_R g580 ( 
.A(n_511),
.Y(n_580)
);

INVx6_ASAP7_75t_L g581 ( 
.A(n_509),
.Y(n_581)
);

INVx2_ASAP7_75t_SL g582 ( 
.A(n_509),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_507),
.Y(n_583)
);

AOI22xp33_ASAP7_75t_SL g584 ( 
.A1(n_516),
.A2(n_488),
.B1(n_483),
.B2(n_452),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_L g585 ( 
.A(n_501),
.B(n_449),
.Y(n_585)
);

BUFx3_ASAP7_75t_L g586 ( 
.A(n_547),
.Y(n_586)
);

INVx3_ASAP7_75t_SL g587 ( 
.A(n_525),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_508),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_508),
.Y(n_589)
);

INVx1_ASAP7_75t_SL g590 ( 
.A(n_491),
.Y(n_590)
);

INVx3_ASAP7_75t_L g591 ( 
.A(n_509),
.Y(n_591)
);

INVx3_ASAP7_75t_SL g592 ( 
.A(n_525),
.Y(n_592)
);

BUFx2_ASAP7_75t_L g593 ( 
.A(n_497),
.Y(n_593)
);

BUFx12f_ASAP7_75t_L g594 ( 
.A(n_541),
.Y(n_594)
);

BUFx12f_ASAP7_75t_L g595 ( 
.A(n_541),
.Y(n_595)
);

AND2x2_ASAP7_75t_L g596 ( 
.A(n_536),
.B(n_490),
.Y(n_596)
);

BUFx12f_ASAP7_75t_L g597 ( 
.A(n_541),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_545),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_545),
.Y(n_599)
);

HB1xp67_ASAP7_75t_L g600 ( 
.A(n_521),
.Y(n_600)
);

CKINVDCx11_ASAP7_75t_R g601 ( 
.A(n_560),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_556),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_556),
.Y(n_603)
);

OAI22xp5_ASAP7_75t_L g604 ( 
.A1(n_585),
.A2(n_505),
.B1(n_525),
.B2(n_485),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_579),
.B(n_519),
.Y(n_605)
);

AOI22xp33_ASAP7_75t_L g606 ( 
.A1(n_584),
.A2(n_485),
.B1(n_480),
.B2(n_492),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_589),
.Y(n_607)
);

BUFx12f_ASAP7_75t_L g608 ( 
.A(n_569),
.Y(n_608)
);

BUFx3_ASAP7_75t_L g609 ( 
.A(n_569),
.Y(n_609)
);

OAI22xp5_ASAP7_75t_L g610 ( 
.A1(n_572),
.A2(n_486),
.B1(n_449),
.B2(n_522),
.Y(n_610)
);

BUFx10_ASAP7_75t_L g611 ( 
.A(n_573),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_557),
.Y(n_612)
);

INVx5_ASAP7_75t_L g613 ( 
.A(n_576),
.Y(n_613)
);

AOI22xp33_ASAP7_75t_L g614 ( 
.A1(n_590),
.A2(n_480),
.B1(n_483),
.B2(n_512),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_589),
.Y(n_615)
);

BUFx12f_ASAP7_75t_L g616 ( 
.A(n_569),
.Y(n_616)
);

BUFx12f_ASAP7_75t_L g617 ( 
.A(n_594),
.Y(n_617)
);

AOI22xp33_ASAP7_75t_SL g618 ( 
.A1(n_580),
.A2(n_512),
.B1(n_550),
.B2(n_500),
.Y(n_618)
);

AOI22xp33_ASAP7_75t_L g619 ( 
.A1(n_596),
.A2(n_512),
.B1(n_479),
.B2(n_484),
.Y(n_619)
);

OAI22xp33_ASAP7_75t_L g620 ( 
.A1(n_587),
.A2(n_484),
.B1(n_528),
.B2(n_523),
.Y(n_620)
);

BUFx2_ASAP7_75t_SL g621 ( 
.A(n_561),
.Y(n_621)
);

INVx1_ASAP7_75t_SL g622 ( 
.A(n_561),
.Y(n_622)
);

AOI22xp33_ASAP7_75t_L g623 ( 
.A1(n_596),
.A2(n_565),
.B1(n_567),
.B2(n_452),
.Y(n_623)
);

AND2x4_ASAP7_75t_L g624 ( 
.A(n_553),
.B(n_521),
.Y(n_624)
);

INVx6_ASAP7_75t_L g625 ( 
.A(n_576),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_557),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_563),
.Y(n_627)
);

OAI22xp5_ASAP7_75t_L g628 ( 
.A1(n_587),
.A2(n_486),
.B1(n_522),
.B2(n_528),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_580),
.Y(n_629)
);

AOI22xp33_ASAP7_75t_L g630 ( 
.A1(n_565),
.A2(n_567),
.B1(n_571),
.B2(n_570),
.Y(n_630)
);

AOI22xp33_ASAP7_75t_L g631 ( 
.A1(n_570),
.A2(n_455),
.B1(n_500),
.B2(n_458),
.Y(n_631)
);

AOI22xp33_ASAP7_75t_L g632 ( 
.A1(n_571),
.A2(n_455),
.B1(n_500),
.B2(n_458),
.Y(n_632)
);

CKINVDCx6p67_ASAP7_75t_R g633 ( 
.A(n_594),
.Y(n_633)
);

CKINVDCx20_ASAP7_75t_R g634 ( 
.A(n_595),
.Y(n_634)
);

HB1xp67_ASAP7_75t_L g635 ( 
.A(n_566),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_575),
.B(n_600),
.Y(n_636)
);

BUFx8_ASAP7_75t_L g637 ( 
.A(n_595),
.Y(n_637)
);

AOI22xp33_ASAP7_75t_L g638 ( 
.A1(n_573),
.A2(n_457),
.B1(n_550),
.B2(n_517),
.Y(n_638)
);

OAI22xp5_ASAP7_75t_L g639 ( 
.A1(n_587),
.A2(n_486),
.B1(n_535),
.B2(n_520),
.Y(n_639)
);

OAI22xp5_ASAP7_75t_L g640 ( 
.A1(n_592),
.A2(n_535),
.B1(n_566),
.B2(n_593),
.Y(n_640)
);

CKINVDCx14_ASAP7_75t_R g641 ( 
.A(n_597),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_563),
.Y(n_642)
);

INVx6_ASAP7_75t_L g643 ( 
.A(n_576),
.Y(n_643)
);

OAI22xp5_ASAP7_75t_L g644 ( 
.A1(n_592),
.A2(n_535),
.B1(n_520),
.B2(n_438),
.Y(n_644)
);

BUFx3_ASAP7_75t_L g645 ( 
.A(n_597),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_605),
.B(n_573),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_602),
.Y(n_647)
);

OAI22xp5_ASAP7_75t_L g648 ( 
.A1(n_623),
.A2(n_592),
.B1(n_593),
.B2(n_555),
.Y(n_648)
);

BUFx3_ASAP7_75t_L g649 ( 
.A(n_645),
.Y(n_649)
);

AOI22xp33_ASAP7_75t_SL g650 ( 
.A1(n_604),
.A2(n_550),
.B1(n_568),
.B2(n_574),
.Y(n_650)
);

AND2x2_ASAP7_75t_L g651 ( 
.A(n_635),
.B(n_583),
.Y(n_651)
);

AOI22xp33_ASAP7_75t_L g652 ( 
.A1(n_606),
.A2(n_614),
.B1(n_632),
.B2(n_631),
.Y(n_652)
);

AOI22xp33_ASAP7_75t_SL g653 ( 
.A1(n_644),
.A2(n_568),
.B1(n_574),
.B2(n_548),
.Y(n_653)
);

OAI22xp33_ASAP7_75t_L g654 ( 
.A1(n_640),
.A2(n_555),
.B1(n_548),
.B2(n_553),
.Y(n_654)
);

AND2x2_ASAP7_75t_L g655 ( 
.A(n_635),
.B(n_583),
.Y(n_655)
);

AOI22xp33_ASAP7_75t_L g656 ( 
.A1(n_606),
.A2(n_573),
.B1(n_548),
.B2(n_457),
.Y(n_656)
);

AOI22xp33_ASAP7_75t_L g657 ( 
.A1(n_614),
.A2(n_554),
.B1(n_534),
.B2(n_586),
.Y(n_657)
);

AOI222xp33_ASAP7_75t_L g658 ( 
.A1(n_623),
.A2(n_436),
.B1(n_432),
.B2(n_446),
.C1(n_451),
.C2(n_443),
.Y(n_658)
);

AOI22xp33_ASAP7_75t_SL g659 ( 
.A1(n_621),
.A2(n_639),
.B1(n_586),
.B2(n_629),
.Y(n_659)
);

AOI22xp33_ASAP7_75t_L g660 ( 
.A1(n_631),
.A2(n_554),
.B1(n_465),
.B2(n_464),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_603),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_612),
.Y(n_662)
);

AOI211xp5_ASAP7_75t_L g663 ( 
.A1(n_620),
.A2(n_476),
.B(n_474),
.C(n_432),
.Y(n_663)
);

AOI22xp33_ASAP7_75t_L g664 ( 
.A1(n_632),
.A2(n_554),
.B1(n_464),
.B2(n_465),
.Y(n_664)
);

OAI21xp33_ASAP7_75t_L g665 ( 
.A1(n_620),
.A2(n_438),
.B(n_472),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_637),
.Y(n_666)
);

AND2x2_ASAP7_75t_L g667 ( 
.A(n_626),
.B(n_588),
.Y(n_667)
);

AOI22xp33_ASAP7_75t_L g668 ( 
.A1(n_618),
.A2(n_471),
.B1(n_473),
.B2(n_454),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_627),
.Y(n_669)
);

OAI22xp5_ASAP7_75t_L g670 ( 
.A1(n_638),
.A2(n_622),
.B1(n_619),
.B2(n_630),
.Y(n_670)
);

NOR2xp33_ASAP7_75t_L g671 ( 
.A(n_601),
.B(n_609),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_607),
.Y(n_672)
);

INVx1_ASAP7_75t_SL g673 ( 
.A(n_636),
.Y(n_673)
);

OAI22xp5_ASAP7_75t_L g674 ( 
.A1(n_638),
.A2(n_555),
.B1(n_477),
.B2(n_526),
.Y(n_674)
);

INVx3_ASAP7_75t_L g675 ( 
.A(n_613),
.Y(n_675)
);

BUFx2_ASAP7_75t_L g676 ( 
.A(n_624),
.Y(n_676)
);

AOI22xp33_ASAP7_75t_L g677 ( 
.A1(n_619),
.A2(n_471),
.B1(n_473),
.B2(n_454),
.Y(n_677)
);

OAI22xp5_ASAP7_75t_L g678 ( 
.A1(n_630),
.A2(n_628),
.B1(n_610),
.B2(n_477),
.Y(n_678)
);

OAI22xp5_ASAP7_75t_L g679 ( 
.A1(n_625),
.A2(n_477),
.B1(n_526),
.B2(n_472),
.Y(n_679)
);

OAI222xp33_ASAP7_75t_L g680 ( 
.A1(n_642),
.A2(n_502),
.B1(n_598),
.B2(n_588),
.C1(n_562),
.C2(n_599),
.Y(n_680)
);

OAI22xp5_ASAP7_75t_L g681 ( 
.A1(n_625),
.A2(n_423),
.B1(n_578),
.B2(n_562),
.Y(n_681)
);

AOI22xp33_ASAP7_75t_L g682 ( 
.A1(n_615),
.A2(n_473),
.B1(n_454),
.B2(n_475),
.Y(n_682)
);

AND2x2_ASAP7_75t_L g683 ( 
.A(n_611),
.B(n_598),
.Y(n_683)
);

OAI21xp33_ASAP7_75t_L g684 ( 
.A1(n_641),
.A2(n_423),
.B(n_463),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_637),
.Y(n_685)
);

CKINVDCx20_ASAP7_75t_R g686 ( 
.A(n_634),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_611),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_625),
.Y(n_688)
);

AOI22xp33_ASAP7_75t_L g689 ( 
.A1(n_624),
.A2(n_475),
.B1(n_543),
.B2(n_599),
.Y(n_689)
);

INVx1_ASAP7_75t_SL g690 ( 
.A(n_608),
.Y(n_690)
);

AOI22xp33_ASAP7_75t_L g691 ( 
.A1(n_643),
.A2(n_475),
.B1(n_542),
.B2(n_463),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_643),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_643),
.B(n_446),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_613),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_613),
.Y(n_695)
);

NOR2xp33_ASAP7_75t_L g696 ( 
.A(n_616),
.B(n_478),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_SL g697 ( 
.A(n_663),
.B(n_613),
.Y(n_697)
);

OAI222xp33_ASAP7_75t_L g698 ( 
.A1(n_652),
.A2(n_670),
.B1(n_650),
.B2(n_673),
.C1(n_646),
.C2(n_657),
.Y(n_698)
);

AOI221xp5_ASAP7_75t_SL g699 ( 
.A1(n_684),
.A2(n_641),
.B1(n_476),
.B2(n_474),
.C(n_451),
.Y(n_699)
);

AOI22xp33_ASAP7_75t_L g700 ( 
.A1(n_658),
.A2(n_540),
.B1(n_433),
.B2(n_549),
.Y(n_700)
);

AOI22xp33_ASAP7_75t_L g701 ( 
.A1(n_668),
.A2(n_549),
.B1(n_437),
.B2(n_499),
.Y(n_701)
);

OAI222xp33_ASAP7_75t_L g702 ( 
.A1(n_656),
.A2(n_502),
.B1(n_562),
.B2(n_443),
.C1(n_441),
.C2(n_447),
.Y(n_702)
);

AOI22xp33_ASAP7_75t_L g703 ( 
.A1(n_660),
.A2(n_527),
.B1(n_530),
.B2(n_546),
.Y(n_703)
);

OAI22xp5_ASAP7_75t_L g704 ( 
.A1(n_664),
.A2(n_659),
.B1(n_648),
.B2(n_691),
.Y(n_704)
);

AOI22xp33_ASAP7_75t_L g705 ( 
.A1(n_665),
.A2(n_524),
.B1(n_498),
.B2(n_453),
.Y(n_705)
);

NAND3xp33_ASAP7_75t_L g706 ( 
.A(n_693),
.B(n_447),
.C(n_453),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_651),
.B(n_591),
.Y(n_707)
);

AOI22xp33_ASAP7_75t_L g708 ( 
.A1(n_653),
.A2(n_496),
.B1(n_493),
.B2(n_509),
.Y(n_708)
);

AOI22xp33_ASAP7_75t_L g709 ( 
.A1(n_677),
.A2(n_532),
.B1(n_441),
.B2(n_544),
.Y(n_709)
);

AOI22xp33_ASAP7_75t_L g710 ( 
.A1(n_678),
.A2(n_529),
.B1(n_531),
.B2(n_424),
.Y(n_710)
);

AOI22xp33_ASAP7_75t_L g711 ( 
.A1(n_689),
.A2(n_424),
.B1(n_617),
.B2(n_633),
.Y(n_711)
);

AOI22xp5_ASAP7_75t_L g712 ( 
.A1(n_696),
.A2(n_436),
.B1(n_577),
.B2(n_578),
.Y(n_712)
);

OAI211xp5_ASAP7_75t_SL g713 ( 
.A1(n_671),
.A2(n_469),
.B(n_478),
.C(n_591),
.Y(n_713)
);

AOI22xp33_ASAP7_75t_L g714 ( 
.A1(n_672),
.A2(n_424),
.B1(n_462),
.B2(n_558),
.Y(n_714)
);

OAI22xp5_ASAP7_75t_L g715 ( 
.A1(n_674),
.A2(n_578),
.B1(n_577),
.B2(n_564),
.Y(n_715)
);

AOI22xp33_ASAP7_75t_L g716 ( 
.A1(n_672),
.A2(n_424),
.B1(n_462),
.B2(n_558),
.Y(n_716)
);

OAI22xp5_ASAP7_75t_L g717 ( 
.A1(n_676),
.A2(n_577),
.B1(n_564),
.B2(n_552),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_651),
.B(n_591),
.Y(n_718)
);

OAI22xp5_ASAP7_75t_L g719 ( 
.A1(n_676),
.A2(n_577),
.B1(n_564),
.B2(n_552),
.Y(n_719)
);

AOI22xp33_ASAP7_75t_SL g720 ( 
.A1(n_681),
.A2(n_444),
.B1(n_436),
.B2(n_551),
.Y(n_720)
);

AOI22xp33_ASAP7_75t_L g721 ( 
.A1(n_683),
.A2(n_469),
.B1(n_470),
.B2(n_421),
.Y(n_721)
);

AND2x2_ASAP7_75t_L g722 ( 
.A(n_662),
.B(n_582),
.Y(n_722)
);

AOI22xp33_ASAP7_75t_L g723 ( 
.A1(n_683),
.A2(n_470),
.B1(n_421),
.B2(n_551),
.Y(n_723)
);

NAND3xp33_ASAP7_75t_L g724 ( 
.A(n_655),
.B(n_582),
.C(n_444),
.Y(n_724)
);

OAI22xp5_ASAP7_75t_L g725 ( 
.A1(n_686),
.A2(n_564),
.B1(n_581),
.B2(n_559),
.Y(n_725)
);

NAND3xp33_ASAP7_75t_L g726 ( 
.A(n_655),
.B(n_252),
.C(n_551),
.Y(n_726)
);

OAI22xp33_ASAP7_75t_L g727 ( 
.A1(n_654),
.A2(n_686),
.B1(n_690),
.B2(n_649),
.Y(n_727)
);

OAI21xp33_ASAP7_75t_L g728 ( 
.A1(n_662),
.A2(n_559),
.B(n_252),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_667),
.B(n_581),
.Y(n_729)
);

AND2x2_ASAP7_75t_L g730 ( 
.A(n_647),
.B(n_581),
.Y(n_730)
);

INVx1_ASAP7_75t_SL g731 ( 
.A(n_649),
.Y(n_731)
);

OAI22xp5_ASAP7_75t_L g732 ( 
.A1(n_666),
.A2(n_564),
.B1(n_581),
.B2(n_559),
.Y(n_732)
);

AOI22xp33_ASAP7_75t_L g733 ( 
.A1(n_682),
.A2(n_564),
.B1(n_537),
.B2(n_538),
.Y(n_733)
);

AOI22xp33_ASAP7_75t_L g734 ( 
.A1(n_667),
.A2(n_669),
.B1(n_661),
.B2(n_687),
.Y(n_734)
);

OAI22xp33_ASAP7_75t_L g735 ( 
.A1(n_688),
.A2(n_537),
.B1(n_538),
.B2(n_487),
.Y(n_735)
);

AOI22xp33_ASAP7_75t_SL g736 ( 
.A1(n_679),
.A2(n_487),
.B1(n_285),
.B2(n_51),
.Y(n_736)
);

AOI22xp33_ASAP7_75t_SL g737 ( 
.A1(n_687),
.A2(n_285),
.B1(n_50),
.B2(n_52),
.Y(n_737)
);

AOI22xp33_ASAP7_75t_L g738 ( 
.A1(n_692),
.A2(n_285),
.B1(n_53),
.B2(n_55),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_722),
.Y(n_739)
);

OAI221xp5_ASAP7_75t_L g740 ( 
.A1(n_699),
.A2(n_688),
.B1(n_692),
.B2(n_695),
.C(n_694),
.Y(n_740)
);

OAI22xp5_ASAP7_75t_L g741 ( 
.A1(n_704),
.A2(n_685),
.B1(n_666),
.B2(n_694),
.Y(n_741)
);

AND2x2_ASAP7_75t_SL g742 ( 
.A(n_734),
.B(n_675),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_722),
.B(n_675),
.Y(n_743)
);

OAI221xp5_ASAP7_75t_L g744 ( 
.A1(n_712),
.A2(n_685),
.B1(n_675),
.B2(n_680),
.C(n_285),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_730),
.B(n_47),
.Y(n_745)
);

AND2x2_ASAP7_75t_L g746 ( 
.A(n_730),
.B(n_56),
.Y(n_746)
);

OAI22xp33_ASAP7_75t_L g747 ( 
.A1(n_712),
.A2(n_285),
.B1(n_59),
.B2(n_60),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_707),
.B(n_58),
.Y(n_748)
);

AND2x2_ASAP7_75t_L g749 ( 
.A(n_718),
.B(n_61),
.Y(n_749)
);

AND2x2_ASAP7_75t_L g750 ( 
.A(n_729),
.B(n_63),
.Y(n_750)
);

AND2x2_ASAP7_75t_L g751 ( 
.A(n_724),
.B(n_64),
.Y(n_751)
);

OA211x2_ASAP7_75t_L g752 ( 
.A1(n_697),
.A2(n_65),
.B(n_66),
.C(n_68),
.Y(n_752)
);

AND2x2_ASAP7_75t_L g753 ( 
.A(n_724),
.B(n_69),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_728),
.Y(n_754)
);

OAI21xp5_ASAP7_75t_SL g755 ( 
.A1(n_698),
.A2(n_70),
.B(n_71),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_731),
.B(n_73),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_697),
.B(n_177),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_727),
.B(n_74),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_705),
.B(n_176),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_720),
.B(n_78),
.Y(n_760)
);

OAI21xp5_ASAP7_75t_L g761 ( 
.A1(n_713),
.A2(n_79),
.B(n_80),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_725),
.B(n_175),
.Y(n_762)
);

OAI21xp5_ASAP7_75t_L g763 ( 
.A1(n_726),
.A2(n_85),
.B(n_86),
.Y(n_763)
);

AOI22xp33_ASAP7_75t_L g764 ( 
.A1(n_700),
.A2(n_87),
.B1(n_88),
.B2(n_91),
.Y(n_764)
);

AOI22xp33_ASAP7_75t_L g765 ( 
.A1(n_706),
.A2(n_174),
.B1(n_94),
.B2(n_95),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_728),
.B(n_703),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_717),
.B(n_93),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_719),
.B(n_732),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_735),
.B(n_172),
.Y(n_769)
);

AOI22xp5_ASAP7_75t_L g770 ( 
.A1(n_755),
.A2(n_708),
.B1(n_711),
.B2(n_715),
.Y(n_770)
);

AOI22xp5_ASAP7_75t_L g771 ( 
.A1(n_755),
.A2(n_736),
.B1(n_737),
.B2(n_701),
.Y(n_771)
);

NOR3xp33_ASAP7_75t_L g772 ( 
.A(n_741),
.B(n_702),
.C(n_738),
.Y(n_772)
);

OAI211xp5_ASAP7_75t_L g773 ( 
.A1(n_761),
.A2(n_710),
.B(n_721),
.C(n_723),
.Y(n_773)
);

AND2x2_ASAP7_75t_L g774 ( 
.A(n_739),
.B(n_716),
.Y(n_774)
);

AND2x2_ASAP7_75t_L g775 ( 
.A(n_739),
.B(n_743),
.Y(n_775)
);

NOR2xp33_ASAP7_75t_L g776 ( 
.A(n_749),
.B(n_97),
.Y(n_776)
);

NAND3xp33_ASAP7_75t_L g777 ( 
.A(n_751),
.B(n_714),
.C(n_709),
.Y(n_777)
);

XNOR2xp5_ASAP7_75t_L g778 ( 
.A(n_742),
.B(n_746),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_754),
.B(n_733),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_754),
.Y(n_780)
);

AND2x2_ASAP7_75t_L g781 ( 
.A(n_742),
.B(n_749),
.Y(n_781)
);

AND2x2_ASAP7_75t_L g782 ( 
.A(n_742),
.B(n_98),
.Y(n_782)
);

OR2x2_ASAP7_75t_L g783 ( 
.A(n_768),
.B(n_99),
.Y(n_783)
);

AOI22xp5_ASAP7_75t_L g784 ( 
.A1(n_744),
.A2(n_101),
.B1(n_102),
.B2(n_103),
.Y(n_784)
);

NAND4xp25_ASAP7_75t_L g785 ( 
.A(n_740),
.B(n_104),
.C(n_106),
.D(n_107),
.Y(n_785)
);

NAND3xp33_ASAP7_75t_L g786 ( 
.A(n_751),
.B(n_753),
.C(n_758),
.Y(n_786)
);

AND2x2_ASAP7_75t_L g787 ( 
.A(n_746),
.B(n_109),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_753),
.Y(n_788)
);

OAI211xp5_ASAP7_75t_SL g789 ( 
.A1(n_760),
.A2(n_110),
.B(n_111),
.C(n_112),
.Y(n_789)
);

NOR2x1_ASAP7_75t_L g790 ( 
.A(n_786),
.B(n_748),
.Y(n_790)
);

NAND4xp75_ASAP7_75t_L g791 ( 
.A(n_782),
.B(n_752),
.C(n_750),
.D(n_757),
.Y(n_791)
);

BUFx6f_ASAP7_75t_L g792 ( 
.A(n_783),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_780),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_788),
.B(n_750),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_SL g795 ( 
.A(n_781),
.B(n_766),
.Y(n_795)
);

XNOR2xp5_ASAP7_75t_L g796 ( 
.A(n_778),
.B(n_787),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_775),
.B(n_745),
.Y(n_797)
);

INVx3_ASAP7_75t_L g798 ( 
.A(n_774),
.Y(n_798)
);

XNOR2xp5_ASAP7_75t_L g799 ( 
.A(n_770),
.B(n_756),
.Y(n_799)
);

XNOR2xp5_ASAP7_75t_L g800 ( 
.A(n_796),
.B(n_771),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_793),
.Y(n_801)
);

XNOR2x2_ASAP7_75t_L g802 ( 
.A(n_790),
.B(n_785),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_790),
.B(n_798),
.Y(n_803)
);

INVxp67_ASAP7_75t_SL g804 ( 
.A(n_798),
.Y(n_804)
);

OAI22x1_ASAP7_75t_L g805 ( 
.A1(n_800),
.A2(n_804),
.B1(n_799),
.B2(n_795),
.Y(n_805)
);

INVx3_ASAP7_75t_L g806 ( 
.A(n_802),
.Y(n_806)
);

AOI22x1_ASAP7_75t_L g807 ( 
.A1(n_804),
.A2(n_792),
.B1(n_763),
.B2(n_791),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_801),
.Y(n_808)
);

OA22x2_ASAP7_75t_L g809 ( 
.A1(n_803),
.A2(n_794),
.B1(n_797),
.B2(n_784),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_801),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_806),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_808),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_810),
.Y(n_813)
);

NAND4xp25_ASAP7_75t_L g814 ( 
.A(n_811),
.B(n_806),
.C(n_772),
.D(n_776),
.Y(n_814)
);

NAND4xp75_ASAP7_75t_L g815 ( 
.A(n_811),
.B(n_805),
.C(n_807),
.D(n_752),
.Y(n_815)
);

OAI22xp5_ASAP7_75t_L g816 ( 
.A1(n_815),
.A2(n_807),
.B1(n_809),
.B2(n_812),
.Y(n_816)
);

AOI22xp33_ASAP7_75t_L g817 ( 
.A1(n_814),
.A2(n_772),
.B1(n_813),
.B2(n_777),
.Y(n_817)
);

AOI22xp5_ASAP7_75t_L g818 ( 
.A1(n_814),
.A2(n_792),
.B1(n_773),
.B2(n_789),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_818),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_817),
.Y(n_820)
);

OAI22xp33_ASAP7_75t_L g821 ( 
.A1(n_816),
.A2(n_792),
.B1(n_759),
.B2(n_762),
.Y(n_821)
);

AOI22xp5_ASAP7_75t_L g822 ( 
.A1(n_818),
.A2(n_773),
.B1(n_789),
.B2(n_779),
.Y(n_822)
);

AO22x2_ASAP7_75t_L g823 ( 
.A1(n_816),
.A2(n_779),
.B1(n_769),
.B2(n_767),
.Y(n_823)
);

NOR2xp33_ASAP7_75t_L g824 ( 
.A(n_818),
.B(n_747),
.Y(n_824)
);

AND2x4_ASAP7_75t_L g825 ( 
.A(n_819),
.B(n_765),
.Y(n_825)
);

INVx2_ASAP7_75t_L g826 ( 
.A(n_823),
.Y(n_826)
);

AOI22xp5_ASAP7_75t_L g827 ( 
.A1(n_822),
.A2(n_764),
.B1(n_115),
.B2(n_121),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_820),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_824),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_821),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_820),
.Y(n_831)
);

AND5x1_ASAP7_75t_L g832 ( 
.A(n_827),
.B(n_113),
.C(n_122),
.D(n_123),
.E(n_124),
.Y(n_832)
);

OAI21xp5_ASAP7_75t_L g833 ( 
.A1(n_829),
.A2(n_125),
.B(n_126),
.Y(n_833)
);

NOR2xp67_ASAP7_75t_L g834 ( 
.A(n_830),
.B(n_127),
.Y(n_834)
);

NOR3xp33_ASAP7_75t_L g835 ( 
.A(n_828),
.B(n_128),
.C(n_130),
.Y(n_835)
);

AND3x4_ASAP7_75t_L g836 ( 
.A(n_825),
.B(n_131),
.C(n_132),
.Y(n_836)
);

AND4x1_ASAP7_75t_L g837 ( 
.A(n_831),
.B(n_133),
.C(n_139),
.D(n_141),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_836),
.Y(n_838)
);

NAND2x1_ASAP7_75t_L g839 ( 
.A(n_834),
.B(n_826),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_833),
.Y(n_840)
);

AOI22xp5_ASAP7_75t_L g841 ( 
.A1(n_835),
.A2(n_825),
.B1(n_837),
.B2(n_832),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_836),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_836),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_840),
.Y(n_844)
);

AO22x2_ASAP7_75t_L g845 ( 
.A1(n_839),
.A2(n_143),
.B1(n_146),
.B2(n_148),
.Y(n_845)
);

NAND4xp25_ASAP7_75t_L g846 ( 
.A(n_838),
.B(n_843),
.C(n_842),
.D(n_841),
.Y(n_846)
);

OAI22xp5_ASAP7_75t_L g847 ( 
.A1(n_838),
.A2(n_149),
.B1(n_150),
.B2(n_151),
.Y(n_847)
);

INVx4_ASAP7_75t_L g848 ( 
.A(n_838),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_844),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_848),
.Y(n_850)
);

OAI22xp5_ASAP7_75t_L g851 ( 
.A1(n_850),
.A2(n_849),
.B1(n_845),
.B2(n_847),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_851),
.Y(n_852)
);

OAI22xp33_ASAP7_75t_L g853 ( 
.A1(n_852),
.A2(n_846),
.B1(n_153),
.B2(n_154),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_853),
.Y(n_854)
);

AOI221xp5_ASAP7_75t_L g855 ( 
.A1(n_854),
.A2(n_152),
.B1(n_155),
.B2(n_156),
.C(n_157),
.Y(n_855)
);

AOI211xp5_ASAP7_75t_L g856 ( 
.A1(n_855),
.A2(n_159),
.B(n_160),
.C(n_161),
.Y(n_856)
);


endmodule