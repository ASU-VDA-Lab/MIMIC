module real_jpeg_32320_n_13 (n_8, n_116, n_0, n_111, n_2, n_114, n_10, n_9, n_12, n_6, n_121, n_11, n_112, n_120, n_7, n_117, n_3, n_119, n_5, n_4, n_115, n_1, n_118, n_113, n_13);

input n_8;
input n_116;
input n_0;
input n_111;
input n_2;
input n_114;
input n_10;
input n_9;
input n_12;
input n_6;
input n_121;
input n_11;
input n_112;
input n_120;
input n_7;
input n_117;
input n_3;
input n_119;
input n_5;
input n_4;
input n_115;
input n_1;
input n_118;
input n_113;

output n_13;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_68;
wire n_78;
wire n_83;
wire n_104;
wire n_64;
wire n_47;
wire n_22;
wire n_87;
wire n_105;
wire n_40;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_44;
wire n_28;
wire n_62;
wire n_106;
wire n_45;
wire n_42;
wire n_18;
wire n_77;
wire n_39;
wire n_94;
wire n_26;
wire n_19;
wire n_17;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_0),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_0),
.B(n_44),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_1),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_1),
.B(n_93),
.Y(n_105)
);

AOI221xp5_ASAP7_75t_L g58 ( 
.A1(n_2),
.A2(n_10),
.B1(n_59),
.B2(n_64),
.C(n_65),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_2),
.B(n_59),
.C(n_64),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_3),
.B(n_50),
.Y(n_49)
);

HAxp5_ASAP7_75t_SL g100 ( 
.A(n_3),
.B(n_101),
.CON(n_100),
.SN(n_100)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_5),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_6),
.Y(n_40)
);

AOI322xp5_ASAP7_75t_L g103 ( 
.A1(n_6),
.A2(n_34),
.A3(n_36),
.B1(n_42),
.B2(n_104),
.C1(n_106),
.C2(n_121),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g16 ( 
.A(n_7),
.B(n_17),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_8),
.B(n_61),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_9),
.Y(n_85)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_10),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g28 ( 
.A(n_11),
.B(n_29),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_11),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g14 ( 
.A1(n_12),
.A2(n_15),
.B1(n_16),
.B2(n_21),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

XOR2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_22),
.Y(n_13)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_17),
.B(n_116),
.Y(n_64)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_19),
.Y(n_96)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_20),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_20),
.Y(n_63)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_20),
.Y(n_90)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

AOI31xp67_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_55),
.A3(n_91),
.B(n_98),
.Y(n_24)
);

NOR3xp33_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_41),
.C(n_49),
.Y(n_25)
);

OAI21xp5_ASAP7_75t_L g98 ( 
.A1(n_26),
.A2(n_99),
.B(n_103),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_34),
.Y(n_26)
);

INVxp67_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NOR3xp33_ASAP7_75t_L g104 ( 
.A(n_28),
.B(n_49),
.C(n_105),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_29),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_31),
.Y(n_29)
);

INVx2_ASAP7_75t_SL g82 ( 
.A(n_31),
.Y(n_82)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_33),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_35),
.B(n_40),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_112),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

OA21x2_ASAP7_75t_SL g99 ( 
.A1(n_41),
.A2(n_100),
.B(n_102),
.Y(n_99)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_43),
.B(n_48),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_46),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

HB1xp67_ASAP7_75t_L g101 ( 
.A(n_50),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_52),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_85),
.C(n_86),
.Y(n_55)
);

AOI21xp5_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_77),
.B(n_84),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_67),
.B1(n_75),
.B2(n_76),
.Y(n_57)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_60),
.B(n_66),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_63),
.Y(n_61)
);

INVx2_ASAP7_75t_SL g66 ( 
.A(n_64),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_70),
.Y(n_68)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_78),
.B(n_83),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_78),
.B(n_83),
.Y(n_84)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_81),
.Y(n_79)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_89),
.Y(n_87)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_92),
.B(n_97),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_95),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

BUFx24_ASAP7_75t_SL g109 ( 
.A(n_100),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_108),
.Y(n_106)
);

CKINVDCx14_ASAP7_75t_R g30 ( 
.A(n_111),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_113),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_114),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_115),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_117),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_118),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_119),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_120),
.Y(n_94)
);


endmodule