module fake_jpeg_2926_n_183 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_183);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_183;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_170;
wire n_162;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_93;
wire n_54;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx5_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

INVx4_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_1),
.B(n_3),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_11),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

INVx11_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

INVx6_ASAP7_75t_SL g27 ( 
.A(n_10),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_21),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_29),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

BUFx2_ASAP7_75t_L g62 ( 
.A(n_30),
.Y(n_62)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_31),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

BUFx2_ASAP7_75t_L g72 ( 
.A(n_32),
.Y(n_72)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_33),
.Y(n_78)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_34),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_35),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_36),
.Y(n_80)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

INVx2_ASAP7_75t_SL g38 ( 
.A(n_13),
.Y(n_38)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_38),
.Y(n_70)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_14),
.B(n_0),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_40),
.B(n_45),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_41),
.Y(n_77)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

BUFx12_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_43),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

BUFx12_ASAP7_75t_L g74 ( 
.A(n_44),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_14),
.B(n_0),
.C(n_2),
.Y(n_45)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_46),
.B(n_49),
.Y(n_54)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_19),
.Y(n_47)
);

OR2x2_ASAP7_75t_L g63 ( 
.A(n_47),
.B(n_48),
.Y(n_63)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_16),
.B(n_2),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_18),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_50),
.B(n_52),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_19),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_51),
.B(n_12),
.Y(n_73)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_22),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_29),
.A2(n_25),
.B1(n_28),
.B2(n_17),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_56),
.A2(n_64),
.B1(n_82),
.B2(n_5),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_47),
.B(n_23),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_58),
.B(n_84),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_38),
.A2(n_25),
.B1(n_15),
.B2(n_24),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_61),
.A2(n_34),
.B1(n_50),
.B2(n_42),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_30),
.A2(n_25),
.B1(n_28),
.B2(n_17),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_36),
.B(n_16),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_68),
.B(n_76),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_73),
.B(n_59),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_48),
.B(n_23),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_75),
.B(n_83),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_36),
.B(n_20),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_35),
.B(n_20),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_79),
.B(n_81),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_41),
.B(n_24),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_32),
.A2(n_24),
.B1(n_15),
.B2(n_4),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_43),
.B(n_15),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_33),
.B(n_2),
.Y(n_84)
);

OAI32xp33_ASAP7_75t_L g85 ( 
.A1(n_58),
.A2(n_51),
.A3(n_44),
.B1(n_39),
.B2(n_37),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_85),
.B(n_89),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_63),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_87),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_84),
.B(n_50),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_90),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_75),
.B(n_3),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_92),
.B(n_96),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_63),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_93),
.B(n_97),
.Y(n_122)
);

AO22x1_ASAP7_75t_L g94 ( 
.A1(n_57),
.A2(n_46),
.B1(n_5),
.B2(n_6),
.Y(n_94)
);

O2A1O1Ixp33_ASAP7_75t_L g108 ( 
.A1(n_94),
.A2(n_78),
.B(n_70),
.C(n_71),
.Y(n_108)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_57),
.Y(n_95)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_95),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_53),
.B(n_4),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_54),
.B(n_4),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_99),
.A2(n_72),
.B1(n_65),
.B2(n_78),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_66),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_100),
.B(n_104),
.Y(n_113)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_62),
.Y(n_101)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_101),
.Y(n_117)
);

AOI22x1_ASAP7_75t_L g102 ( 
.A1(n_62),
.A2(n_5),
.B1(n_7),
.B2(n_9),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_102),
.A2(n_59),
.B1(n_77),
.B2(n_80),
.Y(n_118)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_59),
.Y(n_103)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_103),
.Y(n_125)
);

OR2x2_ASAP7_75t_L g104 ( 
.A(n_67),
.B(n_9),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_82),
.A2(n_9),
.B1(n_11),
.B2(n_55),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_105),
.A2(n_72),
.B1(n_71),
.B2(n_55),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_106),
.Y(n_127)
);

AOI21xp33_ASAP7_75t_L g107 ( 
.A1(n_70),
.A2(n_80),
.B(n_67),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_107),
.B(n_69),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_108),
.B(n_118),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_109),
.B(n_115),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_112),
.B(n_101),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_86),
.B(n_65),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_93),
.A2(n_77),
.B(n_69),
.Y(n_119)
);

NOR3xp33_ASAP7_75t_L g137 ( 
.A(n_119),
.B(n_120),
.C(n_113),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_86),
.A2(n_59),
.B1(n_74),
.B2(n_60),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_121),
.B(n_124),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_89),
.A2(n_85),
.B1(n_87),
.B2(n_106),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_106),
.A2(n_60),
.B1(n_74),
.B2(n_92),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_126),
.B(n_94),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_122),
.B(n_96),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_128),
.B(n_138),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_119),
.A2(n_100),
.B(n_104),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_130),
.Y(n_152)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_110),
.Y(n_131)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_131),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_127),
.B(n_98),
.C(n_95),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_133),
.B(n_127),
.C(n_123),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_135),
.B(n_141),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_136),
.B(n_137),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_123),
.B(n_88),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_117),
.Y(n_139)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_139),
.Y(n_144)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_110),
.Y(n_140)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_140),
.Y(n_146)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_117),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_132),
.A2(n_111),
.B1(n_115),
.B2(n_124),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_143),
.A2(n_130),
.B1(n_114),
.B2(n_121),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_141),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_145),
.A2(n_140),
.B(n_131),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_133),
.B(n_111),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_149),
.B(n_150),
.C(n_126),
.Y(n_156)
);

AO22x1_ASAP7_75t_SL g153 ( 
.A1(n_143),
.A2(n_129),
.B1(n_135),
.B2(n_132),
.Y(n_153)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_153),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_147),
.B(n_134),
.Y(n_154)
);

NAND3xp33_ASAP7_75t_L g164 ( 
.A(n_154),
.B(n_157),
.C(n_158),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_152),
.A2(n_116),
.B1(n_129),
.B2(n_118),
.Y(n_155)
);

HB1xp67_ASAP7_75t_L g163 ( 
.A(n_155),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_156),
.B(n_159),
.C(n_160),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_148),
.A2(n_91),
.B(n_116),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_150),
.B(n_114),
.C(n_125),
.Y(n_160)
);

OA21x2_ASAP7_75t_SL g165 ( 
.A1(n_154),
.A2(n_142),
.B(n_152),
.Y(n_165)
);

OA21x2_ASAP7_75t_SL g168 ( 
.A1(n_165),
.A2(n_166),
.B(n_151),
.Y(n_168)
);

NAND3xp33_ASAP7_75t_L g166 ( 
.A(n_153),
.B(n_97),
.C(n_88),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_161),
.A2(n_147),
.B1(n_149),
.B2(n_109),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_167),
.B(n_170),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_168),
.B(n_169),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_164),
.A2(n_108),
.B(n_146),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_164),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_162),
.B(n_144),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_171),
.B(n_144),
.C(n_146),
.Y(n_172)
);

OAI211xp5_ASAP7_75t_L g176 ( 
.A1(n_172),
.A2(n_175),
.B(n_173),
.C(n_169),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_170),
.B(n_125),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_176),
.B(n_177),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_174),
.A2(n_167),
.B1(n_163),
.B2(n_171),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_175),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_178),
.B(n_102),
.C(n_103),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_179),
.A2(n_102),
.B(n_94),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_181),
.B(n_180),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_182),
.B(n_74),
.Y(n_183)
);


endmodule