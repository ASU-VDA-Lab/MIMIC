module fake_jpeg_17500_n_352 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_352);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_352;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx1_ASAP7_75t_SL g26 ( 
.A(n_8),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_14),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVx11_ASAP7_75t_SL g31 ( 
.A(n_8),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_14),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_8),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_25),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_36),
.B(n_37),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g37 ( 
.A(n_31),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_23),
.B(n_0),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_41),
.B(n_23),
.Y(n_57)
);

OR2x2_ASAP7_75t_L g42 ( 
.A(n_22),
.B(n_0),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_42),
.B(n_49),
.Y(n_66)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

INVx2_ASAP7_75t_SL g44 ( 
.A(n_21),
.Y(n_44)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

BUFx2_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_21),
.Y(n_48)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_26),
.B(n_35),
.Y(n_49)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_16),
.Y(n_50)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_44),
.B(n_21),
.C(n_30),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_51),
.B(n_52),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_27),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_57),
.B(n_70),
.Y(n_84)
);

OAI22xp33_ASAP7_75t_L g60 ( 
.A1(n_39),
.A2(n_31),
.B1(n_26),
.B2(n_16),
.Y(n_60)
);

OAI22xp33_ASAP7_75t_L g97 ( 
.A1(n_60),
.A2(n_50),
.B1(n_47),
.B2(n_44),
.Y(n_97)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g93 ( 
.A(n_61),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_43),
.A2(n_26),
.B1(n_33),
.B2(n_29),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_62),
.A2(n_74),
.B1(n_22),
.B2(n_35),
.Y(n_86)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_68),
.Y(n_85)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_69),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_42),
.B(n_25),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_42),
.B(n_25),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_72),
.B(n_23),
.Y(n_92)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_38),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_73),
.B(n_38),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_39),
.A2(n_33),
.B1(n_29),
.B2(n_28),
.Y(n_74)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_45),
.Y(n_75)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_75),
.Y(n_98)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_56),
.Y(n_76)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_76),
.Y(n_112)
);

OAI32xp33_ASAP7_75t_L g77 ( 
.A1(n_66),
.A2(n_49),
.A3(n_36),
.B1(n_28),
.B2(n_17),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_77),
.A2(n_57),
.B1(n_27),
.B2(n_32),
.Y(n_116)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_78),
.Y(n_126)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_56),
.Y(n_79)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_79),
.Y(n_129)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_54),
.Y(n_80)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_80),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_71),
.B(n_20),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_81),
.B(n_83),
.Y(n_110)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_54),
.Y(n_82)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_82),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_67),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_86),
.B(n_97),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_52),
.B(n_20),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_87),
.B(n_89),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_67),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_63),
.Y(n_90)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_90),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_92),
.B(n_109),
.Y(n_136)
);

INVx2_ASAP7_75t_SL g94 ( 
.A(n_61),
.Y(n_94)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_94),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_58),
.A2(n_22),
.B1(n_24),
.B2(n_35),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_95),
.A2(n_32),
.B1(n_27),
.B2(n_34),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_53),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_96),
.B(n_100),
.Y(n_115)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_61),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g125 ( 
.A(n_99),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_64),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_64),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_101),
.Y(n_121)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_55),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_102),
.B(n_104),
.Y(n_127)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_63),
.Y(n_103)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_103),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_55),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_59),
.B(n_17),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_105),
.B(n_108),
.Y(n_137)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_59),
.Y(n_106)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_106),
.Y(n_123)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_58),
.Y(n_107)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_107),
.Y(n_138)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_68),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_57),
.B(n_32),
.Y(n_109)
);

A2O1A1Ixp33_ASAP7_75t_SL g111 ( 
.A1(n_84),
.A2(n_51),
.B(n_38),
.C(n_60),
.Y(n_111)
);

O2A1O1Ixp33_ASAP7_75t_L g153 ( 
.A1(n_111),
.A2(n_99),
.B(n_88),
.C(n_90),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_113),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_116),
.B(n_11),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_107),
.A2(n_69),
.B1(n_50),
.B2(n_73),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_118),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_91),
.A2(n_75),
.B1(n_65),
.B2(n_40),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_122),
.A2(n_92),
.B1(n_79),
.B2(n_76),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_85),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_124),
.B(n_128),
.Y(n_149)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_93),
.Y(n_128)
);

OAI21xp33_ASAP7_75t_L g130 ( 
.A1(n_109),
.A2(n_13),
.B(n_10),
.Y(n_130)
);

OR2x2_ASAP7_75t_SL g158 ( 
.A(n_130),
.B(n_134),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_91),
.A2(n_65),
.B1(n_40),
.B2(n_44),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_131),
.A2(n_132),
.B1(n_34),
.B2(n_102),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_91),
.A2(n_34),
.B1(n_37),
.B2(n_12),
.Y(n_132)
);

NOR2x1_ASAP7_75t_L g134 ( 
.A(n_77),
.B(n_24),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_115),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_140),
.B(n_160),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_131),
.A2(n_92),
.B(n_85),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_141),
.A2(n_138),
.B(n_139),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_142),
.A2(n_146),
.B1(n_155),
.B2(n_162),
.Y(n_183)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_123),
.Y(n_143)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_143),
.Y(n_175)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_123),
.Y(n_144)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_144),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_145),
.A2(n_161),
.B1(n_138),
.B2(n_120),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_135),
.A2(n_98),
.B1(n_97),
.B2(n_108),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_122),
.B(n_98),
.C(n_93),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_147),
.B(n_151),
.C(n_156),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_136),
.B(n_116),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_148),
.B(n_166),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_136),
.B(n_132),
.C(n_126),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_117),
.Y(n_152)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_152),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_153),
.A2(n_129),
.B(n_112),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_135),
.A2(n_103),
.B1(n_82),
.B2(n_80),
.Y(n_155)
);

MAJx2_ASAP7_75t_L g156 ( 
.A(n_134),
.B(n_106),
.C(n_30),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_117),
.Y(n_157)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_157),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_126),
.B(n_93),
.C(n_88),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_159),
.B(n_169),
.C(n_129),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_119),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_111),
.A2(n_94),
.B1(n_101),
.B2(n_24),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_110),
.B(n_94),
.Y(n_163)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_163),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_137),
.Y(n_164)
);

HB1xp67_ASAP7_75t_L g184 ( 
.A(n_164),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_135),
.A2(n_11),
.B1(n_15),
.B2(n_14),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_165),
.A2(n_10),
.B1(n_15),
.B2(n_13),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_114),
.B(n_21),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_120),
.Y(n_167)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_167),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_124),
.B(n_111),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_168),
.B(n_1),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_111),
.B(n_93),
.C(n_21),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_133),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_170),
.B(n_171),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_119),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_133),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_172),
.B(n_125),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_174),
.B(n_182),
.C(n_197),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_176),
.A2(n_185),
.B1(n_187),
.B2(n_193),
.Y(n_218)
);

OAI21xp33_ASAP7_75t_L g177 ( 
.A1(n_168),
.A2(n_111),
.B(n_112),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_177),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_148),
.B(n_127),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_SL g219 ( 
.A(n_179),
.B(n_181),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_149),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_180),
.B(n_195),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_169),
.B(n_139),
.C(n_125),
.Y(n_182)
);

OAI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_150),
.A2(n_128),
.B1(n_30),
.B2(n_19),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_189),
.A2(n_162),
.B1(n_164),
.B2(n_154),
.Y(n_210)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_190),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_146),
.A2(n_19),
.B1(n_121),
.B2(n_12),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_152),
.Y(n_195)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_196),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_151),
.B(n_121),
.C(n_19),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_141),
.B(n_161),
.Y(n_198)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_198),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_143),
.Y(n_199)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_199),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_145),
.A2(n_11),
.B1(n_10),
.B2(n_3),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_200),
.A2(n_156),
.B1(n_158),
.B2(n_157),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_153),
.B(n_1),
.Y(n_202)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_202),
.Y(n_229)
);

HB1xp67_ASAP7_75t_L g203 ( 
.A(n_144),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_203),
.B(n_205),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_159),
.Y(n_205)
);

INVx1_ASAP7_75t_SL g206 ( 
.A(n_170),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_206),
.B(n_167),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_140),
.B(n_121),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_207),
.B(n_172),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_194),
.B(n_153),
.Y(n_208)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_208),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_210),
.B(n_215),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_191),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_211),
.A2(n_223),
.B(n_226),
.Y(n_245)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_214),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_178),
.B(n_166),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_198),
.A2(n_155),
.B1(n_147),
.B2(n_165),
.Y(n_216)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_216),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_202),
.A2(n_142),
.B1(n_156),
.B2(n_158),
.Y(n_217)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_217),
.Y(n_252)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_222),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_191),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_224),
.Y(n_251)
);

INVx2_ASAP7_75t_SL g225 ( 
.A(n_206),
.Y(n_225)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_225),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_183),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_192),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_227),
.A2(n_228),
.B(n_230),
.Y(n_249)
);

XOR2x2_ASAP7_75t_L g230 ( 
.A(n_173),
.B(n_174),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_184),
.B(n_2),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_231),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_205),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_SL g250 ( 
.A1(n_232),
.A2(n_200),
.B(n_181),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_188),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_233),
.B(n_234),
.Y(n_240)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_192),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_199),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_235),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_229),
.B(n_180),
.Y(n_242)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_242),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_237),
.B(n_230),
.C(n_173),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_243),
.B(n_244),
.C(n_246),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_219),
.B(n_179),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_219),
.B(n_182),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_229),
.B(n_194),
.Y(n_247)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_247),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_237),
.B(n_221),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_248),
.B(n_254),
.C(n_216),
.Y(n_270)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_250),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_211),
.B(n_196),
.Y(n_253)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_253),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_220),
.B(n_197),
.C(n_176),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_220),
.A2(n_185),
.B1(n_175),
.B2(n_186),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_256),
.A2(n_228),
.B1(n_213),
.B2(n_232),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_223),
.B(n_204),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_257),
.B(n_258),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_227),
.B(n_204),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_208),
.A2(n_186),
.B(n_175),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_262),
.A2(n_209),
.B1(n_5),
.B2(n_6),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_238),
.B(n_225),
.Y(n_264)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_264),
.Y(n_286)
);

INVx1_ASAP7_75t_SL g267 ( 
.A(n_256),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_267),
.B(n_280),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_270),
.B(n_273),
.C(n_277),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_263),
.A2(n_218),
.B1(n_213),
.B2(n_225),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_271),
.A2(n_285),
.B1(n_255),
.B2(n_253),
.Y(n_299)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_272),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_243),
.B(n_217),
.C(n_212),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_252),
.A2(n_233),
.B1(n_212),
.B2(n_234),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_275),
.A2(n_241),
.B1(n_252),
.B2(n_263),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_SL g276 ( 
.A(n_244),
.B(n_210),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_276),
.B(n_249),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_248),
.B(n_236),
.C(n_201),
.Y(n_277)
);

CKINVDCx16_ASAP7_75t_R g278 ( 
.A(n_257),
.Y(n_278)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_278),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_246),
.B(n_226),
.C(n_235),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_279),
.B(n_254),
.C(n_261),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_258),
.Y(n_280)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_281),
.Y(n_301)
);

INVxp33_ASAP7_75t_SL g282 ( 
.A(n_255),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g291 ( 
.A(n_282),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_241),
.B(n_209),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_283),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_259),
.B(n_4),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_287),
.B(n_294),
.C(n_295),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_288),
.A2(n_276),
.B1(n_265),
.B2(n_6),
.Y(n_316)
);

AO21x1_ASAP7_75t_L g289 ( 
.A1(n_274),
.A2(n_249),
.B(n_250),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_289),
.B(n_272),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_L g293 ( 
.A1(n_275),
.A2(n_262),
.B(n_261),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_293),
.A2(n_297),
.B(n_269),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_265),
.B(n_240),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_L g297 ( 
.A1(n_268),
.A2(n_242),
.B(n_240),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_299),
.B(n_245),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_270),
.B(n_239),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_302),
.B(n_279),
.C(n_295),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_298),
.A2(n_267),
.B(n_271),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_303),
.A2(n_306),
.B1(n_308),
.B2(n_311),
.Y(n_329)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_305),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_307),
.B(n_309),
.C(n_312),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_291),
.A2(n_283),
.B1(n_266),
.B2(n_284),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_294),
.B(n_277),
.C(n_273),
.Y(n_309)
);

FAx1_ASAP7_75t_SL g310 ( 
.A(n_293),
.B(n_247),
.CI(n_266),
.CON(n_310),
.SN(n_310)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_310),
.B(n_313),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_L g312 ( 
.A1(n_290),
.A2(n_251),
.B(n_245),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_286),
.B(n_251),
.Y(n_313)
);

OR2x2_ASAP7_75t_L g314 ( 
.A(n_296),
.B(n_260),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_314),
.B(n_315),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_300),
.B(n_260),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_316),
.B(n_287),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_301),
.B(n_4),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_317),
.B(n_5),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_SL g318 ( 
.A1(n_303),
.A2(n_291),
.B(n_289),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g338 ( 
.A1(n_318),
.A2(n_308),
.B(n_7),
.Y(n_338)
);

BUFx24_ASAP7_75t_SL g319 ( 
.A(n_310),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_319),
.B(n_323),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_316),
.B(n_302),
.Y(n_323)
);

NAND2xp33_ASAP7_75t_SL g336 ( 
.A(n_325),
.B(n_312),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_314),
.A2(n_297),
.B1(n_288),
.B2(n_292),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_326),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_311),
.B(n_292),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_327),
.B(n_328),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_329),
.B(n_310),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_330),
.B(n_331),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_320),
.B(n_307),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_L g333 ( 
.A1(n_320),
.A2(n_309),
.B(n_304),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g340 ( 
.A(n_333),
.B(n_338),
.Y(n_340)
);

AND2x2_ASAP7_75t_L g339 ( 
.A(n_336),
.B(n_325),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_322),
.B(n_304),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_337),
.B(n_326),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_339),
.B(n_341),
.Y(n_345)
);

AND2x2_ASAP7_75t_L g341 ( 
.A(n_335),
.B(n_321),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_343),
.B(n_344),
.Y(n_347)
);

NAND3xp33_ASAP7_75t_L g344 ( 
.A(n_334),
.B(n_324),
.C(n_329),
.Y(n_344)
);

INVxp67_ASAP7_75t_L g346 ( 
.A(n_342),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_L g348 ( 
.A1(n_346),
.A2(n_332),
.B(n_340),
.Y(n_348)
);

OAI21xp5_ASAP7_75t_SL g349 ( 
.A1(n_348),
.A2(n_332),
.B(n_345),
.Y(n_349)
);

NOR3xp33_ASAP7_75t_L g350 ( 
.A(n_349),
.B(n_347),
.C(n_7),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_350),
.B(n_5),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_351),
.B(n_8),
.Y(n_352)
);


endmodule