module real_jpeg_17435_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_216;
wire n_202;
wire n_128;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_0),
.A2(n_15),
.B1(n_20),
.B2(n_21),
.Y(n_19)
);

INVx5_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_1),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_1),
.B(n_76),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_1),
.B(n_92),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_1),
.B(n_156),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g205 ( 
.A(n_1),
.B(n_206),
.Y(n_205)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_2),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g122 ( 
.A(n_2),
.Y(n_122)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_2),
.Y(n_198)
);

BUFx3_ASAP7_75t_L g272 ( 
.A(n_2),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_3),
.Y(n_101)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_3),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_4),
.B(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_4),
.B(n_98),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_4),
.A2(n_9),
.B1(n_120),
.B2(n_123),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_4),
.B(n_163),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g185 ( 
.A(n_4),
.B(n_186),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_4),
.B(n_231),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_4),
.B(n_256),
.Y(n_255)
);

AND2x2_ASAP7_75t_L g259 ( 
.A(n_4),
.B(n_260),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_4),
.B(n_298),
.Y(n_297)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_5),
.B(n_62),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_5),
.B(n_71),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_5),
.B(n_103),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_5),
.B(n_112),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_5),
.B(n_134),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g201 ( 
.A(n_5),
.B(n_202),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g269 ( 
.A(n_5),
.B(n_270),
.Y(n_269)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_6),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_6),
.Y(n_76)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_6),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_6),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g286 ( 
.A(n_6),
.Y(n_286)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_7),
.B(n_54),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_8),
.B(n_30),
.Y(n_29)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_8),
.B(n_64),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_8),
.B(n_79),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_8),
.B(n_151),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g264 ( 
.A(n_8),
.B(n_53),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_8),
.B(n_267),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_8),
.B(n_281),
.Y(n_280)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_9),
.B(n_115),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_9),
.B(n_139),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_9),
.Y(n_192)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_10),
.Y(n_42)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_10),
.Y(n_204)
);

BUFx4f_ASAP7_75t_L g322 ( 
.A(n_10),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_11),
.B(n_73),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_11),
.B(n_210),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_11),
.B(n_236),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_11),
.B(n_30),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_11),
.B(n_305),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_11),
.B(n_312),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_11),
.B(n_318),
.Y(n_317)
);

AND2x2_ASAP7_75t_L g40 ( 
.A(n_12),
.B(n_41),
.Y(n_40)
);

AND2x2_ASAP7_75t_SL g52 ( 
.A(n_12),
.B(n_53),
.Y(n_52)
);

AND2x4_ASAP7_75t_SL g84 ( 
.A(n_12),
.B(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_12),
.B(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_13),
.Y(n_60)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_14),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_14),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_14),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_14),
.Y(n_148)
);

INVx3_ASAP7_75t_L g234 ( 
.A(n_14),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_16),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_16),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_17),
.B(n_54),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_17),
.B(n_169),
.Y(n_168)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_18),
.Y(n_74)
);

BUFx5_ASAP7_75t_L g112 ( 
.A(n_18),
.Y(n_112)
);

BUFx5_ASAP7_75t_L g165 ( 
.A(n_18),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_216),
.Y(n_21)
);

AOI21xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_175),
.B(n_214),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_24),
.B(n_176),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_107),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_68),
.C(n_90),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_SL g177 ( 
.A(n_26),
.B(n_178),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_45),
.C(n_55),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

XNOR2x2_ASAP7_75t_L g241 ( 
.A(n_28),
.B(n_242),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_35),
.Y(n_28)
);

MAJx2_ASAP7_75t_L g127 ( 
.A(n_29),
.B(n_40),
.C(n_44),
.Y(n_127)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_34),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g158 ( 
.A(n_34),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g35 ( 
.A1(n_36),
.A2(n_40),
.B1(n_43),
.B2(n_44),
.Y(n_35)
);

INVx1_ASAP7_75t_SL g44 ( 
.A(n_36),
.Y(n_44)
);

OR2x2_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_38),
.Y(n_36)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_40),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_42),
.Y(n_116)
);

INVx5_ASAP7_75t_L g170 ( 
.A(n_42),
.Y(n_170)
);

INVx4_ASAP7_75t_L g268 ( 
.A(n_42),
.Y(n_268)
);

HB1xp67_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_46),
.B(n_55),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_52),
.Y(n_46)
);

XOR2xp5_ASAP7_75t_SL g240 ( 
.A(n_47),
.B(n_52),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_51),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_61),
.C(n_63),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_56),
.A2(n_61),
.B1(n_226),
.B2(n_227),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_56),
.Y(n_226)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_61),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_61),
.A2(n_227),
.B1(n_303),
.B2(n_304),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_61),
.B(n_303),
.C(n_307),
.Y(n_329)
);

XOR2x1_ASAP7_75t_L g224 ( 
.A(n_63),
.B(n_225),
.Y(n_224)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_68),
.B(n_90),
.Y(n_178)
);

XOR2x2_ASAP7_75t_SL g68 ( 
.A(n_69),
.B(n_77),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_69),
.B(n_78),
.C(n_88),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_72),
.C(n_75),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_70),
.A2(n_75),
.B1(n_182),
.B2(n_183),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_70),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_70),
.B(n_253),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_SL g180 ( 
.A(n_72),
.B(n_181),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_75),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_84),
.B1(n_88),
.B2(n_89),
.Y(n_77)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_78),
.Y(n_89)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_82),
.Y(n_190)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_84),
.Y(n_88)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_85),
.Y(n_313)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

XOR2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_96),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_91),
.B(n_97),
.C(n_105),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_102),
.B1(n_105),
.B2(n_106),
.Y(n_96)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_97),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx4_ASAP7_75t_L g210 ( 
.A(n_100),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_102),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_102),
.A2(n_105),
.B1(n_235),
.B2(n_291),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_105),
.B(n_230),
.C(n_235),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_108),
.A2(n_144),
.B1(n_173),
.B2(n_174),
.Y(n_107)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_108),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_128),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_118),
.C(n_127),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_110),
.B(n_212),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_113),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_111),
.B(n_114),
.C(n_117),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_117),
.Y(n_113)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_118),
.A2(n_119),
.B1(n_127),
.B2(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_119),
.A2(n_185),
.B(n_191),
.Y(n_184)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_126),
.Y(n_136)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_126),
.Y(n_238)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_127),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_129),
.A2(n_141),
.B1(n_142),
.B2(n_143),
.Y(n_128)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_129),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_131),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_132),
.A2(n_133),
.B1(n_137),
.B2(n_138),
.Y(n_131)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_133),
.B(n_200),
.C(n_208),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_133),
.A2(n_208),
.B1(n_209),
.B2(n_339),
.Y(n_338)
);

INVxp67_ASAP7_75t_L g339 ( 
.A(n_133),
.Y(n_339)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVxp67_ASAP7_75t_R g137 ( 
.A(n_138),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

BUFx2_ASAP7_75t_L g256 ( 
.A(n_140),
.Y(n_256)
);

INVxp67_ASAP7_75t_SL g143 ( 
.A(n_141),
.Y(n_143)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_144),
.Y(n_174)
);

XNOR2x2_ASAP7_75t_SL g144 ( 
.A(n_145),
.B(n_159),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_149),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_155),
.Y(n_149)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

BUFx2_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_161),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_166),
.Y(n_161)
);

INVx1_ASAP7_75t_SL g163 ( 
.A(n_164),
.Y(n_163)
);

INVx8_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_167),
.A2(n_168),
.B1(n_171),
.B2(n_172),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_SL g172 ( 
.A(n_171),
.Y(n_172)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_179),
.C(n_211),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_177),
.B(n_244),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_179),
.B(n_211),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_184),
.C(n_199),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_180),
.B(n_184),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_182),
.B(n_254),
.C(n_255),
.Y(n_288)
);

INVx1_ASAP7_75t_SL g186 ( 
.A(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_193),
.Y(n_191)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_197),
.Y(n_207)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_197),
.Y(n_299)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_199),
.B(n_221),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_200),
.B(n_338),
.Y(n_337)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_205),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_201),
.B(n_205),
.Y(n_279)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_201),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_201),
.A2(n_296),
.B1(n_297),
.B2(n_315),
.Y(n_314)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_204),
.Y(n_263)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_217),
.A2(n_245),
.B(n_352),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_243),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_219),
.B(n_243),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_222),
.C(n_241),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_220),
.B(n_349),
.Y(n_348)
);

HB1xp67_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_223),
.B(n_241),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_SL g223 ( 
.A(n_224),
.B(n_228),
.C(n_239),
.Y(n_223)
);

XOR2x1_ASAP7_75t_L g343 ( 
.A(n_224),
.B(n_344),
.Y(n_343)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_229),
.B(n_240),
.Y(n_344)
);

XOR2x1_ASAP7_75t_L g289 ( 
.A(n_230),
.B(n_290),
.Y(n_289)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx5_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

BUFx3_ASAP7_75t_L g306 ( 
.A(n_234),
.Y(n_306)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_235),
.Y(n_291)
);

INVx4_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

HB1xp67_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_248),
.A2(n_347),
.B(n_351),
.Y(n_247)
);

AOI21x1_ASAP7_75t_L g248 ( 
.A1(n_249),
.A2(n_332),
.B(n_346),
.Y(n_248)
);

OAI21x1_ASAP7_75t_L g249 ( 
.A1(n_250),
.A2(n_292),
.B(n_331),
.Y(n_249)
);

AND2x2_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_275),
.Y(n_250)
);

OR2x2_ASAP7_75t_L g331 ( 
.A(n_251),
.B(n_275),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_257),
.C(n_265),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_SL g326 ( 
.A(n_252),
.B(n_327),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_255),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_257),
.A2(n_258),
.B1(n_265),
.B2(n_328),
.Y(n_327)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_264),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_SL g308 ( 
.A(n_259),
.B(n_264),
.Y(n_308)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_265),
.Y(n_328)
);

AO22x1_ASAP7_75t_SL g265 ( 
.A1(n_266),
.A2(n_269),
.B1(n_273),
.B2(n_274),
.Y(n_265)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_266),
.Y(n_273)
);

INVx3_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_SL g274 ( 
.A(n_269),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_269),
.B(n_273),
.Y(n_277)
);

INVx4_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx3_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_274),
.B(n_317),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_287),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_276),
.B(n_288),
.C(n_289),
.Y(n_345)
);

XOR2x1_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_278),
.Y(n_276)
);

MAJx2_ASAP7_75t_L g341 ( 
.A(n_277),
.B(n_279),
.C(n_280),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_280),
.Y(n_278)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

HB1xp67_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx4_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx3_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx6_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_289),
.Y(n_287)
);

AOI21x1_ASAP7_75t_L g292 ( 
.A1(n_293),
.A2(n_325),
.B(n_330),
.Y(n_292)
);

OAI21x1_ASAP7_75t_SL g293 ( 
.A1(n_294),
.A2(n_309),
.B(n_324),
.Y(n_293)
);

NOR2x1_ASAP7_75t_SL g294 ( 
.A(n_295),
.B(n_300),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_295),
.B(n_300),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_297),
.Y(n_295)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_297),
.Y(n_315)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_301),
.A2(n_302),
.B1(n_307),
.B2(n_308),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

AOI21x1_ASAP7_75t_SL g309 ( 
.A1(n_310),
.A2(n_316),
.B(n_323),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_314),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_311),
.B(n_314),
.Y(n_323)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_326),
.B(n_329),
.Y(n_325)
);

NOR2x1_ASAP7_75t_SL g330 ( 
.A(n_326),
.B(n_329),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_333),
.B(n_345),
.Y(n_332)
);

NOR2x1_ASAP7_75t_L g346 ( 
.A(n_333),
.B(n_345),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_334),
.A2(n_335),
.B1(n_342),
.B2(n_343),
.Y(n_333)
);

INVxp67_ASAP7_75t_SL g334 ( 
.A(n_335),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_336),
.A2(n_337),
.B1(n_340),
.B2(n_341),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_336),
.B(n_341),
.C(n_342),
.Y(n_350)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

NOR2xp67_ASAP7_75t_L g347 ( 
.A(n_348),
.B(n_350),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_348),
.B(n_350),
.Y(n_351)
);

INVxp67_ASAP7_75t_SL g352 ( 
.A(n_353),
.Y(n_352)
);


endmodule