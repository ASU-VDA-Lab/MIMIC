module fake_jpeg_14106_n_25 (n_3, n_2, n_1, n_0, n_4, n_5, n_25);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_25;

wire n_13;
wire n_21;
wire n_10;
wire n_23;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_16;
wire n_24;
wire n_9;
wire n_11;
wire n_17;
wire n_12;
wire n_8;
wire n_15;
wire n_7;

OAI22xp5_ASAP7_75t_L g6 ( 
.A1(n_1),
.A2(n_5),
.B1(n_3),
.B2(n_4),
.Y(n_6)
);

OAI22xp5_ASAP7_75t_SL g7 ( 
.A1(n_0),
.A2(n_1),
.B1(n_2),
.B2(n_5),
.Y(n_7)
);

OAI22xp5_ASAP7_75t_SL g8 ( 
.A1(n_4),
.A2(n_0),
.B1(n_3),
.B2(n_5),
.Y(n_8)
);

NAND2xp5_ASAP7_75t_L g9 ( 
.A(n_3),
.B(n_4),
.Y(n_9)
);

OR2x2_ASAP7_75t_L g10 ( 
.A(n_1),
.B(n_2),
.Y(n_10)
);

INVx2_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

INVx11_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

OAI22xp5_ASAP7_75t_L g13 ( 
.A1(n_9),
.A2(n_0),
.B1(n_1),
.B2(n_10),
.Y(n_13)
);

AOI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_13),
.A2(n_15),
.B1(n_17),
.B2(n_7),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_14),
.B(n_16),
.Y(n_19)
);

O2A1O1Ixp33_ASAP7_75t_L g15 ( 
.A1(n_9),
.A2(n_10),
.B(n_12),
.C(n_8),
.Y(n_15)
);

AND2x2_ASAP7_75t_SL g16 ( 
.A(n_7),
.B(n_8),
.Y(n_16)
);

AND2x2_ASAP7_75t_L g17 ( 
.A(n_10),
.B(n_11),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_13),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_18),
.B(n_16),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_20),
.B(n_6),
.C(n_7),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_21),
.B(n_22),
.C(n_12),
.Y(n_24)
);

O2A1O1Ixp33_ASAP7_75t_SL g23 ( 
.A1(n_21),
.A2(n_20),
.B(n_19),
.C(n_6),
.Y(n_23)
);

OAI31xp67_ASAP7_75t_L g25 ( 
.A1(n_23),
.A2(n_24),
.A3(n_12),
.B(n_11),
.Y(n_25)
);


endmodule