module fake_jpeg_29691_n_174 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_174);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_174;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_120;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_10),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_33),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_13),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_7),
.Y(n_56)
);

INVx13_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

INVx1_ASAP7_75t_SL g58 ( 
.A(n_0),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_9),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_30),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_31),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_15),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_14),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_20),
.Y(n_68)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_34),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_43),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_28),
.Y(n_71)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_4),
.Y(n_72)
);

CKINVDCx14_ASAP7_75t_R g73 ( 
.A(n_51),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_57),
.Y(n_74)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_74),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_58),
.B(n_0),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_75),
.B(n_80),
.Y(n_85)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_67),
.Y(n_76)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_76),
.Y(n_94)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_72),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_77),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_52),
.B(n_1),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_78),
.B(n_83),
.Y(n_93)
);

NAND2x1_ASAP7_75t_SL g79 ( 
.A(n_58),
.B(n_1),
.Y(n_79)
);

OR2x2_ASAP7_75t_L g91 ( 
.A(n_79),
.B(n_82),
.Y(n_91)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_72),
.Y(n_80)
);

INVx11_ASAP7_75t_L g81 ( 
.A(n_63),
.Y(n_81)
);

INVx2_ASAP7_75t_SL g96 ( 
.A(n_81),
.Y(n_96)
);

OR2x4_ASAP7_75t_L g82 ( 
.A(n_56),
.B(n_2),
.Y(n_82)
);

INVx2_ASAP7_75t_SL g83 ( 
.A(n_67),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_79),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_84),
.B(n_86),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_83),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_80),
.A2(n_63),
.B1(n_66),
.B2(n_69),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_87),
.A2(n_64),
.B1(n_60),
.B2(n_68),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_82),
.A2(n_66),
.B1(n_69),
.B2(n_68),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_88),
.A2(n_70),
.B1(n_62),
.B2(n_55),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_74),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_90),
.B(n_92),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_81),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_76),
.B(n_73),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_95),
.B(n_64),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_78),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_98),
.B(n_3),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_99),
.B(n_102),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_91),
.A2(n_71),
.B1(n_54),
.B2(n_59),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_101),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_91),
.A2(n_64),
.B(n_60),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_97),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_103),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_85),
.B(n_93),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_104),
.B(n_113),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_105),
.A2(n_107),
.B1(n_25),
.B2(n_47),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_94),
.A2(n_65),
.B(n_61),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_106),
.B(n_19),
.Y(n_130)
);

OAI21xp33_ASAP7_75t_L g108 ( 
.A1(n_97),
.A2(n_57),
.B(n_53),
.Y(n_108)
);

O2A1O1Ixp33_ASAP7_75t_L g127 ( 
.A1(n_108),
.A2(n_11),
.B(n_12),
.C(n_16),
.Y(n_127)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_89),
.Y(n_109)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_109),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_87),
.B(n_2),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_111),
.B(n_29),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_112),
.B(n_115),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_86),
.B(n_3),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_89),
.B(n_4),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_114),
.B(n_117),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_96),
.B(n_5),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_96),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_116),
.B(n_6),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_98),
.B(n_5),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_108),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_119),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_120),
.A2(n_128),
.B1(n_133),
.B2(n_41),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_122),
.B(n_123),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_100),
.B(n_8),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_110),
.B(n_9),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_124),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_101),
.B(n_10),
.Y(n_125)
);

NOR4xp25_ASAP7_75t_L g151 ( 
.A(n_125),
.B(n_129),
.C(n_121),
.D(n_127),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_127),
.A2(n_32),
.B1(n_37),
.B2(n_38),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_111),
.A2(n_11),
.B1(n_17),
.B2(n_18),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_102),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_130),
.B(n_138),
.Y(n_148)
);

INVx13_ASAP7_75t_L g131 ( 
.A(n_103),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_105),
.A2(n_21),
.B1(n_22),
.B2(n_23),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_100),
.A2(n_24),
.B(n_26),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_136),
.B(n_139),
.C(n_132),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_104),
.B(n_27),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_139),
.B(n_46),
.Y(n_150)
);

HB1xp67_ASAP7_75t_L g140 ( 
.A(n_126),
.Y(n_140)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_140),
.Y(n_157)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_137),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_141),
.B(n_143),
.Y(n_159)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_126),
.Y(n_142)
);

HB1xp67_ASAP7_75t_L g158 ( 
.A(n_142),
.Y(n_158)
);

NAND3xp33_ASAP7_75t_L g163 ( 
.A(n_144),
.B(n_145),
.C(n_149),
.Y(n_163)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_118),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_118),
.A2(n_49),
.B1(n_44),
.B2(n_45),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_146),
.A2(n_151),
.B1(n_155),
.B2(n_147),
.Y(n_162)
);

NOR2xp67_ASAP7_75t_L g149 ( 
.A(n_132),
.B(n_42),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_150),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_153),
.Y(n_161)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_131),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_154),
.A2(n_119),
.B1(n_134),
.B2(n_135),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_160),
.B(n_162),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_161),
.B(n_148),
.C(n_155),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_165),
.B(n_167),
.Y(n_168)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_157),
.Y(n_166)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_166),
.Y(n_169)
);

HB1xp67_ASAP7_75t_L g167 ( 
.A(n_158),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_168),
.B(n_159),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_170),
.A2(n_164),
.B(n_169),
.Y(n_171)
);

NAND2xp33_ASAP7_75t_SL g172 ( 
.A(n_171),
.B(n_163),
.Y(n_172)
);

NAND2x1_ASAP7_75t_L g173 ( 
.A(n_172),
.B(n_156),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_173),
.B(n_152),
.Y(n_174)
);


endmodule