module real_aes_2235_n_77 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_527, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_77);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_527;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_77;
wire n_480;
wire n_113;
wire n_476;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_522;
wire n_485;
wire n_222;
wire n_503;
wire n_287;
wire n_357;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_341;
wire n_232;
wire n_460;
wire n_401;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_320;
wire n_260;
wire n_97;
wire n_186;
wire n_138;
wire n_379;
wire n_453;
wire n_374;
wire n_235;
wire n_399;
wire n_378;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_145;
wire n_415;
wire n_227;
wire n_92;
wire n_519;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_292;
wire n_400;
wire n_116;
wire n_94;
wire n_289;
wire n_462;
wire n_280;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_408;
wire n_184;
wire n_372;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_104;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_506;
wire n_513;
wire n_297;
wire n_383;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_164;
wire n_231;
wire n_102;
wire n_454;
wire n_122;
wire n_443;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_204;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_331;
wire n_93;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_323;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_368;
wire n_505;
wire n_434;
wire n_502;
wire n_250;
wire n_85;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_402;
wire n_87;
wire n_171;
wire n_78;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_501;
wire n_488;
wire n_251;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_158;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_109;
wire n_203;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_155;
wire n_243;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_446;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_180;
wire n_212;
wire n_210;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_103;
wire n_166;
wire n_224;
wire n_151;
wire n_130;
wire n_253;
wire n_459;
wire n_99;
wire n_440;
wire n_525;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_305;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_473;
wire n_465;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_340;
wire n_483;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_206;
wire n_307;
wire n_500;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_264;
wire n_237;
wire n_91;
AO22x2_ASAP7_75t_L g91 ( .A1(n_0), .A2(n_49), .B1(n_88), .B2(n_92), .Y(n_91) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_1), .B(n_164), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_2), .B(n_179), .Y(n_259) );
INVx1_ASAP7_75t_L g152 ( .A(n_3), .Y(n_152) );
OAI22xp5_ASAP7_75t_SL g495 ( .A1(n_4), .A2(n_496), .B1(n_497), .B2(n_498), .Y(n_495) );
INVx1_ASAP7_75t_L g498 ( .A(n_4), .Y(n_498) );
INVx1_ASAP7_75t_L g497 ( .A(n_5), .Y(n_497) );
AO22x2_ASAP7_75t_L g87 ( .A1(n_6), .A2(n_15), .B1(n_88), .B2(n_89), .Y(n_87) );
AND2x2_ASAP7_75t_L g199 ( .A(n_7), .B(n_200), .Y(n_199) );
AND2x2_ASAP7_75t_L g261 ( .A(n_8), .B(n_188), .Y(n_261) );
INVx2_ASAP7_75t_L g185 ( .A(n_9), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_10), .B(n_179), .Y(n_233) );
INVx1_ASAP7_75t_L g488 ( .A(n_11), .Y(n_488) );
NAND2xp5_ASAP7_75t_SL g266 ( .A(n_12), .B(n_164), .Y(n_266) );
INVx1_ASAP7_75t_L g525 ( .A(n_12), .Y(n_525) );
AOI22xp33_ASAP7_75t_L g204 ( .A1(n_13), .A2(n_70), .B1(n_164), .B2(n_205), .Y(n_204) );
INVx1_ASAP7_75t_L g489 ( .A(n_14), .Y(n_489) );
OAI221xp5_ASAP7_75t_L g504 ( .A1(n_15), .A2(n_49), .B1(n_54), .B2(n_505), .C(n_507), .Y(n_504) );
OR2x2_ASAP7_75t_L g186 ( .A(n_16), .B(n_69), .Y(n_186) );
OA21x2_ASAP7_75t_L g189 ( .A1(n_16), .A2(n_69), .B(n_185), .Y(n_189) );
INVx3_ASAP7_75t_L g88 ( .A(n_17), .Y(n_88) );
AO21x2_ASAP7_75t_L g228 ( .A1(n_18), .A2(n_200), .B(n_229), .Y(n_228) );
AOI22xp33_ASAP7_75t_L g111 ( .A1(n_19), .A2(n_44), .B1(n_112), .B2(n_114), .Y(n_111) );
AOI21xp5_ASAP7_75t_L g256 ( .A1(n_20), .A2(n_172), .B(n_257), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_21), .B(n_179), .Y(n_241) );
INVx1_ASAP7_75t_SL g99 ( .A(n_22), .Y(n_99) );
INVx1_ASAP7_75t_L g154 ( .A(n_23), .Y(n_154) );
AND2x2_ASAP7_75t_L g170 ( .A(n_23), .B(n_152), .Y(n_170) );
AND2x2_ASAP7_75t_L g173 ( .A(n_23), .B(n_174), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_24), .B(n_164), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_25), .B(n_179), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_26), .B(n_164), .Y(n_163) );
AOI21xp5_ASAP7_75t_L g194 ( .A1(n_27), .A2(n_172), .B(n_195), .Y(n_194) );
AO22x2_ASAP7_75t_L g94 ( .A1(n_28), .A2(n_54), .B1(n_88), .B2(n_95), .Y(n_94) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_29), .B(n_181), .Y(n_180) );
NAND2xp5_ASAP7_75t_SL g230 ( .A(n_30), .B(n_164), .Y(n_230) );
INVx1_ASAP7_75t_L g167 ( .A(n_31), .Y(n_167) );
INVx1_ASAP7_75t_L g176 ( .A(n_31), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_32), .B(n_179), .Y(n_197) );
AND2x2_ASAP7_75t_L g218 ( .A(n_33), .B(n_183), .Y(n_218) );
INVx1_ASAP7_75t_L g100 ( .A(n_34), .Y(n_100) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_35), .B(n_181), .Y(n_196) );
AOI22xp33_ASAP7_75t_L g130 ( .A1(n_36), .A2(n_65), .B1(n_131), .B2(n_134), .Y(n_130) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_37), .B(n_181), .Y(n_240) );
NAND2xp5_ASAP7_75t_SL g198 ( .A(n_38), .B(n_164), .Y(n_198) );
AOI22xp33_ASAP7_75t_L g115 ( .A1(n_39), .A2(n_63), .B1(n_116), .B2(n_119), .Y(n_115) );
AOI22xp33_ASAP7_75t_L g106 ( .A1(n_40), .A2(n_48), .B1(n_107), .B2(n_108), .Y(n_106) );
NAND2xp5_ASAP7_75t_SL g220 ( .A(n_41), .B(n_164), .Y(n_220) );
AOI21xp5_ASAP7_75t_L g238 ( .A1(n_42), .A2(n_172), .B(n_239), .Y(n_238) );
AND2x2_ASAP7_75t_L g272 ( .A(n_43), .B(n_184), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_45), .B(n_181), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_46), .B(n_181), .Y(n_234) );
AOI22xp5_ASAP7_75t_L g492 ( .A1(n_46), .A2(n_493), .B1(n_494), .B2(n_495), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_46), .Y(n_493) );
AOI22xp5_ASAP7_75t_L g209 ( .A1(n_47), .A2(n_71), .B1(n_172), .B2(n_210), .Y(n_209) );
INVxp33_ASAP7_75t_L g509 ( .A(n_49), .Y(n_509) );
AOI22xp33_ASAP7_75t_SL g122 ( .A1(n_50), .A2(n_66), .B1(n_123), .B2(n_127), .Y(n_122) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_51), .B(n_179), .Y(n_269) );
INVx1_ASAP7_75t_L g169 ( .A(n_52), .Y(n_169) );
INVx1_ASAP7_75t_L g174 ( .A(n_52), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_53), .B(n_181), .Y(n_258) );
INVxp67_ASAP7_75t_L g508 ( .A(n_54), .Y(n_508) );
AOI21xp5_ASAP7_75t_L g221 ( .A1(n_55), .A2(n_172), .B(n_222), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_56), .B(n_144), .Y(n_143) );
AOI21xp5_ASAP7_75t_L g171 ( .A1(n_57), .A2(n_172), .B(n_177), .Y(n_171) );
AOI21xp5_ASAP7_75t_L g231 ( .A1(n_58), .A2(n_172), .B(n_232), .Y(n_231) );
AND2x2_ASAP7_75t_L g243 ( .A(n_59), .B(n_184), .Y(n_243) );
AOI22xp5_ASAP7_75t_L g79 ( .A1(n_60), .A2(n_80), .B1(n_147), .B2(n_148), .Y(n_79) );
CKINVDCx20_ASAP7_75t_R g147 ( .A(n_60), .Y(n_147) );
AOI22xp33_ASAP7_75t_L g139 ( .A1(n_61), .A2(n_67), .B1(n_140), .B2(n_141), .Y(n_139) );
NAND2xp5_ASAP7_75t_SL g202 ( .A(n_62), .B(n_183), .Y(n_202) );
AND2x2_ASAP7_75t_L g187 ( .A(n_64), .B(n_188), .Y(n_187) );
AOI22xp33_ASAP7_75t_L g83 ( .A1(n_68), .A2(n_73), .B1(n_84), .B2(n_101), .Y(n_83) );
AOI21xp5_ASAP7_75t_L g267 ( .A1(n_72), .A2(n_172), .B(n_268), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_74), .B(n_179), .Y(n_178) );
BUFx2_ASAP7_75t_L g271 ( .A(n_75), .Y(n_271) );
BUFx2_ASAP7_75t_SL g506 ( .A(n_76), .Y(n_506) );
AOI221xp5_ASAP7_75t_L g77 ( .A1(n_78), .A2(n_149), .B1(n_155), .B2(n_483), .C(n_484), .Y(n_77) );
INVxp67_ASAP7_75t_L g78 ( .A(n_79), .Y(n_78) );
CKINVDCx20_ASAP7_75t_R g148 ( .A(n_80), .Y(n_148) );
OAI222xp33_ASAP7_75t_L g484 ( .A1(n_80), .A2(n_148), .B1(n_485), .B2(n_517), .C1(n_520), .C2(n_525), .Y(n_484) );
HB1xp67_ASAP7_75t_L g80 ( .A(n_81), .Y(n_80) );
NOR3xp33_ASAP7_75t_L g81 ( .A(n_82), .B(n_121), .C(n_138), .Y(n_81) );
NAND4xp25_ASAP7_75t_L g82 ( .A(n_83), .B(n_106), .C(n_111), .D(n_115), .Y(n_82) );
AND2x6_ASAP7_75t_L g84 ( .A(n_85), .B(n_93), .Y(n_84) );
AND2x2_ASAP7_75t_L g112 ( .A(n_85), .B(n_113), .Y(n_112) );
AND2x4_ASAP7_75t_L g118 ( .A(n_85), .B(n_102), .Y(n_118) );
AND2x2_ASAP7_75t_L g146 ( .A(n_85), .B(n_137), .Y(n_146) );
AND2x4_ASAP7_75t_L g85 ( .A(n_86), .B(n_90), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_87), .Y(n_86) );
INVx1_ASAP7_75t_L g105 ( .A(n_87), .Y(n_105) );
AND2x2_ASAP7_75t_L g110 ( .A(n_87), .B(n_91), .Y(n_110) );
AND2x4_ASAP7_75t_L g120 ( .A(n_87), .B(n_90), .Y(n_120) );
INVx2_ASAP7_75t_L g89 ( .A(n_88), .Y(n_89) );
INVx1_ASAP7_75t_L g92 ( .A(n_88), .Y(n_92) );
INVx1_ASAP7_75t_L g95 ( .A(n_88), .Y(n_95) );
OAI22x1_ASAP7_75t_L g97 ( .A1(n_88), .A2(n_98), .B1(n_99), .B2(n_100), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_88), .Y(n_98) );
INVxp67_ASAP7_75t_L g142 ( .A(n_90), .Y(n_142) );
INVx2_ASAP7_75t_L g90 ( .A(n_91), .Y(n_90) );
AND2x2_ASAP7_75t_L g104 ( .A(n_91), .B(n_105), .Y(n_104) );
AND2x2_ASAP7_75t_L g107 ( .A(n_93), .B(n_104), .Y(n_107) );
AND2x2_ASAP7_75t_L g140 ( .A(n_93), .B(n_120), .Y(n_140) );
AND2x2_ASAP7_75t_L g93 ( .A(n_94), .B(n_96), .Y(n_93) );
INVx2_ASAP7_75t_L g103 ( .A(n_94), .Y(n_103) );
BUFx2_ASAP7_75t_L g109 ( .A(n_94), .Y(n_109) );
AND2x2_ASAP7_75t_L g137 ( .A(n_94), .B(n_97), .Y(n_137) );
AND2x4_ASAP7_75t_L g102 ( .A(n_96), .B(n_103), .Y(n_102) );
INVx2_ASAP7_75t_L g96 ( .A(n_97), .Y(n_96) );
AND2x2_ASAP7_75t_L g113 ( .A(n_97), .B(n_103), .Y(n_113) );
HB1xp67_ASAP7_75t_L g126 ( .A(n_97), .Y(n_126) );
AND2x6_ASAP7_75t_L g101 ( .A(n_102), .B(n_104), .Y(n_101) );
AND2x4_ASAP7_75t_L g114 ( .A(n_102), .B(n_110), .Y(n_114) );
AND2x4_ASAP7_75t_L g119 ( .A(n_102), .B(n_120), .Y(n_119) );
AND2x2_ASAP7_75t_L g133 ( .A(n_104), .B(n_113), .Y(n_133) );
HB1xp67_ASAP7_75t_L g136 ( .A(n_105), .Y(n_136) );
AND2x4_ASAP7_75t_L g108 ( .A(n_109), .B(n_110), .Y(n_108) );
AND2x2_ASAP7_75t_L g125 ( .A(n_110), .B(n_126), .Y(n_125) );
AND2x2_ASAP7_75t_L g129 ( .A(n_113), .B(n_120), .Y(n_129) );
INVx3_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
INVx8_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
NAND2xp5_ASAP7_75t_L g121 ( .A(n_122), .B(n_130), .Y(n_121) );
INVx2_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
INVx3_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
INVx2_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
INVx2_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
INVx4_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
INVx3_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
AND2x2_ASAP7_75t_L g134 ( .A(n_135), .B(n_137), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
AND2x2_ASAP7_75t_L g141 ( .A(n_137), .B(n_142), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g138 ( .A(n_139), .B(n_143), .Y(n_138) );
INVx4_ASAP7_75t_SL g144 ( .A(n_145), .Y(n_144) );
INVx6_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx2_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
OR2x2_ASAP7_75t_SL g150 ( .A(n_151), .B(n_153), .Y(n_150) );
AND2x2_ASAP7_75t_L g206 ( .A(n_151), .B(n_207), .Y(n_206) );
INVx1_ASAP7_75t_L g510 ( .A(n_151), .Y(n_510) );
HB1xp67_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
AND2x2_ASAP7_75t_L g175 ( .A(n_152), .B(n_176), .Y(n_175) );
AND3x1_ASAP7_75t_SL g503 ( .A(n_153), .B(n_504), .C(n_510), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_153), .B(n_516), .Y(n_515) );
INVx1_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
NOR2x1p5_ASAP7_75t_L g211 ( .A(n_154), .B(n_212), .Y(n_211) );
INVx3_ASAP7_75t_SL g155 ( .A(n_156), .Y(n_155) );
AND2x4_ASAP7_75t_SL g156 ( .A(n_157), .B(n_379), .Y(n_156) );
NOR3xp33_ASAP7_75t_SL g157 ( .A(n_158), .B(n_288), .C(n_320), .Y(n_157) );
OAI221xp5_ASAP7_75t_L g158 ( .A1(n_159), .A2(n_214), .B1(n_244), .B2(n_262), .C(n_273), .Y(n_158) );
OR2x2_ASAP7_75t_L g159 ( .A(n_160), .B(n_190), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
AND2x2_ASAP7_75t_L g250 ( .A(n_161), .B(n_191), .Y(n_250) );
INVx4_ASAP7_75t_L g279 ( .A(n_161), .Y(n_279) );
AND2x4_ASAP7_75t_SL g319 ( .A(n_161), .B(n_252), .Y(n_319) );
BUFx2_ASAP7_75t_L g329 ( .A(n_161), .Y(n_329) );
NOR2x1_ASAP7_75t_L g395 ( .A(n_161), .B(n_334), .Y(n_395) );
AND2x2_ASAP7_75t_L g404 ( .A(n_161), .B(n_332), .Y(n_404) );
OR2x2_ASAP7_75t_L g412 ( .A(n_161), .B(n_413), .Y(n_412) );
AND2x2_ASAP7_75t_L g438 ( .A(n_161), .B(n_277), .Y(n_438) );
AND2x4_ASAP7_75t_L g457 ( .A(n_161), .B(n_458), .Y(n_457) );
OR2x6_ASAP7_75t_L g161 ( .A(n_162), .B(n_187), .Y(n_161) );
AOI21xp5_ASAP7_75t_L g162 ( .A1(n_163), .A2(n_171), .B(n_183), .Y(n_162) );
HB1xp67_ASAP7_75t_L g483 ( .A(n_164), .Y(n_483) );
AND2x4_ASAP7_75t_L g164 ( .A(n_165), .B(n_170), .Y(n_164) );
AND2x4_ASAP7_75t_L g165 ( .A(n_166), .B(n_168), .Y(n_165) );
AND2x6_ASAP7_75t_L g181 ( .A(n_166), .B(n_174), .Y(n_181) );
INVx2_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
AND2x4_ASAP7_75t_L g179 ( .A(n_168), .B(n_176), .Y(n_179) );
INVx2_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
INVx5_ASAP7_75t_L g182 ( .A(n_170), .Y(n_182) );
AND2x6_ASAP7_75t_L g172 ( .A(n_173), .B(n_175), .Y(n_172) );
BUFx3_ASAP7_75t_L g208 ( .A(n_173), .Y(n_208) );
INVx2_ASAP7_75t_L g213 ( .A(n_174), .Y(n_213) );
AND2x4_ASAP7_75t_L g210 ( .A(n_175), .B(n_211), .Y(n_210) );
INVx2_ASAP7_75t_L g207 ( .A(n_176), .Y(n_207) );
AOI21xp5_ASAP7_75t_L g177 ( .A1(n_178), .A2(n_180), .B(n_182), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_181), .B(n_271), .Y(n_270) );
AOI21xp5_ASAP7_75t_L g195 ( .A1(n_182), .A2(n_196), .B(n_197), .Y(n_195) );
AOI21xp5_ASAP7_75t_L g222 ( .A1(n_182), .A2(n_223), .B(n_224), .Y(n_222) );
AOI21xp5_ASAP7_75t_L g232 ( .A1(n_182), .A2(n_233), .B(n_234), .Y(n_232) );
AOI21xp5_ASAP7_75t_L g239 ( .A1(n_182), .A2(n_240), .B(n_241), .Y(n_239) );
AOI21xp5_ASAP7_75t_L g257 ( .A1(n_182), .A2(n_258), .B(n_259), .Y(n_257) );
AOI21xp5_ASAP7_75t_L g268 ( .A1(n_182), .A2(n_269), .B(n_270), .Y(n_268) );
AO21x2_ASAP7_75t_L g203 ( .A1(n_183), .A2(n_204), .B(n_209), .Y(n_203) );
CKINVDCx5p33_ASAP7_75t_R g254 ( .A(n_183), .Y(n_254) );
BUFx6f_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
AND2x2_ASAP7_75t_SL g184 ( .A(n_185), .B(n_186), .Y(n_184) );
AND2x4_ASAP7_75t_L g225 ( .A(n_185), .B(n_186), .Y(n_225) );
AOI21xp5_ASAP7_75t_L g265 ( .A1(n_188), .A2(n_266), .B(n_267), .Y(n_265) );
BUFx4f_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
INVx3_ASAP7_75t_L g192 ( .A(n_189), .Y(n_192) );
INVx2_ASAP7_75t_SL g370 ( .A(n_190), .Y(n_370) );
OR2x2_ASAP7_75t_L g190 ( .A(n_191), .B(n_201), .Y(n_190) );
AND2x2_ASAP7_75t_L g277 ( .A(n_191), .B(n_253), .Y(n_277) );
INVx2_ASAP7_75t_L g304 ( .A(n_191), .Y(n_304) );
INVx2_ASAP7_75t_L g334 ( .A(n_191), .Y(n_334) );
AND2x2_ASAP7_75t_L g348 ( .A(n_191), .B(n_252), .Y(n_348) );
AO21x2_ASAP7_75t_L g191 ( .A1(n_192), .A2(n_193), .B(n_199), .Y(n_191) );
INVx4_ASAP7_75t_L g200 ( .A(n_192), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_194), .B(n_198), .Y(n_193) );
INVx3_ASAP7_75t_L g236 ( .A(n_200), .Y(n_236) );
AND2x2_ASAP7_75t_L g278 ( .A(n_201), .B(n_279), .Y(n_278) );
INVx2_ASAP7_75t_L g301 ( .A(n_201), .Y(n_301) );
BUFx3_ASAP7_75t_L g315 ( .A(n_201), .Y(n_315) );
AND2x2_ASAP7_75t_L g344 ( .A(n_201), .B(n_345), .Y(n_344) );
AND2x4_ASAP7_75t_L g201 ( .A(n_202), .B(n_203), .Y(n_201) );
AND2x4_ASAP7_75t_L g248 ( .A(n_202), .B(n_203), .Y(n_248) );
AND2x4_ASAP7_75t_L g205 ( .A(n_206), .B(n_208), .Y(n_205) );
HB1xp67_ASAP7_75t_L g524 ( .A(n_207), .Y(n_524) );
HB1xp67_ASAP7_75t_L g523 ( .A(n_211), .Y(n_523) );
INVx3_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
INVx1_ASAP7_75t_L g350 ( .A(n_214), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_215), .B(n_226), .Y(n_214) );
OR2x2_ASAP7_75t_L g461 ( .A(n_215), .B(n_262), .Y(n_461) );
INVx2_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
AND2x2_ASAP7_75t_L g317 ( .A(n_216), .B(n_318), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_216), .B(n_226), .Y(n_378) );
OR2x2_ASAP7_75t_L g476 ( .A(n_216), .B(n_398), .Y(n_476) );
INVx2_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
AND2x2_ASAP7_75t_L g287 ( .A(n_217), .B(n_263), .Y(n_287) );
OR2x2_ASAP7_75t_SL g297 ( .A(n_217), .B(n_298), .Y(n_297) );
INVx4_ASAP7_75t_L g308 ( .A(n_217), .Y(n_308) );
HB1xp67_ASAP7_75t_L g359 ( .A(n_217), .Y(n_359) );
NAND2x1_ASAP7_75t_L g365 ( .A(n_217), .B(n_264), .Y(n_365) );
AND2x2_ASAP7_75t_L g390 ( .A(n_217), .B(n_228), .Y(n_390) );
OR2x2_ASAP7_75t_L g411 ( .A(n_217), .B(n_294), .Y(n_411) );
OR2x6_ASAP7_75t_L g217 ( .A(n_218), .B(n_219), .Y(n_217) );
AOI21xp5_ASAP7_75t_L g219 ( .A1(n_220), .A2(n_221), .B(n_225), .Y(n_219) );
AOI21xp5_ASAP7_75t_L g229 ( .A1(n_225), .A2(n_230), .B(n_231), .Y(n_229) );
INVx1_ASAP7_75t_L g306 ( .A(n_226), .Y(n_306) );
O2A1O1Ixp33_ASAP7_75t_L g399 ( .A1(n_226), .A2(n_400), .B(n_403), .C(n_405), .Y(n_399) );
AND2x2_ASAP7_75t_L g472 ( .A(n_226), .B(n_247), .Y(n_472) );
AND2x2_ASAP7_75t_L g226 ( .A(n_227), .B(n_235), .Y(n_226) );
INVx1_ASAP7_75t_L g339 ( .A(n_227), .Y(n_339) );
AND2x2_ASAP7_75t_L g409 ( .A(n_227), .B(n_264), .Y(n_409) );
INVx2_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
INVx1_ASAP7_75t_L g283 ( .A(n_228), .Y(n_283) );
OR2x2_ASAP7_75t_L g298 ( .A(n_228), .B(n_264), .Y(n_298) );
INVx1_ASAP7_75t_L g314 ( .A(n_228), .Y(n_314) );
AND2x2_ASAP7_75t_L g326 ( .A(n_228), .B(n_235), .Y(n_326) );
HB1xp67_ASAP7_75t_L g432 ( .A(n_228), .Y(n_432) );
NOR2x1_ASAP7_75t_SL g263 ( .A(n_235), .B(n_264), .Y(n_263) );
AO21x1_ASAP7_75t_SL g235 ( .A1(n_236), .A2(n_237), .B(n_243), .Y(n_235) );
AO21x2_ASAP7_75t_L g295 ( .A1(n_236), .A2(n_237), .B(n_243), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_238), .B(n_242), .Y(n_237) );
INVxp67_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
AND2x2_ASAP7_75t_L g245 ( .A(n_246), .B(n_249), .Y(n_245) );
OR2x2_ASAP7_75t_L g396 ( .A(n_246), .B(n_331), .Y(n_396) );
INVx2_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_247), .B(n_414), .Y(n_413) );
OR2x2_ASAP7_75t_L g478 ( .A(n_247), .B(n_375), .Y(n_478) );
INVx3_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
AND2x2_ASAP7_75t_L g323 ( .A(n_248), .B(n_304), .Y(n_323) );
AND2x2_ASAP7_75t_L g419 ( .A(n_248), .B(n_332), .Y(n_419) );
INVx1_ASAP7_75t_L g336 ( .A(n_249), .Y(n_336) );
AND2x2_ASAP7_75t_L g249 ( .A(n_250), .B(n_251), .Y(n_249) );
INVx1_ASAP7_75t_L g386 ( .A(n_250), .Y(n_386) );
INVx2_ASAP7_75t_L g353 ( .A(n_251), .Y(n_353) );
HB1xp67_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
AND2x2_ASAP7_75t_L g303 ( .A(n_252), .B(n_304), .Y(n_303) );
INVx2_ASAP7_75t_L g333 ( .A(n_252), .Y(n_333) );
INVx1_ASAP7_75t_L g458 ( .A(n_252), .Y(n_458) );
INVx3_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
HB1xp67_ASAP7_75t_L g415 ( .A(n_253), .Y(n_415) );
AOI21x1_ASAP7_75t_L g253 ( .A1(n_254), .A2(n_255), .B(n_261), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_256), .B(n_260), .Y(n_255) );
OR2x2_ASAP7_75t_L g429 ( .A(n_262), .B(n_430), .Y(n_429) );
INVx2_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
INVx2_ASAP7_75t_SL g284 ( .A(n_264), .Y(n_284) );
OR2x2_ASAP7_75t_L g307 ( .A(n_264), .B(n_308), .Y(n_307) );
AND2x2_ASAP7_75t_L g318 ( .A(n_264), .B(n_294), .Y(n_318) );
AND2x2_ASAP7_75t_L g392 ( .A(n_264), .B(n_308), .Y(n_392) );
BUFx2_ASAP7_75t_L g475 ( .A(n_264), .Y(n_475) );
OR2x6_ASAP7_75t_L g264 ( .A(n_265), .B(n_272), .Y(n_264) );
CKINVDCx16_ASAP7_75t_R g511 ( .A(n_271), .Y(n_511) );
AOI22xp5_ASAP7_75t_L g517 ( .A1(n_271), .A2(n_503), .B1(n_518), .B2(n_519), .Y(n_517) );
AOI21xp5_ASAP7_75t_L g273 ( .A1(n_274), .A2(n_280), .B(n_285), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_276), .B(n_278), .Y(n_275) );
AND2x2_ASAP7_75t_L g427 ( .A(n_276), .B(n_349), .Y(n_427) );
BUFx2_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
AND2x2_ASAP7_75t_L g286 ( .A(n_277), .B(n_279), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_278), .B(n_348), .Y(n_449) );
INVx1_ASAP7_75t_L g479 ( .A(n_278), .Y(n_479) );
NAND2x1p5_ASAP7_75t_L g375 ( .A(n_279), .B(n_376), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_279), .B(n_415), .Y(n_452) );
INVxp67_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_282), .B(n_284), .Y(n_281) );
AND2x4_ASAP7_75t_SL g316 ( .A(n_282), .B(n_317), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_282), .B(n_310), .Y(n_463) );
INVx3_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
NOR2xp33_ASAP7_75t_L g421 ( .A(n_283), .B(n_365), .Y(n_421) );
AND2x2_ASAP7_75t_L g439 ( .A(n_283), .B(n_392), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_284), .B(n_326), .Y(n_342) );
A2O1A1Ixp33_ASAP7_75t_L g371 ( .A1(n_284), .A2(n_330), .B(n_372), .C(n_377), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_284), .B(n_402), .Y(n_401) );
AND2x2_ASAP7_75t_L g285 ( .A(n_286), .B(n_287), .Y(n_285) );
AOI221xp5_ASAP7_75t_L g466 ( .A1(n_286), .A2(n_359), .B1(n_467), .B2(n_473), .C(n_477), .Y(n_466) );
INVx1_ASAP7_75t_SL g454 ( .A(n_287), .Y(n_454) );
OAI221xp5_ASAP7_75t_L g288 ( .A1(n_289), .A2(n_299), .B1(n_305), .B2(n_309), .C(n_527), .Y(n_288) );
INVx2_ASAP7_75t_SL g289 ( .A(n_290), .Y(n_289) );
AND2x4_ASAP7_75t_L g290 ( .A(n_291), .B(n_296), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
INVx1_ASAP7_75t_L g364 ( .A(n_293), .Y(n_364) );
HB1xp67_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
AND2x2_ASAP7_75t_L g338 ( .A(n_294), .B(n_339), .Y(n_338) );
AND2x2_ASAP7_75t_L g369 ( .A(n_294), .B(n_314), .Y(n_369) );
INVx2_ASAP7_75t_L g402 ( .A(n_294), .Y(n_402) );
INVx3_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
INVx2_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
OAI32xp33_ASAP7_75t_L g453 ( .A1(n_297), .A2(n_344), .A3(n_375), .B1(n_454), .B2(n_455), .Y(n_453) );
OR2x2_ASAP7_75t_L g424 ( .A(n_298), .B(n_411), .Y(n_424) );
INVx1_ASAP7_75t_L g434 ( .A(n_299), .Y(n_434) );
OR2x2_ASAP7_75t_L g299 ( .A(n_300), .B(n_302), .Y(n_299) );
INVx2_ASAP7_75t_L g349 ( .A(n_300), .Y(n_349) );
AND2x2_ASAP7_75t_L g420 ( .A(n_300), .B(n_395), .Y(n_420) );
OR2x2_ASAP7_75t_L g451 ( .A(n_300), .B(n_452), .Y(n_451) );
INVx2_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_301), .B(n_356), .Y(n_355) );
INVx1_ASAP7_75t_SL g302 ( .A(n_303), .Y(n_302) );
INVx1_ASAP7_75t_L g345 ( .A(n_304), .Y(n_345) );
OR2x2_ASAP7_75t_L g305 ( .A(n_306), .B(n_307), .Y(n_305) );
INVx2_ASAP7_75t_SL g310 ( .A(n_307), .Y(n_310) );
OR2x2_ASAP7_75t_L g397 ( .A(n_307), .B(n_398), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_308), .B(n_326), .Y(n_325) );
NOR2xp67_ASAP7_75t_L g431 ( .A(n_308), .B(n_432), .Y(n_431) );
BUFx2_ASAP7_75t_L g444 ( .A(n_308), .Y(n_444) );
A2O1A1Ixp33_ASAP7_75t_L g309 ( .A1(n_310), .A2(n_311), .B(n_316), .C(n_319), .Y(n_309) );
AND2x2_ASAP7_75t_L g459 ( .A(n_311), .B(n_460), .Y(n_459) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
OR2x2_ASAP7_75t_L g312 ( .A(n_313), .B(n_315), .Y(n_312) );
BUFx2_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
OR2x2_ASAP7_75t_L g385 ( .A(n_315), .B(n_386), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_315), .B(n_319), .Y(n_406) );
AND2x2_ASAP7_75t_L g437 ( .A(n_315), .B(n_438), .Y(n_437) );
O2A1O1Ixp33_ASAP7_75t_L g447 ( .A1(n_317), .A2(n_448), .B(n_450), .C(n_453), .Y(n_447) );
AOI222xp33_ASAP7_75t_L g321 ( .A1(n_318), .A2(n_322), .B1(n_324), .B2(n_327), .C1(n_335), .C2(n_337), .Y(n_321) );
AND2x2_ASAP7_75t_L g389 ( .A(n_318), .B(n_390), .Y(n_389) );
AND2x2_ASAP7_75t_L g322 ( .A(n_319), .B(n_323), .Y(n_322) );
INVx2_ASAP7_75t_SL g343 ( .A(n_319), .Y(n_343) );
NAND4xp25_ASAP7_75t_L g320 ( .A(n_321), .B(n_340), .C(n_361), .D(n_371), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_323), .B(n_329), .Y(n_383) );
INVx1_ASAP7_75t_SL g324 ( .A(n_325), .Y(n_324) );
AND2x2_ASAP7_75t_L g391 ( .A(n_326), .B(n_392), .Y(n_391) );
INVx2_ASAP7_75t_SL g398 ( .A(n_326), .Y(n_398) );
AND2x2_ASAP7_75t_L g327 ( .A(n_328), .B(n_330), .Y(n_327) );
A2O1A1Ixp33_ASAP7_75t_L g361 ( .A1(n_328), .A2(n_362), .B(n_366), .C(n_370), .Y(n_361) );
INVx2_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_329), .B(n_344), .Y(n_465) );
OR2x2_ASAP7_75t_L g469 ( .A(n_329), .B(n_355), .Y(n_469) );
INVx1_ASAP7_75t_L g442 ( .A(n_330), .Y(n_442) );
INVx2_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
AND2x2_ASAP7_75t_L g332 ( .A(n_333), .B(n_334), .Y(n_332) );
INVx1_ASAP7_75t_SL g376 ( .A(n_333), .Y(n_376) );
INVx1_ASAP7_75t_L g356 ( .A(n_334), .Y(n_356) );
INVx2_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_336), .B(n_373), .Y(n_372) );
BUFx2_ASAP7_75t_SL g337 ( .A(n_338), .Y(n_337) );
INVx1_ASAP7_75t_L g360 ( .A(n_338), .Y(n_360) );
AOI322xp5_ASAP7_75t_L g340 ( .A1(n_341), .A2(n_343), .A3(n_344), .B1(n_346), .B2(n_350), .C1(n_351), .C2(n_357), .Y(n_340) );
INVxp67_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
O2A1O1Ixp33_ASAP7_75t_SL g422 ( .A1(n_343), .A2(n_423), .B(n_424), .C(n_425), .Y(n_422) );
INVx1_ASAP7_75t_L g445 ( .A(n_344), .Y(n_445) );
NOR2xp67_ASAP7_75t_L g346 ( .A(n_347), .B(n_349), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
AND2x2_ASAP7_75t_L g403 ( .A(n_349), .B(n_404), .Y(n_403) );
AND2x2_ASAP7_75t_L g351 ( .A(n_352), .B(n_354), .Y(n_351) );
INVx2_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx2_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
HB1xp67_ASAP7_75t_L g425 ( .A(n_355), .Y(n_425) );
INVx2_ASAP7_75t_SL g357 ( .A(n_358), .Y(n_357) );
OR2x2_ASAP7_75t_L g358 ( .A(n_359), .B(n_360), .Y(n_358) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
OR2x2_ASAP7_75t_L g363 ( .A(n_364), .B(n_365), .Y(n_363) );
INVx3_ASAP7_75t_L g368 ( .A(n_365), .Y(n_368) );
OR2x2_ASAP7_75t_L g436 ( .A(n_365), .B(n_398), .Y(n_436) );
NOR2xp33_ASAP7_75t_L g481 ( .A(n_365), .B(n_482), .Y(n_481) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_368), .B(n_369), .Y(n_367) );
INVx1_ASAP7_75t_SL g468 ( .A(n_369), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_370), .B(n_374), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
NAND3xp33_ASAP7_75t_SL g473 ( .A(n_378), .B(n_474), .C(n_476), .Y(n_473) );
NOR3xp33_ASAP7_75t_SL g379 ( .A(n_380), .B(n_417), .C(n_446), .Y(n_379) );
NAND2xp5_ASAP7_75t_SL g380 ( .A(n_381), .B(n_399), .Y(n_380) );
O2A1O1Ixp33_ASAP7_75t_L g381 ( .A1(n_382), .A2(n_384), .B(n_387), .C(n_393), .Y(n_381) );
OAI31xp33_ASAP7_75t_L g426 ( .A1(n_382), .A2(n_404), .A3(n_427), .B(n_428), .Y(n_426) );
INVx1_ASAP7_75t_SL g382 ( .A(n_383), .Y(n_382) );
INVx1_ASAP7_75t_SL g384 ( .A(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
NOR2xp33_ASAP7_75t_L g388 ( .A(n_389), .B(n_391), .Y(n_388) );
INVx2_ASAP7_75t_L g441 ( .A(n_389), .Y(n_441) );
INVx1_ASAP7_75t_L g416 ( .A(n_391), .Y(n_416) );
AOI21xp5_ASAP7_75t_L g393 ( .A1(n_394), .A2(n_396), .B(n_397), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
OR2x2_ASAP7_75t_L g443 ( .A(n_401), .B(n_444), .Y(n_443) );
INVxp67_ASAP7_75t_L g482 ( .A(n_402), .Y(n_482) );
OAI22xp33_ASAP7_75t_SL g405 ( .A1(n_406), .A2(n_407), .B1(n_412), .B2(n_416), .Y(n_405) );
INVx3_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
AND2x4_ASAP7_75t_L g408 ( .A(n_409), .B(n_410), .Y(n_408) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
HB1xp67_ASAP7_75t_L g423 ( .A(n_411), .Y(n_423) );
OR2x2_ASAP7_75t_L g474 ( .A(n_411), .B(n_475), .Y(n_474) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
NAND3xp33_ASAP7_75t_SL g417 ( .A(n_418), .B(n_426), .C(n_433), .Y(n_417) );
O2A1O1Ixp33_ASAP7_75t_L g418 ( .A1(n_419), .A2(n_420), .B(n_421), .C(n_422), .Y(n_418) );
INVx2_ASAP7_75t_L g455 ( .A(n_419), .Y(n_455) );
INVx1_ASAP7_75t_SL g428 ( .A(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
AOI221xp5_ASAP7_75t_L g433 ( .A1(n_434), .A2(n_435), .B1(n_437), .B2(n_439), .C(n_440), .Y(n_433) );
INVx2_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
OAI22xp33_ASAP7_75t_L g440 ( .A1(n_441), .A2(n_442), .B1(n_443), .B2(n_445), .Y(n_440) );
NAND3xp33_ASAP7_75t_SL g446 ( .A(n_447), .B(n_456), .C(n_466), .Y(n_446) );
INVxp33_ASAP7_75t_SL g448 ( .A(n_449), .Y(n_448) );
INVx1_ASAP7_75t_SL g450 ( .A(n_451), .Y(n_450) );
AOI22xp5_ASAP7_75t_L g456 ( .A1(n_457), .A2(n_459), .B1(n_462), .B2(n_464), .Y(n_456) );
INVx2_ASAP7_75t_L g470 ( .A(n_457), .Y(n_470) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx1_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
OAI22xp5_ASAP7_75t_L g467 ( .A1(n_468), .A2(n_469), .B1(n_470), .B2(n_471), .Y(n_467) );
INVx1_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
OAI22xp33_ASAP7_75t_SL g477 ( .A1(n_476), .A2(n_478), .B1(n_479), .B2(n_480), .Y(n_477) );
INVx1_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
AOI22xp33_ASAP7_75t_L g485 ( .A1(n_486), .A2(n_501), .B1(n_511), .B2(n_512), .Y(n_485) );
CKINVDCx20_ASAP7_75t_R g518 ( .A(n_486), .Y(n_518) );
AOI22xp5_ASAP7_75t_L g486 ( .A1(n_487), .A2(n_492), .B1(n_499), .B2(n_500), .Y(n_486) );
CKINVDCx20_ASAP7_75t_R g499 ( .A(n_487), .Y(n_499) );
AOI22xp5_ASAP7_75t_L g487 ( .A1(n_488), .A2(n_489), .B1(n_490), .B2(n_491), .Y(n_487) );
INVx1_ASAP7_75t_L g490 ( .A(n_488), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_489), .Y(n_491) );
INVx1_ASAP7_75t_L g500 ( .A(n_492), .Y(n_500) );
INVx1_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
INVx1_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
CKINVDCx20_ASAP7_75t_R g501 ( .A(n_502), .Y(n_501) );
CKINVDCx20_ASAP7_75t_R g502 ( .A(n_503), .Y(n_502) );
INVxp67_ASAP7_75t_L g516 ( .A(n_504), .Y(n_516) );
CKINVDCx8_ASAP7_75t_R g505 ( .A(n_506), .Y(n_505) );
NOR2xp33_ASAP7_75t_L g507 ( .A(n_508), .B(n_509), .Y(n_507) );
CKINVDCx16_ASAP7_75t_R g514 ( .A(n_510), .Y(n_514) );
AO21x1_ASAP7_75t_SL g522 ( .A1(n_510), .A2(n_523), .B(n_524), .Y(n_522) );
CKINVDCx20_ASAP7_75t_R g512 ( .A(n_513), .Y(n_512) );
CKINVDCx20_ASAP7_75t_R g519 ( .A(n_513), .Y(n_519) );
OR2x2_ASAP7_75t_L g513 ( .A(n_514), .B(n_515), .Y(n_513) );
CKINVDCx20_ASAP7_75t_R g520 ( .A(n_521), .Y(n_520) );
CKINVDCx20_ASAP7_75t_R g521 ( .A(n_522), .Y(n_521) );
endmodule