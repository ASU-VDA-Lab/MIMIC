module fake_jpeg_15893_n_244 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_244);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_244;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx11_ASAP7_75t_SL g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx16f_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx6f_ASAP7_75t_SL g21 ( 
.A(n_8),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx4f_ASAP7_75t_SL g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_10),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_12),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_5),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_16),
.B(n_0),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_36),
.B(n_45),
.Y(n_51)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_16),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_42),
.B(n_46),
.Y(n_55)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_25),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_25),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_47),
.B(n_35),
.Y(n_67)
);

HB1xp67_ASAP7_75t_L g48 ( 
.A(n_20),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_48),
.B(n_18),
.Y(n_66)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_49),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_17),
.B(n_0),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_50),
.B(n_35),
.Y(n_59)
);

NAND2x1_ASAP7_75t_SL g53 ( 
.A(n_40),
.B(n_20),
.Y(n_53)
);

NAND2xp67_ASAP7_75t_L g80 ( 
.A(n_53),
.B(n_40),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_39),
.A2(n_34),
.B1(n_28),
.B2(n_19),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_56),
.A2(n_64),
.B1(n_30),
.B2(n_44),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_59),
.B(n_67),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_37),
.B(n_29),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_60),
.B(n_69),
.Y(n_88)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_63),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_39),
.A2(n_28),
.B1(n_34),
.B2(n_33),
.Y(n_64)
);

AOI21xp33_ASAP7_75t_SL g65 ( 
.A1(n_48),
.A2(n_20),
.B(n_19),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_65),
.B(n_23),
.C(n_31),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_66),
.B(n_18),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_37),
.B(n_29),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_55),
.A2(n_38),
.B1(n_44),
.B2(n_34),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_71),
.A2(n_79),
.B1(n_83),
.B2(n_86),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_72),
.B(n_74),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_59),
.B(n_36),
.Y(n_74)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_62),
.Y(n_75)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_75),
.Y(n_115)
);

AOI32xp33_ASAP7_75t_L g76 ( 
.A1(n_51),
.A2(n_44),
.A3(n_49),
.B1(n_20),
.B2(n_50),
.Y(n_76)
);

AOI32xp33_ASAP7_75t_L g111 ( 
.A1(n_76),
.A2(n_100),
.A3(n_52),
.B1(n_23),
.B2(n_70),
.Y(n_111)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_62),
.Y(n_77)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_77),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_60),
.B(n_42),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_78),
.B(n_81),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_65),
.A2(n_38),
.B1(n_24),
.B2(n_33),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_80),
.B(n_105),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_69),
.B(n_42),
.Y(n_81)
);

HB1xp67_ASAP7_75t_L g82 ( 
.A(n_54),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_82),
.B(n_87),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_64),
.A2(n_22),
.B1(n_17),
.B2(n_27),
.Y(n_83)
);

CKINVDCx6p67_ASAP7_75t_R g84 ( 
.A(n_68),
.Y(n_84)
);

INVx1_ASAP7_75t_SL g124 ( 
.A(n_84),
.Y(n_124)
);

BUFx8_ASAP7_75t_L g85 ( 
.A(n_53),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_85),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_55),
.A2(n_22),
.B1(n_27),
.B2(n_24),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_54),
.Y(n_87)
);

INVx13_ASAP7_75t_L g89 ( 
.A(n_53),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_89),
.B(n_93),
.Y(n_118)
);

O2A1O1Ixp33_ASAP7_75t_SL g90 ( 
.A1(n_55),
.A2(n_47),
.B(n_46),
.C(n_43),
.Y(n_90)
);

O2A1O1Ixp33_ASAP7_75t_L g113 ( 
.A1(n_90),
.A2(n_103),
.B(n_104),
.C(n_23),
.Y(n_113)
);

BUFx24_ASAP7_75t_L g91 ( 
.A(n_61),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_91),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_61),
.A2(n_43),
.B1(n_49),
.B2(n_30),
.Y(n_92)
);

OR2x2_ASAP7_75t_L g122 ( 
.A(n_92),
.B(n_101),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_68),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_94),
.B(n_95),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_67),
.B(n_47),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_70),
.A2(n_45),
.B1(n_41),
.B2(n_46),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_96),
.A2(n_31),
.B1(n_2),
.B2(n_3),
.Y(n_128)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_57),
.Y(n_97)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_97),
.Y(n_114)
);

BUFx2_ASAP7_75t_L g98 ( 
.A(n_58),
.Y(n_98)
);

INVx5_ASAP7_75t_L g117 ( 
.A(n_98),
.Y(n_117)
);

NAND2xp33_ASAP7_75t_SL g100 ( 
.A(n_63),
.B(n_45),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_68),
.Y(n_101)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_52),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_102),
.B(n_52),
.Y(n_116)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_58),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_67),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_57),
.B(n_1),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_SL g112 ( 
.A(n_106),
.B(n_23),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_111),
.B(n_80),
.Y(n_132)
);

CKINVDCx14_ASAP7_75t_R g139 ( 
.A(n_112),
.Y(n_139)
);

CKINVDCx14_ASAP7_75t_R g144 ( 
.A(n_113),
.Y(n_144)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_116),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_88),
.B(n_41),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_120),
.B(n_127),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_106),
.B(n_18),
.C(n_26),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_125),
.B(n_85),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_88),
.B(n_73),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_128),
.A2(n_129),
.B1(n_71),
.B2(n_102),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_88),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_115),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_131),
.A2(n_132),
.B(n_140),
.Y(n_155)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_116),
.Y(n_134)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_134),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_114),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_135),
.B(n_142),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_136),
.B(n_1),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_118),
.A2(n_120),
.B1(n_127),
.B2(n_123),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_138),
.A2(n_141),
.B1(n_143),
.B2(n_146),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_123),
.A2(n_89),
.B1(n_93),
.B2(n_100),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_109),
.B(n_108),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_111),
.A2(n_130),
.B1(n_128),
.B2(n_125),
.Y(n_143)
);

AOI322xp5_ASAP7_75t_L g145 ( 
.A1(n_126),
.A2(n_85),
.A3(n_90),
.B1(n_105),
.B2(n_98),
.C1(n_26),
.C2(n_96),
.Y(n_145)
);

A2O1A1O1Ixp25_ASAP7_75t_L g151 ( 
.A1(n_145),
.A2(n_126),
.B(n_122),
.C(n_130),
.D(n_129),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_113),
.A2(n_99),
.B1(n_103),
.B2(n_97),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_115),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_147),
.A2(n_124),
.B(n_107),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_108),
.B(n_105),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_148),
.A2(n_122),
.B(n_119),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_110),
.B(n_77),
.Y(n_149)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_149),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_138),
.B(n_112),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_150),
.B(n_154),
.C(n_156),
.Y(n_170)
);

AOI221xp5_ASAP7_75t_L g173 ( 
.A1(n_151),
.A2(n_158),
.B1(n_143),
.B2(n_141),
.C(n_144),
.Y(n_173)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_149),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_153),
.B(n_162),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_138),
.B(n_126),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_139),
.B(n_140),
.C(n_137),
.Y(n_156)
);

AO21x1_ASAP7_75t_L g172 ( 
.A1(n_157),
.A2(n_159),
.B(n_160),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_132),
.A2(n_122),
.B(n_119),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_139),
.A2(n_124),
.B(n_121),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_133),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_163),
.A2(n_164),
.B(n_145),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_144),
.A2(n_121),
.B(n_117),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_133),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_165),
.B(n_167),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_134),
.Y(n_167)
);

INVx5_ASAP7_75t_L g171 ( 
.A(n_157),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_171),
.B(n_177),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_SL g197 ( 
.A(n_173),
.B(n_26),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_150),
.B(n_137),
.C(n_148),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_174),
.B(n_178),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_161),
.A2(n_142),
.B1(n_146),
.B2(n_136),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_175),
.A2(n_176),
.B1(n_185),
.B2(n_184),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_160),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_176),
.B(n_179),
.Y(n_188)
);

INVx13_ASAP7_75t_L g177 ( 
.A(n_152),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_156),
.B(n_147),
.C(n_131),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_166),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_181),
.A2(n_172),
.B1(n_178),
.B2(n_174),
.Y(n_199)
);

OR2x2_ASAP7_75t_L g182 ( 
.A(n_161),
.B(n_75),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_182),
.B(n_185),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_154),
.B(n_114),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_183),
.B(n_151),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_168),
.A2(n_99),
.B1(n_117),
.B2(n_84),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_184),
.A2(n_158),
.B1(n_163),
.B2(n_168),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_164),
.Y(n_185)
);

CKINVDCx16_ASAP7_75t_R g186 ( 
.A(n_169),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_186),
.B(n_189),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_180),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_187),
.B(n_182),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_189),
.A2(n_190),
.B1(n_198),
.B2(n_172),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_171),
.A2(n_163),
.B1(n_159),
.B2(n_155),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_170),
.B(n_155),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_193),
.B(n_196),
.Y(n_201)
);

INVx13_ASAP7_75t_L g195 ( 
.A(n_177),
.Y(n_195)
);

BUFx2_ASAP7_75t_L g204 ( 
.A(n_195),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_197),
.B(n_199),
.Y(n_205)
);

O2A1O1Ixp33_ASAP7_75t_L g200 ( 
.A1(n_191),
.A2(n_172),
.B(n_179),
.C(n_175),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_200),
.A2(n_208),
.B1(n_209),
.B2(n_211),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_SL g213 ( 
.A(n_202),
.B(n_198),
.Y(n_213)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_188),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_203),
.A2(n_210),
.B(n_84),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_193),
.B(n_194),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_206),
.B(n_207),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_194),
.B(n_170),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_190),
.B(n_183),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_192),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_213),
.B(n_218),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_200),
.A2(n_181),
.B1(n_197),
.B2(n_196),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_214),
.B(n_220),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_206),
.B(n_195),
.C(n_91),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_215),
.B(n_216),
.C(n_217),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_205),
.B(n_91),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_207),
.B(n_101),
.C(n_84),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_205),
.B(n_201),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_201),
.A2(n_15),
.B1(n_4),
.B2(n_5),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_221),
.A2(n_204),
.B(n_4),
.Y(n_225)
);

OA21x2_ASAP7_75t_SL g222 ( 
.A1(n_219),
.A2(n_204),
.B(n_15),
.Y(n_222)
);

OR2x2_ASAP7_75t_L g233 ( 
.A(n_222),
.B(n_223),
.Y(n_233)
);

HB1xp67_ASAP7_75t_L g223 ( 
.A(n_217),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_225),
.B(n_10),
.Y(n_232)
);

OA21x2_ASAP7_75t_SL g227 ( 
.A1(n_215),
.A2(n_2),
.B(n_6),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_227),
.A2(n_7),
.B(n_9),
.Y(n_229)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_229),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_224),
.A2(n_216),
.B(n_218),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_230),
.B(n_231),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_224),
.A2(n_226),
.B(n_228),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_232),
.B(n_10),
.Y(n_235)
);

AOI322xp5_ASAP7_75t_L g238 ( 
.A1(n_235),
.A2(n_237),
.A3(n_228),
.B1(n_213),
.B2(n_14),
.C1(n_13),
.C2(n_11),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_233),
.B(n_226),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_238),
.B(n_13),
.Y(n_241)
);

O2A1O1Ixp33_ASAP7_75t_SL g239 ( 
.A1(n_236),
.A2(n_234),
.B(n_212),
.C(n_14),
.Y(n_239)
);

NOR2xp67_ASAP7_75t_L g240 ( 
.A(n_239),
.B(n_11),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_240),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_242),
.A2(n_241),
.B(n_212),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_243),
.B(n_14),
.Y(n_244)
);


endmodule