module real_aes_7921_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_666;
wire n_537;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_369;
wire n_343;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_725;
wire n_504;
wire n_310;
wire n_455;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_502;
wire n_434;
wire n_527;
wire n_600;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_249;
wire n_623;
wire n_721;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_717;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_418;
wire n_140;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_639;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g108 ( .A(n_0), .Y(n_108) );
INVx1_ASAP7_75t_L g455 ( .A(n_1), .Y(n_455) );
INVx1_ASAP7_75t_L g259 ( .A(n_2), .Y(n_259) );
AOI22xp33_ASAP7_75t_L g530 ( .A1(n_3), .A2(n_36), .B1(n_209), .B2(n_494), .Y(n_530) );
AOI21xp33_ASAP7_75t_L g220 ( .A1(n_4), .A2(n_142), .B(n_221), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_5), .B(n_164), .Y(n_480) );
AND2x6_ASAP7_75t_L g147 ( .A(n_6), .B(n_148), .Y(n_147) );
AOI21xp5_ASAP7_75t_L g140 ( .A1(n_7), .A2(n_141), .B(n_149), .Y(n_140) );
INVx1_ASAP7_75t_L g105 ( .A(n_8), .Y(n_105) );
NOR2xp33_ASAP7_75t_L g123 ( .A(n_8), .B(n_37), .Y(n_123) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_9), .B(n_207), .Y(n_206) );
INVx1_ASAP7_75t_L g226 ( .A(n_10), .Y(n_226) );
INVx1_ASAP7_75t_L g139 ( .A(n_11), .Y(n_139) );
INVx1_ASAP7_75t_L g449 ( .A(n_12), .Y(n_449) );
INVx1_ASAP7_75t_L g159 ( .A(n_13), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_14), .B(n_233), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_15), .B(n_165), .Y(n_482) );
AO32x2_ASAP7_75t_L g528 ( .A1(n_16), .A2(n_164), .A3(n_180), .B1(n_468), .B2(n_529), .Y(n_528) );
NAND2xp5_ASAP7_75t_SL g514 ( .A(n_17), .B(n_209), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_18), .B(n_176), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_19), .B(n_165), .Y(n_458) );
AOI22xp33_ASAP7_75t_L g531 ( .A1(n_20), .A2(n_48), .B1(n_209), .B2(n_494), .Y(n_531) );
NAND2xp5_ASAP7_75t_SL g169 ( .A(n_21), .B(n_142), .Y(n_169) );
AOI22xp33_ASAP7_75t_SL g495 ( .A1(n_22), .A2(n_74), .B1(n_209), .B2(n_233), .Y(n_495) );
NAND2xp5_ASAP7_75t_SL g504 ( .A(n_23), .B(n_209), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_24), .B(n_219), .Y(n_249) );
A2O1A1Ixp33_ASAP7_75t_L g155 ( .A1(n_25), .A2(n_156), .B(n_158), .C(n_160), .Y(n_155) );
BUFx6f_ASAP7_75t_L g146 ( .A(n_26), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_27), .B(n_135), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_28), .B(n_191), .Y(n_260) );
AOI222xp33_ASAP7_75t_SL g125 ( .A1(n_29), .A2(n_88), .B1(n_126), .B2(n_714), .C1(n_715), .C2(n_718), .Y(n_125) );
INVx1_ASAP7_75t_L g714 ( .A(n_29), .Y(n_714) );
INVx1_ASAP7_75t_L g238 ( .A(n_30), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_31), .B(n_135), .Y(n_506) );
INVx2_ASAP7_75t_L g145 ( .A(n_32), .Y(n_145) );
NAND2xp5_ASAP7_75t_SL g463 ( .A(n_33), .B(n_209), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_34), .B(n_135), .Y(n_516) );
A2O1A1Ixp33_ASAP7_75t_L g170 ( .A1(n_35), .A2(n_147), .B(n_152), .C(n_171), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g104 ( .A(n_37), .B(n_105), .Y(n_104) );
INVx1_ASAP7_75t_L g236 ( .A(n_38), .Y(n_236) );
NAND2xp5_ASAP7_75t_SL g190 ( .A(n_39), .B(n_191), .Y(n_190) );
CKINVDCx20_ASAP7_75t_R g124 ( .A(n_40), .Y(n_124) );
NAND2xp5_ASAP7_75t_SL g475 ( .A(n_41), .B(n_209), .Y(n_475) );
AOI22xp33_ASAP7_75t_L g493 ( .A1(n_42), .A2(n_84), .B1(n_161), .B2(n_494), .Y(n_493) );
NAND2xp5_ASAP7_75t_SL g478 ( .A(n_43), .B(n_209), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_44), .B(n_209), .Y(n_450) );
CKINVDCx16_ASAP7_75t_R g239 ( .A(n_45), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_46), .B(n_454), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_47), .B(n_142), .Y(n_210) );
AOI22xp33_ASAP7_75t_SL g486 ( .A1(n_49), .A2(n_59), .B1(n_209), .B2(n_233), .Y(n_486) );
AOI22xp33_ASAP7_75t_L g99 ( .A1(n_50), .A2(n_100), .B1(n_113), .B2(n_729), .Y(n_99) );
AOI22xp5_ASAP7_75t_L g232 ( .A1(n_51), .A2(n_152), .B1(n_233), .B2(n_235), .Y(n_232) );
CKINVDCx20_ASAP7_75t_R g182 ( .A(n_52), .Y(n_182) );
NAND2xp5_ASAP7_75t_SL g467 ( .A(n_53), .B(n_209), .Y(n_467) );
CKINVDCx16_ASAP7_75t_R g256 ( .A(n_54), .Y(n_256) );
NAND2xp5_ASAP7_75t_SL g510 ( .A(n_55), .B(n_209), .Y(n_510) );
A2O1A1Ixp33_ASAP7_75t_L g223 ( .A1(n_56), .A2(n_224), .B(n_225), .C(n_227), .Y(n_223) );
CKINVDCx20_ASAP7_75t_R g195 ( .A(n_57), .Y(n_195) );
INVx1_ASAP7_75t_L g222 ( .A(n_58), .Y(n_222) );
INVx1_ASAP7_75t_L g148 ( .A(n_60), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_61), .B(n_209), .Y(n_456) );
INVx1_ASAP7_75t_L g138 ( .A(n_62), .Y(n_138) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_63), .Y(n_117) );
AO32x2_ASAP7_75t_L g491 ( .A1(n_64), .A2(n_164), .A3(n_201), .B1(n_468), .B2(n_492), .Y(n_491) );
INVx1_ASAP7_75t_L g466 ( .A(n_65), .Y(n_466) );
INVx1_ASAP7_75t_L g501 ( .A(n_66), .Y(n_501) );
A2O1A1Ixp33_ASAP7_75t_SL g246 ( .A1(n_67), .A2(n_176), .B(n_227), .C(n_247), .Y(n_246) );
INVxp67_ASAP7_75t_L g248 ( .A(n_68), .Y(n_248) );
NAND2xp5_ASAP7_75t_SL g502 ( .A(n_69), .B(n_233), .Y(n_502) );
INVx1_ASAP7_75t_L g112 ( .A(n_70), .Y(n_112) );
CKINVDCx20_ASAP7_75t_R g241 ( .A(n_71), .Y(n_241) );
INVx1_ASAP7_75t_L g186 ( .A(n_72), .Y(n_186) );
OAI22xp5_ASAP7_75t_L g725 ( .A1(n_73), .A2(n_128), .B1(n_716), .B2(n_726), .Y(n_725) );
CKINVDCx20_ASAP7_75t_R g726 ( .A(n_73), .Y(n_726) );
A2O1A1Ixp33_ASAP7_75t_L g188 ( .A1(n_75), .A2(n_147), .B(n_152), .C(n_189), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_76), .B(n_494), .Y(n_515) );
NAND2xp5_ASAP7_75t_SL g505 ( .A(n_77), .B(n_233), .Y(n_505) );
NAND2xp5_ASAP7_75t_SL g172 ( .A(n_78), .B(n_173), .Y(n_172) );
INVx2_ASAP7_75t_L g136 ( .A(n_79), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_80), .B(n_176), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_81), .B(n_233), .Y(n_476) );
A2O1A1Ixp33_ASAP7_75t_L g257 ( .A1(n_82), .A2(n_147), .B(n_152), .C(n_258), .Y(n_257) );
INVx2_ASAP7_75t_L g109 ( .A(n_83), .Y(n_109) );
OR2x2_ASAP7_75t_L g120 ( .A(n_83), .B(n_121), .Y(n_120) );
OR2x2_ASAP7_75t_L g127 ( .A(n_83), .B(n_122), .Y(n_127) );
AOI22xp33_ASAP7_75t_L g485 ( .A1(n_85), .A2(n_98), .B1(n_233), .B2(n_234), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_86), .B(n_135), .Y(n_228) );
CKINVDCx20_ASAP7_75t_R g263 ( .A(n_87), .Y(n_263) );
A2O1A1Ixp33_ASAP7_75t_L g203 ( .A1(n_89), .A2(n_147), .B(n_152), .C(n_204), .Y(n_203) );
CKINVDCx20_ASAP7_75t_R g212 ( .A(n_90), .Y(n_212) );
INVx1_ASAP7_75t_L g245 ( .A(n_91), .Y(n_245) );
CKINVDCx16_ASAP7_75t_R g150 ( .A(n_92), .Y(n_150) );
NAND2xp5_ASAP7_75t_SL g205 ( .A(n_93), .B(n_173), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_94), .B(n_233), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_95), .B(n_164), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_96), .B(n_112), .Y(n_111) );
AOI21xp5_ASAP7_75t_L g243 ( .A1(n_97), .A2(n_142), .B(n_244), .Y(n_243) );
CKINVDCx20_ASAP7_75t_R g100 ( .A(n_101), .Y(n_100) );
CKINVDCx16_ASAP7_75t_R g101 ( .A(n_102), .Y(n_101) );
INVx2_ASAP7_75t_L g729 ( .A(n_102), .Y(n_729) );
AND2x2_ASAP7_75t_L g102 ( .A(n_103), .B(n_106), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
CKINVDCx14_ASAP7_75t_R g106 ( .A(n_107), .Y(n_106) );
NAND3xp33_ASAP7_75t_SL g107 ( .A(n_108), .B(n_109), .C(n_110), .Y(n_107) );
AND2x2_ASAP7_75t_L g122 ( .A(n_108), .B(n_123), .Y(n_122) );
OR2x2_ASAP7_75t_L g438 ( .A(n_109), .B(n_122), .Y(n_438) );
NOR2x2_ASAP7_75t_L g720 ( .A(n_109), .B(n_121), .Y(n_720) );
INVx1_ASAP7_75t_SL g110 ( .A(n_111), .Y(n_110) );
AOI22x1_ASAP7_75t_L g113 ( .A1(n_114), .A2(n_125), .B1(n_721), .B2(n_724), .Y(n_113) );
NOR2xp33_ASAP7_75t_L g114 ( .A(n_115), .B(n_118), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
INVx2_ASAP7_75t_L g723 ( .A(n_117), .Y(n_723) );
AOI21xp5_ASAP7_75t_L g724 ( .A1(n_118), .A2(n_725), .B(n_727), .Y(n_724) );
NOR2xp33_ASAP7_75t_SL g118 ( .A(n_119), .B(n_124), .Y(n_118) );
HB1xp67_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx1_ASAP7_75t_SL g728 ( .A(n_120), .Y(n_728) );
INVx2_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
OAI22xp5_ASAP7_75t_L g126 ( .A1(n_127), .A2(n_128), .B1(n_436), .B2(n_439), .Y(n_126) );
OAI22xp5_ASAP7_75t_SL g715 ( .A1(n_127), .A2(n_438), .B1(n_716), .B2(n_717), .Y(n_715) );
INVx2_ASAP7_75t_SL g716 ( .A(n_128), .Y(n_716) );
OR4x2_ASAP7_75t_L g128 ( .A(n_129), .B(n_332), .C(n_391), .D(n_418), .Y(n_128) );
NAND3xp33_ASAP7_75t_SL g129 ( .A(n_130), .B(n_274), .C(n_299), .Y(n_129) );
O2A1O1Ixp33_ASAP7_75t_L g130 ( .A1(n_131), .A2(n_197), .B(n_217), .C(n_250), .Y(n_130) );
AOI211xp5_ASAP7_75t_SL g422 ( .A1(n_131), .A2(n_423), .B(n_425), .C(n_428), .Y(n_422) );
AND2x2_ASAP7_75t_L g131 ( .A(n_132), .B(n_166), .Y(n_131) );
INVx1_ASAP7_75t_L g297 ( .A(n_132), .Y(n_297) );
INVx1_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
OR2x2_ASAP7_75t_L g272 ( .A(n_133), .B(n_273), .Y(n_272) );
INVx2_ASAP7_75t_L g304 ( .A(n_133), .Y(n_304) );
AND2x2_ASAP7_75t_L g359 ( .A(n_133), .B(n_328), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_133), .B(n_215), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_133), .B(n_216), .Y(n_417) );
INVx2_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
INVx1_ASAP7_75t_L g278 ( .A(n_134), .Y(n_278) );
AND2x2_ASAP7_75t_L g321 ( .A(n_134), .B(n_184), .Y(n_321) );
AND2x2_ASAP7_75t_L g339 ( .A(n_134), .B(n_216), .Y(n_339) );
OA21x2_ASAP7_75t_L g134 ( .A1(n_135), .A2(n_140), .B(n_163), .Y(n_134) );
INVx1_ASAP7_75t_L g196 ( .A(n_135), .Y(n_196) );
INVx2_ASAP7_75t_L g201 ( .A(n_135), .Y(n_201) );
OA21x2_ASAP7_75t_L g498 ( .A1(n_135), .A2(n_499), .B(n_506), .Y(n_498) );
OA21x2_ASAP7_75t_L g507 ( .A1(n_135), .A2(n_508), .B(n_516), .Y(n_507) );
AND2x2_ASAP7_75t_SL g135 ( .A(n_136), .B(n_137), .Y(n_135) );
AND2x2_ASAP7_75t_L g165 ( .A(n_136), .B(n_137), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_138), .B(n_139), .Y(n_137) );
BUFx2_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
AND2x4_ASAP7_75t_L g142 ( .A(n_143), .B(n_147), .Y(n_142) );
NAND2x1p5_ASAP7_75t_L g187 ( .A(n_143), .B(n_147), .Y(n_187) );
AND2x2_ASAP7_75t_L g143 ( .A(n_144), .B(n_146), .Y(n_143) );
INVx1_ASAP7_75t_L g454 ( .A(n_144), .Y(n_454) );
INVx1_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx2_ASAP7_75t_L g153 ( .A(n_145), .Y(n_153) );
INVx1_ASAP7_75t_L g234 ( .A(n_145), .Y(n_234) );
INVx1_ASAP7_75t_L g154 ( .A(n_146), .Y(n_154) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_146), .Y(n_157) );
INVx3_ASAP7_75t_L g174 ( .A(n_146), .Y(n_174) );
INVx1_ASAP7_75t_L g176 ( .A(n_146), .Y(n_176) );
BUFx6f_ASAP7_75t_L g191 ( .A(n_146), .Y(n_191) );
INVx4_ASAP7_75t_SL g162 ( .A(n_147), .Y(n_162) );
OAI21xp5_ASAP7_75t_L g447 ( .A1(n_147), .A2(n_448), .B(n_452), .Y(n_447) );
BUFx3_ASAP7_75t_L g468 ( .A(n_147), .Y(n_468) );
OAI21xp5_ASAP7_75t_L g473 ( .A1(n_147), .A2(n_474), .B(n_477), .Y(n_473) );
OAI21xp5_ASAP7_75t_L g499 ( .A1(n_147), .A2(n_500), .B(n_503), .Y(n_499) );
OAI21xp5_ASAP7_75t_L g508 ( .A1(n_147), .A2(n_509), .B(n_513), .Y(n_508) );
O2A1O1Ixp33_ASAP7_75t_L g149 ( .A1(n_150), .A2(n_151), .B(n_155), .C(n_162), .Y(n_149) );
O2A1O1Ixp33_ASAP7_75t_L g221 ( .A1(n_151), .A2(n_162), .B(n_222), .C(n_223), .Y(n_221) );
O2A1O1Ixp33_ASAP7_75t_L g244 ( .A1(n_151), .A2(n_162), .B(n_245), .C(n_246), .Y(n_244) );
INVx5_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
AND2x6_ASAP7_75t_L g152 ( .A(n_153), .B(n_154), .Y(n_152) );
BUFx3_ASAP7_75t_L g161 ( .A(n_153), .Y(n_161) );
BUFx6f_ASAP7_75t_L g209 ( .A(n_153), .Y(n_209) );
INVx1_ASAP7_75t_L g494 ( .A(n_153), .Y(n_494) );
NOR2xp33_ASAP7_75t_L g158 ( .A(n_156), .B(n_159), .Y(n_158) );
INVx1_ASAP7_75t_L g451 ( .A(n_156), .Y(n_451) );
AOI21xp5_ASAP7_75t_L g503 ( .A1(n_156), .A2(n_504), .B(n_505), .Y(n_503) );
INVx4_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
OAI22xp5_ASAP7_75t_SL g235 ( .A1(n_157), .A2(n_236), .B1(n_237), .B2(n_238), .Y(n_235) );
INVx2_ASAP7_75t_L g237 ( .A(n_157), .Y(n_237) );
INVx1_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx2_ASAP7_75t_L g178 ( .A(n_161), .Y(n_178) );
OAI22xp33_ASAP7_75t_L g231 ( .A1(n_162), .A2(n_187), .B1(n_232), .B2(n_239), .Y(n_231) );
INVx4_ASAP7_75t_L g183 ( .A(n_164), .Y(n_183) );
OA21x2_ASAP7_75t_L g242 ( .A1(n_164), .A2(n_243), .B(n_249), .Y(n_242) );
OA21x2_ASAP7_75t_L g472 ( .A1(n_164), .A2(n_473), .B(n_480), .Y(n_472) );
BUFx6f_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
INVx1_ASAP7_75t_L g180 ( .A(n_165), .Y(n_180) );
INVx4_ASAP7_75t_L g271 ( .A(n_166), .Y(n_271) );
OAI21xp5_ASAP7_75t_L g326 ( .A1(n_166), .A2(n_327), .B(n_329), .Y(n_326) );
AND2x2_ASAP7_75t_L g407 ( .A(n_166), .B(n_408), .Y(n_407) );
AND2x2_ASAP7_75t_L g166 ( .A(n_167), .B(n_184), .Y(n_166) );
INVx1_ASAP7_75t_L g214 ( .A(n_167), .Y(n_214) );
AND2x2_ASAP7_75t_L g276 ( .A(n_167), .B(n_216), .Y(n_276) );
OR2x2_ASAP7_75t_L g305 ( .A(n_167), .B(n_306), .Y(n_305) );
INVx2_ASAP7_75t_L g319 ( .A(n_167), .Y(n_319) );
INVx3_ASAP7_75t_L g328 ( .A(n_167), .Y(n_328) );
AND2x2_ASAP7_75t_L g338 ( .A(n_167), .B(n_339), .Y(n_338) );
AND2x2_ASAP7_75t_L g371 ( .A(n_167), .B(n_277), .Y(n_371) );
AND2x2_ASAP7_75t_L g395 ( .A(n_167), .B(n_351), .Y(n_395) );
OR2x6_ASAP7_75t_L g167 ( .A(n_168), .B(n_181), .Y(n_167) );
AOI21xp5_ASAP7_75t_SL g168 ( .A1(n_169), .A2(n_170), .B(n_179), .Y(n_168) );
AOI21xp5_ASAP7_75t_L g171 ( .A1(n_172), .A2(n_175), .B(n_177), .Y(n_171) );
O2A1O1Ixp33_ASAP7_75t_L g258 ( .A1(n_173), .A2(n_259), .B(n_260), .C(n_261), .Y(n_258) );
INVx2_ASAP7_75t_L g457 ( .A(n_173), .Y(n_457) );
AOI21xp5_ASAP7_75t_L g462 ( .A1(n_173), .A2(n_463), .B(n_464), .Y(n_462) );
AOI21xp5_ASAP7_75t_L g474 ( .A1(n_173), .A2(n_475), .B(n_476), .Y(n_474) );
O2A1O1Ixp5_ASAP7_75t_SL g500 ( .A1(n_173), .A2(n_227), .B(n_501), .C(n_502), .Y(n_500) );
INVx5_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
NOR2xp33_ASAP7_75t_L g225 ( .A(n_174), .B(n_226), .Y(n_225) );
NOR2xp33_ASAP7_75t_L g247 ( .A(n_174), .B(n_248), .Y(n_247) );
OAI22xp5_ASAP7_75t_SL g492 ( .A1(n_174), .A2(n_191), .B1(n_493), .B2(n_495), .Y(n_492) );
INVx1_ASAP7_75t_L g512 ( .A(n_176), .Y(n_512) );
AOI21xp5_ASAP7_75t_L g189 ( .A1(n_177), .A2(n_190), .B(n_192), .Y(n_189) );
INVx2_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
INVx1_ASAP7_75t_L g193 ( .A(n_179), .Y(n_193) );
OA21x2_ASAP7_75t_L g446 ( .A1(n_179), .A2(n_447), .B(n_458), .Y(n_446) );
OA21x2_ASAP7_75t_L g460 ( .A1(n_179), .A2(n_461), .B(n_469), .Y(n_460) );
INVx2_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
AO21x2_ASAP7_75t_L g230 ( .A1(n_180), .A2(n_231), .B(n_240), .Y(n_230) );
NOR2xp33_ASAP7_75t_L g240 ( .A(n_180), .B(n_241), .Y(n_240) );
AO21x2_ASAP7_75t_L g254 ( .A1(n_180), .A2(n_255), .B(n_262), .Y(n_254) );
NOR2xp33_ASAP7_75t_SL g181 ( .A(n_182), .B(n_183), .Y(n_181) );
INVx3_ASAP7_75t_L g219 ( .A(n_183), .Y(n_219) );
NAND3xp33_ASAP7_75t_L g483 ( .A(n_183), .B(n_468), .C(n_484), .Y(n_483) );
AO21x1_ASAP7_75t_L g562 ( .A1(n_183), .A2(n_484), .B(n_563), .Y(n_562) );
INVx2_ASAP7_75t_L g216 ( .A(n_184), .Y(n_216) );
AND2x2_ASAP7_75t_L g431 ( .A(n_184), .B(n_273), .Y(n_431) );
AO21x2_ASAP7_75t_L g184 ( .A1(n_185), .A2(n_193), .B(n_194), .Y(n_184) );
OAI21xp5_ASAP7_75t_L g185 ( .A1(n_186), .A2(n_187), .B(n_188), .Y(n_185) );
OAI21xp5_ASAP7_75t_L g255 ( .A1(n_187), .A2(n_256), .B(n_257), .Y(n_255) );
INVx4_ASAP7_75t_L g207 ( .A(n_191), .Y(n_207) );
INVx2_ASAP7_75t_L g224 ( .A(n_191), .Y(n_224) );
OAI22xp5_ASAP7_75t_L g484 ( .A1(n_191), .A2(n_457), .B1(n_485), .B2(n_486), .Y(n_484) );
OAI22xp5_ASAP7_75t_L g529 ( .A1(n_191), .A2(n_457), .B1(n_530), .B2(n_531), .Y(n_529) );
NOR2xp33_ASAP7_75t_L g194 ( .A(n_195), .B(n_196), .Y(n_194) );
NOR2xp33_ASAP7_75t_L g211 ( .A(n_196), .B(n_212), .Y(n_211) );
NOR2xp33_ASAP7_75t_L g262 ( .A(n_196), .B(n_263), .Y(n_262) );
AND2x2_ASAP7_75t_L g197 ( .A(n_198), .B(n_213), .Y(n_197) );
INVx1_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
NOR2xp33_ASAP7_75t_L g327 ( .A(n_199), .B(n_328), .Y(n_327) );
AND2x2_ASAP7_75t_L g351 ( .A(n_199), .B(n_339), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_199), .B(n_328), .Y(n_413) );
INVx1_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
INVx2_ASAP7_75t_L g273 ( .A(n_200), .Y(n_273) );
AND2x2_ASAP7_75t_L g277 ( .A(n_200), .B(n_278), .Y(n_277) );
AND2x2_ASAP7_75t_L g318 ( .A(n_200), .B(n_319), .Y(n_318) );
AO21x2_ASAP7_75t_L g200 ( .A1(n_201), .A2(n_202), .B(n_211), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_203), .B(n_210), .Y(n_202) );
AOI21xp5_ASAP7_75t_L g204 ( .A1(n_205), .A2(n_206), .B(n_208), .Y(n_204) );
HB1xp67_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
INVx3_ASAP7_75t_L g227 ( .A(n_209), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_213), .B(n_314), .Y(n_336) );
INVx1_ASAP7_75t_L g375 ( .A(n_213), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_213), .B(n_302), .Y(n_419) );
AND2x2_ASAP7_75t_L g213 ( .A(n_214), .B(n_215), .Y(n_213) );
AND2x2_ASAP7_75t_L g282 ( .A(n_214), .B(n_277), .Y(n_282) );
INVx2_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_216), .B(n_273), .Y(n_306) );
INVx1_ASAP7_75t_L g385 ( .A(n_216), .Y(n_385) );
AOI322xp5_ASAP7_75t_L g409 ( .A1(n_217), .A2(n_324), .A3(n_384), .B1(n_410), .B2(n_412), .C1(n_414), .C2(n_416), .Y(n_409) );
AND2x2_ASAP7_75t_SL g217 ( .A(n_218), .B(n_229), .Y(n_217) );
AND2x2_ASAP7_75t_L g264 ( .A(n_218), .B(n_242), .Y(n_264) );
INVx1_ASAP7_75t_SL g267 ( .A(n_218), .Y(n_267) );
AND2x2_ASAP7_75t_L g269 ( .A(n_218), .B(n_230), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_218), .B(n_286), .Y(n_292) );
INVx2_ASAP7_75t_L g311 ( .A(n_218), .Y(n_311) );
AND2x2_ASAP7_75t_L g324 ( .A(n_218), .B(n_325), .Y(n_324) );
OR2x2_ASAP7_75t_L g362 ( .A(n_218), .B(n_286), .Y(n_362) );
BUFx2_ASAP7_75t_L g379 ( .A(n_218), .Y(n_379) );
AND2x2_ASAP7_75t_L g393 ( .A(n_218), .B(n_253), .Y(n_393) );
OA21x2_ASAP7_75t_L g218 ( .A1(n_219), .A2(n_220), .B(n_228), .Y(n_218) );
O2A1O1Ixp5_ASAP7_75t_L g465 ( .A1(n_224), .A2(n_453), .B(n_466), .C(n_467), .Y(n_465) );
AOI21xp5_ASAP7_75t_L g513 ( .A1(n_224), .A2(n_514), .B(n_515), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_229), .B(n_281), .Y(n_308) );
AND2x2_ASAP7_75t_L g435 ( .A(n_229), .B(n_311), .Y(n_435) );
AND2x2_ASAP7_75t_L g229 ( .A(n_230), .B(n_242), .Y(n_229) );
OR2x2_ASAP7_75t_L g280 ( .A(n_230), .B(n_281), .Y(n_280) );
INVx3_ASAP7_75t_L g286 ( .A(n_230), .Y(n_286) );
AND2x2_ASAP7_75t_L g331 ( .A(n_230), .B(n_254), .Y(n_331) );
NOR2xp33_ASAP7_75t_L g378 ( .A(n_230), .B(n_379), .Y(n_378) );
HB1xp67_ASAP7_75t_L g415 ( .A(n_230), .Y(n_415) );
INVx2_ASAP7_75t_L g261 ( .A(n_233), .Y(n_261) );
INVx3_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
AND2x2_ASAP7_75t_L g266 ( .A(n_242), .B(n_267), .Y(n_266) );
INVx1_ASAP7_75t_L g288 ( .A(n_242), .Y(n_288) );
BUFx2_ASAP7_75t_L g294 ( .A(n_242), .Y(n_294) );
AND2x2_ASAP7_75t_L g313 ( .A(n_242), .B(n_286), .Y(n_313) );
INVx3_ASAP7_75t_L g325 ( .A(n_242), .Y(n_325) );
OR2x2_ASAP7_75t_L g335 ( .A(n_242), .B(n_286), .Y(n_335) );
AOI31xp33_ASAP7_75t_SL g250 ( .A1(n_251), .A2(n_265), .A3(n_268), .B(n_270), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_252), .B(n_264), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_252), .B(n_287), .Y(n_298) );
OR2x2_ASAP7_75t_L g322 ( .A(n_252), .B(n_292), .Y(n_322) );
INVx1_ASAP7_75t_SL g252 ( .A(n_253), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_253), .B(n_266), .Y(n_265) );
OR2x2_ASAP7_75t_L g343 ( .A(n_253), .B(n_335), .Y(n_343) );
NOR2xp33_ASAP7_75t_L g353 ( .A(n_253), .B(n_325), .Y(n_353) );
AND2x2_ASAP7_75t_L g360 ( .A(n_253), .B(n_361), .Y(n_360) );
NAND2x1_ASAP7_75t_L g388 ( .A(n_253), .B(n_324), .Y(n_388) );
NOR2xp33_ASAP7_75t_L g389 ( .A(n_253), .B(n_379), .Y(n_389) );
AND2x2_ASAP7_75t_L g401 ( .A(n_253), .B(n_286), .Y(n_401) );
INVx3_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
INVx3_ASAP7_75t_L g281 ( .A(n_254), .Y(n_281) );
O2A1O1Ixp33_ASAP7_75t_L g448 ( .A1(n_261), .A2(n_449), .B(n_450), .C(n_451), .Y(n_448) );
INVx1_ASAP7_75t_L g347 ( .A(n_264), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_264), .B(n_401), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_266), .B(n_342), .Y(n_376) );
AND2x4_ASAP7_75t_L g287 ( .A(n_267), .B(n_288), .Y(n_287) );
CKINVDCx16_ASAP7_75t_R g268 ( .A(n_269), .Y(n_268) );
OR2x2_ASAP7_75t_L g270 ( .A(n_271), .B(n_272), .Y(n_270) );
INVx2_ASAP7_75t_L g366 ( .A(n_272), .Y(n_366) );
NOR2xp33_ASAP7_75t_L g383 ( .A(n_272), .B(n_384), .Y(n_383) );
AND2x2_ASAP7_75t_L g314 ( .A(n_273), .B(n_304), .Y(n_314) );
AND2x2_ASAP7_75t_L g408 ( .A(n_273), .B(n_278), .Y(n_408) );
INVx1_ASAP7_75t_L g433 ( .A(n_273), .Y(n_433) );
AOI221xp5_ASAP7_75t_L g274 ( .A1(n_275), .A2(n_279), .B1(n_282), .B2(n_283), .C(n_289), .Y(n_274) );
CKINVDCx14_ASAP7_75t_R g295 ( .A(n_275), .Y(n_295) );
AND2x2_ASAP7_75t_L g275 ( .A(n_276), .B(n_277), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_276), .B(n_297), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_279), .B(n_330), .Y(n_349) );
INVx3_ASAP7_75t_SL g279 ( .A(n_280), .Y(n_279) );
OR2x2_ASAP7_75t_L g398 ( .A(n_280), .B(n_294), .Y(n_398) );
AND2x2_ASAP7_75t_L g312 ( .A(n_281), .B(n_313), .Y(n_312) );
INVx1_ASAP7_75t_L g342 ( .A(n_281), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_281), .B(n_325), .Y(n_370) );
NOR3xp33_ASAP7_75t_L g412 ( .A(n_281), .B(n_382), .C(n_413), .Y(n_412) );
AOI211xp5_ASAP7_75t_SL g345 ( .A1(n_282), .A2(n_346), .B(n_348), .C(n_356), .Y(n_345) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
OAI22xp33_ASAP7_75t_L g334 ( .A1(n_284), .A2(n_335), .B1(n_336), .B2(n_337), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_285), .B(n_287), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_285), .B(n_324), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_285), .B(n_369), .Y(n_368) );
BUFx2_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
AND2x2_ASAP7_75t_L g427 ( .A(n_287), .B(n_401), .Y(n_427) );
OAI22xp5_ASAP7_75t_L g289 ( .A1(n_290), .A2(n_295), .B1(n_296), .B2(n_298), .Y(n_289) );
NOR2xp33_ASAP7_75t_SL g290 ( .A(n_291), .B(n_293), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_293), .B(n_342), .Y(n_373) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
OAI22xp5_ASAP7_75t_L g425 ( .A1(n_296), .A2(n_388), .B1(n_419), .B2(n_426), .Y(n_425) );
AOI221xp5_ASAP7_75t_L g299 ( .A1(n_300), .A2(n_307), .B1(n_309), .B2(n_314), .C(n_315), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
OR2x2_ASAP7_75t_L g301 ( .A(n_302), .B(n_305), .Y(n_301) );
HB1xp67_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
INVxp67_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
OAI221xp5_ASAP7_75t_L g315 ( .A1(n_305), .A2(n_316), .B1(n_322), .B2(n_323), .C(n_326), .Y(n_315) );
INVx1_ASAP7_75t_L g358 ( .A(n_306), .Y(n_358) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_311), .B(n_312), .Y(n_310) );
INVx1_ASAP7_75t_SL g330 ( .A(n_311), .Y(n_330) );
OR2x2_ASAP7_75t_L g403 ( .A(n_311), .B(n_335), .Y(n_403) );
AND2x2_ASAP7_75t_L g405 ( .A(n_311), .B(n_313), .Y(n_405) );
INVx1_ASAP7_75t_L g344 ( .A(n_314), .Y(n_344) );
OR2x2_ASAP7_75t_L g316 ( .A(n_317), .B(n_320), .Y(n_316) );
AOI21xp33_ASAP7_75t_SL g374 ( .A1(n_317), .A2(n_375), .B(n_376), .Y(n_374) );
OR2x2_ASAP7_75t_L g381 ( .A(n_317), .B(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
AND2x2_ASAP7_75t_L g355 ( .A(n_318), .B(n_339), .Y(n_355) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
NAND2xp33_ASAP7_75t_SL g372 ( .A(n_323), .B(n_373), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_324), .B(n_342), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_325), .B(n_361), .Y(n_424) );
O2A1O1Ixp33_ASAP7_75t_L g340 ( .A1(n_328), .A2(n_341), .B(n_343), .C(n_344), .Y(n_340) );
NAND2x1_ASAP7_75t_SL g365 ( .A(n_328), .B(n_366), .Y(n_365) );
AOI22xp5_ASAP7_75t_L g377 ( .A1(n_329), .A2(n_378), .B1(n_380), .B2(n_383), .Y(n_377) );
AND2x2_ASAP7_75t_L g329 ( .A(n_330), .B(n_331), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_331), .B(n_421), .Y(n_420) );
NAND5xp2_ASAP7_75t_L g332 ( .A(n_333), .B(n_345), .C(n_363), .D(n_377), .E(n_386), .Y(n_332) );
NOR2xp33_ASAP7_75t_L g333 ( .A(n_334), .B(n_340), .Y(n_333) );
INVx1_ASAP7_75t_L g390 ( .A(n_336), .Y(n_390) );
INVx1_ASAP7_75t_SL g337 ( .A(n_338), .Y(n_337) );
AOI221xp5_ASAP7_75t_L g396 ( .A1(n_338), .A2(n_357), .B1(n_397), .B2(n_399), .C(n_402), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_339), .B(n_433), .Y(n_432) );
NOR2xp33_ASAP7_75t_L g346 ( .A(n_342), .B(n_347), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_342), .B(n_408), .Y(n_411) );
OAI22xp5_ASAP7_75t_L g348 ( .A1(n_349), .A2(n_350), .B1(n_352), .B2(n_354), .Y(n_348) );
INVx1_ASAP7_75t_SL g350 ( .A(n_351), .Y(n_350) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
AND2x2_ASAP7_75t_L g356 ( .A(n_357), .B(n_360), .Y(n_356) );
AND2x2_ASAP7_75t_L g357 ( .A(n_358), .B(n_359), .Y(n_357) );
AND2x2_ASAP7_75t_L g430 ( .A(n_359), .B(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
AOI221xp5_ASAP7_75t_L g363 ( .A1(n_364), .A2(n_367), .B1(n_371), .B2(n_372), .C(n_374), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
AND2x2_ASAP7_75t_L g414 ( .A(n_369), .B(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVx1_ASAP7_75t_SL g421 ( .A(n_379), .Y(n_421) );
INVx1_ASAP7_75t_SL g380 ( .A(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
OAI21xp5_ASAP7_75t_SL g386 ( .A1(n_387), .A2(n_389), .B(n_390), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
OAI211xp5_ASAP7_75t_SL g391 ( .A1(n_392), .A2(n_394), .B(n_396), .C(n_409), .Y(n_391) );
INVx1_ASAP7_75t_SL g392 ( .A(n_393), .Y(n_392) );
A2O1A1Ixp33_ASAP7_75t_L g418 ( .A1(n_394), .A2(n_419), .B(n_420), .C(n_422), .Y(n_418) );
INVx1_ASAP7_75t_SL g394 ( .A(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
NAND2xp5_ASAP7_75t_SL g399 ( .A(n_398), .B(n_400), .Y(n_399) );
AOI21xp33_ASAP7_75t_L g402 ( .A1(n_403), .A2(n_404), .B(n_406), .Y(n_402) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx2_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
AOI21xp33_ASAP7_75t_L g428 ( .A1(n_429), .A2(n_432), .B(n_434), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx2_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx2_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx1_ASAP7_75t_L g717 ( .A(n_439), .Y(n_717) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx2_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
OR5x1_ASAP7_75t_L g441 ( .A(n_442), .B(n_605), .C(n_663), .D(n_699), .E(n_706), .Y(n_441) );
NAND3xp33_ASAP7_75t_SL g442 ( .A(n_443), .B(n_551), .C(n_575), .Y(n_442) );
AOI221xp5_ASAP7_75t_L g443 ( .A1(n_444), .A2(n_487), .B1(n_517), .B2(n_522), .C(n_532), .Y(n_443) );
OAI21xp5_ASAP7_75t_SL g685 ( .A1(n_444), .A2(n_686), .B(n_688), .Y(n_685) );
AND2x2_ASAP7_75t_L g444 ( .A(n_445), .B(n_470), .Y(n_444) );
NAND2x1p5_ASAP7_75t_L g675 ( .A(n_445), .B(n_676), .Y(n_675) );
AND2x2_ASAP7_75t_L g445 ( .A(n_446), .B(n_459), .Y(n_445) );
INVx2_ASAP7_75t_L g521 ( .A(n_446), .Y(n_521) );
AND2x2_ASAP7_75t_L g534 ( .A(n_446), .B(n_472), .Y(n_534) );
AND2x2_ASAP7_75t_L g588 ( .A(n_446), .B(n_471), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_446), .B(n_460), .Y(n_603) );
O2A1O1Ixp33_ASAP7_75t_L g452 ( .A1(n_453), .A2(n_455), .B(n_456), .C(n_457), .Y(n_452) );
INVx2_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
AOI21xp5_ASAP7_75t_L g477 ( .A1(n_457), .A2(n_478), .B(n_479), .Y(n_477) );
AND2x2_ASAP7_75t_L g621 ( .A(n_459), .B(n_562), .Y(n_621) );
AND2x2_ASAP7_75t_L g654 ( .A(n_459), .B(n_472), .Y(n_654) );
INVx2_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
OR2x2_ASAP7_75t_L g561 ( .A(n_460), .B(n_562), .Y(n_561) );
AND2x2_ASAP7_75t_L g574 ( .A(n_460), .B(n_472), .Y(n_574) );
AND2x2_ASAP7_75t_L g581 ( .A(n_460), .B(n_562), .Y(n_581) );
HB1xp67_ASAP7_75t_L g590 ( .A(n_460), .Y(n_590) );
AND2x2_ASAP7_75t_L g597 ( .A(n_460), .B(n_471), .Y(n_597) );
INVx1_ASAP7_75t_L g628 ( .A(n_460), .Y(n_628) );
OAI21xp5_ASAP7_75t_L g461 ( .A1(n_462), .A2(n_465), .B(n_468), .Y(n_461) );
INVx1_ASAP7_75t_L g604 ( .A(n_470), .Y(n_604) );
AND2x2_ASAP7_75t_L g470 ( .A(n_471), .B(n_481), .Y(n_470) );
INVx2_ASAP7_75t_L g560 ( .A(n_471), .Y(n_560) );
AND2x2_ASAP7_75t_L g582 ( .A(n_471), .B(n_521), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_471), .B(n_628), .Y(n_633) );
INVx3_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_472), .B(n_521), .Y(n_520) );
AND2x2_ASAP7_75t_L g705 ( .A(n_472), .B(n_669), .Y(n_705) );
INVx2_ASAP7_75t_L g519 ( .A(n_481), .Y(n_519) );
INVx3_ASAP7_75t_L g620 ( .A(n_481), .Y(n_620) );
OR2x2_ASAP7_75t_L g650 ( .A(n_481), .B(n_651), .Y(n_650) );
NOR2x1_ASAP7_75t_L g676 ( .A(n_481), .B(n_560), .Y(n_676) );
AND2x4_ASAP7_75t_L g481 ( .A(n_482), .B(n_483), .Y(n_481) );
INVx1_ASAP7_75t_L g563 ( .A(n_482), .Y(n_563) );
AOI33xp33_ASAP7_75t_L g696 ( .A1(n_487), .A2(n_534), .A3(n_548), .B1(n_620), .B2(n_697), .B3(n_698), .Y(n_696) );
INVx1_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
OR2x2_ASAP7_75t_L g488 ( .A(n_489), .B(n_496), .Y(n_488) );
OR2x2_ASAP7_75t_L g549 ( .A(n_489), .B(n_550), .Y(n_549) );
NOR2xp33_ASAP7_75t_L g608 ( .A(n_489), .B(n_546), .Y(n_608) );
OR2x2_ASAP7_75t_L g661 ( .A(n_489), .B(n_662), .Y(n_661) );
INVx2_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
AND2x2_ASAP7_75t_L g587 ( .A(n_490), .B(n_588), .Y(n_587) );
OR2x2_ASAP7_75t_L g612 ( .A(n_490), .B(n_496), .Y(n_612) );
AND2x2_ASAP7_75t_L g679 ( .A(n_490), .B(n_524), .Y(n_679) );
AOI21xp5_ASAP7_75t_L g704 ( .A1(n_490), .A2(n_579), .B(n_705), .Y(n_704) );
BUFx6f_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
INVx1_ASAP7_75t_L g526 ( .A(n_491), .Y(n_526) );
INVx1_ASAP7_75t_L g539 ( .A(n_491), .Y(n_539) );
AND2x2_ASAP7_75t_L g558 ( .A(n_491), .B(n_528), .Y(n_558) );
AND2x2_ASAP7_75t_L g607 ( .A(n_491), .B(n_527), .Y(n_607) );
INVx2_ASAP7_75t_SL g649 ( .A(n_496), .Y(n_649) );
OR2x2_ASAP7_75t_L g496 ( .A(n_497), .B(n_507), .Y(n_496) );
INVx2_ASAP7_75t_L g569 ( .A(n_497), .Y(n_569) );
INVx1_ASAP7_75t_L g700 ( .A(n_497), .Y(n_700) );
AND2x2_ASAP7_75t_L g713 ( .A(n_497), .B(n_594), .Y(n_713) );
INVx2_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
INVx2_ASAP7_75t_L g540 ( .A(n_498), .Y(n_540) );
OR2x2_ASAP7_75t_L g546 ( .A(n_498), .B(n_547), .Y(n_546) );
HB1xp67_ASAP7_75t_L g557 ( .A(n_498), .Y(n_557) );
HB1xp67_ASAP7_75t_L g524 ( .A(n_507), .Y(n_524) );
AND2x2_ASAP7_75t_L g541 ( .A(n_507), .B(n_527), .Y(n_541) );
INVx1_ASAP7_75t_L g547 ( .A(n_507), .Y(n_547) );
INVx1_ASAP7_75t_L g554 ( .A(n_507), .Y(n_554) );
AND2x2_ASAP7_75t_L g579 ( .A(n_507), .B(n_528), .Y(n_579) );
INVx2_ASAP7_75t_L g595 ( .A(n_507), .Y(n_595) );
AND2x2_ASAP7_75t_L g688 ( .A(n_507), .B(n_689), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_507), .B(n_569), .Y(n_709) );
AOI21xp5_ASAP7_75t_L g509 ( .A1(n_510), .A2(n_511), .B(n_512), .Y(n_509) );
INVx1_ASAP7_75t_SL g517 ( .A(n_518), .Y(n_517) );
OR2x2_ASAP7_75t_L g518 ( .A(n_519), .B(n_520), .Y(n_518) );
INVx2_ASAP7_75t_L g543 ( .A(n_519), .Y(n_543) );
INVx1_ASAP7_75t_L g572 ( .A(n_519), .Y(n_572) );
NOR2xp33_ASAP7_75t_L g669 ( .A(n_519), .B(n_603), .Y(n_669) );
INVx1_ASAP7_75t_SL g629 ( .A(n_520), .Y(n_629) );
INVx2_ASAP7_75t_L g550 ( .A(n_521), .Y(n_550) );
AND2x2_ASAP7_75t_L g619 ( .A(n_521), .B(n_620), .Y(n_619) );
AND2x2_ASAP7_75t_L g635 ( .A(n_521), .B(n_636), .Y(n_635) );
AND2x2_ASAP7_75t_L g522 ( .A(n_523), .B(n_525), .Y(n_522) );
INVx1_ASAP7_75t_L g697 ( .A(n_523), .Y(n_697) );
INVx1_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
AND2x2_ASAP7_75t_L g552 ( .A(n_525), .B(n_553), .Y(n_552) );
AND2x2_ASAP7_75t_L g655 ( .A(n_525), .B(n_645), .Y(n_655) );
AOI21xp5_ASAP7_75t_L g707 ( .A1(n_525), .A2(n_666), .B(n_708), .Y(n_707) );
AND2x2_ASAP7_75t_L g525 ( .A(n_526), .B(n_527), .Y(n_525) );
AND2x2_ASAP7_75t_L g568 ( .A(n_526), .B(n_569), .Y(n_568) );
BUFx2_ASAP7_75t_L g593 ( .A(n_526), .Y(n_593) );
INVx1_ASAP7_75t_L g617 ( .A(n_526), .Y(n_617) );
OR2x2_ASAP7_75t_L g681 ( .A(n_527), .B(n_540), .Y(n_681) );
NOR2xp67_ASAP7_75t_L g689 ( .A(n_527), .B(n_690), .Y(n_689) );
INVx2_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
AND2x2_ASAP7_75t_L g594 ( .A(n_528), .B(n_595), .Y(n_594) );
BUFx2_ASAP7_75t_L g601 ( .A(n_528), .Y(n_601) );
OAI22xp5_ASAP7_75t_L g532 ( .A1(n_533), .A2(n_535), .B1(n_542), .B2(n_544), .Y(n_532) );
OR2x2_ASAP7_75t_L g611 ( .A(n_533), .B(n_561), .Y(n_611) );
INVx1_ASAP7_75t_SL g533 ( .A(n_534), .Y(n_533) );
AOI222xp33_ASAP7_75t_L g652 ( .A1(n_534), .A2(n_653), .B1(n_655), .B2(n_656), .C1(n_657), .C2(n_660), .Y(n_652) );
INVx1_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
AND2x2_ASAP7_75t_L g536 ( .A(n_537), .B(n_541), .Y(n_536) );
INVx1_ASAP7_75t_SL g537 ( .A(n_538), .Y(n_537) );
OR2x2_ASAP7_75t_L g599 ( .A(n_538), .B(n_600), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_539), .B(n_540), .Y(n_538) );
AND2x2_ASAP7_75t_SL g553 ( .A(n_540), .B(n_554), .Y(n_553) );
HB1xp67_ASAP7_75t_L g624 ( .A(n_540), .Y(n_624) );
AND2x2_ASAP7_75t_L g672 ( .A(n_540), .B(n_541), .Y(n_672) );
INVx1_ASAP7_75t_L g690 ( .A(n_540), .Y(n_690) );
INVx1_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
AND2x2_ASAP7_75t_L g656 ( .A(n_543), .B(n_582), .Y(n_656) );
AND2x2_ASAP7_75t_L g698 ( .A(n_543), .B(n_574), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_545), .B(n_548), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_545), .B(n_593), .Y(n_680) );
INVx2_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
NAND2xp5_ASAP7_75t_SL g577 ( .A(n_546), .B(n_578), .Y(n_577) );
INVx1_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
AND2x2_ASAP7_75t_L g573 ( .A(n_550), .B(n_574), .Y(n_573) );
INVx3_ASAP7_75t_L g641 ( .A(n_550), .Y(n_641) );
O2A1O1Ixp33_ASAP7_75t_L g551 ( .A1(n_552), .A2(n_555), .B(n_559), .C(n_564), .Y(n_551) );
INVxp67_ASAP7_75t_L g565 ( .A(n_552), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_553), .B(n_617), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_553), .B(n_600), .Y(n_695) );
BUFx3_ASAP7_75t_L g659 ( .A(n_554), .Y(n_659) );
INVx1_ASAP7_75t_L g566 ( .A(n_555), .Y(n_566) );
AND2x2_ASAP7_75t_L g555 ( .A(n_556), .B(n_558), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
AND2x2_ASAP7_75t_L g585 ( .A(n_557), .B(n_579), .Y(n_585) );
INVx1_ASAP7_75t_SL g625 ( .A(n_558), .Y(n_625) );
NOR2xp33_ASAP7_75t_L g559 ( .A(n_560), .B(n_561), .Y(n_559) );
INVx1_ASAP7_75t_L g615 ( .A(n_560), .Y(n_615) );
AND2x2_ASAP7_75t_L g638 ( .A(n_560), .B(n_621), .Y(n_638) );
INVx1_ASAP7_75t_SL g609 ( .A(n_561), .Y(n_609) );
INVx1_ASAP7_75t_L g636 ( .A(n_562), .Y(n_636) );
AOI31xp33_ASAP7_75t_L g564 ( .A1(n_565), .A2(n_566), .A3(n_567), .B(n_570), .Y(n_564) );
INVx1_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
AND2x2_ASAP7_75t_L g657 ( .A(n_568), .B(n_658), .Y(n_657) );
INVx1_ASAP7_75t_L g631 ( .A(n_569), .Y(n_631) );
BUFx2_ASAP7_75t_L g645 ( .A(n_569), .Y(n_645) );
AND2x2_ASAP7_75t_L g673 ( .A(n_569), .B(n_594), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_571), .B(n_573), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
INVx1_ASAP7_75t_SL g646 ( .A(n_573), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_574), .B(n_641), .Y(n_687) );
AND2x2_ASAP7_75t_L g694 ( .A(n_574), .B(n_620), .Y(n_694) );
AOI211xp5_ASAP7_75t_L g575 ( .A1(n_576), .A2(n_580), .B(n_583), .C(n_598), .Y(n_575) );
INVxp67_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
INVx2_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
AOI221xp5_ASAP7_75t_L g606 ( .A1(n_580), .A2(n_607), .B1(n_608), .B2(n_609), .C(n_610), .Y(n_606) );
AND2x2_ASAP7_75t_L g580 ( .A(n_581), .B(n_582), .Y(n_580) );
AND2x2_ASAP7_75t_L g614 ( .A(n_581), .B(n_615), .Y(n_614) );
INVx2_ASAP7_75t_L g651 ( .A(n_582), .Y(n_651) );
OAI32xp33_ASAP7_75t_L g583 ( .A1(n_584), .A2(n_586), .A3(n_589), .B1(n_591), .B2(n_596), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
O2A1O1Ixp33_ASAP7_75t_L g637 ( .A1(n_585), .A2(n_638), .B(n_639), .C(n_642), .Y(n_637) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
AND2x2_ASAP7_75t_L g592 ( .A(n_593), .B(n_594), .Y(n_592) );
OAI21xp5_ASAP7_75t_SL g701 ( .A1(n_593), .A2(n_702), .B(n_703), .Y(n_701) );
INVx1_ASAP7_75t_L g662 ( .A(n_594), .Y(n_662) );
INVxp67_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
NOR2xp33_ASAP7_75t_L g598 ( .A(n_599), .B(n_602), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_600), .B(n_631), .Y(n_630) );
AND2x2_ASAP7_75t_L g648 ( .A(n_600), .B(n_649), .Y(n_648) );
INVx2_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
INVx1_ASAP7_75t_L g665 ( .A(n_602), .Y(n_665) );
OR2x2_ASAP7_75t_L g602 ( .A(n_603), .B(n_604), .Y(n_602) );
NAND4xp25_ASAP7_75t_SL g605 ( .A(n_606), .B(n_618), .C(n_637), .D(n_652), .Y(n_605) );
AND2x2_ASAP7_75t_L g644 ( .A(n_607), .B(n_645), .Y(n_644) );
AND2x4_ASAP7_75t_L g666 ( .A(n_607), .B(n_659), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_609), .B(n_641), .Y(n_640) );
OAI22xp5_ASAP7_75t_L g610 ( .A1(n_611), .A2(n_612), .B1(n_613), .B2(n_616), .Y(n_610) );
OAI22xp5_ASAP7_75t_L g692 ( .A1(n_611), .A2(n_662), .B1(n_693), .B2(n_695), .Y(n_692) );
O2A1O1Ixp33_ASAP7_75t_L g699 ( .A1(n_611), .A2(n_700), .B(n_701), .C(n_704), .Y(n_699) );
INVx2_ASAP7_75t_L g670 ( .A(n_612), .Y(n_670) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
AOI222xp33_ASAP7_75t_L g664 ( .A1(n_614), .A2(n_648), .B1(n_665), .B2(n_666), .C1(n_667), .C2(n_670), .Y(n_664) );
O2A1O1Ixp33_ASAP7_75t_L g618 ( .A1(n_619), .A2(n_621), .B(n_622), .C(n_626), .Y(n_618) );
INVx1_ASAP7_75t_L g684 ( .A(n_619), .Y(n_684) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
OAI22xp33_ASAP7_75t_L g626 ( .A1(n_623), .A2(n_627), .B1(n_630), .B2(n_632), .Y(n_626) );
OR2x2_ASAP7_75t_L g623 ( .A(n_624), .B(n_625), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_628), .B(n_629), .Y(n_627) );
OR2x2_ASAP7_75t_L g632 ( .A(n_633), .B(n_634), .Y(n_632) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
AND2x2_ASAP7_75t_L g653 ( .A(n_635), .B(n_654), .Y(n_653) );
INVx1_ASAP7_75t_L g711 ( .A(n_638), .Y(n_711) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
OAI22xp33_ASAP7_75t_L g642 ( .A1(n_643), .A2(n_646), .B1(n_647), .B2(n_650), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_645), .B(n_679), .Y(n_678) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
INVx1_ASAP7_75t_L g702 ( .A(n_650), .Y(n_702) );
INVx1_ASAP7_75t_L g683 ( .A(n_654), .Y(n_683) );
CKINVDCx16_ASAP7_75t_R g710 ( .A(n_656), .Y(n_710) );
INVxp67_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
NAND5xp2_ASAP7_75t_L g663 ( .A(n_664), .B(n_671), .C(n_685), .D(n_691), .E(n_696), .Y(n_663) );
INVx1_ASAP7_75t_SL g667 ( .A(n_668), .Y(n_667) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
O2A1O1Ixp33_ASAP7_75t_L g671 ( .A1(n_672), .A2(n_673), .B(n_674), .C(n_677), .Y(n_671) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
AOI31xp33_ASAP7_75t_L g677 ( .A1(n_678), .A2(n_680), .A3(n_681), .B(n_682), .Y(n_677) );
INVx1_ASAP7_75t_L g703 ( .A(n_679), .Y(n_703) );
OR2x2_ASAP7_75t_L g682 ( .A(n_683), .B(n_684), .Y(n_682) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
OAI222xp33_ASAP7_75t_L g706 ( .A1(n_693), .A2(n_695), .B1(n_707), .B2(n_710), .C1(n_711), .C2(n_712), .Y(n_706) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
INVx2_ASAP7_75t_SL g712 ( .A(n_713), .Y(n_712) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVx2_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx1_ASAP7_75t_SL g721 ( .A(n_722), .Y(n_721) );
BUFx2_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
endmodule