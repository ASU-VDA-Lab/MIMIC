module fake_jpeg_30023_n_475 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_475);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_475;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_292;
wire n_213;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx14_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx8_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_3),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

CKINVDCx16_ASAP7_75t_R g28 ( 
.A(n_11),
.Y(n_28)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx8_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_1),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

BUFx12_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

CKINVDCx5p33_ASAP7_75t_R g42 ( 
.A(n_11),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_13),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_2),
.Y(n_45)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_15),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_2),
.Y(n_47)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_2),
.Y(n_48)
);

CKINVDCx16_ASAP7_75t_R g49 ( 
.A(n_8),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_37),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_50),
.B(n_52),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_24),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_51),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_30),
.B(n_7),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_42),
.B(n_8),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_53),
.B(n_66),
.Y(n_108)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_54),
.Y(n_124)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_55),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_24),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_56),
.Y(n_133)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_57),
.Y(n_112)
);

BUFx2_ASAP7_75t_L g58 ( 
.A(n_23),
.Y(n_58)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_58),
.Y(n_151)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_59),
.Y(n_117)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_48),
.Y(n_60)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_60),
.Y(n_126)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_20),
.Y(n_61)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_61),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_62),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_30),
.B(n_15),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_63),
.B(n_85),
.Y(n_131)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_64),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_24),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_65),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_42),
.B(n_15),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_24),
.Y(n_67)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_67),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_68),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_17),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_69),
.B(n_71),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_40),
.Y(n_70)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_70),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_18),
.Y(n_71)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_72),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_40),
.Y(n_73)
);

INVx6_ASAP7_75t_L g137 ( 
.A(n_73),
.Y(n_137)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_41),
.Y(n_74)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_74),
.Y(n_104)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_20),
.Y(n_75)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_75),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_17),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_76),
.B(n_78),
.Y(n_127)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_18),
.Y(n_77)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_77),
.Y(n_130)
);

BUFx4f_ASAP7_75t_SL g78 ( 
.A(n_42),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_28),
.B(n_14),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_79),
.B(n_80),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_23),
.B(n_33),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_40),
.Y(n_81)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_81),
.Y(n_107)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_41),
.Y(n_82)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_82),
.Y(n_123)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_27),
.Y(n_83)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_83),
.Y(n_134)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_18),
.Y(n_84)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_84),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_23),
.B(n_14),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_45),
.Y(n_86)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_86),
.Y(n_145)
);

INVx3_ASAP7_75t_SL g87 ( 
.A(n_31),
.Y(n_87)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_87),
.Y(n_140)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_45),
.Y(n_88)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_88),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_31),
.Y(n_89)
);

INVx5_ASAP7_75t_L g132 ( 
.A(n_89),
.Y(n_132)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_27),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_90),
.Y(n_125)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_46),
.Y(n_91)
);

NAND2xp33_ASAP7_75t_SL g102 ( 
.A(n_91),
.B(n_17),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_31),
.Y(n_92)
);

INVx5_ASAP7_75t_L g143 ( 
.A(n_92),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_23),
.B(n_14),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_93),
.B(n_33),
.Y(n_139)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_45),
.Y(n_94)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_94),
.Y(n_138)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_41),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_95),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_32),
.Y(n_96)
);

BUFx12f_ASAP7_75t_L g144 ( 
.A(n_96),
.Y(n_144)
);

OR2x2_ASAP7_75t_L g97 ( 
.A(n_43),
.B(n_14),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_97),
.B(n_98),
.Y(n_105)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_46),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g190 ( 
.A(n_102),
.B(n_112),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_97),
.A2(n_46),
.B1(n_32),
.B2(n_43),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_106),
.A2(n_115),
.B1(n_118),
.B2(n_120),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_89),
.A2(n_96),
.B1(n_92),
.B2(n_70),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g179 ( 
.A1(n_109),
.A2(n_121),
.B1(n_150),
.B2(n_29),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_87),
.A2(n_32),
.B1(n_41),
.B2(n_21),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_111),
.A2(n_113),
.B1(n_136),
.B2(n_148),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_59),
.A2(n_21),
.B1(n_22),
.B2(n_45),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_51),
.A2(n_21),
.B1(n_34),
.B2(n_26),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_86),
.A2(n_34),
.B1(n_25),
.B2(n_26),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_56),
.A2(n_25),
.B1(n_28),
.B2(n_49),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_65),
.A2(n_49),
.B1(n_22),
.B2(n_16),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_60),
.A2(n_47),
.B1(n_44),
.B2(n_39),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g198 ( 
.A(n_139),
.B(n_0),
.Y(n_198)
);

A2O1A1Ixp33_ASAP7_75t_L g142 ( 
.A1(n_78),
.A2(n_44),
.B(n_39),
.C(n_35),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_142),
.B(n_147),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_88),
.A2(n_16),
.B1(n_35),
.B2(n_47),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_146),
.A2(n_81),
.B1(n_73),
.B2(n_68),
.Y(n_167)
);

A2O1A1Ixp33_ASAP7_75t_L g147 ( 
.A1(n_78),
.A2(n_33),
.B(n_23),
.C(n_10),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_64),
.A2(n_47),
.B1(n_33),
.B2(n_10),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_67),
.A2(n_29),
.B1(n_19),
.B2(n_33),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_116),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_155),
.B(n_156),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_116),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_131),
.B(n_93),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_157),
.B(n_158),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_114),
.B(n_85),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_128),
.B(n_94),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_160),
.B(n_162),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_105),
.B(n_71),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_140),
.A2(n_58),
.B1(n_54),
.B2(n_62),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_163),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_134),
.A2(n_95),
.B1(n_82),
.B2(n_72),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_165),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_141),
.B(n_80),
.C(n_74),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_166),
.B(n_180),
.C(n_135),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_167),
.A2(n_201),
.B1(n_122),
.B2(n_137),
.Y(n_211)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_145),
.Y(n_168)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_168),
.Y(n_205)
);

INVx1_ASAP7_75t_SL g169 ( 
.A(n_151),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_169),
.B(n_189),
.Y(n_216)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_153),
.Y(n_170)
);

INVx1_ASAP7_75t_SL g236 ( 
.A(n_170),
.Y(n_236)
);

NOR2x1_ASAP7_75t_L g171 ( 
.A(n_118),
.B(n_47),
.Y(n_171)
);

OR2x2_ASAP7_75t_L g226 ( 
.A(n_171),
.B(n_184),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_100),
.B(n_47),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_172),
.B(n_185),
.Y(n_229)
);

HB1xp67_ASAP7_75t_L g173 ( 
.A(n_153),
.Y(n_173)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_173),
.Y(n_212)
);

HB1xp67_ASAP7_75t_L g174 ( 
.A(n_124),
.Y(n_174)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_174),
.Y(n_206)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_145),
.Y(n_175)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_175),
.Y(n_210)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_138),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g223 ( 
.A(n_176),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_127),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_177),
.B(n_183),
.Y(n_214)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_152),
.Y(n_178)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_178),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_179),
.A2(n_99),
.B1(n_107),
.B2(n_129),
.Y(n_237)
);

OR2x2_ASAP7_75t_SL g180 ( 
.A(n_147),
.B(n_142),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_102),
.A2(n_13),
.B(n_12),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_181),
.A2(n_159),
.B(n_190),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_132),
.A2(n_143),
.B1(n_130),
.B2(n_135),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_182),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_110),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_146),
.A2(n_29),
.B1(n_19),
.B2(n_38),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_108),
.B(n_38),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_151),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_186),
.B(n_187),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_125),
.B(n_12),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_138),
.Y(n_188)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_188),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_130),
.A2(n_19),
.B1(n_38),
.B2(n_12),
.Y(n_189)
);

AND2x2_ASAP7_75t_L g239 ( 
.A(n_190),
.B(n_198),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_112),
.B(n_9),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_191),
.B(n_129),
.Y(n_227)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_117),
.Y(n_192)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_192),
.Y(n_228)
);

OA22x2_ASAP7_75t_L g193 ( 
.A1(n_101),
.A2(n_38),
.B1(n_1),
.B2(n_2),
.Y(n_193)
);

O2A1O1Ixp33_ASAP7_75t_SL g235 ( 
.A1(n_193),
.A2(n_144),
.B(n_107),
.C(n_99),
.Y(n_235)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_117),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_194),
.B(n_196),
.Y(n_220)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_152),
.Y(n_195)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_195),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_149),
.B(n_123),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_132),
.A2(n_9),
.B1(n_38),
.B2(n_3),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_197),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_126),
.B(n_0),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_199),
.B(n_200),
.Y(n_233)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_126),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_101),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_201)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_144),
.Y(n_202)
);

INVx2_ASAP7_75t_SL g208 ( 
.A(n_202),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_211),
.A2(n_164),
.B1(n_161),
.B2(n_184),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_215),
.A2(n_190),
.B(n_181),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_196),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_221),
.B(n_183),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_222),
.B(n_240),
.C(n_215),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_159),
.A2(n_122),
.B1(n_137),
.B2(n_119),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_224),
.A2(n_225),
.B1(n_234),
.B2(n_189),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_L g225 ( 
.A1(n_167),
.A2(n_119),
.B1(n_154),
.B2(n_133),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_227),
.B(n_171),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_171),
.A2(n_143),
.B1(n_154),
.B2(n_133),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_235),
.A2(n_237),
.B1(n_231),
.B2(n_190),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_SL g238 ( 
.A(n_180),
.B(n_103),
.C(n_144),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_238),
.A2(n_169),
.B(n_193),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_166),
.B(n_124),
.C(n_123),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_240),
.B(n_158),
.C(n_198),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_227),
.B(n_160),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_241),
.B(n_242),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_207),
.B(n_191),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_243),
.A2(n_226),
.B1(n_234),
.B2(n_216),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_244),
.A2(n_264),
.B1(n_269),
.B2(n_218),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_245),
.B(n_246),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_214),
.B(n_177),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_207),
.B(n_199),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_247),
.B(n_254),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_SL g287 ( 
.A1(n_248),
.A2(n_274),
.B(n_216),
.Y(n_287)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_228),
.Y(n_249)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_249),
.Y(n_278)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_228),
.Y(n_250)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_250),
.Y(n_284)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_219),
.Y(n_251)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_251),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_252),
.B(n_256),
.C(n_257),
.Y(n_275)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_219),
.Y(n_253)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_253),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_221),
.B(n_198),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_204),
.Y(n_255)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_255),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_222),
.B(n_157),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_239),
.B(n_185),
.C(n_180),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_204),
.Y(n_258)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_258),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_214),
.B(n_172),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_259),
.B(n_271),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_SL g294 ( 
.A(n_260),
.B(n_268),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_261),
.B(n_239),
.C(n_229),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_233),
.B(n_187),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_262),
.B(n_267),
.Y(n_286)
);

INVx8_ASAP7_75t_L g263 ( 
.A(n_209),
.Y(n_263)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_263),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_226),
.A2(n_211),
.B1(n_235),
.B2(n_238),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_235),
.A2(n_164),
.B1(n_201),
.B2(n_193),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_265),
.A2(n_243),
.B1(n_267),
.B2(n_226),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_209),
.Y(n_266)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_266),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_233),
.B(n_193),
.Y(n_267)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_212),
.Y(n_270)
);

CKINVDCx16_ASAP7_75t_R g305 ( 
.A(n_270),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_220),
.B(n_162),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_209),
.Y(n_272)
);

AOI22xp33_ASAP7_75t_SL g300 ( 
.A1(n_272),
.A2(n_236),
.B1(n_208),
.B2(n_169),
.Y(n_300)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_212),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_273),
.B(n_223),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_L g274 ( 
.A1(n_239),
.A2(n_193),
.B(n_200),
.Y(n_274)
);

AOI32xp33_ASAP7_75t_L g276 ( 
.A1(n_274),
.A2(n_268),
.A3(n_264),
.B1(n_252),
.B2(n_248),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_SL g312 ( 
.A(n_276),
.B(n_261),
.C(n_259),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_256),
.B(n_257),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_277),
.B(n_288),
.C(n_301),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_279),
.A2(n_282),
.B1(n_292),
.B2(n_302),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_245),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_280),
.B(n_305),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_244),
.A2(n_237),
.B1(n_216),
.B2(n_230),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_283),
.B(n_289),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g329 ( 
.A(n_287),
.Y(n_329)
);

XNOR2x1_ASAP7_75t_SL g291 ( 
.A(n_254),
.B(n_239),
.Y(n_291)
);

XNOR2x1_ASAP7_75t_SL g311 ( 
.A(n_291),
.B(n_241),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_269),
.A2(n_216),
.B1(n_232),
.B2(n_217),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_297),
.B(n_304),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_SL g326 ( 
.A1(n_300),
.A2(n_236),
.B(n_208),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_256),
.B(n_229),
.C(n_203),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_265),
.A2(n_224),
.B1(n_225),
.B2(n_203),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_255),
.B(n_220),
.Y(n_304)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_298),
.Y(n_307)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_307),
.Y(n_338)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_298),
.Y(n_308)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_308),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_L g310 ( 
.A1(n_279),
.A2(n_258),
.B(n_260),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g351 ( 
.A(n_310),
.Y(n_351)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_311),
.B(n_294),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_SL g341 ( 
.A(n_312),
.B(n_316),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_280),
.B(n_242),
.Y(n_315)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_315),
.Y(n_347)
);

NOR2xp67_ASAP7_75t_SL g316 ( 
.A(n_294),
.B(n_246),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_299),
.B(n_304),
.Y(n_317)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_317),
.Y(n_360)
);

CKINVDCx16_ASAP7_75t_R g318 ( 
.A(n_289),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_318),
.B(n_320),
.Y(n_342)
);

CKINVDCx16_ASAP7_75t_R g320 ( 
.A(n_290),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_299),
.B(n_247),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_321),
.B(n_330),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_275),
.B(n_261),
.C(n_271),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_322),
.B(n_301),
.C(n_287),
.Y(n_344)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_278),
.Y(n_323)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_323),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_282),
.A2(n_262),
.B1(n_217),
.B2(n_270),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_324),
.A2(n_328),
.B1(n_306),
.B2(n_192),
.Y(n_358)
);

CKINVDCx16_ASAP7_75t_R g325 ( 
.A(n_290),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_325),
.B(n_326),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_277),
.B(n_273),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_327),
.B(n_335),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_302),
.A2(n_249),
.B1(n_250),
.B2(n_251),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_296),
.B(n_253),
.Y(n_330)
);

NAND3xp33_ASAP7_75t_L g331 ( 
.A(n_285),
.B(n_223),
.C(n_156),
.Y(n_331)
);

INVxp33_ASAP7_75t_L g362 ( 
.A(n_331),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_SL g332 ( 
.A(n_285),
.B(n_155),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_332),
.Y(n_355)
);

OAI22x1_ASAP7_75t_L g333 ( 
.A1(n_276),
.A2(n_208),
.B1(n_236),
.B2(n_263),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_L g340 ( 
.A1(n_333),
.A2(n_283),
.B1(n_297),
.B2(n_292),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_334),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_275),
.B(n_174),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_281),
.B(n_266),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_336),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_SL g375 ( 
.A(n_337),
.B(n_324),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_340),
.A2(n_316),
.B1(n_326),
.B2(n_311),
.Y(n_383)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_327),
.B(n_288),
.Y(n_343)
);

XOR2xp5_ASAP7_75t_L g366 ( 
.A(n_343),
.B(n_335),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_344),
.B(n_346),
.C(n_348),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_333),
.A2(n_286),
.B1(n_305),
.B2(n_303),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_345),
.A2(n_357),
.B1(n_314),
.B2(n_308),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_319),
.B(n_281),
.C(n_286),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_319),
.B(n_296),
.C(n_291),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_L g349 ( 
.A1(n_313),
.A2(n_295),
.B1(n_293),
.B2(n_284),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_L g374 ( 
.A1(n_349),
.A2(n_328),
.B1(n_309),
.B2(n_325),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_322),
.B(n_284),
.C(n_278),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_352),
.B(n_312),
.C(n_310),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_333),
.A2(n_303),
.B1(n_295),
.B2(n_293),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_358),
.A2(n_363),
.B1(n_318),
.B2(n_307),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_L g363 ( 
.A1(n_313),
.A2(n_306),
.B1(n_266),
.B2(n_263),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_317),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_364),
.B(n_320),
.Y(n_367)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_338),
.Y(n_365)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_365),
.Y(n_391)
);

XOR2xp5_ASAP7_75t_L g395 ( 
.A(n_366),
.B(n_375),
.Y(n_395)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_367),
.Y(n_400)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_338),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_368),
.B(n_376),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_SL g404 ( 
.A1(n_369),
.A2(n_377),
.B1(n_383),
.B2(n_359),
.Y(n_404)
);

CKINVDCx16_ASAP7_75t_R g370 ( 
.A(n_342),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_SL g408 ( 
.A(n_370),
.B(n_373),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_372),
.B(n_378),
.C(n_388),
.Y(n_401)
);

OAI21xp5_ASAP7_75t_SL g373 ( 
.A1(n_354),
.A2(n_329),
.B(n_351),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g392 ( 
.A1(n_374),
.A2(n_382),
.B1(n_358),
.B2(n_360),
.Y(n_392)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_339),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_351),
.A2(n_330),
.B1(n_309),
.B2(n_314),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_352),
.B(n_344),
.C(n_343),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_356),
.B(n_332),
.Y(n_379)
);

CKINVDCx14_ASAP7_75t_R g402 ( 
.A(n_379),
.Y(n_402)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_339),
.Y(n_380)
);

OR2x2_ASAP7_75t_L g406 ( 
.A(n_380),
.B(n_387),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_355),
.B(n_336),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_381),
.B(n_389),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_SL g384 ( 
.A(n_337),
.B(n_315),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g399 ( 
.A(n_384),
.B(n_386),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_L g385 ( 
.A1(n_355),
.A2(n_321),
.B1(n_323),
.B2(n_272),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_L g396 ( 
.A1(n_385),
.A2(n_347),
.B1(n_361),
.B2(n_350),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_SL g386 ( 
.A(n_341),
.B(n_206),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_360),
.Y(n_387)
);

XOR2xp5_ASAP7_75t_L g388 ( 
.A(n_353),
.B(n_173),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_356),
.B(n_206),
.Y(n_389)
);

OAI322xp33_ASAP7_75t_L g390 ( 
.A1(n_367),
.A2(n_341),
.A3(n_362),
.B1(n_364),
.B2(n_348),
.C1(n_346),
.C2(n_350),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_390),
.B(n_188),
.Y(n_425)
);

XOR2xp5_ASAP7_75t_L g421 ( 
.A(n_392),
.B(n_375),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_382),
.A2(n_363),
.B1(n_347),
.B2(n_361),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_SL g422 ( 
.A1(n_393),
.A2(n_403),
.B1(n_384),
.B2(n_388),
.Y(n_422)
);

OAI21xp5_ASAP7_75t_L g394 ( 
.A1(n_383),
.A2(n_345),
.B(n_357),
.Y(n_394)
);

AO21x1_ASAP7_75t_L g410 ( 
.A1(n_394),
.A2(n_381),
.B(n_377),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_L g413 ( 
.A1(n_396),
.A2(n_404),
.B1(n_400),
.B2(n_407),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_L g403 ( 
.A1(n_387),
.A2(n_359),
.B1(n_353),
.B2(n_208),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_SL g411 ( 
.A(n_404),
.B(n_386),
.Y(n_411)
);

BUFx24_ASAP7_75t_SL g405 ( 
.A(n_373),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_405),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_SL g407 ( 
.A1(n_369),
.A2(n_194),
.B1(n_210),
.B2(n_205),
.Y(n_407)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_407),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_L g436 ( 
.A(n_410),
.B(n_411),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_402),
.B(n_365),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_412),
.B(n_416),
.Y(n_433)
);

XOR2xp5_ASAP7_75t_L g434 ( 
.A(n_413),
.B(n_421),
.Y(n_434)
);

AOI21xp5_ASAP7_75t_L g414 ( 
.A1(n_394),
.A2(n_368),
.B(n_380),
.Y(n_414)
);

AOI21xp5_ASAP7_75t_L g429 ( 
.A1(n_414),
.A2(n_425),
.B(n_398),
.Y(n_429)
);

CKINVDCx16_ASAP7_75t_R g416 ( 
.A(n_406),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_401),
.B(n_378),
.C(n_371),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_417),
.B(n_418),
.C(n_420),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_401),
.B(n_371),
.C(n_366),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_406),
.B(n_376),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_419),
.B(n_423),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_403),
.B(n_372),
.C(n_395),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g437 ( 
.A(n_422),
.B(n_399),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_L g423 ( 
.A1(n_408),
.A2(n_213),
.B1(n_210),
.B2(n_205),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_400),
.A2(n_213),
.B1(n_170),
.B2(n_176),
.Y(n_424)
);

INVxp67_ASAP7_75t_L g426 ( 
.A(n_424),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_SL g427 ( 
.A(n_415),
.B(n_417),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_427),
.B(n_428),
.Y(n_450)
);

CKINVDCx16_ASAP7_75t_R g428 ( 
.A(n_419),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_SL g442 ( 
.A(n_429),
.B(n_437),
.Y(n_442)
);

AND2x2_ASAP7_75t_L g430 ( 
.A(n_425),
.B(n_393),
.Y(n_430)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_430),
.Y(n_445)
);

OAI21xp5_ASAP7_75t_L g432 ( 
.A1(n_420),
.A2(n_397),
.B(n_391),
.Y(n_432)
);

AOI21xp5_ASAP7_75t_L g446 ( 
.A1(n_432),
.A2(n_433),
.B(n_439),
.Y(n_446)
);

AOI21xp5_ASAP7_75t_L g435 ( 
.A1(n_412),
.A2(n_397),
.B(n_391),
.Y(n_435)
);

OAI21xp5_ASAP7_75t_SL g441 ( 
.A1(n_435),
.A2(n_409),
.B(n_410),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_418),
.B(n_395),
.C(n_392),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_438),
.B(n_421),
.C(n_422),
.Y(n_448)
);

INVxp67_ASAP7_75t_L g439 ( 
.A(n_414),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_439),
.B(n_436),
.Y(n_451)
);

AOI21xp5_ASAP7_75t_L g459 ( 
.A1(n_441),
.A2(n_449),
.B(n_202),
.Y(n_459)
);

BUFx3_ASAP7_75t_L g443 ( 
.A(n_434),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_443),
.B(n_446),
.Y(n_458)
);

NOR2xp67_ASAP7_75t_SL g444 ( 
.A(n_431),
.B(n_411),
.Y(n_444)
);

OAI21xp5_ASAP7_75t_L g461 ( 
.A1(n_444),
.A2(n_195),
.B(n_178),
.Y(n_461)
);

INVxp67_ASAP7_75t_L g447 ( 
.A(n_434),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_447),
.B(n_448),
.Y(n_460)
);

AOI21xp5_ASAP7_75t_L g449 ( 
.A1(n_430),
.A2(n_413),
.B(n_409),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_451),
.B(n_452),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_SL g452 ( 
.A1(n_426),
.A2(n_424),
.B1(n_399),
.B2(n_170),
.Y(n_452)
);

AOI21xp33_ASAP7_75t_L g453 ( 
.A1(n_450),
.A2(n_440),
.B(n_431),
.Y(n_453)
);

BUFx24_ASAP7_75t_SL g462 ( 
.A(n_453),
.Y(n_462)
);

OAI21xp5_ASAP7_75t_SL g455 ( 
.A1(n_442),
.A2(n_438),
.B(n_426),
.Y(n_455)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_455),
.Y(n_465)
);

NAND2x1p5_ASAP7_75t_L g456 ( 
.A(n_445),
.B(n_436),
.Y(n_456)
);

AOI22xp5_ASAP7_75t_SL g467 ( 
.A1(n_456),
.A2(n_175),
.B1(n_168),
.B2(n_104),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_443),
.B(n_437),
.Y(n_457)
);

XOR2xp5_ASAP7_75t_L g463 ( 
.A(n_457),
.B(n_459),
.Y(n_463)
);

OAI21xp5_ASAP7_75t_L g464 ( 
.A1(n_461),
.A2(n_449),
.B(n_452),
.Y(n_464)
);

AO21x1_ASAP7_75t_L g470 ( 
.A1(n_464),
.A2(n_466),
.B(n_467),
.Y(n_470)
);

OAI21xp5_ASAP7_75t_L g466 ( 
.A1(n_458),
.A2(n_448),
.B(n_447),
.Y(n_466)
);

A2O1A1O1Ixp25_ASAP7_75t_L g468 ( 
.A1(n_462),
.A2(n_460),
.B(n_456),
.C(n_454),
.D(n_104),
.Y(n_468)
);

NOR3xp33_ASAP7_75t_L g471 ( 
.A(n_468),
.B(n_469),
.C(n_465),
.Y(n_471)
);

OAI21x1_ASAP7_75t_L g469 ( 
.A1(n_463),
.A2(n_103),
.B(n_4),
.Y(n_469)
);

AOI321xp33_ASAP7_75t_L g473 ( 
.A1(n_471),
.A2(n_472),
.A3(n_4),
.B1(n_5),
.B2(n_6),
.C(n_416),
.Y(n_473)
);

OAI321xp33_ASAP7_75t_L g472 ( 
.A1(n_470),
.A2(n_3),
.A3(n_4),
.B1(n_5),
.B2(n_6),
.C(n_450),
.Y(n_472)
);

OAI21xp5_ASAP7_75t_SL g474 ( 
.A1(n_473),
.A2(n_4),
.B(n_5),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_SL g475 ( 
.A(n_474),
.B(n_5),
.Y(n_475)
);


endmodule