module fake_jpeg_14364_n_643 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_643);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_643;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_511;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_384;
wire n_296;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_538;
wire n_47;
wire n_312;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx13_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx16f_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

BUFx4f_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

BUFx8_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_4),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_16),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_6),
.Y(n_42)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_5),
.Y(n_44)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_8),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_9),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_9),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_12),
.Y(n_50)
);

BUFx10_ASAP7_75t_L g51 ( 
.A(n_0),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_7),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_7),
.Y(n_53)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_8),
.Y(n_54)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_15),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_10),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_11),
.Y(n_57)
);

BUFx12_ASAP7_75t_L g58 ( 
.A(n_3),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_4),
.Y(n_59)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_12),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_16),
.Y(n_61)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_60),
.Y(n_62)
);

INVx5_ASAP7_75t_L g153 ( 
.A(n_62),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_61),
.B(n_9),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_63),
.B(n_71),
.Y(n_197)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_64),
.Y(n_130)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_33),
.Y(n_65)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_65),
.Y(n_136)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_24),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_66),
.Y(n_134)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_67),
.Y(n_164)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_22),
.Y(n_68)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_68),
.Y(n_141)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_60),
.Y(n_69)
);

BUFx5_ASAP7_75t_L g161 ( 
.A(n_69),
.Y(n_161)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_22),
.Y(n_70)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_70),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_61),
.B(n_10),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_19),
.B(n_32),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_72),
.B(n_95),
.Y(n_157)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_40),
.Y(n_73)
);

INVx5_ASAP7_75t_L g204 ( 
.A(n_73),
.Y(n_204)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_37),
.Y(n_74)
);

INVx5_ASAP7_75t_L g181 ( 
.A(n_74),
.Y(n_181)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_35),
.Y(n_75)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_75),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_31),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_76),
.Y(n_137)
);

INVx2_ASAP7_75t_SL g77 ( 
.A(n_42),
.Y(n_77)
);

INVx4_ASAP7_75t_SL g205 ( 
.A(n_77),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_31),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_78),
.Y(n_158)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_20),
.Y(n_79)
);

INVx5_ASAP7_75t_L g182 ( 
.A(n_79),
.Y(n_182)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_35),
.Y(n_80)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_80),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_31),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_81),
.Y(n_159)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_24),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_82),
.Y(n_176)
);

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_37),
.Y(n_83)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_83),
.Y(n_144)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_33),
.Y(n_84)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_84),
.Y(n_184)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_33),
.Y(n_85)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_85),
.Y(n_190)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_40),
.Y(n_86)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_86),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_24),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_87),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_26),
.Y(n_88)
);

INVx6_ASAP7_75t_L g173 ( 
.A(n_88),
.Y(n_173)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_47),
.Y(n_89)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_89),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_26),
.Y(n_90)
);

INVx6_ASAP7_75t_L g189 ( 
.A(n_90),
.Y(n_189)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_26),
.Y(n_91)
);

INVx6_ASAP7_75t_L g198 ( 
.A(n_91),
.Y(n_198)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_35),
.Y(n_92)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_92),
.Y(n_149)
);

NOR2xp67_ASAP7_75t_L g93 ( 
.A(n_25),
.B(n_10),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_93),
.B(n_116),
.Y(n_135)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_34),
.Y(n_94)
);

INVx8_ASAP7_75t_L g148 ( 
.A(n_94),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_19),
.B(n_7),
.Y(n_95)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_20),
.Y(n_96)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_96),
.Y(n_145)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_34),
.Y(n_97)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_97),
.Y(n_152)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_47),
.Y(n_98)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_98),
.Y(n_160)
);

INVx2_ASAP7_75t_SL g99 ( 
.A(n_42),
.Y(n_99)
);

BUFx12f_ASAP7_75t_SL g175 ( 
.A(n_99),
.Y(n_175)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_39),
.Y(n_100)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_100),
.Y(n_192)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_25),
.Y(n_101)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_101),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_34),
.Y(n_102)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_102),
.Y(n_162)
);

BUFx12f_ASAP7_75t_L g103 ( 
.A(n_37),
.Y(n_103)
);

INVx2_ASAP7_75t_SL g140 ( 
.A(n_103),
.Y(n_140)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_33),
.Y(n_104)
);

INVx2_ASAP7_75t_SL g165 ( 
.A(n_104),
.Y(n_165)
);

BUFx12f_ASAP7_75t_L g105 ( 
.A(n_37),
.Y(n_105)
);

INVx2_ASAP7_75t_SL g212 ( 
.A(n_105),
.Y(n_212)
);

INVx11_ASAP7_75t_L g106 ( 
.A(n_45),
.Y(n_106)
);

BUFx10_ASAP7_75t_L g191 ( 
.A(n_106),
.Y(n_191)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_46),
.Y(n_107)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_107),
.Y(n_163)
);

CKINVDCx9p33_ASAP7_75t_R g108 ( 
.A(n_51),
.Y(n_108)
);

INVx5_ASAP7_75t_SL g156 ( 
.A(n_108),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_50),
.Y(n_109)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_109),
.Y(n_168)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_47),
.Y(n_110)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_110),
.Y(n_183)
);

BUFx5_ASAP7_75t_L g111 ( 
.A(n_39),
.Y(n_111)
);

CKINVDCx6p67_ASAP7_75t_R g131 ( 
.A(n_111),
.Y(n_131)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_46),
.Y(n_112)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_112),
.Y(n_185)
);

INVx8_ASAP7_75t_L g113 ( 
.A(n_44),
.Y(n_113)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_113),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_32),
.B(n_11),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g195 ( 
.A(n_114),
.B(n_119),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_50),
.Y(n_115)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_115),
.Y(n_193)
);

BUFx12f_ASAP7_75t_SL g116 ( 
.A(n_49),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_50),
.Y(n_117)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_117),
.Y(n_209)
);

INVx2_ASAP7_75t_SL g118 ( 
.A(n_42),
.Y(n_118)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_118),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_41),
.B(n_11),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g120 ( 
.A(n_44),
.Y(n_120)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_120),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_27),
.Y(n_121)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_121),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_27),
.Y(n_122)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_122),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_27),
.Y(n_123)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_123),
.Y(n_206)
);

BUFx3_ASAP7_75t_L g124 ( 
.A(n_36),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_124),
.B(n_125),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_41),
.B(n_17),
.Y(n_125)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_36),
.Y(n_126)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_126),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_30),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_127),
.B(n_128),
.Y(n_143)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_52),
.Y(n_128)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_36),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_129),
.B(n_47),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_L g132 ( 
.A1(n_66),
.A2(n_30),
.B1(n_55),
.B2(n_52),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_132),
.A2(n_150),
.B1(n_167),
.B2(n_177),
.Y(n_219)
);

OAI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_87),
.A2(n_51),
.B1(n_54),
.B2(n_45),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_139),
.A2(n_172),
.B1(n_174),
.B2(n_6),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_146),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_74),
.A2(n_49),
.B1(n_51),
.B2(n_42),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_63),
.B(n_56),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_151),
.B(n_178),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_72),
.B(n_56),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_154),
.B(n_155),
.Y(n_222)
);

AOI21xp33_ASAP7_75t_L g155 ( 
.A1(n_71),
.A2(n_38),
.B(n_53),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_95),
.B(n_57),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_166),
.B(n_169),
.Y(n_244)
);

AO22x1_ASAP7_75t_SL g167 ( 
.A1(n_82),
.A2(n_51),
.B1(n_54),
.B2(n_43),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_114),
.B(n_57),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_119),
.B(n_29),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_171),
.B(n_180),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_125),
.A2(n_55),
.B1(n_30),
.B2(n_38),
.Y(n_172)
);

OAI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_88),
.A2(n_90),
.B1(n_102),
.B2(n_109),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_83),
.A2(n_51),
.B1(n_55),
.B2(n_54),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_77),
.B(n_53),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_103),
.B(n_29),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_99),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_188),
.B(n_210),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_118),
.B(n_23),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_196),
.B(n_0),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_105),
.A2(n_48),
.B1(n_43),
.B2(n_59),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_200),
.A2(n_203),
.B1(n_113),
.B2(n_48),
.Y(n_217)
);

AND2x2_ASAP7_75t_SL g201 ( 
.A(n_79),
.B(n_48),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g223 ( 
.A(n_201),
.B(n_123),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_62),
.A2(n_48),
.B1(n_43),
.B2(n_59),
.Y(n_203)
);

OR2x2_ASAP7_75t_L g210 ( 
.A(n_96),
.B(n_28),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_L g213 ( 
.A1(n_91),
.A2(n_94),
.B1(n_97),
.B2(n_81),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_213),
.A2(n_58),
.B1(n_1),
.B2(n_2),
.Y(n_235)
);

AO22x2_ASAP7_75t_L g214 ( 
.A1(n_167),
.A2(n_76),
.B1(n_78),
.B2(n_115),
.Y(n_214)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_214),
.Y(n_290)
);

INVx6_ASAP7_75t_L g215 ( 
.A(n_202),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g307 ( 
.A(n_215),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_217),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_156),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_218),
.B(n_220),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_156),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_192),
.A2(n_23),
.B1(n_28),
.B2(n_117),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_221),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g340 ( 
.A(n_223),
.Y(n_340)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_152),
.Y(n_224)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_224),
.Y(n_295)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_130),
.Y(n_225)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_225),
.Y(n_299)
);

AOI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_192),
.A2(n_127),
.B1(n_122),
.B2(n_121),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g350 ( 
.A(n_226),
.Y(n_350)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_133),
.Y(n_227)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_227),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_229),
.B(n_265),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_195),
.A2(n_21),
.B1(n_58),
.B2(n_12),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g314 ( 
.A1(n_230),
.A2(n_237),
.B(n_257),
.Y(n_314)
);

A2O1A1Ixp33_ASAP7_75t_L g231 ( 
.A1(n_195),
.A2(n_21),
.B(n_13),
.C(n_18),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g310 ( 
.A(n_231),
.B(n_161),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_141),
.B(n_21),
.C(n_58),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_232),
.B(n_280),
.C(n_287),
.Y(n_309)
);

INVx1_ASAP7_75t_SL g233 ( 
.A(n_179),
.Y(n_233)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_233),
.Y(n_304)
);

AOI22xp33_ASAP7_75t_L g234 ( 
.A1(n_174),
.A2(n_58),
.B1(n_18),
.B2(n_17),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_234),
.A2(n_254),
.B1(n_263),
.B2(n_278),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_235),
.A2(n_236),
.B1(n_255),
.B2(n_258),
.Y(n_296)
);

OAI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_210),
.A2(n_18),
.B1(n_17),
.B2(n_15),
.Y(n_236)
);

O2A1O1Ixp33_ASAP7_75t_L g237 ( 
.A1(n_201),
.A2(n_0),
.B(n_1),
.C(n_2),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_147),
.Y(n_238)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_238),
.Y(n_306)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_149),
.Y(n_239)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_239),
.Y(n_317)
);

HAxp5_ASAP7_75t_SL g240 ( 
.A(n_157),
.B(n_18),
.CON(n_240),
.SN(n_240)
);

BUFx8_ASAP7_75t_L g347 ( 
.A(n_240),
.Y(n_347)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_162),
.Y(n_241)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_241),
.Y(n_312)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_142),
.Y(n_242)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_242),
.Y(n_321)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_168),
.Y(n_243)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_243),
.Y(n_332)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_150),
.Y(n_245)
);

HB1xp67_ASAP7_75t_L g311 ( 
.A(n_245),
.Y(n_311)
);

INVx2_ASAP7_75t_SL g247 ( 
.A(n_186),
.Y(n_247)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_247),
.Y(n_335)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_170),
.Y(n_248)
);

INVx2_ASAP7_75t_SL g348 ( 
.A(n_248),
.Y(n_348)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_199),
.Y(n_249)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_249),
.Y(n_334)
);

INVx6_ASAP7_75t_L g250 ( 
.A(n_202),
.Y(n_250)
);

INVx4_ASAP7_75t_L g315 ( 
.A(n_250),
.Y(n_315)
);

AOI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_211),
.A2(n_14),
.B1(n_13),
.B2(n_2),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_SL g300 ( 
.A1(n_251),
.A2(n_277),
.B1(n_181),
.B2(n_144),
.Y(n_300)
);

INVx11_ASAP7_75t_L g253 ( 
.A(n_191),
.Y(n_253)
);

INVx11_ASAP7_75t_L g302 ( 
.A(n_253),
.Y(n_302)
);

AOI22xp33_ASAP7_75t_L g254 ( 
.A1(n_132),
.A2(n_14),
.B1(n_1),
.B2(n_2),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_213),
.A2(n_143),
.B1(n_138),
.B2(n_135),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_193),
.Y(n_256)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_256),
.Y(n_336)
);

NAND2x1_ASAP7_75t_SL g257 ( 
.A(n_175),
.B(n_205),
.Y(n_257)
);

OAI22xp33_ASAP7_75t_SL g258 ( 
.A1(n_177),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_258)
);

CKINVDCx14_ASAP7_75t_R g259 ( 
.A(n_205),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_259),
.B(n_285),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_197),
.B(n_3),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_260),
.B(n_284),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_203),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_261),
.A2(n_269),
.B1(n_273),
.B2(n_275),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_157),
.B(n_207),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_SL g331 ( 
.A(n_262),
.B(n_274),
.Y(n_331)
);

INVx11_ASAP7_75t_L g264 ( 
.A(n_191),
.Y(n_264)
);

BUFx2_ASAP7_75t_L g303 ( 
.A(n_264),
.Y(n_303)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_206),
.Y(n_265)
);

INVx5_ASAP7_75t_L g266 ( 
.A(n_181),
.Y(n_266)
);

INVx3_ASAP7_75t_L g291 ( 
.A(n_266),
.Y(n_291)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_163),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_267),
.B(n_271),
.Y(n_343)
);

INVx6_ASAP7_75t_L g268 ( 
.A(n_137),
.Y(n_268)
);

INVx4_ASAP7_75t_L g326 ( 
.A(n_268),
.Y(n_326)
);

OAI22xp33_ASAP7_75t_L g269 ( 
.A1(n_200),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_209),
.Y(n_270)
);

INVx3_ASAP7_75t_L g337 ( 
.A(n_270),
.Y(n_337)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_185),
.Y(n_271)
);

INVx3_ASAP7_75t_L g272 ( 
.A(n_204),
.Y(n_272)
);

INVx4_ASAP7_75t_L g346 ( 
.A(n_272),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_198),
.A2(n_173),
.B1(n_189),
.B2(n_134),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_165),
.B(n_5),
.Y(n_274)
);

OAI22xp33_ASAP7_75t_SL g275 ( 
.A1(n_139),
.A2(n_176),
.B1(n_134),
.B2(n_158),
.Y(n_275)
);

INVx1_ASAP7_75t_SL g276 ( 
.A(n_208),
.Y(n_276)
);

CKINVDCx16_ASAP7_75t_R g328 ( 
.A(n_276),
.Y(n_328)
);

AOI22xp33_ASAP7_75t_SL g277 ( 
.A1(n_145),
.A2(n_187),
.B1(n_182),
.B2(n_153),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_198),
.A2(n_173),
.B1(n_189),
.B2(n_176),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g279 ( 
.A(n_137),
.Y(n_279)
);

INVx8_ASAP7_75t_L g298 ( 
.A(n_279),
.Y(n_298)
);

AND2x2_ASAP7_75t_L g280 ( 
.A(n_164),
.B(n_194),
.Y(n_280)
);

BUFx2_ASAP7_75t_SL g281 ( 
.A(n_131),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_281),
.Y(n_308)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_160),
.Y(n_282)
);

INVx3_ASAP7_75t_L g342 ( 
.A(n_282),
.Y(n_342)
);

OAI22xp33_ASAP7_75t_SL g283 ( 
.A1(n_158),
.A2(n_159),
.B1(n_145),
.B2(n_184),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_283),
.A2(n_140),
.B1(n_212),
.B2(n_153),
.Y(n_320)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_183),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_160),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_165),
.B(n_136),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_SL g333 ( 
.A(n_286),
.B(n_220),
.Y(n_333)
);

AND2x2_ASAP7_75t_L g287 ( 
.A(n_190),
.B(n_144),
.Y(n_287)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_148),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_288),
.B(n_131),
.Y(n_327)
);

HB1xp67_ASAP7_75t_L g289 ( 
.A(n_140),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_289),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_229),
.B(n_148),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_293),
.B(n_294),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_260),
.B(n_216),
.Y(n_294)
);

INVxp67_ASAP7_75t_L g393 ( 
.A(n_300),
.Y(n_393)
);

OR2x2_ASAP7_75t_L g366 ( 
.A(n_310),
.B(n_349),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_216),
.B(n_159),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_313),
.B(n_330),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_320),
.A2(n_323),
.B1(n_325),
.B2(n_329),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_L g323 ( 
.A1(n_263),
.A2(n_245),
.B1(n_228),
.B2(n_222),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_257),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_324),
.B(n_287),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_L g325 ( 
.A1(n_228),
.A2(n_182),
.B1(n_191),
.B2(n_212),
.Y(n_325)
);

INVxp67_ASAP7_75t_L g396 ( 
.A(n_327),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_L g329 ( 
.A1(n_214),
.A2(n_131),
.B1(n_230),
.B2(n_252),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_231),
.B(n_242),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_333),
.B(n_344),
.Y(n_351)
);

MAJx2_ASAP7_75t_L g338 ( 
.A(n_246),
.B(n_244),
.C(n_255),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_338),
.B(n_271),
.C(n_239),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_248),
.B(n_233),
.Y(n_344)
);

OAI21xp5_ASAP7_75t_L g345 ( 
.A1(n_257),
.A2(n_237),
.B(n_223),
.Y(n_345)
);

A2O1A1O1Ixp25_ASAP7_75t_L g354 ( 
.A1(n_345),
.A2(n_314),
.B(n_330),
.C(n_340),
.D(n_309),
.Y(n_354)
);

AOI22xp33_ASAP7_75t_SL g349 ( 
.A1(n_219),
.A2(n_235),
.B1(n_265),
.B2(n_249),
.Y(n_349)
);

AND2x2_ASAP7_75t_L g352 ( 
.A(n_324),
.B(n_223),
.Y(n_352)
);

CKINVDCx14_ASAP7_75t_R g434 ( 
.A(n_352),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_297),
.A2(n_261),
.B1(n_232),
.B2(n_240),
.Y(n_353)
);

OAI21xp5_ASAP7_75t_L g410 ( 
.A1(n_353),
.A2(n_354),
.B(n_361),
.Y(n_410)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_321),
.Y(n_355)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_355),
.Y(n_403)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_334),
.Y(n_357)
);

HB1xp67_ASAP7_75t_L g401 ( 
.A(n_357),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_319),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_358),
.B(n_368),
.Y(n_408)
);

HB1xp67_ASAP7_75t_L g359 ( 
.A(n_346),
.Y(n_359)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_359),
.Y(n_407)
);

AOI21xp5_ASAP7_75t_L g360 ( 
.A1(n_311),
.A2(n_269),
.B(n_218),
.Y(n_360)
);

AOI21xp5_ASAP7_75t_L g422 ( 
.A1(n_360),
.A2(n_379),
.B(n_350),
.Y(n_422)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_321),
.Y(n_362)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_362),
.Y(n_409)
);

AND2x2_ASAP7_75t_L g363 ( 
.A(n_345),
.B(n_280),
.Y(n_363)
);

CKINVDCx16_ASAP7_75t_R g425 ( 
.A(n_363),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_290),
.A2(n_214),
.B1(n_247),
.B2(n_267),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_364),
.A2(n_377),
.B1(n_385),
.B2(n_390),
.Y(n_427)
);

INVx1_ASAP7_75t_SL g365 ( 
.A(n_304),
.Y(n_365)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_365),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_331),
.B(n_276),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_334),
.Y(n_369)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_369),
.Y(n_414)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_348),
.Y(n_370)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_370),
.Y(n_420)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_348),
.Y(n_372)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_372),
.Y(n_428)
);

MAJx3_ASAP7_75t_L g373 ( 
.A(n_314),
.B(n_280),
.C(n_287),
.Y(n_373)
);

OAI21xp5_ASAP7_75t_L g415 ( 
.A1(n_373),
.A2(n_375),
.B(n_395),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_294),
.B(n_214),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_374),
.B(n_383),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_297),
.A2(n_288),
.B1(n_214),
.B2(n_278),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g418 ( 
.A(n_376),
.B(n_398),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_L g377 ( 
.A1(n_290),
.A2(n_215),
.B1(n_268),
.B2(n_250),
.Y(n_377)
);

BUFx6f_ASAP7_75t_L g378 ( 
.A(n_298),
.Y(n_378)
);

BUFx6f_ASAP7_75t_L g406 ( 
.A(n_378),
.Y(n_406)
);

AOI21xp5_ASAP7_75t_L g379 ( 
.A1(n_305),
.A2(n_266),
.B(n_285),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_348),
.Y(n_380)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_380),
.Y(n_429)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_335),
.Y(n_381)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_381),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_SL g382 ( 
.A(n_339),
.B(n_225),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_SL g405 ( 
.A(n_382),
.B(n_389),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_292),
.B(n_227),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_292),
.B(n_238),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_384),
.B(n_391),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_L g385 ( 
.A1(n_341),
.A2(n_247),
.B1(n_279),
.B2(n_273),
.Y(n_385)
);

INVx3_ASAP7_75t_L g386 ( 
.A(n_346),
.Y(n_386)
);

AOI22xp33_ASAP7_75t_SL g404 ( 
.A1(n_386),
.A2(n_388),
.B1(n_308),
.B2(n_303),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_318),
.A2(n_241),
.B1(n_243),
.B2(n_270),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_SL g435 ( 
.A1(n_387),
.A2(n_392),
.B1(n_317),
.B2(n_304),
.Y(n_435)
);

INVx3_ASAP7_75t_L g388 ( 
.A(n_315),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_335),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_341),
.A2(n_224),
.B1(n_256),
.B2(n_279),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_299),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_L g392 ( 
.A1(n_340),
.A2(n_284),
.B1(n_272),
.B2(n_282),
.Y(n_392)
);

CKINVDCx16_ASAP7_75t_R g394 ( 
.A(n_322),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_394),
.B(n_397),
.Y(n_438)
);

OAI21xp33_ASAP7_75t_SL g395 ( 
.A1(n_305),
.A2(n_253),
.B(n_264),
.Y(n_395)
);

OR2x2_ASAP7_75t_L g397 ( 
.A(n_310),
.B(n_347),
.Y(n_397)
);

AND2x2_ASAP7_75t_L g398 ( 
.A(n_309),
.B(n_343),
.Y(n_398)
);

XOR2xp5_ASAP7_75t_L g399 ( 
.A(n_398),
.B(n_313),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_399),
.B(n_402),
.C(n_411),
.Y(n_469)
);

AOI32xp33_ASAP7_75t_L g400 ( 
.A1(n_366),
.A2(n_354),
.A3(n_371),
.B1(n_358),
.B2(n_393),
.Y(n_400)
);

OAI21xp5_ASAP7_75t_SL g445 ( 
.A1(n_400),
.A2(n_422),
.B(n_397),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_398),
.B(n_356),
.C(n_376),
.Y(n_402)
);

BUFx3_ASAP7_75t_L g470 ( 
.A(n_404),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_356),
.B(n_338),
.C(n_293),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_352),
.B(n_301),
.C(n_306),
.Y(n_417)
);

XOR2xp5_ASAP7_75t_L g451 ( 
.A(n_417),
.B(n_423),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_371),
.B(n_299),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_419),
.B(n_436),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_351),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_421),
.B(n_431),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_352),
.B(n_306),
.C(n_301),
.Y(n_423)
);

AOI22xp33_ASAP7_75t_SL g424 ( 
.A1(n_393),
.A2(n_350),
.B1(n_308),
.B2(n_303),
.Y(n_424)
);

CKINVDCx16_ASAP7_75t_R g453 ( 
.A(n_424),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_383),
.B(n_317),
.C(n_316),
.Y(n_426)
);

XOR2xp5_ASAP7_75t_L g463 ( 
.A(n_426),
.B(n_430),
.Y(n_463)
);

XOR2xp5_ASAP7_75t_L g430 ( 
.A(n_384),
.B(n_296),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_392),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_L g433 ( 
.A1(n_385),
.A2(n_364),
.B1(n_374),
.B2(n_390),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_SL g446 ( 
.A1(n_433),
.A2(n_353),
.B1(n_360),
.B2(n_396),
.Y(n_446)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_435),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_391),
.B(n_296),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_355),
.B(n_316),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_437),
.B(n_380),
.Y(n_457)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_436),
.A2(n_366),
.B1(n_363),
.B2(n_367),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_L g502 ( 
.A1(n_440),
.A2(n_448),
.B1(n_473),
.B2(n_428),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_SL g443 ( 
.A(n_405),
.B(n_419),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_443),
.B(n_447),
.Y(n_482)
);

OAI22xp5_ASAP7_75t_L g444 ( 
.A1(n_433),
.A2(n_375),
.B1(n_367),
.B2(n_387),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_L g481 ( 
.A1(n_444),
.A2(n_446),
.B1(n_475),
.B2(n_434),
.Y(n_481)
);

A2O1A1Ixp33_ASAP7_75t_L g479 ( 
.A1(n_445),
.A2(n_400),
.B(n_410),
.C(n_415),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_401),
.Y(n_447)
);

AOI22xp5_ASAP7_75t_L g448 ( 
.A1(n_430),
.A2(n_363),
.B1(n_396),
.B2(n_362),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_437),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_449),
.B(n_455),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_421),
.B(n_291),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_SL g480 ( 
.A(n_450),
.B(n_456),
.Y(n_480)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_432),
.Y(n_452)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_452),
.Y(n_476)
);

FAx1_ASAP7_75t_SL g454 ( 
.A(n_413),
.B(n_411),
.CI(n_410),
.CON(n_454),
.SN(n_454)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_454),
.B(n_464),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_408),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_438),
.B(n_291),
.Y(n_456)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_457),
.Y(n_488)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_432),
.Y(n_458)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_458),
.Y(n_494)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_403),
.Y(n_459)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_459),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_405),
.B(n_389),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_460),
.B(n_462),
.Y(n_495)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_403),
.Y(n_461)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_461),
.Y(n_509)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_409),
.Y(n_462)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_414),
.Y(n_464)
);

XOR2xp5_ASAP7_75t_L g465 ( 
.A(n_418),
.B(n_373),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_465),
.B(n_468),
.C(n_402),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_SL g466 ( 
.A(n_416),
.B(n_372),
.Y(n_466)
);

XNOR2xp5_ASAP7_75t_SL g487 ( 
.A(n_466),
.B(n_441),
.Y(n_487)
);

AND2x2_ASAP7_75t_L g467 ( 
.A(n_415),
.B(n_379),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g486 ( 
.A(n_467),
.Y(n_486)
);

XOR2xp5_ASAP7_75t_L g468 ( 
.A(n_418),
.B(n_373),
.Y(n_468)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_409),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_471),
.B(n_472),
.Y(n_498)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_420),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_420),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_416),
.B(n_381),
.Y(n_474)
);

CKINVDCx20_ASAP7_75t_R g497 ( 
.A(n_474),
.Y(n_497)
);

OAI22xp5_ASAP7_75t_SL g475 ( 
.A1(n_413),
.A2(n_365),
.B1(n_370),
.B2(n_369),
.Y(n_475)
);

XNOR2x1_ASAP7_75t_L g520 ( 
.A(n_477),
.B(n_478),
.Y(n_520)
);

XNOR2x1_ASAP7_75t_L g478 ( 
.A(n_465),
.B(n_399),
.Y(n_478)
);

AOI21xp5_ASAP7_75t_L g514 ( 
.A1(n_479),
.A2(n_467),
.B(n_460),
.Y(n_514)
);

OAI22xp5_ASAP7_75t_SL g510 ( 
.A1(n_481),
.A2(n_491),
.B1(n_496),
.B2(n_507),
.Y(n_510)
);

XNOR2xp5_ASAP7_75t_L g484 ( 
.A(n_451),
.B(n_426),
.Y(n_484)
);

XOR2xp5_ASAP7_75t_L g517 ( 
.A(n_484),
.B(n_485),
.Y(n_517)
);

XOR2xp5_ASAP7_75t_L g485 ( 
.A(n_463),
.B(n_451),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_487),
.B(n_504),
.Y(n_536)
);

OAI22xp5_ASAP7_75t_SL g489 ( 
.A1(n_439),
.A2(n_422),
.B1(n_427),
.B2(n_431),
.Y(n_489)
);

AOI22xp5_ASAP7_75t_L g518 ( 
.A1(n_489),
.A2(n_501),
.B1(n_502),
.B2(n_473),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_469),
.B(n_463),
.C(n_468),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_490),
.B(n_500),
.C(n_503),
.Y(n_526)
);

AOI22xp5_ASAP7_75t_L g491 ( 
.A1(n_439),
.A2(n_435),
.B1(n_425),
.B2(n_427),
.Y(n_491)
);

XOR2xp5_ASAP7_75t_L g493 ( 
.A(n_469),
.B(n_417),
.Y(n_493)
);

XOR2xp5_ASAP7_75t_L g531 ( 
.A(n_493),
.B(n_347),
.Y(n_531)
);

AOI22xp5_ASAP7_75t_L g496 ( 
.A1(n_444),
.A2(n_425),
.B1(n_423),
.B2(n_429),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_448),
.B(n_412),
.C(n_429),
.Y(n_500)
);

OAI22xp5_ASAP7_75t_SL g501 ( 
.A1(n_440),
.A2(n_428),
.B1(n_412),
.B2(n_407),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_446),
.B(n_407),
.C(n_414),
.Y(n_503)
);

CKINVDCx16_ASAP7_75t_R g504 ( 
.A(n_457),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_445),
.B(n_386),
.C(n_357),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g537 ( 
.A(n_505),
.B(n_508),
.C(n_302),
.Y(n_537)
);

AOI21xp33_ASAP7_75t_L g506 ( 
.A1(n_455),
.A2(n_467),
.B(n_442),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_SL g525 ( 
.A(n_506),
.B(n_461),
.Y(n_525)
);

AOI22xp5_ASAP7_75t_L g507 ( 
.A1(n_449),
.A2(n_406),
.B1(n_378),
.B2(n_388),
.Y(n_507)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_474),
.B(n_342),
.C(n_295),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_497),
.B(n_466),
.Y(n_511)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_511),
.Y(n_547)
);

XNOR2xp5_ASAP7_75t_L g512 ( 
.A(n_493),
.B(n_442),
.Y(n_512)
);

MAJx2_ASAP7_75t_L g551 ( 
.A(n_512),
.B(n_516),
.C(n_522),
.Y(n_551)
);

OAI22xp5_ASAP7_75t_SL g513 ( 
.A1(n_481),
.A2(n_441),
.B1(n_453),
.B2(n_443),
.Y(n_513)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_513),
.Y(n_543)
);

OAI21xp5_ASAP7_75t_SL g545 ( 
.A1(n_514),
.A2(n_503),
.B(n_505),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_492),
.B(n_475),
.Y(n_515)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_515),
.Y(n_557)
);

XNOR2xp5_ASAP7_75t_L g516 ( 
.A(n_484),
.B(n_454),
.Y(n_516)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_518),
.Y(n_563)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_492),
.Y(n_519)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_519),
.Y(n_560)
);

OAI22xp5_ASAP7_75t_SL g521 ( 
.A1(n_496),
.A2(n_453),
.B1(n_470),
.B2(n_454),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_521),
.B(n_528),
.Y(n_550)
);

XNOR2xp5_ASAP7_75t_L g522 ( 
.A(n_485),
.B(n_472),
.Y(n_522)
);

XNOR2xp5_ASAP7_75t_L g523 ( 
.A(n_490),
.B(n_471),
.Y(n_523)
);

XNOR2xp5_ASAP7_75t_L g541 ( 
.A(n_523),
.B(n_537),
.Y(n_541)
);

CKINVDCx20_ASAP7_75t_R g524 ( 
.A(n_482),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_SL g549 ( 
.A(n_524),
.B(n_527),
.Y(n_549)
);

AO21x1_ASAP7_75t_L g552 ( 
.A1(n_525),
.A2(n_534),
.B(n_507),
.Y(n_552)
);

CKINVDCx20_ASAP7_75t_R g527 ( 
.A(n_482),
.Y(n_527)
);

AOI22xp5_ASAP7_75t_L g528 ( 
.A1(n_489),
.A2(n_470),
.B1(n_462),
.B2(n_459),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_498),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g556 ( 
.A(n_529),
.B(n_532),
.Y(n_556)
);

OAI22xp5_ASAP7_75t_SL g530 ( 
.A1(n_491),
.A2(n_452),
.B1(n_458),
.B2(n_447),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_530),
.B(n_533),
.Y(n_553)
);

MAJIxp5_ASAP7_75t_L g542 ( 
.A(n_531),
.B(n_539),
.C(n_478),
.Y(n_542)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_495),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_495),
.Y(n_533)
);

AOI22xp5_ASAP7_75t_L g534 ( 
.A1(n_501),
.A2(n_464),
.B1(n_406),
.B2(n_378),
.Y(n_534)
);

INVx1_ASAP7_75t_SL g535 ( 
.A(n_509),
.Y(n_535)
);

INVx11_ASAP7_75t_L g562 ( 
.A(n_535),
.Y(n_562)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_476),
.Y(n_538)
);

CKINVDCx20_ASAP7_75t_R g544 ( 
.A(n_538),
.Y(n_544)
);

MAJIxp5_ASAP7_75t_L g539 ( 
.A(n_477),
.B(n_342),
.C(n_295),
.Y(n_539)
);

AOI21xp5_ASAP7_75t_L g540 ( 
.A1(n_514),
.A2(n_486),
.B(n_483),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_540),
.B(n_546),
.Y(n_585)
);

XOR2xp5_ASAP7_75t_L g572 ( 
.A(n_542),
.B(n_548),
.Y(n_572)
);

XNOR2xp5_ASAP7_75t_L g567 ( 
.A(n_545),
.B(n_555),
.Y(n_567)
);

MAJIxp5_ASAP7_75t_L g546 ( 
.A(n_523),
.B(n_500),
.C(n_508),
.Y(n_546)
);

XNOR2xp5_ASAP7_75t_SL g548 ( 
.A(n_516),
.B(n_520),
.Y(n_548)
);

OAI22xp5_ASAP7_75t_L g566 ( 
.A1(n_552),
.A2(n_528),
.B1(n_518),
.B2(n_534),
.Y(n_566)
);

XNOR2xp5_ASAP7_75t_SL g554 ( 
.A(n_520),
.B(n_487),
.Y(n_554)
);

XOR2xp5_ASAP7_75t_L g583 ( 
.A(n_554),
.B(n_559),
.Y(n_583)
);

XNOR2xp5_ASAP7_75t_L g555 ( 
.A(n_526),
.B(n_488),
.Y(n_555)
);

XNOR2xp5_ASAP7_75t_L g558 ( 
.A(n_526),
.B(n_522),
.Y(n_558)
);

XNOR2xp5_ASAP7_75t_L g580 ( 
.A(n_558),
.B(n_561),
.Y(n_580)
);

XOR2xp5_ASAP7_75t_L g559 ( 
.A(n_517),
.B(n_488),
.Y(n_559)
);

XNOR2xp5_ASAP7_75t_L g561 ( 
.A(n_512),
.B(n_479),
.Y(n_561)
);

MAJIxp5_ASAP7_75t_L g564 ( 
.A(n_517),
.B(n_509),
.C(n_499),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_SL g575 ( 
.A(n_564),
.B(n_530),
.Y(n_575)
);

NAND2xp33_ASAP7_75t_L g565 ( 
.A(n_547),
.B(n_511),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_565),
.B(n_568),
.Y(n_588)
);

AOI22xp5_ASAP7_75t_L g598 ( 
.A1(n_566),
.A2(n_569),
.B1(n_584),
.B2(n_563),
.Y(n_598)
);

OAI22xp5_ASAP7_75t_L g568 ( 
.A1(n_552),
.A2(n_515),
.B1(n_536),
.B2(n_480),
.Y(n_568)
);

OAI22xp5_ASAP7_75t_SL g569 ( 
.A1(n_550),
.A2(n_521),
.B1(n_510),
.B2(n_513),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_549),
.Y(n_570)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_570),
.Y(n_596)
);

MAJIxp5_ASAP7_75t_L g571 ( 
.A(n_541),
.B(n_539),
.C(n_537),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_SL g602 ( 
.A(n_571),
.B(n_575),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_556),
.B(n_535),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_573),
.B(n_578),
.Y(n_593)
);

NOR2xp33_ASAP7_75t_L g574 ( 
.A(n_564),
.B(n_555),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_SL g590 ( 
.A(n_574),
.B(n_545),
.Y(n_590)
);

MAJIxp5_ASAP7_75t_L g576 ( 
.A(n_541),
.B(n_510),
.C(n_531),
.Y(n_576)
);

MAJIxp5_ASAP7_75t_L g589 ( 
.A(n_576),
.B(n_577),
.C(n_579),
.Y(n_589)
);

MAJIxp5_ASAP7_75t_L g577 ( 
.A(n_558),
.B(n_499),
.C(n_494),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_560),
.Y(n_578)
);

MAJIxp5_ASAP7_75t_L g579 ( 
.A(n_546),
.B(n_494),
.C(n_476),
.Y(n_579)
);

MAJIxp5_ASAP7_75t_L g581 ( 
.A(n_559),
.B(n_406),
.C(n_312),
.Y(n_581)
);

MAJIxp5_ASAP7_75t_L g592 ( 
.A(n_581),
.B(n_582),
.C(n_562),
.Y(n_592)
);

MAJIxp5_ASAP7_75t_L g582 ( 
.A(n_542),
.B(n_332),
.C(n_336),
.Y(n_582)
);

OAI22xp5_ASAP7_75t_SL g584 ( 
.A1(n_550),
.A2(n_307),
.B1(n_298),
.B2(n_326),
.Y(n_584)
);

AOI21xp5_ASAP7_75t_L g586 ( 
.A1(n_573),
.A2(n_540),
.B(n_553),
.Y(n_586)
);

OAI21xp5_ASAP7_75t_SL g607 ( 
.A1(n_586),
.A2(n_580),
.B(n_572),
.Y(n_607)
);

NOR2x1_ASAP7_75t_SL g587 ( 
.A(n_569),
.B(n_561),
.Y(n_587)
);

OR2x2_ASAP7_75t_L g613 ( 
.A(n_587),
.B(n_595),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_SL g609 ( 
.A(n_590),
.B(n_328),
.Y(n_609)
);

HB1xp67_ASAP7_75t_L g591 ( 
.A(n_577),
.Y(n_591)
);

AOI22xp33_ASAP7_75t_L g608 ( 
.A1(n_591),
.A2(n_580),
.B1(n_326),
.B2(n_315),
.Y(n_608)
);

HB1xp67_ASAP7_75t_L g615 ( 
.A(n_592),
.Y(n_615)
);

XNOR2xp5_ASAP7_75t_L g594 ( 
.A(n_579),
.B(n_551),
.Y(n_594)
);

NOR2xp67_ASAP7_75t_SL g606 ( 
.A(n_594),
.B(n_599),
.Y(n_606)
);

OAI21xp5_ASAP7_75t_L g595 ( 
.A1(n_585),
.A2(n_543),
.B(n_557),
.Y(n_595)
);

OAI21xp5_ASAP7_75t_L g597 ( 
.A1(n_576),
.A2(n_543),
.B(n_553),
.Y(n_597)
);

AOI22xp5_ASAP7_75t_L g603 ( 
.A1(n_597),
.A2(n_601),
.B1(n_584),
.B2(n_583),
.Y(n_603)
);

XOR2xp5_ASAP7_75t_L g616 ( 
.A(n_598),
.B(n_595),
.Y(n_616)
);

MAJIxp5_ASAP7_75t_L g599 ( 
.A(n_571),
.B(n_563),
.C(n_551),
.Y(n_599)
);

MAJIxp5_ASAP7_75t_L g600 ( 
.A(n_567),
.B(n_548),
.C(n_554),
.Y(n_600)
);

MAJIxp5_ASAP7_75t_L g610 ( 
.A(n_600),
.B(n_337),
.C(n_312),
.Y(n_610)
);

OAI22xp5_ASAP7_75t_SL g601 ( 
.A1(n_581),
.A2(n_544),
.B1(n_562),
.B2(n_307),
.Y(n_601)
);

INVxp67_ASAP7_75t_L g621 ( 
.A(n_603),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_L g604 ( 
.A(n_602),
.B(n_567),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_SL g622 ( 
.A(n_604),
.B(n_611),
.Y(n_622)
);

AOI22xp5_ASAP7_75t_L g605 ( 
.A1(n_588),
.A2(n_583),
.B1(n_572),
.B2(n_582),
.Y(n_605)
);

XOR2xp5_ASAP7_75t_L g626 ( 
.A(n_605),
.B(n_608),
.Y(n_626)
);

AOI21xp5_ASAP7_75t_L g617 ( 
.A1(n_607),
.A2(n_609),
.B(n_612),
.Y(n_617)
);

XNOR2xp5_ASAP7_75t_L g619 ( 
.A(n_610),
.B(n_594),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_L g611 ( 
.A(n_589),
.B(n_332),
.Y(n_611)
);

MAJIxp5_ASAP7_75t_L g612 ( 
.A(n_589),
.B(n_302),
.C(n_336),
.Y(n_612)
);

MAJIxp5_ASAP7_75t_L g614 ( 
.A(n_599),
.B(n_337),
.C(n_347),
.Y(n_614)
);

AOI21xp5_ASAP7_75t_L g618 ( 
.A1(n_614),
.A2(n_592),
.B(n_600),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_L g624 ( 
.A(n_616),
.B(n_598),
.Y(n_624)
);

OAI21x1_ASAP7_75t_L g632 ( 
.A1(n_618),
.A2(n_624),
.B(n_613),
.Y(n_632)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_619),
.Y(n_630)
);

AOI21xp5_ASAP7_75t_L g620 ( 
.A1(n_606),
.A2(n_597),
.B(n_586),
.Y(n_620)
);

AOI21xp5_ASAP7_75t_L g633 ( 
.A1(n_620),
.A2(n_623),
.B(n_603),
.Y(n_633)
);

OAI21xp5_ASAP7_75t_SL g623 ( 
.A1(n_613),
.A2(n_587),
.B(n_596),
.Y(n_623)
);

XNOR2xp5_ASAP7_75t_L g625 ( 
.A(n_610),
.B(n_601),
.Y(n_625)
);

AND2x2_ASAP7_75t_L g629 ( 
.A(n_625),
.B(n_612),
.Y(n_629)
);

INVxp67_ASAP7_75t_L g627 ( 
.A(n_622),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_627),
.B(n_628),
.Y(n_634)
);

MAJIxp5_ASAP7_75t_L g628 ( 
.A(n_621),
.B(n_615),
.C(n_616),
.Y(n_628)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_629),
.Y(n_635)
);

NOR2xp33_ASAP7_75t_L g631 ( 
.A(n_621),
.B(n_593),
.Y(n_631)
);

AOI21xp5_ASAP7_75t_SL g636 ( 
.A1(n_631),
.A2(n_632),
.B(n_633),
.Y(n_636)
);

INVxp67_ASAP7_75t_L g637 ( 
.A(n_631),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_SL g639 ( 
.A(n_637),
.B(n_626),
.Y(n_639)
);

AO21x1_ASAP7_75t_L g638 ( 
.A1(n_635),
.A2(n_630),
.B(n_593),
.Y(n_638)
);

OAI21xp5_ASAP7_75t_SL g640 ( 
.A1(n_638),
.A2(n_639),
.B(n_636),
.Y(n_640)
);

AOI21x1_ASAP7_75t_L g641 ( 
.A1(n_640),
.A2(n_634),
.B(n_617),
.Y(n_641)
);

XOR2xp5_ASAP7_75t_L g642 ( 
.A(n_641),
.B(n_626),
.Y(n_642)
);

AOI21xp5_ASAP7_75t_L g643 ( 
.A1(n_642),
.A2(n_605),
.B(n_614),
.Y(n_643)
);


endmodule