module fake_jpeg_22371_n_58 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_58);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_58;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_43;
wire n_37;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

INVx2_ASAP7_75t_L g8 ( 
.A(n_3),
.Y(n_8)
);

INVx13_ASAP7_75t_L g9 ( 
.A(n_3),
.Y(n_9)
);

BUFx12_ASAP7_75t_L g10 ( 
.A(n_4),
.Y(n_10)
);

BUFx12f_ASAP7_75t_L g11 ( 
.A(n_3),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

BUFx3_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

HB1xp67_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_12),
.B(n_0),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_17),
.B(n_15),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

AND2x2_ASAP7_75t_SL g24 ( 
.A(n_18),
.B(n_19),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

BUFx24_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

OR2x4_ASAP7_75t_L g21 ( 
.A(n_20),
.B(n_14),
.Y(n_21)
);

OAI22xp33_ASAP7_75t_SL g28 ( 
.A1(n_21),
.A2(n_25),
.B1(n_9),
.B2(n_20),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_22),
.B(n_7),
.Y(n_26)
);

OA22x2_ASAP7_75t_L g25 ( 
.A1(n_20),
.A2(n_9),
.B1(n_13),
.B2(n_8),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_26),
.B(n_27),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g27 ( 
.A1(n_25),
.A2(n_8),
.B1(n_13),
.B2(n_18),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_28),
.A2(n_10),
.B1(n_1),
.B2(n_2),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_24),
.B(n_19),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_29),
.B(n_30),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_24),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_23),
.B(n_10),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_31),
.B(n_32),
.Y(n_38)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

CKINVDCx12_ASAP7_75t_R g34 ( 
.A(n_33),
.Y(n_34)
);

AOI21xp5_ASAP7_75t_L g35 ( 
.A1(n_30),
.A2(n_16),
.B(n_18),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_35),
.B(n_39),
.Y(n_41)
);

AND2x6_ASAP7_75t_L g39 ( 
.A(n_29),
.B(n_18),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_40),
.A2(n_27),
.B1(n_32),
.B2(n_26),
.Y(n_43)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_38),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_42),
.A2(n_44),
.B1(n_45),
.B2(n_36),
.Y(n_46)
);

OAI21xp5_ASAP7_75t_L g48 ( 
.A1(n_43),
.A2(n_32),
.B(n_10),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_34),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

OAI21xp5_ASAP7_75t_L g50 ( 
.A1(n_46),
.A2(n_47),
.B(n_48),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_45),
.A2(n_39),
.B1(n_40),
.B2(n_31),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_47),
.B(n_41),
.C(n_42),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_49),
.B(n_43),
.Y(n_52)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_50),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_51),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_SL g54 ( 
.A1(n_52),
.A2(n_51),
.B(n_2),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_53),
.B(n_54),
.C(n_0),
.Y(n_55)
);

BUFx24_ASAP7_75t_SL g56 ( 
.A(n_55),
.Y(n_56)
);

XOR2xp5_ASAP7_75t_L g57 ( 
.A(n_56),
.B(n_6),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_57),
.B(n_7),
.Y(n_58)
);


endmodule