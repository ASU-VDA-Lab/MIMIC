module fake_jpeg_20299_n_261 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_261);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_261;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

BUFx10_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_14),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_8),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx16f_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_6),
.Y(n_32)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_15),
.B(n_0),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_34),
.B(n_41),
.Y(n_56)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

INVx3_ASAP7_75t_SL g60 ( 
.A(n_36),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_20),
.B(n_14),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_16),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_42),
.B(n_43),
.Y(n_65)
);

INVx4_ASAP7_75t_SL g43 ( 
.A(n_28),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_15),
.B(n_30),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_45),
.B(n_15),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g48 ( 
.A(n_45),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_48),
.B(n_67),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_42),
.B(n_15),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_49),
.B(n_15),
.Y(n_83)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_52),
.Y(n_70)
);

OAI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_35),
.A2(n_32),
.B1(n_29),
.B2(n_23),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_53),
.A2(n_24),
.B1(n_17),
.B2(n_22),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g54 ( 
.A1(n_34),
.A2(n_40),
.B(n_33),
.Y(n_54)
);

A2O1A1Ixp33_ASAP7_75t_L g93 ( 
.A1(n_54),
.A2(n_36),
.B(n_39),
.C(n_17),
.Y(n_93)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_57),
.Y(n_104)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_58),
.Y(n_71)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_59),
.Y(n_72)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_62),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_43),
.A2(n_32),
.B1(n_29),
.B2(n_23),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_63),
.A2(n_66),
.B1(n_22),
.B2(n_16),
.Y(n_105)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_64),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_43),
.A2(n_21),
.B1(n_20),
.B2(n_18),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_56),
.B(n_41),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_68),
.B(n_73),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_49),
.B(n_18),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_52),
.Y(n_74)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_74),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_65),
.B(n_54),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_75),
.B(n_76),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_60),
.B(n_21),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_61),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_77),
.B(n_78),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_51),
.B(n_30),
.Y(n_78)
);

OR2x2_ASAP7_75t_L g114 ( 
.A(n_79),
.B(n_100),
.Y(n_114)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_61),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_80),
.B(n_82),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_51),
.B(n_25),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_83),
.B(n_92),
.Y(n_107)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_61),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_85),
.B(n_86),
.Y(n_115)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_58),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_59),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_87),
.B(n_88),
.Y(n_121)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_62),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_51),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_89),
.B(n_96),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_64),
.A2(n_40),
.B1(n_43),
.B2(n_36),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_90),
.A2(n_26),
.B1(n_19),
.B2(n_3),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_51),
.B(n_44),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_91),
.B(n_95),
.C(n_103),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_46),
.B(n_38),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_93),
.A2(n_0),
.B(n_1),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_46),
.A2(n_39),
.B1(n_36),
.B2(n_38),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_94),
.A2(n_97),
.B1(n_105),
.B2(n_103),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_55),
.B(n_44),
.C(n_30),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_55),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_47),
.A2(n_44),
.B1(n_25),
.B2(n_24),
.Y(n_97)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_57),
.Y(n_98)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_98),
.Y(n_117)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_47),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_99),
.B(n_102),
.Y(n_131)
);

INVx1_ASAP7_75t_SL g100 ( 
.A(n_60),
.Y(n_100)
);

CKINVDCx5p33_ASAP7_75t_R g101 ( 
.A(n_60),
.Y(n_101)
);

OR2x2_ASAP7_75t_L g129 ( 
.A(n_101),
.B(n_27),
.Y(n_129)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_50),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_50),
.B(n_44),
.Y(n_103)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_61),
.Y(n_106)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_106),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_100),
.A2(n_30),
.B1(n_1),
.B2(n_2),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_108),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_71),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_111),
.B(n_112),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_101),
.Y(n_112)
);

CKINVDCx14_ASAP7_75t_R g164 ( 
.A(n_118),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_83),
.B(n_31),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_120),
.B(n_122),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_93),
.B(n_27),
.Y(n_122)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_98),
.Y(n_123)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_123),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_69),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_124),
.B(n_104),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_92),
.B(n_27),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_126),
.B(n_136),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_127),
.A2(n_137),
.B1(n_80),
.B2(n_102),
.Y(n_157)
);

NOR3xp33_ASAP7_75t_L g128 ( 
.A(n_79),
.B(n_26),
.C(n_19),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_128),
.B(n_133),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_129),
.Y(n_156)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_91),
.Y(n_133)
);

A2O1A1O1Ixp25_ASAP7_75t_L g134 ( 
.A1(n_103),
.A2(n_26),
.B(n_19),
.C(n_3),
.D(n_4),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_SL g142 ( 
.A(n_134),
.B(n_10),
.C(n_11),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_135),
.A2(n_94),
.B1(n_84),
.B2(n_81),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_72),
.B(n_1),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_97),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_95),
.B(n_7),
.Y(n_138)
);

OAI21xp33_ASAP7_75t_L g140 ( 
.A1(n_138),
.A2(n_10),
.B(n_11),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_140),
.B(n_137),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_142),
.B(n_143),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_116),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_146),
.A2(n_149),
.B1(n_157),
.B2(n_135),
.Y(n_182)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_116),
.Y(n_147)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_147),
.Y(n_166)
);

OAI22x1_ASAP7_75t_SL g149 ( 
.A1(n_122),
.A2(n_90),
.B1(n_91),
.B2(n_77),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_115),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_150),
.B(n_152),
.Y(n_175)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_131),
.Y(n_151)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_151),
.Y(n_169)
);

INVx5_ASAP7_75t_L g152 ( 
.A(n_130),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_113),
.B(n_70),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_153),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_107),
.B(n_74),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_154),
.B(n_158),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_110),
.B(n_70),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_155),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_107),
.B(n_104),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_121),
.Y(n_159)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_159),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_160),
.Y(n_178)
);

BUFx24_ASAP7_75t_SL g161 ( 
.A(n_125),
.Y(n_161)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_161),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_125),
.B(n_10),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_162),
.B(n_163),
.Y(n_172)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_132),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_158),
.B(n_120),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_173),
.B(n_183),
.Y(n_197)
);

MAJx3_ASAP7_75t_L g174 ( 
.A(n_149),
.B(n_133),
.C(n_118),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_SL g192 ( 
.A(n_174),
.B(n_180),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_164),
.A2(n_114),
.B(n_109),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_177),
.A2(n_181),
.B(n_156),
.Y(n_199)
);

OR2x2_ASAP7_75t_L g179 ( 
.A(n_144),
.B(n_111),
.Y(n_179)
);

OA22x2_ASAP7_75t_L g196 ( 
.A1(n_179),
.A2(n_182),
.B1(n_114),
.B2(n_129),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_145),
.A2(n_127),
.B(n_112),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_148),
.B(n_126),
.Y(n_183)
);

BUFx2_ASAP7_75t_L g184 ( 
.A(n_165),
.Y(n_184)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_184),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_148),
.B(n_154),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_185),
.B(n_186),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_144),
.B(n_136),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_174),
.A2(n_157),
.B1(n_145),
.B2(n_141),
.Y(n_190)
);

CKINVDCx14_ASAP7_75t_R g221 ( 
.A(n_190),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_171),
.B(n_150),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_191),
.B(n_193),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_171),
.B(n_152),
.Y(n_193)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_184),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_194),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_174),
.A2(n_156),
.B1(n_146),
.B2(n_151),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_195),
.A2(n_198),
.B1(n_202),
.B2(n_205),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g215 ( 
.A(n_196),
.B(n_182),
.Y(n_215)
);

INVx2_ASAP7_75t_SL g198 ( 
.A(n_184),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_199),
.A2(n_179),
.B(n_167),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_SL g200 ( 
.A(n_177),
.B(n_119),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_200),
.B(n_201),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_SL g201 ( 
.A(n_185),
.B(n_119),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_178),
.A2(n_139),
.B1(n_143),
.B2(n_114),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_SL g203 ( 
.A(n_180),
.B(n_142),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_203),
.B(n_204),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_170),
.B(n_124),
.Y(n_204)
);

CKINVDCx16_ASAP7_75t_R g205 ( 
.A(n_175),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_170),
.B(n_159),
.C(n_147),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_206),
.B(n_178),
.C(n_176),
.Y(n_209)
);

AND3x1_ASAP7_75t_L g207 ( 
.A(n_196),
.B(n_181),
.C(n_179),
.Y(n_207)
);

AOI31xp67_ASAP7_75t_L g224 ( 
.A1(n_207),
.A2(n_196),
.A3(n_204),
.B(n_197),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_209),
.B(n_214),
.C(n_206),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_192),
.B(n_173),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_211),
.B(n_220),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_213),
.A2(n_215),
.B(n_12),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_200),
.B(n_183),
.C(n_186),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_192),
.A2(n_169),
.B1(n_168),
.B2(n_195),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_216),
.A2(n_218),
.B1(n_198),
.B2(n_188),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_203),
.A2(n_169),
.B1(n_168),
.B2(n_166),
.Y(n_218)
);

AOI322xp5_ASAP7_75t_L g219 ( 
.A1(n_189),
.A2(n_166),
.A3(n_172),
.B1(n_187),
.B2(n_134),
.C1(n_129),
.C2(n_138),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_219),
.B(n_138),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_201),
.B(n_172),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_223),
.B(n_208),
.C(n_209),
.Y(n_243)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_224),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_225),
.B(n_226),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_217),
.B(n_187),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_227),
.B(n_228),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_221),
.A2(n_163),
.B(n_194),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_212),
.Y(n_229)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_229),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_215),
.A2(n_165),
.B1(n_117),
.B2(n_123),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_230),
.A2(n_234),
.B1(n_210),
.B2(n_214),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_213),
.A2(n_132),
.B1(n_117),
.B2(n_13),
.Y(n_232)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_232),
.Y(n_242)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_207),
.B(n_11),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_233),
.B(n_12),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_235),
.A2(n_231),
.B1(n_222),
.B2(n_208),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_237),
.A2(n_234),
.B1(n_224),
.B2(n_230),
.Y(n_245)
);

BUFx24_ASAP7_75t_SL g241 ( 
.A(n_223),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_241),
.B(n_243),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_243),
.B(n_231),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_244),
.B(n_245),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_235),
.A2(n_233),
.B1(n_220),
.B2(n_211),
.Y(n_246)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_246),
.B(n_240),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_247),
.B(n_248),
.C(n_239),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_236),
.B(n_222),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_250),
.B(n_248),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_244),
.B(n_238),
.C(n_242),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_251),
.B(n_253),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_SL g254 ( 
.A1(n_252),
.A2(n_249),
.B(n_246),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_254),
.B(n_255),
.C(n_12),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_256),
.Y(n_257)
);

BUFx24_ASAP7_75t_SL g259 ( 
.A(n_257),
.Y(n_259)
);

BUFx24_ASAP7_75t_SL g260 ( 
.A(n_259),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_260),
.B(n_258),
.Y(n_261)
);


endmodule