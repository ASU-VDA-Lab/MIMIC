module fake_jpeg_19625_n_251 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_251);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_251;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_12),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_15),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

INVx6_ASAP7_75t_SL g27 ( 
.A(n_15),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx4f_ASAP7_75t_SL g31 ( 
.A(n_2),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_5),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_13),
.Y(n_33)
);

INVx13_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

BUFx4f_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx2_ASAP7_75t_SL g38 ( 
.A(n_35),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_38),
.B(n_39),
.Y(n_62)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_42),
.B(n_44),
.Y(n_75)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_43),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_24),
.B(n_0),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_20),
.B(n_16),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_46),
.B(n_18),
.Y(n_63)
);

BUFx24_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

OR2x2_ASAP7_75t_L g50 ( 
.A(n_47),
.B(n_24),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_21),
.Y(n_48)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_39),
.B(n_42),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_49),
.B(n_51),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_50),
.B(n_37),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_44),
.B(n_35),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_41),
.A2(n_24),
.B1(n_25),
.B2(n_30),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_54),
.A2(n_57),
.B1(n_65),
.B2(n_29),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_44),
.A2(n_20),
.B1(n_32),
.B2(n_22),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_55),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_38),
.A2(n_25),
.B1(n_30),
.B2(n_32),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_56),
.A2(n_29),
.B1(n_23),
.B2(n_40),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_38),
.A2(n_30),
.B1(n_22),
.B2(n_33),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_58),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_46),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_61),
.B(n_63),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_47),
.A2(n_17),
.B1(n_18),
.B2(n_33),
.Y(n_65)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_66),
.Y(n_98)
);

NAND2xp33_ASAP7_75t_SL g67 ( 
.A(n_45),
.B(n_35),
.Y(n_67)
);

NAND2xp33_ASAP7_75t_SL g87 ( 
.A(n_67),
.B(n_35),
.Y(n_87)
);

OR2x2_ASAP7_75t_L g68 ( 
.A(n_45),
.B(n_17),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_68),
.Y(n_93)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_37),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_69),
.Y(n_91)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_36),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_70),
.Y(n_102)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_71),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_48),
.B(n_26),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_72),
.B(n_31),
.Y(n_78)
);

BUFx2_ASAP7_75t_L g76 ( 
.A(n_74),
.Y(n_76)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_76),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_78),
.B(n_84),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_80),
.A2(n_96),
.B(n_101),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_61),
.B(n_26),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_81),
.B(n_88),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_82),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_51),
.A2(n_40),
.B1(n_27),
.B2(n_43),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_83),
.A2(n_85),
.B1(n_86),
.B2(n_95),
.Y(n_129)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_66),
.Y(n_84)
);

OAI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_49),
.A2(n_52),
.B1(n_53),
.B2(n_55),
.Y(n_85)
);

AND2x2_ASAP7_75t_SL g111 ( 
.A(n_87),
.B(n_74),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_62),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_68),
.B(n_23),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_89),
.B(n_92),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_60),
.A2(n_27),
.B1(n_21),
.B2(n_35),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_90),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_62),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_68),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_94),
.B(n_100),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_50),
.A2(n_27),
.B1(n_48),
.B2(n_31),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_75),
.B(n_31),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_50),
.A2(n_31),
.B1(n_34),
.B2(n_2),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_97),
.A2(n_106),
.B1(n_53),
.B2(n_69),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_75),
.B(n_34),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_99),
.B(n_64),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_58),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_60),
.A2(n_34),
.B1(n_1),
.B2(n_2),
.Y(n_101)
);

AO22x1_ASAP7_75t_L g105 ( 
.A1(n_67),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_105)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_105),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_52),
.A2(n_0),
.B1(n_1),
.B2(n_4),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_111),
.A2(n_80),
.B(n_87),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_79),
.B(n_71),
.C(n_64),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_113),
.B(n_114),
.C(n_127),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_79),
.B(n_92),
.C(n_88),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_104),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_115),
.B(n_117),
.Y(n_148)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_91),
.Y(n_116)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_116),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_104),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_119),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_77),
.B(n_14),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_120),
.B(n_131),
.Y(n_138)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_91),
.Y(n_124)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_124),
.Y(n_140)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_91),
.Y(n_126)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_126),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_93),
.B(n_64),
.C(n_70),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_86),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_128),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_130),
.A2(n_73),
.B1(n_107),
.B2(n_94),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_100),
.B(n_16),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_76),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_132),
.Y(n_147)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_76),
.Y(n_133)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_133),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_118),
.A2(n_111),
.B(n_125),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_134),
.A2(n_136),
.B(n_144),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_137),
.A2(n_154),
.B1(n_128),
.B2(n_117),
.Y(n_164)
);

BUFx2_ASAP7_75t_L g139 ( 
.A(n_133),
.Y(n_139)
);

CKINVDCx14_ASAP7_75t_R g160 ( 
.A(n_139),
.Y(n_160)
);

INVx2_ASAP7_75t_SL g141 ( 
.A(n_116),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_141),
.B(n_145),
.Y(n_180)
);

AND2x4_ASAP7_75t_L g144 ( 
.A(n_111),
.B(n_80),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_122),
.B(n_96),
.Y(n_145)
);

OAI21xp33_ASAP7_75t_SL g146 ( 
.A1(n_129),
.A2(n_93),
.B(n_105),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_146),
.A2(n_153),
.B(n_155),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_121),
.B(n_110),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_150),
.B(n_152),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_110),
.B(n_96),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_112),
.B(n_105),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_129),
.A2(n_107),
.B1(n_73),
.B2(n_83),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_118),
.A2(n_102),
.B(n_97),
.Y(n_155)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_124),
.Y(n_157)
);

BUFx2_ASAP7_75t_L g174 ( 
.A(n_157),
.Y(n_174)
);

A2O1A1Ixp33_ASAP7_75t_L g158 ( 
.A1(n_112),
.A2(n_95),
.B(n_102),
.C(n_103),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_158),
.B(n_153),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_114),
.B(n_103),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_159),
.B(n_108),
.Y(n_175)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_148),
.Y(n_161)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_161),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_148),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_163),
.B(n_167),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_164),
.B(n_166),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_142),
.B(n_115),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_135),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_168),
.A2(n_173),
.B(n_155),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_159),
.B(n_113),
.C(n_127),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_169),
.B(n_175),
.C(n_182),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_156),
.B(n_125),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_170),
.B(n_171),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_156),
.B(n_109),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_153),
.B(n_130),
.Y(n_172)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_172),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_136),
.A2(n_123),
.B(n_132),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_134),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_177),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_158),
.B(n_126),
.Y(n_178)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_178),
.Y(n_197)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_135),
.Y(n_179)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_179),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_151),
.B(n_108),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_181),
.B(n_163),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_144),
.B(n_84),
.C(n_98),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_183),
.B(n_195),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_176),
.B(n_138),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_185),
.B(n_13),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_186),
.A2(n_190),
.B(n_173),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_165),
.A2(n_144),
.B(n_151),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_169),
.B(n_144),
.C(n_154),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_194),
.B(n_198),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_181),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_172),
.A2(n_123),
.B1(n_147),
.B2(n_149),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_196),
.A2(n_141),
.B1(n_143),
.B2(n_174),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_170),
.B(n_149),
.C(n_140),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_174),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_199),
.B(n_139),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_184),
.A2(n_178),
.B1(n_161),
.B2(n_168),
.Y(n_201)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_201),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_202),
.A2(n_205),
.B1(n_194),
.B2(n_190),
.Y(n_216)
);

AOI321xp33_ASAP7_75t_L g204 ( 
.A1(n_192),
.A2(n_165),
.A3(n_162),
.B1(n_171),
.B2(n_175),
.C(n_180),
.Y(n_204)
);

AOI31xp67_ASAP7_75t_L g223 ( 
.A1(n_204),
.A2(n_187),
.A3(n_210),
.B(n_205),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_186),
.A2(n_162),
.B(n_182),
.Y(n_205)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_206),
.Y(n_224)
);

AOI322xp5_ASAP7_75t_L g207 ( 
.A1(n_197),
.A2(n_180),
.A3(n_164),
.B1(n_166),
.B2(n_179),
.C1(n_167),
.C2(n_140),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_207),
.B(n_212),
.Y(n_217)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_208),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_184),
.A2(n_160),
.B1(n_141),
.B2(n_157),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_209),
.B(n_211),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_193),
.A2(n_143),
.B(n_5),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_197),
.A2(n_174),
.B1(n_59),
.B2(n_98),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_213),
.B(n_196),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_193),
.A2(n_4),
.B(n_6),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_214),
.B(n_198),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_216),
.B(n_202),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_203),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_219),
.B(n_221),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_220),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_210),
.B(n_187),
.C(n_192),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_222),
.B(n_189),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_223),
.A2(n_222),
.B1(n_216),
.B2(n_204),
.Y(n_232)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_224),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_228),
.B(n_231),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_229),
.B(n_232),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_215),
.A2(n_191),
.B(n_201),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_230),
.A2(n_227),
.B(n_226),
.Y(n_237)
);

A2O1A1Ixp33_ASAP7_75t_L g231 ( 
.A1(n_218),
.A2(n_191),
.B(n_189),
.C(n_188),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_233),
.B(n_217),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_234),
.A2(n_237),
.B(n_239),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_230),
.A2(n_209),
.B1(n_220),
.B2(n_215),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_236),
.A2(n_235),
.B1(n_237),
.B2(n_238),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_229),
.B(n_225),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_240),
.B(n_241),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_238),
.A2(n_231),
.B1(n_200),
.B2(n_211),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_239),
.A2(n_200),
.B(n_213),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_243),
.A2(n_199),
.B(n_242),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_245),
.A2(n_246),
.B(n_8),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_240),
.A2(n_4),
.B(n_7),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_247),
.B(n_248),
.C(n_59),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_244),
.A2(n_8),
.B(n_9),
.Y(n_248)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_249),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_250),
.A2(n_8),
.B(n_9),
.Y(n_251)
);


endmodule