module fake_jpeg_29698_n_174 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_174);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_174;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_7),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_27),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_14),
.Y(n_51)
);

INVx13_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_1),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_28),
.Y(n_54)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_6),
.Y(n_55)
);

BUFx16f_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_23),
.B(n_13),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_4),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_20),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_29),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_22),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_9),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_15),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_10),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_17),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_33),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_24),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_16),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_10),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_70),
.B(n_72),
.Y(n_81)
);

INVx3_ASAP7_75t_SL g71 ( 
.A(n_56),
.Y(n_71)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_71),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_58),
.B(n_0),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_50),
.Y(n_73)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_73),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_56),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_74),
.B(n_76),
.Y(n_84)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_52),
.Y(n_75)
);

INVx11_ASAP7_75t_L g78 ( 
.A(n_75),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_57),
.Y(n_76)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_52),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_77),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_73),
.A2(n_60),
.B1(n_50),
.B2(n_54),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_82),
.A2(n_47),
.B1(n_53),
.B2(n_60),
.Y(n_96)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_75),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_83),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_74),
.A2(n_47),
.B1(n_53),
.B2(n_68),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_86),
.A2(n_68),
.B1(n_54),
.B2(n_63),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_71),
.B(n_62),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_87),
.B(n_89),
.Y(n_92)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_77),
.Y(n_88)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_88),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_70),
.B(n_64),
.Y(n_89)
);

OR2x2_ASAP7_75t_L g90 ( 
.A(n_71),
.B(n_69),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_90),
.B(n_48),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_85),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_91),
.B(n_98),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_90),
.B(n_69),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_93),
.B(n_97),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_96),
.A2(n_106),
.B1(n_107),
.B2(n_108),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_81),
.B(n_49),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_79),
.Y(n_98)
);

INVx1_ASAP7_75t_SL g99 ( 
.A(n_79),
.Y(n_99)
);

OR2x2_ASAP7_75t_L g120 ( 
.A(n_99),
.B(n_102),
.Y(n_120)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_83),
.Y(n_100)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_100),
.Y(n_112)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_79),
.Y(n_101)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_101),
.Y(n_128)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_80),
.Y(n_103)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_103),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_84),
.B(n_51),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_104),
.B(n_105),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_82),
.B(n_59),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_86),
.A2(n_63),
.B1(n_48),
.B2(n_61),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_80),
.A2(n_67),
.B1(n_65),
.B2(n_66),
.Y(n_108)
);

AOI32xp33_ASAP7_75t_L g111 ( 
.A1(n_108),
.A2(n_26),
.A3(n_31),
.B1(n_46),
.B2(n_44),
.Y(n_111)
);

OR2x2_ASAP7_75t_SL g133 ( 
.A(n_111),
.B(n_25),
.Y(n_133)
);

OAI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_91),
.A2(n_55),
.B1(n_78),
.B2(n_21),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_115),
.A2(n_127),
.B1(n_129),
.B2(n_11),
.Y(n_142)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_95),
.Y(n_116)
);

INVxp67_ASAP7_75t_SL g144 ( 
.A(n_116),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_92),
.B(n_55),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_118),
.B(n_122),
.Y(n_139)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_94),
.Y(n_119)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_119),
.Y(n_146)
);

OR2x2_ASAP7_75t_L g121 ( 
.A(n_99),
.B(n_78),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_121),
.B(n_125),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_95),
.B(n_0),
.Y(n_122)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_98),
.Y(n_123)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_123),
.Y(n_136)
);

O2A1O1Ixp33_ASAP7_75t_L g124 ( 
.A1(n_105),
.A2(n_19),
.B(n_41),
.C(n_40),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_124),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_108),
.Y(n_125)
);

BUFx24_ASAP7_75t_SL g126 ( 
.A(n_97),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_126),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_105),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_105),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_114),
.B(n_30),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_131),
.B(n_11),
.C(n_12),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_110),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_132),
.B(n_138),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_133),
.A2(n_140),
.B1(n_148),
.B2(n_123),
.Y(n_149)
);

INVx13_ASAP7_75t_L g135 ( 
.A(n_128),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_135),
.B(n_142),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_120),
.A2(n_5),
.B(n_6),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_137),
.B(n_141),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_113),
.B(n_5),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_L g140 ( 
.A1(n_117),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_120),
.B(n_8),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_121),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_145),
.Y(n_156)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_112),
.Y(n_147)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_147),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_116),
.A2(n_34),
.B1(n_39),
.B2(n_38),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_149),
.B(n_150),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_134),
.A2(n_124),
.B(n_115),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_145),
.A2(n_132),
.B(n_143),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_151),
.B(n_154),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_131),
.B(n_109),
.Y(n_154)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_158),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_151),
.A2(n_157),
.B1(n_156),
.B2(n_152),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_161),
.A2(n_163),
.B1(n_153),
.B2(n_136),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_155),
.A2(n_139),
.B1(n_148),
.B2(n_146),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_164),
.B(n_165),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_160),
.B(n_154),
.C(n_158),
.Y(n_165)
);

BUFx2_ASAP7_75t_L g166 ( 
.A(n_161),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_167),
.B(n_162),
.Y(n_168)
);

AOI322xp5_ASAP7_75t_L g169 ( 
.A1(n_168),
.A2(n_159),
.A3(n_166),
.B1(n_135),
.B2(n_133),
.C1(n_144),
.C2(n_36),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_169),
.B(n_37),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_170),
.A2(n_130),
.B1(n_32),
.B2(n_18),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_171),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_172),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_173),
.B(n_166),
.Y(n_174)
);


endmodule