module fake_aes_12453_n_655 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_71, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_72, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_655);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_71;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_72;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_655;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_73;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_490;
wire n_247;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_423;
wire n_342;
wire n_420;
wire n_621;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_78;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_75;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_445;
wire n_398;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_74;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_487;
wire n_451;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_99;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g73 ( .A(n_58), .Y(n_73) );
CKINVDCx14_ASAP7_75t_R g74 ( .A(n_4), .Y(n_74) );
BUFx2_ASAP7_75t_L g75 ( .A(n_69), .Y(n_75) );
INVx2_ASAP7_75t_L g76 ( .A(n_15), .Y(n_76) );
CKINVDCx20_ASAP7_75t_R g77 ( .A(n_55), .Y(n_77) );
BUFx2_ASAP7_75t_L g78 ( .A(n_56), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_51), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_30), .Y(n_80) );
INVxp33_ASAP7_75t_L g81 ( .A(n_62), .Y(n_81) );
CKINVDCx20_ASAP7_75t_R g82 ( .A(n_67), .Y(n_82) );
CKINVDCx5p33_ASAP7_75t_R g83 ( .A(n_70), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_65), .Y(n_84) );
CKINVDCx5p33_ASAP7_75t_R g85 ( .A(n_19), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_66), .Y(n_86) );
INVx2_ASAP7_75t_L g87 ( .A(n_71), .Y(n_87) );
CKINVDCx5p33_ASAP7_75t_R g88 ( .A(n_61), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_24), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_32), .Y(n_90) );
CKINVDCx5p33_ASAP7_75t_R g91 ( .A(n_63), .Y(n_91) );
CKINVDCx16_ASAP7_75t_R g92 ( .A(n_54), .Y(n_92) );
INVx2_ASAP7_75t_L g93 ( .A(n_68), .Y(n_93) );
CKINVDCx20_ASAP7_75t_R g94 ( .A(n_9), .Y(n_94) );
CKINVDCx5p33_ASAP7_75t_R g95 ( .A(n_15), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_50), .Y(n_96) );
INVx2_ASAP7_75t_L g97 ( .A(n_47), .Y(n_97) );
CKINVDCx5p33_ASAP7_75t_R g98 ( .A(n_33), .Y(n_98) );
CKINVDCx14_ASAP7_75t_R g99 ( .A(n_4), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_49), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_35), .Y(n_101) );
INVx2_ASAP7_75t_L g102 ( .A(n_57), .Y(n_102) );
NOR2xp67_ASAP7_75t_L g103 ( .A(n_64), .B(n_26), .Y(n_103) );
CKINVDCx5p33_ASAP7_75t_R g104 ( .A(n_52), .Y(n_104) );
INVx2_ASAP7_75t_SL g105 ( .A(n_53), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_59), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g107 ( .A(n_60), .Y(n_107) );
CKINVDCx5p33_ASAP7_75t_R g108 ( .A(n_48), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_28), .Y(n_109) );
INVxp67_ASAP7_75t_SL g110 ( .A(n_13), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_37), .Y(n_111) );
HB1xp67_ASAP7_75t_L g112 ( .A(n_27), .Y(n_112) );
INVxp67_ASAP7_75t_L g113 ( .A(n_44), .Y(n_113) );
BUFx6f_ASAP7_75t_L g114 ( .A(n_87), .Y(n_114) );
BUFx2_ASAP7_75t_L g115 ( .A(n_74), .Y(n_115) );
INVx2_ASAP7_75t_L g116 ( .A(n_87), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_73), .Y(n_117) );
BUFx6f_ASAP7_75t_L g118 ( .A(n_93), .Y(n_118) );
INVx2_ASAP7_75t_SL g119 ( .A(n_75), .Y(n_119) );
CKINVDCx5p33_ASAP7_75t_R g120 ( .A(n_92), .Y(n_120) );
BUFx3_ASAP7_75t_L g121 ( .A(n_75), .Y(n_121) );
INVx2_ASAP7_75t_L g122 ( .A(n_93), .Y(n_122) );
AND2x2_ASAP7_75t_SL g123 ( .A(n_78), .B(n_20), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_73), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_79), .Y(n_125) );
AOI22x1_ASAP7_75t_SL g126 ( .A1(n_94), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_79), .Y(n_127) );
CKINVDCx5p33_ASAP7_75t_R g128 ( .A(n_92), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g129 ( .A(n_78), .B(n_0), .Y(n_129) );
BUFx6f_ASAP7_75t_L g130 ( .A(n_97), .Y(n_130) );
INVx2_ASAP7_75t_L g131 ( .A(n_97), .Y(n_131) );
OAI21x1_ASAP7_75t_L g132 ( .A1(n_102), .A2(n_40), .B(n_72), .Y(n_132) );
AND2x4_ASAP7_75t_L g133 ( .A(n_105), .B(n_1), .Y(n_133) );
INVx2_ASAP7_75t_L g134 ( .A(n_114), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_114), .Y(n_135) );
INVx2_ASAP7_75t_L g136 ( .A(n_114), .Y(n_136) );
INVx2_ASAP7_75t_L g137 ( .A(n_114), .Y(n_137) );
BUFx3_ASAP7_75t_L g138 ( .A(n_133), .Y(n_138) );
BUFx3_ASAP7_75t_L g139 ( .A(n_133), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_114), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_114), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_114), .Y(n_142) );
INVx1_ASAP7_75t_SL g143 ( .A(n_115), .Y(n_143) );
INVx2_ASAP7_75t_L g144 ( .A(n_118), .Y(n_144) );
INVx1_ASAP7_75t_SL g145 ( .A(n_115), .Y(n_145) );
NAND2xp33_ASAP7_75t_SL g146 ( .A(n_120), .B(n_77), .Y(n_146) );
OR2x6_ASAP7_75t_L g147 ( .A(n_129), .B(n_112), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g148 ( .A(n_121), .B(n_105), .Y(n_148) );
INVx2_ASAP7_75t_SL g149 ( .A(n_117), .Y(n_149) );
NAND2xp33_ASAP7_75t_L g150 ( .A(n_119), .B(n_83), .Y(n_150) );
NAND2xp33_ASAP7_75t_L g151 ( .A(n_119), .B(n_85), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_118), .Y(n_152) );
INVx2_ASAP7_75t_L g153 ( .A(n_118), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_121), .B(n_102), .Y(n_154) );
BUFx6f_ASAP7_75t_L g155 ( .A(n_132), .Y(n_155) );
AND2x4_ASAP7_75t_L g156 ( .A(n_121), .B(n_76), .Y(n_156) );
CKINVDCx16_ASAP7_75t_R g157 ( .A(n_119), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_118), .Y(n_158) );
INVx4_ASAP7_75t_L g159 ( .A(n_133), .Y(n_159) );
AND2x2_ASAP7_75t_SL g160 ( .A(n_123), .B(n_80), .Y(n_160) );
BUFx3_ASAP7_75t_L g161 ( .A(n_133), .Y(n_161) );
INVx2_ASAP7_75t_SL g162 ( .A(n_117), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_118), .Y(n_163) );
INVx3_ASAP7_75t_L g164 ( .A(n_133), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_148), .B(n_129), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_156), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_156), .Y(n_167) );
AOI22xp5_ASAP7_75t_L g168 ( .A1(n_160), .A2(n_123), .B1(n_128), .B2(n_99), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_148), .B(n_124), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_154), .B(n_124), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_156), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_156), .Y(n_172) );
AND2x6_ASAP7_75t_SL g173 ( .A(n_147), .B(n_126), .Y(n_173) );
INVx1_ASAP7_75t_SL g174 ( .A(n_143), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_154), .B(n_125), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_156), .Y(n_176) );
AOI22xp5_ASAP7_75t_L g177 ( .A1(n_160), .A2(n_123), .B1(n_82), .B2(n_95), .Y(n_177) );
NAND2xp5_ASAP7_75t_SL g178 ( .A(n_149), .B(n_123), .Y(n_178) );
INVx4_ASAP7_75t_L g179 ( .A(n_159), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_138), .Y(n_180) );
NAND2xp5_ASAP7_75t_SL g181 ( .A(n_149), .B(n_125), .Y(n_181) );
OAI221xp5_ASAP7_75t_L g182 ( .A1(n_147), .A2(n_127), .B1(n_110), .B2(n_76), .C(n_116), .Y(n_182) );
INVx1_ASAP7_75t_L g183 ( .A(n_138), .Y(n_183) );
INVx2_ASAP7_75t_L g184 ( .A(n_164), .Y(n_184) );
NAND2xp5_ASAP7_75t_SL g185 ( .A(n_149), .B(n_127), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_164), .Y(n_186) );
NAND2xp5_ASAP7_75t_SL g187 ( .A(n_162), .B(n_80), .Y(n_187) );
INVx2_ASAP7_75t_L g188 ( .A(n_164), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_164), .Y(n_189) );
INVx4_ASAP7_75t_L g190 ( .A(n_159), .Y(n_190) );
NOR2xp67_ASAP7_75t_L g191 ( .A(n_159), .B(n_116), .Y(n_191) );
INVx2_ASAP7_75t_L g192 ( .A(n_159), .Y(n_192) );
INVx2_ASAP7_75t_L g193 ( .A(n_138), .Y(n_193) );
INVx2_ASAP7_75t_L g194 ( .A(n_139), .Y(n_194) );
NAND3xp33_ASAP7_75t_L g195 ( .A(n_150), .B(n_126), .C(n_84), .Y(n_195) );
NOR2xp33_ASAP7_75t_L g196 ( .A(n_157), .B(n_81), .Y(n_196) );
OR2x6_ASAP7_75t_L g197 ( .A(n_147), .B(n_132), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_162), .B(n_88), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_139), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_162), .B(n_91), .Y(n_200) );
NOR2x2_ASAP7_75t_L g201 ( .A(n_147), .B(n_116), .Y(n_201) );
NAND3xp33_ASAP7_75t_SL g202 ( .A(n_143), .B(n_108), .C(n_107), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_147), .B(n_98), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_147), .B(n_104), .Y(n_204) );
INVx2_ASAP7_75t_L g205 ( .A(n_139), .Y(n_205) );
NOR2xp33_ASAP7_75t_L g206 ( .A(n_157), .B(n_113), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_160), .B(n_122), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_165), .B(n_145), .Y(n_208) );
AOI22xp5_ASAP7_75t_L g209 ( .A1(n_178), .A2(n_145), .B1(n_151), .B2(n_146), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_169), .B(n_161), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_170), .B(n_161), .Y(n_211) );
AOI22xp33_ASAP7_75t_L g212 ( .A1(n_178), .A2(n_161), .B1(n_155), .B2(n_131), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_175), .B(n_196), .Y(n_213) );
OR2x6_ASAP7_75t_L g214 ( .A(n_179), .B(n_155), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_166), .Y(n_215) );
AOI21x1_ASAP7_75t_L g216 ( .A1(n_197), .A2(n_132), .B(n_158), .Y(n_216) );
CKINVDCx5p33_ASAP7_75t_R g217 ( .A(n_174), .Y(n_217) );
OAI22xp5_ASAP7_75t_L g218 ( .A1(n_177), .A2(n_155), .B1(n_131), .B2(n_122), .Y(n_218) );
OAI21x1_ASAP7_75t_L g219 ( .A1(n_187), .A2(n_136), .B(n_137), .Y(n_219) );
OAI21xp5_ASAP7_75t_L g220 ( .A1(n_186), .A2(n_163), .B(n_158), .Y(n_220) );
INVx2_ASAP7_75t_SL g221 ( .A(n_203), .Y(n_221) );
AOI21xp5_ASAP7_75t_L g222 ( .A1(n_181), .A2(n_155), .B(n_163), .Y(n_222) );
NAND2xp5_ASAP7_75t_SL g223 ( .A(n_179), .B(n_155), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_206), .B(n_155), .Y(n_224) );
OAI21xp5_ASAP7_75t_L g225 ( .A1(n_186), .A2(n_141), .B(n_140), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_204), .B(n_155), .Y(n_226) );
AOI21xp5_ASAP7_75t_L g227 ( .A1(n_181), .A2(n_140), .B(n_152), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_167), .B(n_122), .Y(n_228) );
NAND2xp5_ASAP7_75t_SL g229 ( .A(n_179), .B(n_84), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_171), .B(n_131), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_172), .B(n_176), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_189), .Y(n_232) );
AO21x1_ASAP7_75t_L g233 ( .A1(n_187), .A2(n_86), .B(n_109), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_189), .Y(n_234) );
NAND2xp5_ASAP7_75t_SL g235 ( .A(n_190), .B(n_86), .Y(n_235) );
O2A1O1Ixp33_ASAP7_75t_L g236 ( .A1(n_182), .A2(n_111), .B(n_90), .C(n_96), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_190), .B(n_89), .Y(n_237) );
NOR2x1_ASAP7_75t_L g238 ( .A(n_202), .B(n_89), .Y(n_238) );
NAND2xp5_ASAP7_75t_SL g239 ( .A(n_190), .B(n_90), .Y(n_239) );
A2O1A1Ixp33_ASAP7_75t_L g240 ( .A1(n_207), .A2(n_96), .B(n_100), .C(n_101), .Y(n_240) );
NAND2xp5_ASAP7_75t_SL g241 ( .A(n_184), .B(n_100), .Y(n_241) );
NOR2x1p5_ASAP7_75t_SL g242 ( .A(n_184), .B(n_134), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_192), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_208), .B(n_168), .Y(n_244) );
OAI21x1_ASAP7_75t_L g245 ( .A1(n_216), .A2(n_188), .B(n_185), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_237), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_213), .B(n_191), .Y(n_247) );
AOI21xp5_ASAP7_75t_L g248 ( .A1(n_223), .A2(n_185), .B(n_197), .Y(n_248) );
BUFx3_ASAP7_75t_L g249 ( .A(n_217), .Y(n_249) );
AOI21xp5_ASAP7_75t_L g250 ( .A1(n_223), .A2(n_197), .B(n_188), .Y(n_250) );
AO31x2_ASAP7_75t_L g251 ( .A1(n_240), .A2(n_152), .A3(n_142), .B(n_135), .Y(n_251) );
OAI21xp5_ASAP7_75t_L g252 ( .A1(n_226), .A2(n_197), .B(n_180), .Y(n_252) );
INVx3_ASAP7_75t_L g253 ( .A(n_214), .Y(n_253) );
AOI22xp5_ASAP7_75t_L g254 ( .A1(n_221), .A2(n_195), .B1(n_199), .B2(n_183), .Y(n_254) );
AOI21xp5_ASAP7_75t_L g255 ( .A1(n_222), .A2(n_200), .B(n_198), .Y(n_255) );
INVx6_ASAP7_75t_SL g256 ( .A(n_214), .Y(n_256) );
OAI21x1_ASAP7_75t_L g257 ( .A1(n_219), .A2(n_193), .B(n_194), .Y(n_257) );
AOI21xp5_ASAP7_75t_L g258 ( .A1(n_224), .A2(n_192), .B(n_205), .Y(n_258) );
INVx2_ASAP7_75t_L g259 ( .A(n_214), .Y(n_259) );
NAND2xp5_ASAP7_75t_SL g260 ( .A(n_212), .B(n_193), .Y(n_260) );
A2O1A1Ixp33_ASAP7_75t_L g261 ( .A1(n_236), .A2(n_205), .B(n_194), .C(n_103), .Y(n_261) );
AO32x2_ASAP7_75t_L g262 ( .A1(n_218), .A2(n_201), .A3(n_118), .B1(n_130), .B2(n_173), .Y(n_262) );
OR2x6_ASAP7_75t_L g263 ( .A(n_214), .B(n_201), .Y(n_263) );
AO31x2_ASAP7_75t_L g264 ( .A1(n_240), .A2(n_142), .A3(n_141), .B(n_135), .Y(n_264) );
AO21x2_ASAP7_75t_L g265 ( .A1(n_233), .A2(n_103), .B(n_101), .Y(n_265) );
INVxp67_ASAP7_75t_L g266 ( .A(n_229), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_228), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_267), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_244), .B(n_215), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_246), .Y(n_270) );
AOI21xp5_ASAP7_75t_L g271 ( .A1(n_255), .A2(n_219), .B(n_241), .Y(n_271) );
AOI22xp5_ASAP7_75t_L g272 ( .A1(n_263), .A2(n_209), .B1(n_238), .B2(n_229), .Y(n_272) );
OAI21xp5_ASAP7_75t_L g273 ( .A1(n_258), .A2(n_241), .B(n_234), .Y(n_273) );
OA21x2_ASAP7_75t_L g274 ( .A1(n_257), .A2(n_225), .B(n_220), .Y(n_274) );
OAI21xp5_ASAP7_75t_L g275 ( .A1(n_261), .A2(n_232), .B(n_230), .Y(n_275) );
OAI21x1_ASAP7_75t_L g276 ( .A1(n_245), .A2(n_227), .B(n_235), .Y(n_276) );
AO21x1_ASAP7_75t_L g277 ( .A1(n_252), .A2(n_235), .B(n_239), .Y(n_277) );
CKINVDCx5p33_ASAP7_75t_R g278 ( .A(n_249), .Y(n_278) );
AOI21x1_ASAP7_75t_L g279 ( .A1(n_250), .A2(n_239), .B(n_134), .Y(n_279) );
OA21x2_ASAP7_75t_L g280 ( .A1(n_248), .A2(n_137), .B(n_134), .Y(n_280) );
AO21x2_ASAP7_75t_L g281 ( .A1(n_265), .A2(n_231), .B(n_109), .Y(n_281) );
AND2x2_ASAP7_75t_L g282 ( .A(n_263), .B(n_210), .Y(n_282) );
NOR2x1_ASAP7_75t_L g283 ( .A(n_263), .B(n_106), .Y(n_283) );
INVx2_ASAP7_75t_L g284 ( .A(n_259), .Y(n_284) );
BUFx2_ASAP7_75t_L g285 ( .A(n_256), .Y(n_285) );
AOI21xp5_ASAP7_75t_L g286 ( .A1(n_260), .A2(n_211), .B(n_243), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_247), .B(n_242), .Y(n_287) );
OAI21x1_ASAP7_75t_L g288 ( .A1(n_253), .A2(n_153), .B(n_144), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_251), .Y(n_289) );
INVx2_ASAP7_75t_L g290 ( .A(n_280), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_269), .B(n_251), .Y(n_291) );
AO21x2_ASAP7_75t_L g292 ( .A1(n_271), .A2(n_265), .B(n_261), .Y(n_292) );
INVx2_ASAP7_75t_L g293 ( .A(n_280), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_284), .Y(n_294) );
NOR2x1_ASAP7_75t_R g295 ( .A(n_278), .B(n_249), .Y(n_295) );
INVx2_ASAP7_75t_L g296 ( .A(n_280), .Y(n_296) );
AND2x2_ASAP7_75t_L g297 ( .A(n_268), .B(n_262), .Y(n_297) );
INVx2_ASAP7_75t_L g298 ( .A(n_280), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_269), .B(n_251), .Y(n_299) );
OA21x2_ASAP7_75t_L g300 ( .A1(n_271), .A2(n_259), .B(n_266), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_284), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_284), .Y(n_302) );
AO21x2_ASAP7_75t_L g303 ( .A1(n_281), .A2(n_254), .B(n_106), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_289), .Y(n_304) );
CKINVDCx20_ASAP7_75t_R g305 ( .A(n_285), .Y(n_305) );
OAI21xp5_ASAP7_75t_L g306 ( .A1(n_275), .A2(n_266), .B(n_253), .Y(n_306) );
AND2x4_ASAP7_75t_L g307 ( .A(n_282), .B(n_251), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_289), .Y(n_308) );
INVx3_ASAP7_75t_L g309 ( .A(n_288), .Y(n_309) );
HB1xp67_ASAP7_75t_L g310 ( .A(n_268), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_270), .Y(n_311) );
INVx2_ASAP7_75t_L g312 ( .A(n_281), .Y(n_312) );
OR2x2_ASAP7_75t_L g313 ( .A(n_270), .B(n_264), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_287), .Y(n_314) );
AND2x2_ASAP7_75t_L g315 ( .A(n_282), .B(n_262), .Y(n_315) );
HB1xp67_ASAP7_75t_L g316 ( .A(n_283), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_287), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_281), .Y(n_318) );
BUFx6f_ASAP7_75t_L g319 ( .A(n_288), .Y(n_319) );
OR2x6_ASAP7_75t_L g320 ( .A(n_283), .B(n_256), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_281), .Y(n_321) );
INVx2_ASAP7_75t_L g322 ( .A(n_279), .Y(n_322) );
AOI22xp5_ASAP7_75t_L g323 ( .A1(n_314), .A2(n_272), .B1(n_277), .B2(n_275), .Y(n_323) );
INVx2_ASAP7_75t_L g324 ( .A(n_290), .Y(n_324) );
HB1xp67_ASAP7_75t_L g325 ( .A(n_310), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_304), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_304), .Y(n_327) );
INVx3_ASAP7_75t_L g328 ( .A(n_319), .Y(n_328) );
INVx2_ASAP7_75t_L g329 ( .A(n_294), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_308), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_308), .Y(n_331) );
AND2x2_ASAP7_75t_L g332 ( .A(n_307), .B(n_262), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_311), .B(n_272), .Y(n_333) );
HB1xp67_ASAP7_75t_L g334 ( .A(n_294), .Y(n_334) );
AND2x4_ASAP7_75t_L g335 ( .A(n_307), .B(n_279), .Y(n_335) );
INVx3_ASAP7_75t_L g336 ( .A(n_319), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_314), .B(n_277), .Y(n_337) );
AND2x2_ASAP7_75t_L g338 ( .A(n_307), .B(n_262), .Y(n_338) );
AND2x2_ASAP7_75t_L g339 ( .A(n_307), .B(n_264), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_317), .Y(n_340) );
INVx2_ASAP7_75t_L g341 ( .A(n_290), .Y(n_341) );
INVx2_ASAP7_75t_L g342 ( .A(n_290), .Y(n_342) );
OR2x2_ASAP7_75t_L g343 ( .A(n_317), .B(n_264), .Y(n_343) );
INVx2_ASAP7_75t_L g344 ( .A(n_293), .Y(n_344) );
INVx3_ASAP7_75t_L g345 ( .A(n_319), .Y(n_345) );
AND2x2_ASAP7_75t_L g346 ( .A(n_297), .B(n_264), .Y(n_346) );
AND2x2_ASAP7_75t_L g347 ( .A(n_297), .B(n_111), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_313), .Y(n_348) );
CKINVDCx5p33_ASAP7_75t_R g349 ( .A(n_305), .Y(n_349) );
NAND2x1p5_ASAP7_75t_SL g350 ( .A(n_312), .B(n_136), .Y(n_350) );
NOR2x1_ASAP7_75t_L g351 ( .A(n_320), .B(n_273), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_313), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_301), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_302), .Y(n_354) );
OR2x2_ASAP7_75t_L g355 ( .A(n_291), .B(n_273), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_302), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_291), .Y(n_357) );
INVxp67_ASAP7_75t_L g358 ( .A(n_295), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_299), .Y(n_359) );
NOR2xp33_ASAP7_75t_L g360 ( .A(n_295), .B(n_320), .Y(n_360) );
AND2x2_ASAP7_75t_L g361 ( .A(n_315), .B(n_274), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_299), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_318), .Y(n_363) );
AND2x2_ASAP7_75t_L g364 ( .A(n_315), .B(n_274), .Y(n_364) );
INVx2_ASAP7_75t_L g365 ( .A(n_293), .Y(n_365) );
OR2x6_ASAP7_75t_L g366 ( .A(n_320), .B(n_286), .Y(n_366) );
BUFx2_ASAP7_75t_L g367 ( .A(n_309), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_318), .Y(n_368) );
AND2x2_ASAP7_75t_L g369 ( .A(n_321), .B(n_274), .Y(n_369) );
AND2x4_ASAP7_75t_L g370 ( .A(n_309), .B(n_276), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_316), .B(n_118), .Y(n_371) );
INVx2_ASAP7_75t_L g372 ( .A(n_293), .Y(n_372) );
AND2x2_ASAP7_75t_L g373 ( .A(n_321), .B(n_274), .Y(n_373) );
INVx3_ASAP7_75t_L g374 ( .A(n_319), .Y(n_374) );
HB1xp67_ASAP7_75t_L g375 ( .A(n_320), .Y(n_375) );
HB1xp67_ASAP7_75t_L g376 ( .A(n_320), .Y(n_376) );
NOR2x1p5_ASAP7_75t_L g377 ( .A(n_349), .B(n_312), .Y(n_377) );
BUFx3_ASAP7_75t_L g378 ( .A(n_325), .Y(n_378) );
AND2x2_ASAP7_75t_L g379 ( .A(n_339), .B(n_300), .Y(n_379) );
AND2x2_ASAP7_75t_L g380 ( .A(n_339), .B(n_300), .Y(n_380) );
OR2x2_ASAP7_75t_L g381 ( .A(n_357), .B(n_312), .Y(n_381) );
AND2x4_ASAP7_75t_SL g382 ( .A(n_376), .B(n_309), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_347), .B(n_306), .Y(n_383) );
AND2x2_ASAP7_75t_L g384 ( .A(n_361), .B(n_300), .Y(n_384) );
AND2x4_ASAP7_75t_SL g385 ( .A(n_375), .B(n_309), .Y(n_385) );
INVx2_ASAP7_75t_L g386 ( .A(n_324), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_357), .B(n_359), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_326), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_326), .Y(n_389) );
INVx2_ASAP7_75t_L g390 ( .A(n_324), .Y(n_390) );
INVx2_ASAP7_75t_L g391 ( .A(n_324), .Y(n_391) );
HB1xp67_ASAP7_75t_L g392 ( .A(n_334), .Y(n_392) );
INVx2_ASAP7_75t_L g393 ( .A(n_341), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_327), .Y(n_394) );
AND2x4_ASAP7_75t_L g395 ( .A(n_335), .B(n_296), .Y(n_395) );
OR2x2_ASAP7_75t_L g396 ( .A(n_359), .B(n_300), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_330), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_362), .B(n_303), .Y(n_398) );
INVx2_ASAP7_75t_L g399 ( .A(n_341), .Y(n_399) );
AND2x2_ASAP7_75t_L g400 ( .A(n_361), .B(n_300), .Y(n_400) );
OR2x2_ASAP7_75t_L g401 ( .A(n_362), .B(n_292), .Y(n_401) );
INVx2_ASAP7_75t_L g402 ( .A(n_341), .Y(n_402) );
INVx2_ASAP7_75t_L g403 ( .A(n_342), .Y(n_403) );
NOR2xp33_ASAP7_75t_L g404 ( .A(n_358), .B(n_2), .Y(n_404) );
NAND2x1p5_ASAP7_75t_L g405 ( .A(n_351), .B(n_319), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_331), .Y(n_406) );
AND2x2_ASAP7_75t_L g407 ( .A(n_364), .B(n_292), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_331), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_353), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_353), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_340), .B(n_303), .Y(n_411) );
AND2x2_ASAP7_75t_L g412 ( .A(n_364), .B(n_332), .Y(n_412) );
INVx2_ASAP7_75t_L g413 ( .A(n_342), .Y(n_413) );
AND2x2_ASAP7_75t_L g414 ( .A(n_332), .B(n_292), .Y(n_414) );
AND2x2_ASAP7_75t_L g415 ( .A(n_338), .B(n_292), .Y(n_415) );
AND2x4_ASAP7_75t_SL g416 ( .A(n_360), .B(n_319), .Y(n_416) );
INVx4_ASAP7_75t_L g417 ( .A(n_366), .Y(n_417) );
AND2x2_ASAP7_75t_L g418 ( .A(n_338), .B(n_296), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_354), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_356), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_356), .Y(n_421) );
AND2x2_ASAP7_75t_L g422 ( .A(n_346), .B(n_296), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_363), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_363), .Y(n_424) );
INVx2_ASAP7_75t_L g425 ( .A(n_342), .Y(n_425) );
AOI33xp33_ASAP7_75t_L g426 ( .A1(n_348), .A2(n_298), .A3(n_322), .B1(n_153), .B2(n_144), .B3(n_137), .Y(n_426) );
HB1xp67_ASAP7_75t_L g427 ( .A(n_329), .Y(n_427) );
AND2x2_ASAP7_75t_L g428 ( .A(n_352), .B(n_298), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_340), .B(n_352), .Y(n_429) );
OR2x2_ASAP7_75t_L g430 ( .A(n_337), .B(n_298), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_368), .Y(n_431) );
INVx2_ASAP7_75t_L g432 ( .A(n_344), .Y(n_432) );
AND3x1_ASAP7_75t_L g433 ( .A(n_323), .B(n_3), .C(n_5), .Y(n_433) );
AND2x2_ASAP7_75t_L g434 ( .A(n_369), .B(n_322), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_368), .Y(n_435) );
OR2x2_ASAP7_75t_L g436 ( .A(n_355), .B(n_303), .Y(n_436) );
AND2x2_ASAP7_75t_L g437 ( .A(n_369), .B(n_373), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_344), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_333), .B(n_322), .Y(n_439) );
BUFx2_ASAP7_75t_L g440 ( .A(n_367), .Y(n_440) );
AND2x2_ASAP7_75t_L g441 ( .A(n_373), .B(n_130), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_343), .Y(n_442) );
HB1xp67_ASAP7_75t_L g443 ( .A(n_372), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_323), .B(n_3), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_355), .B(n_5), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_343), .Y(n_446) );
AND2x2_ASAP7_75t_L g447 ( .A(n_344), .B(n_130), .Y(n_447) );
AND2x2_ASAP7_75t_L g448 ( .A(n_365), .B(n_130), .Y(n_448) );
INVx3_ASAP7_75t_L g449 ( .A(n_365), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_365), .Y(n_450) );
INVx2_ASAP7_75t_L g451 ( .A(n_449), .Y(n_451) );
NAND2x1_ASAP7_75t_L g452 ( .A(n_417), .B(n_367), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_392), .Y(n_453) );
NOR2xp33_ASAP7_75t_L g454 ( .A(n_378), .B(n_371), .Y(n_454) );
AND2x2_ASAP7_75t_L g455 ( .A(n_437), .B(n_335), .Y(n_455) );
INVx2_ASAP7_75t_L g456 ( .A(n_386), .Y(n_456) );
INVx2_ASAP7_75t_L g457 ( .A(n_386), .Y(n_457) );
HB1xp67_ASAP7_75t_L g458 ( .A(n_443), .Y(n_458) );
AND2x2_ASAP7_75t_L g459 ( .A(n_412), .B(n_370), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_412), .B(n_350), .Y(n_460) );
AND2x2_ASAP7_75t_L g461 ( .A(n_418), .B(n_366), .Y(n_461) );
AND2x2_ASAP7_75t_L g462 ( .A(n_418), .B(n_366), .Y(n_462) );
NOR2xp33_ASAP7_75t_L g463 ( .A(n_445), .B(n_366), .Y(n_463) );
AND2x2_ASAP7_75t_L g464 ( .A(n_379), .B(n_370), .Y(n_464) );
INVx2_ASAP7_75t_L g465 ( .A(n_390), .Y(n_465) );
OAI21xp33_ASAP7_75t_SL g466 ( .A1(n_377), .A2(n_366), .B(n_345), .Y(n_466) );
AND2x2_ASAP7_75t_L g467 ( .A(n_379), .B(n_370), .Y(n_467) );
OR2x2_ASAP7_75t_L g468 ( .A(n_427), .B(n_350), .Y(n_468) );
INVx2_ASAP7_75t_L g469 ( .A(n_390), .Y(n_469) );
AND2x2_ASAP7_75t_L g470 ( .A(n_380), .B(n_370), .Y(n_470) );
NOR2x1p5_ASAP7_75t_L g471 ( .A(n_417), .B(n_328), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_394), .Y(n_472) );
INVx2_ASAP7_75t_L g473 ( .A(n_391), .Y(n_473) );
AND2x2_ASAP7_75t_L g474 ( .A(n_380), .B(n_328), .Y(n_474) );
INVx2_ASAP7_75t_L g475 ( .A(n_391), .Y(n_475) );
INVx2_ASAP7_75t_L g476 ( .A(n_393), .Y(n_476) );
AND2x2_ASAP7_75t_L g477 ( .A(n_414), .B(n_328), .Y(n_477) );
AOI22xp5_ASAP7_75t_L g478 ( .A1(n_433), .A2(n_374), .B1(n_345), .B2(n_336), .Y(n_478) );
NAND2x1_ASAP7_75t_L g479 ( .A(n_417), .B(n_328), .Y(n_479) );
AND2x2_ASAP7_75t_L g480 ( .A(n_422), .B(n_336), .Y(n_480) );
AND2x2_ASAP7_75t_L g481 ( .A(n_422), .B(n_336), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_442), .B(n_336), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_406), .Y(n_483) );
NOR2xp33_ASAP7_75t_L g484 ( .A(n_404), .B(n_6), .Y(n_484) );
AND2x2_ASAP7_75t_L g485 ( .A(n_441), .B(n_374), .Y(n_485) );
NOR2xp33_ASAP7_75t_L g486 ( .A(n_444), .B(n_6), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_406), .Y(n_487) );
AND2x2_ASAP7_75t_L g488 ( .A(n_414), .B(n_374), .Y(n_488) );
AND2x2_ASAP7_75t_L g489 ( .A(n_415), .B(n_345), .Y(n_489) );
AND2x2_ASAP7_75t_L g490 ( .A(n_415), .B(n_345), .Y(n_490) );
NOR2xp33_ASAP7_75t_L g491 ( .A(n_387), .B(n_7), .Y(n_491) );
NAND2xp5_ASAP7_75t_SL g492 ( .A(n_426), .B(n_130), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_388), .Y(n_493) );
NAND2x1_ASAP7_75t_L g494 ( .A(n_440), .B(n_130), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_446), .B(n_7), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_429), .B(n_8), .Y(n_496) );
BUFx3_ASAP7_75t_L g497 ( .A(n_382), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_389), .Y(n_498) );
OAI21xp33_ASAP7_75t_L g499 ( .A1(n_407), .A2(n_130), .B(n_136), .Y(n_499) );
AND2x2_ASAP7_75t_L g500 ( .A(n_384), .B(n_400), .Y(n_500) );
NAND2x1p5_ASAP7_75t_L g501 ( .A(n_440), .B(n_276), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_397), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_408), .Y(n_503) );
HB1xp67_ASAP7_75t_L g504 ( .A(n_438), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_423), .Y(n_505) );
OR2x2_ASAP7_75t_L g506 ( .A(n_381), .B(n_8), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_409), .B(n_9), .Y(n_507) );
NAND2x1_ASAP7_75t_L g508 ( .A(n_395), .B(n_10), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_410), .B(n_10), .Y(n_509) );
AND2x4_ASAP7_75t_SL g510 ( .A(n_395), .B(n_11), .Y(n_510) );
AND2x2_ASAP7_75t_L g511 ( .A(n_384), .B(n_11), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_423), .Y(n_512) );
AND2x2_ASAP7_75t_L g513 ( .A(n_400), .B(n_12), .Y(n_513) );
INVx2_ASAP7_75t_L g514 ( .A(n_399), .Y(n_514) );
INVx1_ASAP7_75t_SL g515 ( .A(n_428), .Y(n_515) );
XNOR2xp5_ASAP7_75t_L g516 ( .A(n_407), .B(n_13), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_419), .B(n_14), .Y(n_517) );
AND2x2_ASAP7_75t_L g518 ( .A(n_434), .B(n_14), .Y(n_518) );
AND2x2_ASAP7_75t_L g519 ( .A(n_434), .B(n_16), .Y(n_519) );
INVx2_ASAP7_75t_L g520 ( .A(n_402), .Y(n_520) );
INVx2_ASAP7_75t_L g521 ( .A(n_402), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_420), .B(n_16), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_424), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_453), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_511), .B(n_431), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_458), .Y(n_526) );
AND2x2_ASAP7_75t_L g527 ( .A(n_500), .B(n_416), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_513), .B(n_431), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_458), .B(n_435), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_504), .B(n_435), .Y(n_530) );
OR2x2_ASAP7_75t_L g531 ( .A(n_515), .B(n_430), .Y(n_531) );
NOR2xp33_ASAP7_75t_L g532 ( .A(n_516), .B(n_383), .Y(n_532) );
AND2x2_ASAP7_75t_L g533 ( .A(n_455), .B(n_416), .Y(n_533) );
AND2x4_ASAP7_75t_L g534 ( .A(n_497), .B(n_382), .Y(n_534) );
HB1xp67_ASAP7_75t_L g535 ( .A(n_504), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_513), .B(n_436), .Y(n_536) );
AND2x2_ASAP7_75t_L g537 ( .A(n_455), .B(n_395), .Y(n_537) );
AND2x2_ASAP7_75t_L g538 ( .A(n_459), .B(n_385), .Y(n_538) );
NAND3xp33_ASAP7_75t_L g539 ( .A(n_491), .B(n_411), .C(n_398), .Y(n_539) );
OAI222xp33_ASAP7_75t_L g540 ( .A1(n_518), .A2(n_421), .B1(n_405), .B2(n_401), .C1(n_396), .C2(n_450), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_493), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_518), .B(n_428), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_519), .B(n_396), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_498), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_502), .Y(n_545) );
AND2x2_ASAP7_75t_L g546 ( .A(n_459), .B(n_385), .Y(n_546) );
INVx2_ASAP7_75t_L g547 ( .A(n_456), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_503), .Y(n_548) );
AOI21xp5_ASAP7_75t_L g549 ( .A1(n_494), .A2(n_405), .B(n_439), .Y(n_549) );
INVx1_ASAP7_75t_SL g550 ( .A(n_497), .Y(n_550) );
AND2x2_ASAP7_75t_L g551 ( .A(n_464), .B(n_438), .Y(n_551) );
AND2x2_ASAP7_75t_L g552 ( .A(n_464), .B(n_405), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_472), .B(n_447), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_483), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_487), .Y(n_555) );
OR2x2_ASAP7_75t_L g556 ( .A(n_460), .B(n_432), .Y(n_556) );
NAND2x1p5_ASAP7_75t_L g557 ( .A(n_508), .B(n_448), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_505), .B(n_448), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_512), .B(n_447), .Y(n_559) );
AND2x4_ASAP7_75t_L g560 ( .A(n_471), .B(n_425), .Y(n_560) );
NAND3xp33_ASAP7_75t_L g561 ( .A(n_491), .B(n_413), .C(n_403), .Y(n_561) );
AND2x2_ASAP7_75t_L g562 ( .A(n_467), .B(n_17), .Y(n_562) );
INVxp67_ASAP7_75t_L g563 ( .A(n_454), .Y(n_563) );
AND2x2_ASAP7_75t_L g564 ( .A(n_470), .B(n_17), .Y(n_564) );
AND2x2_ASAP7_75t_L g565 ( .A(n_461), .B(n_18), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_523), .B(n_18), .Y(n_566) );
HB1xp67_ASAP7_75t_L g567 ( .A(n_474), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_482), .Y(n_568) );
INVx2_ASAP7_75t_SL g569 ( .A(n_510), .Y(n_569) );
NAND2x1p5_ASAP7_75t_L g570 ( .A(n_452), .B(n_21), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_456), .B(n_22), .Y(n_571) );
OR2x2_ASAP7_75t_L g572 ( .A(n_477), .B(n_23), .Y(n_572) );
AND2x2_ASAP7_75t_L g573 ( .A(n_462), .B(n_25), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_457), .B(n_29), .Y(n_574) );
OR2x2_ASAP7_75t_L g575 ( .A(n_477), .B(n_31), .Y(n_575) );
INVx1_ASAP7_75t_SL g576 ( .A(n_510), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_506), .Y(n_577) );
AND2x4_ASAP7_75t_L g578 ( .A(n_488), .B(n_34), .Y(n_578) );
INVx2_ASAP7_75t_L g579 ( .A(n_535), .Y(n_579) );
NAND4xp75_ASAP7_75t_L g580 ( .A(n_569), .B(n_466), .C(n_484), .D(n_463), .Y(n_580) );
AOI221xp5_ASAP7_75t_SL g581 ( .A1(n_563), .A2(n_484), .B1(n_463), .B2(n_486), .C(n_495), .Y(n_581) );
OAI21xp5_ASAP7_75t_L g582 ( .A1(n_561), .A2(n_492), .B(n_454), .Y(n_582) );
AND3x1_ASAP7_75t_L g583 ( .A(n_532), .B(n_486), .C(n_478), .Y(n_583) );
INVx3_ASAP7_75t_L g584 ( .A(n_534), .Y(n_584) );
OAI21xp5_ASAP7_75t_SL g585 ( .A1(n_576), .A2(n_499), .B(n_496), .Y(n_585) );
AOI22xp33_ASAP7_75t_SL g586 ( .A1(n_576), .A2(n_489), .B1(n_490), .B2(n_481), .Y(n_586) );
AOI22xp5_ASAP7_75t_L g587 ( .A1(n_539), .A2(n_489), .B1(n_490), .B2(n_480), .Y(n_587) );
OAI22xp33_ASAP7_75t_L g588 ( .A1(n_550), .A2(n_479), .B1(n_468), .B2(n_501), .Y(n_588) );
INVx3_ASAP7_75t_L g589 ( .A(n_534), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_568), .B(n_465), .Y(n_590) );
OR2x2_ASAP7_75t_L g591 ( .A(n_531), .B(n_469), .Y(n_591) );
OAI21xp33_ASAP7_75t_SL g592 ( .A1(n_550), .A2(n_485), .B(n_521), .Y(n_592) );
OAI221xp5_ASAP7_75t_L g593 ( .A1(n_539), .A2(n_522), .B1(n_507), .B2(n_517), .C(n_509), .Y(n_593) );
INVxp67_ASAP7_75t_L g594 ( .A(n_524), .Y(n_594) );
AOI22xp5_ASAP7_75t_L g595 ( .A1(n_561), .A2(n_451), .B1(n_514), .B2(n_475), .Y(n_595) );
NOR2xp33_ASAP7_75t_L g596 ( .A(n_577), .B(n_520), .Y(n_596) );
AOI21xp33_ASAP7_75t_L g597 ( .A1(n_566), .A2(n_562), .B(n_564), .Y(n_597) );
INVx2_ASAP7_75t_L g598 ( .A(n_547), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_529), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_526), .B(n_520), .Y(n_600) );
OAI31xp33_ASAP7_75t_SL g601 ( .A1(n_527), .A2(n_476), .A3(n_475), .B(n_473), .Y(n_601) );
OR2x2_ASAP7_75t_L g602 ( .A(n_556), .B(n_469), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_529), .Y(n_603) );
INVxp67_ASAP7_75t_L g604 ( .A(n_541), .Y(n_604) );
NAND4xp25_ASAP7_75t_L g605 ( .A(n_565), .B(n_36), .C(n_38), .D(n_39), .Y(n_605) );
OAI21xp33_ASAP7_75t_L g606 ( .A1(n_567), .A2(n_41), .B(n_42), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_530), .Y(n_607) );
INVxp67_ASAP7_75t_L g608 ( .A(n_544), .Y(n_608) );
INVx1_ASAP7_75t_SL g609 ( .A(n_551), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_536), .B(n_43), .Y(n_610) );
AOI22xp33_ASAP7_75t_L g611 ( .A1(n_584), .A2(n_552), .B1(n_543), .B2(n_578), .Y(n_611) );
AOI22xp5_ASAP7_75t_L g612 ( .A1(n_583), .A2(n_525), .B1(n_528), .B2(n_542), .Y(n_612) );
INVxp67_ASAP7_75t_L g613 ( .A(n_596), .Y(n_613) );
OAI31xp33_ASAP7_75t_L g614 ( .A1(n_588), .A2(n_540), .A3(n_557), .B(n_570), .Y(n_614) );
AOI21xp5_ASAP7_75t_L g615 ( .A1(n_592), .A2(n_570), .B(n_549), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_599), .B(n_548), .Y(n_616) );
AOI221xp5_ASAP7_75t_SL g617 ( .A1(n_592), .A2(n_545), .B1(n_537), .B2(n_533), .C(n_538), .Y(n_617) );
NOR2xp33_ASAP7_75t_L g618 ( .A(n_584), .B(n_546), .Y(n_618) );
BUFx2_ASAP7_75t_L g619 ( .A(n_589), .Y(n_619) );
AOI221xp5_ASAP7_75t_L g620 ( .A1(n_581), .A2(n_597), .B1(n_594), .B2(n_604), .C(n_608), .Y(n_620) );
NAND4xp25_ASAP7_75t_SL g621 ( .A(n_586), .B(n_573), .C(n_575), .D(n_572), .Y(n_621) );
AOI211xp5_ASAP7_75t_L g622 ( .A1(n_585), .A2(n_582), .B(n_601), .C(n_605), .Y(n_622) );
AOI22xp5_ASAP7_75t_L g623 ( .A1(n_580), .A2(n_578), .B1(n_555), .B2(n_554), .Y(n_623) );
AOI21xp5_ASAP7_75t_L g624 ( .A1(n_606), .A2(n_560), .B(n_574), .Y(n_624) );
OAI211xp5_ASAP7_75t_L g625 ( .A1(n_587), .A2(n_559), .B(n_558), .C(n_553), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_603), .B(n_607), .Y(n_626) );
OAI22xp33_ASAP7_75t_L g627 ( .A1(n_609), .A2(n_571), .B1(n_45), .B2(n_46), .Y(n_627) );
AOI21x1_ASAP7_75t_L g628 ( .A1(n_579), .A2(n_600), .B(n_590), .Y(n_628) );
NAND4xp75_ASAP7_75t_L g629 ( .A(n_610), .B(n_595), .C(n_598), .D(n_591), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_602), .B(n_599), .Y(n_630) );
AOI221xp5_ASAP7_75t_L g631 ( .A1(n_583), .A2(n_581), .B1(n_593), .B2(n_592), .C(n_597), .Y(n_631) );
NAND4xp25_ASAP7_75t_L g632 ( .A(n_581), .B(n_576), .C(n_582), .D(n_484), .Y(n_632) );
NAND3xp33_ASAP7_75t_SL g633 ( .A(n_582), .B(n_550), .C(n_576), .Y(n_633) );
INVx1_ASAP7_75t_L g634 ( .A(n_626), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_616), .Y(n_635) );
NAND5xp2_ASAP7_75t_L g636 ( .A(n_614), .B(n_631), .C(n_622), .D(n_623), .E(n_617), .Y(n_636) );
NAND4xp25_ASAP7_75t_SL g637 ( .A(n_615), .B(n_620), .C(n_612), .D(n_611), .Y(n_637) );
OAI22xp5_ASAP7_75t_L g638 ( .A1(n_619), .A2(n_629), .B1(n_613), .B2(n_618), .Y(n_638) );
NOR2xp33_ASAP7_75t_L g639 ( .A(n_632), .B(n_633), .Y(n_639) );
INVx2_ASAP7_75t_L g640 ( .A(n_635), .Y(n_640) );
NOR2x1_ASAP7_75t_L g641 ( .A(n_636), .B(n_621), .Y(n_641) );
NAND2xp5_ASAP7_75t_SL g642 ( .A(n_638), .B(n_628), .Y(n_642) );
AND2x2_ASAP7_75t_L g643 ( .A(n_639), .B(n_630), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_640), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_643), .B(n_634), .Y(n_645) );
AND2x2_ASAP7_75t_L g646 ( .A(n_641), .B(n_625), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_646), .B(n_642), .Y(n_647) );
AOI21x1_ASAP7_75t_L g648 ( .A1(n_646), .A2(n_637), .B(n_624), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_647), .Y(n_649) );
INVx3_ASAP7_75t_L g650 ( .A(n_648), .Y(n_650) );
AOI21xp33_ASAP7_75t_L g651 ( .A1(n_649), .A2(n_650), .B(n_644), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_651), .Y(n_652) );
OAI21xp5_ASAP7_75t_L g653 ( .A1(n_652), .A2(n_649), .B(n_650), .Y(n_653) );
AOI21xp5_ASAP7_75t_SL g654 ( .A1(n_653), .A2(n_645), .B(n_650), .Y(n_654) );
AOI21xp33_ASAP7_75t_SL g655 ( .A1(n_654), .A2(n_650), .B(n_627), .Y(n_655) );
endmodule