module fake_jpeg_28636_n_118 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_118);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_118;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_32),
.B(n_8),
.Y(n_39)
);

CKINVDCx14_ASAP7_75t_R g40 ( 
.A(n_26),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_14),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

OR2x2_ASAP7_75t_L g43 ( 
.A(n_21),
.B(n_10),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_22),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_6),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_10),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_2),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_44),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_51),
.A2(n_58),
.B1(n_53),
.B2(n_49),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_38),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_52)
);

O2A1O1Ixp33_ASAP7_75t_L g61 ( 
.A1(n_52),
.A2(n_50),
.B(n_49),
.C(n_48),
.Y(n_61)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_53),
.Y(n_62)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_47),
.Y(n_54)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_54),
.Y(n_63)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_47),
.Y(n_55)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_55),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_43),
.B(n_3),
.Y(n_56)
);

OR2x2_ASAP7_75t_L g70 ( 
.A(n_56),
.B(n_4),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_38),
.B(n_18),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_57),
.B(n_39),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_42),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_56),
.B(n_43),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_59),
.B(n_66),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_61),
.A2(n_54),
.B1(n_46),
.B2(n_45),
.Y(n_80)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_55),
.Y(n_64)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_64),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_65),
.A2(n_51),
.B1(n_58),
.B2(n_53),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_57),
.B(n_50),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_55),
.Y(n_67)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_67),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_57),
.B(n_41),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_68),
.B(n_71),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_69),
.B(n_7),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_70),
.B(n_5),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_52),
.B(n_41),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_72),
.A2(n_17),
.B(n_19),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_67),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_73),
.B(n_76),
.Y(n_86)
);

A2O1A1O1Ixp25_ASAP7_75t_L g74 ( 
.A1(n_69),
.A2(n_40),
.B(n_45),
.C(n_42),
.D(n_46),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_SL g94 ( 
.A(n_74),
.B(n_15),
.C(n_16),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_63),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_77),
.B(n_12),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_80),
.B(n_29),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g81 ( 
.A(n_61),
.B(n_54),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_L g90 ( 
.A(n_81),
.B(n_62),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_60),
.A2(n_54),
.B1(n_8),
.B2(n_9),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_83),
.A2(n_63),
.B1(n_9),
.B2(n_11),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_84),
.B(n_85),
.Y(n_91)
);

HB1xp67_ASAP7_75t_L g85 ( 
.A(n_60),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_87),
.A2(n_96),
.B1(n_99),
.B2(n_74),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_SL g88 ( 
.A1(n_78),
.A2(n_70),
.B(n_11),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_88),
.B(n_89),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_84),
.B(n_7),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_90),
.B(n_98),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_92),
.B(n_97),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_75),
.B(n_12),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_93),
.B(n_95),
.Y(n_107)
);

XNOR2x2_ASAP7_75t_L g105 ( 
.A(n_94),
.B(n_98),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_81),
.B(n_62),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_76),
.A2(n_20),
.B(n_23),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_73),
.A2(n_25),
.B(n_28),
.Y(n_98)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_86),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_101),
.B(n_102),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_105),
.Y(n_110)
);

FAx1_ASAP7_75t_L g106 ( 
.A(n_90),
.B(n_82),
.CI(n_79),
.CON(n_106),
.SN(n_106)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_106),
.B(n_91),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_109),
.B(n_111),
.C(n_107),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_100),
.A2(n_87),
.B1(n_33),
.B2(n_34),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_108),
.A2(n_100),
.B(n_103),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_112),
.A2(n_113),
.B(n_104),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_114),
.B(n_109),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_115),
.Y(n_116)
);

AOI321xp33_ASAP7_75t_L g117 ( 
.A1(n_116),
.A2(n_110),
.A3(n_106),
.B1(n_111),
.B2(n_35),
.C(n_30),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_117),
.B(n_37),
.Y(n_118)
);


endmodule