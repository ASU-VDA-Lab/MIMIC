module fake_jpeg_13831_n_56 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_56);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_56;

wire n_13;
wire n_21;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_44;
wire n_26;
wire n_38;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

NAND2xp5_ASAP7_75t_SL g8 ( 
.A(n_0),
.B(n_1),
.Y(n_8)
);

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_0),
.Y(n_9)
);

INVx3_ASAP7_75t_L g10 ( 
.A(n_7),
.Y(n_10)
);

CKINVDCx14_ASAP7_75t_R g11 ( 
.A(n_0),
.Y(n_11)
);

INVx11_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_2),
.Y(n_13)
);

INVx5_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

INVx3_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVx8_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_SL g18 ( 
.A1(n_11),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_18)
);

OAI21xp5_ASAP7_75t_L g25 ( 
.A1(n_18),
.A2(n_20),
.B(n_21),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_8),
.B(n_4),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_19),
.B(n_6),
.Y(n_26)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_8),
.A2(n_2),
.B(n_5),
.Y(n_20)
);

AO22x1_ASAP7_75t_L g21 ( 
.A1(n_12),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_22),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_20),
.B(n_16),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g31 ( 
.A(n_23),
.B(n_16),
.C(n_15),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_26),
.B(n_27),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_21),
.B(n_13),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_22),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_29),
.B(n_17),
.Y(n_37)
);

OA21x2_ASAP7_75t_L g30 ( 
.A1(n_23),
.A2(n_18),
.B(n_21),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_30),
.B(n_31),
.Y(n_42)
);

HB1xp67_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

HB1xp67_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

OAI22xp33_ASAP7_75t_L g34 ( 
.A1(n_24),
.A2(n_22),
.B1(n_16),
.B2(n_15),
.Y(n_34)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

INVx1_ASAP7_75t_SL g35 ( 
.A(n_28),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_35),
.Y(n_40)
);

NOR2x1_ASAP7_75t_L g36 ( 
.A(n_25),
.B(n_12),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_36),
.B(n_37),
.C(n_25),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_41),
.A2(n_36),
.B1(n_30),
.B2(n_10),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_10),
.C(n_15),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_43),
.B(n_10),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_44),
.B(n_45),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_42),
.A2(n_39),
.B1(n_34),
.B2(n_40),
.Y(n_46)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_46),
.Y(n_48)
);

INVxp33_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_47),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_48),
.A2(n_47),
.B1(n_42),
.B2(n_35),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_51),
.B(n_52),
.C(n_50),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_48),
.B(n_28),
.C(n_13),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_53),
.B(n_49),
.Y(n_54)
);

AOI31xp33_ASAP7_75t_L g55 ( 
.A1(n_54),
.A2(n_11),
.A3(n_14),
.B(n_9),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_55),
.A2(n_9),
.B1(n_14),
.B2(n_27),
.Y(n_56)
);


endmodule