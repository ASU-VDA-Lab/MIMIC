module fake_jpeg_8910_n_341 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_341);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_341;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_11),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx12_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx8_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

INVx1_ASAP7_75t_SL g34 ( 
.A(n_5),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_34),
.B(n_0),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_36),
.B(n_48),
.Y(n_69)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

BUFx4f_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

INVx1_ASAP7_75t_SL g38 ( 
.A(n_21),
.Y(n_38)
);

INVx2_ASAP7_75t_SL g75 ( 
.A(n_38),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g39 ( 
.A1(n_27),
.A2(n_14),
.B(n_13),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_39),
.B(n_43),
.Y(n_65)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_40),
.Y(n_72)
);

BUFx12_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_16),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_21),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_45),
.B(n_47),
.Y(n_58)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_24),
.Y(n_46)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_21),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_21),
.Y(n_49)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_49),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_46),
.Y(n_50)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_50),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_53),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_42),
.A2(n_34),
.B1(n_16),
.B2(n_23),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_54),
.A2(n_57),
.B1(n_60),
.B2(n_61),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_55),
.Y(n_96)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_56),
.B(n_62),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_37),
.A2(n_24),
.B1(n_33),
.B2(n_19),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_40),
.A2(n_33),
.B1(n_19),
.B2(n_20),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_39),
.A2(n_16),
.B1(n_23),
.B2(n_20),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_38),
.A2(n_33),
.B1(n_20),
.B2(n_22),
.Y(n_64)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_64),
.A2(n_68),
.B(n_70),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_48),
.A2(n_22),
.B1(n_17),
.B2(n_29),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_66),
.A2(n_32),
.B1(n_31),
.B2(n_18),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_49),
.A2(n_22),
.B1(n_17),
.B2(n_29),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_49),
.A2(n_25),
.B1(n_26),
.B2(n_28),
.Y(n_70)
);

BUFx16f_ASAP7_75t_L g71 ( 
.A(n_41),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g112 ( 
.A(n_71),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_74),
.Y(n_79)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_41),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_76),
.B(n_41),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_36),
.B(n_28),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_77),
.B(n_25),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_71),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_78),
.B(n_80),
.Y(n_123)
);

OR2x2_ASAP7_75t_L g80 ( 
.A(n_65),
.B(n_43),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_77),
.B(n_13),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_81),
.B(n_82),
.Y(n_143)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_58),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_73),
.A2(n_28),
.B1(n_26),
.B2(n_25),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_83),
.A2(n_104),
.B1(n_75),
.B2(n_32),
.Y(n_131)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_58),
.Y(n_84)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_84),
.Y(n_119)
);

BUFx12_ASAP7_75t_L g85 ( 
.A(n_71),
.Y(n_85)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_85),
.Y(n_124)
);

OAI22xp33_ASAP7_75t_L g87 ( 
.A1(n_73),
.A2(n_45),
.B1(n_35),
.B2(n_31),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_87),
.A2(n_110),
.B1(n_67),
.B2(n_52),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_90),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_66),
.B(n_18),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_91),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_51),
.B(n_18),
.Y(n_92)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_92),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_65),
.B(n_31),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_94),
.B(n_95),
.Y(n_125)
);

BUFx24_ASAP7_75t_L g97 ( 
.A(n_59),
.Y(n_97)
);

CKINVDCx5p33_ASAP7_75t_R g144 ( 
.A(n_97),
.Y(n_144)
);

AND2x4_ASAP7_75t_L g98 ( 
.A(n_69),
.B(n_32),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_98),
.A2(n_32),
.B(n_30),
.Y(n_146)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_72),
.Y(n_99)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_99),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_51),
.B(n_18),
.Y(n_100)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_100),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_69),
.B(n_26),
.Y(n_101)
);

AOI21xp33_ASAP7_75t_L g137 ( 
.A1(n_101),
.A2(n_114),
.B(n_95),
.Y(n_137)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_60),
.Y(n_102)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_102),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_72),
.A2(n_10),
.B1(n_12),
.B2(n_14),
.Y(n_104)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_59),
.Y(n_105)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_105),
.Y(n_136)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_57),
.Y(n_106)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_106),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_53),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_107),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_108),
.A2(n_32),
.B1(n_35),
.B2(n_18),
.Y(n_138)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_69),
.Y(n_109)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_109),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_56),
.A2(n_35),
.B1(n_21),
.B2(n_30),
.Y(n_110)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_59),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_111),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_74),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_113),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_62),
.B(n_52),
.Y(n_114)
);

BUFx12f_ASAP7_75t_L g115 ( 
.A(n_76),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_115),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_116),
.A2(n_126),
.B1(n_130),
.B2(n_139),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_106),
.A2(n_67),
.B1(n_75),
.B2(n_63),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_103),
.A2(n_63),
.B1(n_75),
.B2(n_55),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_128),
.A2(n_131),
.B1(n_138),
.B2(n_99),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_109),
.A2(n_98),
.B1(n_101),
.B2(n_88),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_103),
.A2(n_41),
.B(n_18),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_132),
.A2(n_137),
.B(n_146),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_98),
.A2(n_50),
.B1(n_35),
.B2(n_30),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_114),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_142),
.B(n_145),
.Y(n_170)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_89),
.Y(n_145)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_126),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_148),
.B(n_149),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_144),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_125),
.B(n_94),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_150),
.B(n_158),
.C(n_172),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_130),
.A2(n_88),
.B1(n_108),
.B2(n_98),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_151),
.A2(n_157),
.B1(n_169),
.B2(n_124),
.Y(n_211)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_116),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_153),
.B(n_154),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_144),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_139),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_155),
.B(n_162),
.Y(n_203)
);

OAI21xp33_ASAP7_75t_SL g184 ( 
.A1(n_156),
.A2(n_118),
.B(n_120),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_134),
.A2(n_80),
.B1(n_111),
.B2(n_105),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_125),
.B(n_110),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_146),
.B(n_141),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_159),
.A2(n_121),
.B(n_120),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_140),
.A2(n_93),
.B1(n_87),
.B2(n_96),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_160),
.A2(n_166),
.B1(n_180),
.B2(n_118),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_142),
.B(n_79),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_161),
.B(n_167),
.Y(n_191)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_123),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_140),
.A2(n_132),
.B1(n_135),
.B2(n_134),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_163),
.A2(n_133),
.B1(n_122),
.B2(n_145),
.Y(n_181)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_129),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_164),
.B(n_165),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_144),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_135),
.A2(n_93),
.B1(n_96),
.B2(n_86),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_123),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_128),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_168),
.B(n_171),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_141),
.A2(n_86),
.B1(n_97),
.B2(n_107),
.Y(n_169)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_143),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_137),
.B(n_97),
.C(n_112),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_129),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_173),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_131),
.A2(n_117),
.B(n_133),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_174),
.A2(n_127),
.B(n_112),
.Y(n_198)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_143),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_175),
.B(n_177),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_119),
.B(n_112),
.Y(n_176)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_176),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_119),
.B(n_79),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_121),
.B(n_115),
.Y(n_178)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_178),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_138),
.Y(n_179)
);

HB1xp67_ASAP7_75t_L g188 ( 
.A(n_179),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_122),
.A2(n_30),
.B1(n_21),
.B2(n_115),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_181),
.B(n_197),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_150),
.B(n_152),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_183),
.B(n_190),
.C(n_214),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_184),
.A2(n_211),
.B1(n_160),
.B2(n_180),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_L g219 ( 
.A1(n_186),
.A2(n_155),
.B1(n_167),
.B2(n_162),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_187),
.A2(n_192),
.B(n_198),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_152),
.B(n_85),
.Y(n_190)
);

OA21x2_ASAP7_75t_L g192 ( 
.A1(n_168),
.A2(n_136),
.B(n_30),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_161),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_195),
.B(n_199),
.Y(n_218)
);

AO22x1_ASAP7_75t_L g196 ( 
.A1(n_153),
.A2(n_124),
.B1(n_30),
.B2(n_136),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_196),
.B(n_0),
.Y(n_234)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_177),
.Y(n_197)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_164),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_174),
.A2(n_127),
.B(n_1),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_200),
.A2(n_207),
.B(n_210),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_170),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_202),
.B(n_212),
.Y(n_220)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_166),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_204),
.B(n_206),
.Y(n_237)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_169),
.Y(n_206)
);

OA21x2_ASAP7_75t_L g207 ( 
.A1(n_148),
.A2(n_0),
.B(n_1),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_158),
.B(n_172),
.Y(n_209)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_209),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_179),
.A2(n_85),
.B(n_124),
.Y(n_210)
);

INVx2_ASAP7_75t_SL g212 ( 
.A(n_173),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_151),
.B(n_11),
.Y(n_214)
);

NAND3xp33_ASAP7_75t_L g216 ( 
.A(n_208),
.B(n_157),
.C(n_175),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_216),
.B(n_225),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_183),
.B(n_147),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_217),
.B(n_226),
.C(n_229),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_219),
.A2(n_224),
.B1(n_186),
.B2(n_204),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_208),
.Y(n_221)
);

OR2x2_ASAP7_75t_L g256 ( 
.A(n_221),
.B(n_228),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_205),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_213),
.B(n_147),
.C(n_159),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_191),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_213),
.B(n_159),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_203),
.B(n_171),
.Y(n_231)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_231),
.Y(n_247)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_191),
.Y(n_232)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_232),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_211),
.A2(n_165),
.B1(n_154),
.B2(n_149),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_233),
.A2(n_242),
.B1(n_207),
.B2(n_212),
.Y(n_252)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_234),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_189),
.B(n_11),
.Y(n_235)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_235),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_201),
.B(n_10),
.Y(n_236)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_236),
.Y(n_264)
);

OR2x2_ASAP7_75t_L g238 ( 
.A(n_193),
.B(n_1),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g260 ( 
.A1(n_238),
.A2(n_234),
.B(n_231),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_209),
.B(n_2),
.C(n_3),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_239),
.B(n_196),
.C(n_3),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_193),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_240),
.A2(n_197),
.B1(n_182),
.B2(n_207),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_194),
.B(n_10),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_241),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_206),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_242)
);

CKINVDCx14_ASAP7_75t_R g266 ( 
.A(n_243),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_227),
.A2(n_185),
.B1(n_200),
.B2(n_182),
.Y(n_244)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_244),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_246),
.B(n_259),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_226),
.B(n_229),
.C(n_230),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_249),
.B(n_250),
.C(n_251),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_230),
.B(n_190),
.C(n_198),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_223),
.B(n_214),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_252),
.A2(n_240),
.B1(n_228),
.B2(n_225),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_217),
.B(n_187),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_254),
.B(n_257),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_223),
.B(n_210),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_232),
.B(n_192),
.C(n_188),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_258),
.B(n_239),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_220),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_L g274 ( 
.A1(n_260),
.A2(n_238),
.B(n_221),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_237),
.A2(n_192),
.B1(n_196),
.B2(n_199),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_261),
.A2(n_2),
.B1(n_6),
.B2(n_7),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g276 ( 
.A(n_263),
.B(n_238),
.Y(n_276)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_261),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_268),
.B(n_272),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_245),
.B(n_212),
.Y(n_269)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_269),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_255),
.A2(n_227),
.B1(n_237),
.B2(n_224),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_270),
.A2(n_278),
.B1(n_281),
.B2(n_265),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_271),
.B(n_276),
.Y(n_288)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_255),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_SL g273 ( 
.A1(n_252),
.A2(n_215),
.B(n_233),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_273),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_SL g297 ( 
.A(n_274),
.B(n_283),
.Y(n_297)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_256),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_279),
.A2(n_282),
.B1(n_246),
.B2(n_263),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_256),
.B(n_218),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_280),
.B(n_264),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_258),
.A2(n_215),
.B(n_222),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_265),
.A2(n_222),
.B1(n_242),
.B2(n_7),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_249),
.B(n_6),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_284),
.B(n_262),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_277),
.B(n_248),
.C(n_275),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_286),
.B(n_291),
.Y(n_305)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_287),
.Y(n_304)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_290),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_277),
.B(n_248),
.C(n_257),
.Y(n_291)
);

INVx13_ASAP7_75t_L g292 ( 
.A(n_280),
.Y(n_292)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_292),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_275),
.B(n_250),
.C(n_254),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_293),
.B(n_295),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_284),
.B(n_251),
.C(n_253),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_271),
.B(n_260),
.C(n_247),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_298),
.B(n_301),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_299),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_300),
.B(n_278),
.Y(n_302)
);

INVx13_ASAP7_75t_L g301 ( 
.A(n_272),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_302),
.B(n_306),
.Y(n_318)
);

AOI21x1_ASAP7_75t_SL g303 ( 
.A1(n_297),
.A2(n_273),
.B(n_268),
.Y(n_303)
);

AND2x2_ASAP7_75t_L g322 ( 
.A(n_303),
.B(n_309),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_293),
.B(n_281),
.Y(n_306)
);

NOR2xp67_ASAP7_75t_SL g309 ( 
.A(n_294),
.B(n_267),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_300),
.B(n_296),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_310),
.A2(n_313),
.B(n_290),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_296),
.B(n_274),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_L g315 ( 
.A1(n_307),
.A2(n_285),
.B1(n_266),
.B2(n_292),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_315),
.B(n_319),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_303),
.A2(n_304),
.B1(n_312),
.B2(n_308),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_316),
.B(n_320),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_305),
.B(n_286),
.C(n_291),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_317),
.B(n_314),
.C(n_306),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_SL g319 ( 
.A(n_311),
.B(n_288),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_310),
.B(n_289),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_302),
.B(n_301),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_321),
.A2(n_297),
.B1(n_283),
.B2(n_282),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_323),
.A2(n_288),
.B1(n_295),
.B2(n_299),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_322),
.A2(n_313),
.B1(n_279),
.B2(n_298),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_324),
.B(n_328),
.Y(n_334)
);

AND2x2_ASAP7_75t_L g333 ( 
.A(n_326),
.B(n_330),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_329),
.B(n_318),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_317),
.B(n_6),
.C(n_7),
.Y(n_330)
);

AOI21xp5_ASAP7_75t_SL g331 ( 
.A1(n_327),
.A2(n_322),
.B(n_318),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_L g336 ( 
.A1(n_331),
.A2(n_332),
.B(n_329),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_334),
.B(n_326),
.C(n_325),
.Y(n_335)
);

O2A1O1Ixp33_ASAP7_75t_SL g337 ( 
.A1(n_335),
.A2(n_336),
.B(n_333),
.C(n_330),
.Y(n_337)
);

NOR2xp67_ASAP7_75t_SL g338 ( 
.A(n_337),
.B(n_6),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_338),
.B(n_8),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_L g340 ( 
.A1(n_339),
.A2(n_8),
.B(n_9),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_SL g341 ( 
.A1(n_340),
.A2(n_9),
.B(n_334),
.Y(n_341)
);


endmodule