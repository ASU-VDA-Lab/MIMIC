module fake_jpeg_25085_n_328 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_328);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_328;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_12),
.Y(n_17)
);

BUFx2_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_0),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_0),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_4),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_9),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

INVx3_ASAP7_75t_SL g56 ( 
.A(n_35),
.Y(n_56)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_36),
.B(n_30),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_25),
.B(n_15),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_37),
.B(n_40),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_25),
.B(n_15),
.Y(n_40)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx1_ASAP7_75t_SL g72 ( 
.A(n_46),
.Y(n_72)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

BUFx2_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_53),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_55),
.B(n_57),
.Y(n_66)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_58),
.Y(n_83)
);

INVx2_ASAP7_75t_SL g59 ( 
.A(n_39),
.Y(n_59)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_59),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_60),
.Y(n_64)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_61),
.Y(n_90)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_63),
.Y(n_78)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_65),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_54),
.B(n_40),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_70),
.B(n_81),
.Y(n_101)
);

OR2x2_ASAP7_75t_L g71 ( 
.A(n_54),
.B(n_38),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_71),
.B(n_79),
.Y(n_102)
);

OAI21xp33_ASAP7_75t_L g73 ( 
.A1(n_47),
.A2(n_37),
.B(n_25),
.Y(n_73)
);

XOR2x1_ASAP7_75t_SL g93 ( 
.A(n_73),
.B(n_18),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_62),
.A2(n_42),
.B1(n_36),
.B2(n_30),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_74),
.A2(n_76),
.B1(n_88),
.B2(n_56),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_47),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_75),
.B(n_59),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_62),
.A2(n_41),
.B1(n_44),
.B2(n_19),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_52),
.B(n_38),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_77),
.B(n_91),
.C(n_63),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_53),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_49),
.A2(n_41),
.B1(n_26),
.B2(n_34),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_80),
.A2(n_56),
.B1(n_50),
.B2(n_61),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_52),
.B(n_44),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_60),
.B(n_44),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_82),
.B(n_84),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_51),
.B(n_38),
.Y(n_84)
);

BUFx4f_ASAP7_75t_L g85 ( 
.A(n_49),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_85),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_48),
.Y(n_86)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_86),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_51),
.A2(n_22),
.B1(n_32),
.B2(n_19),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_48),
.B(n_38),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_89),
.B(n_46),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_45),
.B(n_38),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_93),
.B(n_100),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_70),
.B(n_19),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_95),
.B(n_96),
.Y(n_120)
);

FAx1_ASAP7_75t_SL g96 ( 
.A(n_71),
.B(n_43),
.CI(n_18),
.CON(n_96),
.SN(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_67),
.Y(n_97)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_97),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_71),
.A2(n_0),
.B(n_1),
.Y(n_98)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_98),
.Y(n_138)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_81),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_99),
.B(n_110),
.Y(n_137)
);

OAI22x1_ASAP7_75t_L g103 ( 
.A1(n_77),
.A2(n_31),
.B1(n_26),
.B2(n_18),
.Y(n_103)
);

AOI22x1_ASAP7_75t_SL g121 ( 
.A1(n_103),
.A2(n_85),
.B1(n_31),
.B2(n_64),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_105),
.B(n_115),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_106),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_107),
.A2(n_68),
.B1(n_83),
.B2(n_79),
.Y(n_128)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_83),
.Y(n_108)
);

INVxp33_ASAP7_75t_SL g146 ( 
.A(n_108),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_84),
.B(n_26),
.C(n_58),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_109),
.B(n_90),
.C(n_64),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_66),
.B(n_17),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_111),
.B(n_112),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_82),
.B(n_22),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_77),
.A2(n_0),
.B(n_1),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_113),
.B(n_117),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_76),
.A2(n_32),
.B1(n_22),
.B2(n_34),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_114),
.A2(n_88),
.B1(n_27),
.B2(n_29),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_74),
.B(n_89),
.Y(n_115)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_91),
.Y(n_117)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_67),
.Y(n_118)
);

HB1xp67_ASAP7_75t_L g136 ( 
.A(n_118),
.Y(n_136)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_91),
.Y(n_119)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_119),
.Y(n_122)
);

OAI21xp33_ASAP7_75t_SL g156 ( 
.A1(n_121),
.A2(n_148),
.B(n_108),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_93),
.A2(n_103),
.B1(n_100),
.B2(n_115),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_123),
.A2(n_126),
.B1(n_144),
.B2(n_20),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_124),
.B(n_119),
.Y(n_150)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_111),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_125),
.B(n_139),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_128),
.A2(n_132),
.B1(n_134),
.B2(n_114),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_115),
.A2(n_90),
.B1(n_68),
.B2(n_87),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_130),
.A2(n_133),
.B1(n_142),
.B2(n_116),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_104),
.A2(n_78),
.B1(n_69),
.B2(n_87),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_99),
.A2(n_72),
.B1(n_78),
.B2(n_69),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_101),
.A2(n_72),
.B1(n_21),
.B2(n_17),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_101),
.B(n_104),
.C(n_105),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_135),
.B(n_147),
.C(n_95),
.Y(n_152)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_112),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_102),
.A2(n_85),
.B1(n_32),
.B2(n_23),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_L g144 ( 
.A1(n_98),
.A2(n_21),
.B1(n_65),
.B2(n_33),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_109),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_145),
.B(n_124),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_102),
.B(n_86),
.C(n_28),
.Y(n_147)
);

NAND2xp33_ASAP7_75t_SL g148 ( 
.A(n_96),
.B(n_31),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_133),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_149),
.A2(n_160),
.B(n_161),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_150),
.B(n_162),
.C(n_152),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_152),
.B(n_153),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_127),
.A2(n_117),
.B(n_116),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_154),
.A2(n_167),
.B(n_173),
.Y(n_203)
);

INVxp33_ASAP7_75t_SL g155 ( 
.A(n_146),
.Y(n_155)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_155),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_156),
.A2(n_157),
.B1(n_165),
.B2(n_168),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_136),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_158),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_159),
.Y(n_205)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_132),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_130),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_135),
.B(n_96),
.C(n_113),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_141),
.B(n_110),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_SL g195 ( 
.A(n_163),
.B(n_171),
.Y(n_195)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_140),
.Y(n_164)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_164),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_140),
.B(n_97),
.Y(n_166)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_166),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_121),
.A2(n_92),
.B1(n_94),
.B2(n_118),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_137),
.A2(n_27),
.B1(n_29),
.B2(n_33),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_125),
.B(n_92),
.Y(n_169)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_169),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_137),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_170),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_141),
.B(n_24),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_129),
.Y(n_172)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_172),
.Y(n_200)
);

OAI21xp33_ASAP7_75t_SL g173 ( 
.A1(n_138),
.A2(n_20),
.B(n_28),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_129),
.Y(n_174)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_174),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_139),
.B(n_23),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g199 ( 
.A(n_175),
.Y(n_199)
);

INVxp33_ASAP7_75t_L g176 ( 
.A(n_143),
.Y(n_176)
);

INVx1_ASAP7_75t_SL g196 ( 
.A(n_176),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_127),
.A2(n_94),
.B1(n_24),
.B2(n_9),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_177),
.A2(n_120),
.B1(n_122),
.B2(n_145),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_120),
.B(n_24),
.Y(n_178)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_178),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_147),
.Y(n_179)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_179),
.Y(n_209)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_142),
.Y(n_180)
);

OA21x2_ASAP7_75t_L g187 ( 
.A1(n_180),
.A2(n_149),
.B(n_161),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_126),
.A2(n_15),
.B1(n_14),
.B2(n_13),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_181),
.A2(n_131),
.B1(n_148),
.B2(n_14),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_182),
.B(n_210),
.C(n_151),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_186),
.A2(n_189),
.B1(n_191),
.B2(n_180),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_187),
.B(n_169),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_160),
.A2(n_127),
.B1(n_122),
.B2(n_131),
.Y(n_188)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_188),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_153),
.A2(n_131),
.B(n_2),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_190),
.A2(n_1),
.B(n_3),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_157),
.A2(n_14),
.B1(n_13),
.B2(n_11),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_150),
.B(n_13),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_194),
.B(n_207),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_162),
.B(n_11),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_171),
.B(n_10),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_208),
.B(n_211),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_164),
.B(n_10),
.C(n_2),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_154),
.B(n_10),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_198),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_212),
.B(n_218),
.Y(n_239)
);

OAI21xp33_ASAP7_75t_L g213 ( 
.A1(n_190),
.A2(n_170),
.B(n_177),
.Y(n_213)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_213),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_SL g214 ( 
.A(n_195),
.B(n_163),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_214),
.B(n_217),
.Y(n_240)
);

AOI21xp33_ASAP7_75t_L g215 ( 
.A1(n_203),
.A2(n_179),
.B(n_151),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_215),
.A2(n_216),
.B1(n_226),
.B2(n_227),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_195),
.B(n_178),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_204),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_219),
.B(n_235),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_SL g220 ( 
.A(n_208),
.B(n_166),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_220),
.B(n_186),
.Y(n_251)
);

HB1xp67_ASAP7_75t_L g221 ( 
.A(n_202),
.Y(n_221)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_221),
.Y(n_247)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_222),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_199),
.B(n_159),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_225),
.B(n_230),
.Y(n_243)
);

AOI22x1_ASAP7_75t_L g226 ( 
.A1(n_205),
.A2(n_158),
.B1(n_3),
.B2(n_4),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_182),
.B(n_1),
.C(n_3),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_228),
.B(n_189),
.C(n_211),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_203),
.A2(n_3),
.B(n_4),
.Y(n_229)
);

CKINVDCx16_ASAP7_75t_R g249 ( 
.A(n_229),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_192),
.B(n_5),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_183),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_231),
.B(n_232),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_193),
.B(n_5),
.Y(n_232)
);

INVx3_ASAP7_75t_SL g233 ( 
.A(n_196),
.Y(n_233)
);

INVx1_ASAP7_75t_SL g255 ( 
.A(n_233),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_210),
.B(n_5),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_200),
.Y(n_236)
);

BUFx3_ASAP7_75t_L g242 ( 
.A(n_236),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_207),
.B(n_6),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_237),
.B(n_191),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_238),
.B(n_257),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_219),
.B(n_185),
.C(n_209),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_245),
.B(n_246),
.C(n_248),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_220),
.B(n_185),
.C(n_209),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_223),
.B(n_188),
.C(n_194),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_251),
.B(n_224),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_223),
.B(n_197),
.C(n_206),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_254),
.B(n_256),
.C(n_258),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_217),
.B(n_187),
.C(n_183),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_224),
.B(n_187),
.C(n_201),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_SL g279 ( 
.A(n_259),
.B(n_248),
.Y(n_279)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_239),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_260),
.B(n_261),
.Y(n_280)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_242),
.Y(n_261)
);

INVxp67_ASAP7_75t_SL g262 ( 
.A(n_244),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_262),
.B(n_265),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_240),
.B(n_214),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_263),
.B(n_271),
.Y(n_281)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_243),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_246),
.B(n_234),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_268),
.B(n_269),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_245),
.B(n_234),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_242),
.B(n_230),
.Y(n_270)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_270),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_240),
.B(n_222),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_254),
.B(n_258),
.C(n_251),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_272),
.B(n_249),
.C(n_227),
.Y(n_290)
);

CKINVDCx16_ASAP7_75t_R g273 ( 
.A(n_250),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_273),
.Y(n_277)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_255),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_274),
.B(n_275),
.Y(n_287)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_255),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_264),
.B(n_247),
.C(n_256),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_276),
.B(n_284),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_266),
.A2(n_241),
.B(n_231),
.Y(n_278)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_278),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_279),
.B(n_286),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_264),
.B(n_238),
.C(n_253),
.Y(n_284)
);

AND2x2_ASAP7_75t_L g285 ( 
.A(n_271),
.B(n_226),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g302 ( 
.A1(n_285),
.A2(n_196),
.B(n_283),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_259),
.B(n_252),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_263),
.B(n_228),
.Y(n_288)
);

AND2x2_ASAP7_75t_L g301 ( 
.A(n_288),
.B(n_232),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_SL g296 ( 
.A(n_290),
.B(n_268),
.Y(n_296)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_280),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_292),
.B(n_298),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_277),
.B(n_287),
.Y(n_293)
);

OR2x2_ASAP7_75t_L g307 ( 
.A(n_293),
.B(n_294),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_285),
.A2(n_205),
.B1(n_233),
.B2(n_269),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_282),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_295),
.B(n_297),
.Y(n_311)
);

AND2x2_ASAP7_75t_L g305 ( 
.A(n_296),
.B(n_288),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_289),
.A2(n_184),
.B1(n_226),
.B2(n_267),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_290),
.A2(n_267),
.B1(n_272),
.B2(n_229),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_301),
.B(n_279),
.C(n_8),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_302),
.B(n_281),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_286),
.B(n_6),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_303),
.B(n_6),
.Y(n_304)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_304),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_305),
.B(n_306),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_297),
.B(n_281),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_308),
.B(n_309),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_299),
.B(n_8),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_SL g314 ( 
.A(n_310),
.B(n_291),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_314),
.B(n_315),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_SL g315 ( 
.A(n_307),
.B(n_298),
.Y(n_315)
);

NOR2xp67_ASAP7_75t_SL g316 ( 
.A(n_312),
.B(n_300),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_316),
.B(n_300),
.Y(n_322)
);

OAI21x1_ASAP7_75t_L g317 ( 
.A1(n_306),
.A2(n_301),
.B(n_294),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_317),
.B(n_311),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_321),
.B(n_322),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_323),
.B(n_320),
.C(n_313),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_SL g325 ( 
.A1(n_324),
.A2(n_319),
.B(n_318),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_325),
.B(n_321),
.Y(n_326)
);

BUFx24_ASAP7_75t_SL g327 ( 
.A(n_326),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_327),
.B(n_304),
.C(n_8),
.Y(n_328)
);


endmodule