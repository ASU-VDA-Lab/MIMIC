module fake_jpeg_4620_n_228 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_228);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_228;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_152;
wire n_73;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_127;
wire n_76;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVxp67_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_4),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

INVx13_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

INVx5_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_23),
.B(n_0),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_32),
.B(n_35),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_17),
.B(n_0),
.Y(n_34)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_34),
.Y(n_64)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_24),
.B(n_1),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_37),
.B(n_39),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_24),
.B(n_1),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

BUFx16f_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

BUFx4f_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_41),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_17),
.Y(n_42)
);

CKINVDCx12_ASAP7_75t_R g53 ( 
.A(n_42),
.Y(n_53)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_45),
.B(n_57),
.Y(n_78)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_46),
.A2(n_28),
.B1(n_24),
.B2(n_16),
.Y(n_71)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_50),
.B(n_61),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_35),
.A2(n_31),
.B1(n_18),
.B2(n_19),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_51),
.A2(n_52),
.B1(n_60),
.B2(n_28),
.Y(n_80)
);

OA22x2_ASAP7_75t_L g52 ( 
.A1(n_32),
.A2(n_31),
.B1(n_29),
.B2(n_27),
.Y(n_52)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_56),
.Y(n_69)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

BUFx16f_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_58),
.Y(n_76)
);

OAI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_35),
.A2(n_31),
.B1(n_18),
.B2(n_19),
.Y(n_60)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_33),
.Y(n_61)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_62),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_63),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_44),
.B(n_32),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_65),
.B(n_30),
.Y(n_99)
);

INVx13_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_66),
.B(n_80),
.Y(n_94)
);

AND2x4_ASAP7_75t_SL g67 ( 
.A(n_52),
.B(n_36),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_67),
.A2(n_77),
.B(n_79),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_53),
.B(n_42),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_68),
.B(n_82),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_52),
.A2(n_15),
.B1(n_22),
.B2(n_26),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_70),
.A2(n_75),
.B1(n_84),
.B2(n_21),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_71),
.A2(n_48),
.B1(n_3),
.B2(n_4),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_59),
.B(n_16),
.C(n_25),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_72),
.B(n_20),
.Y(n_87)
);

OA22x2_ASAP7_75t_L g75 ( 
.A1(n_58),
.A2(n_49),
.B1(n_60),
.B2(n_51),
.Y(n_75)
);

NAND2xp33_ASAP7_75t_SL g77 ( 
.A(n_59),
.B(n_26),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_SL g79 ( 
.A1(n_64),
.A2(n_39),
.B(n_37),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_43),
.B(n_22),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_54),
.B(n_28),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_83),
.B(n_29),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_54),
.A2(n_21),
.B1(n_25),
.B2(n_48),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_78),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_86),
.B(n_91),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_87),
.B(n_95),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_88),
.B(n_89),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_SL g89 ( 
.A(n_65),
.B(n_20),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_78),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_92),
.B(n_93),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_68),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_67),
.B(n_20),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_83),
.B(n_47),
.Y(n_96)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_96),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_97),
.B(n_101),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_99),
.B(n_100),
.Y(n_124)
);

NAND3xp33_ASAP7_75t_L g100 ( 
.A(n_77),
.B(n_30),
.C(n_3),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_85),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_85),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_102),
.B(n_81),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_82),
.B(n_29),
.Y(n_103)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_103),
.Y(n_118)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_74),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_104),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_67),
.B(n_30),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_105),
.B(n_75),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_79),
.B(n_82),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_106),
.B(n_108),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_74),
.Y(n_107)
);

INVxp33_ASAP7_75t_L g126 ( 
.A(n_107),
.Y(n_126)
);

NOR3xp33_ASAP7_75t_L g108 ( 
.A(n_75),
.B(n_2),
.C(n_5),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_99),
.B(n_106),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_110),
.B(n_114),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_94),
.A2(n_75),
.B1(n_67),
.B2(n_70),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_112),
.A2(n_117),
.B1(n_127),
.B2(n_130),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_98),
.B(n_86),
.Y(n_114)
);

CKINVDCx14_ASAP7_75t_R g115 ( 
.A(n_97),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_115),
.B(n_119),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_98),
.A2(n_75),
.B1(n_81),
.B2(n_74),
.Y(n_117)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_107),
.Y(n_119)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_107),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_123),
.B(n_129),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_125),
.B(n_93),
.Y(n_136)
);

INVx13_ASAP7_75t_L g129 ( 
.A(n_102),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_88),
.A2(n_72),
.B1(n_63),
.B2(n_56),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_120),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_131),
.B(n_134),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_110),
.B(n_92),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_133),
.B(n_144),
.Y(n_155)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_125),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_136),
.B(n_138),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_121),
.A2(n_105),
.B1(n_95),
.B2(n_90),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_137),
.A2(n_149),
.B1(n_118),
.B2(n_124),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_111),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_116),
.B(n_90),
.Y(n_141)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_141),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_128),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_142),
.B(n_143),
.Y(n_160)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_117),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_114),
.B(n_121),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_130),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_145),
.B(n_146),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_121),
.B(n_109),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_118),
.A2(n_95),
.B1(n_105),
.B2(n_89),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_147),
.A2(n_76),
.B(n_27),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_SL g148 ( 
.A(n_109),
.B(n_87),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_148),
.B(n_29),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_112),
.A2(n_87),
.B1(n_104),
.B2(n_76),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_116),
.B(n_122),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_150),
.B(n_151),
.Y(n_168)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_127),
.Y(n_151)
);

OAI21xp33_ASAP7_75t_L g152 ( 
.A1(n_144),
.A2(n_122),
.B(n_129),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_152),
.B(n_159),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_153),
.A2(n_154),
.B(n_164),
.Y(n_176)
);

NOR3xp33_ASAP7_75t_L g154 ( 
.A(n_131),
.B(n_124),
.C(n_129),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_157),
.B(n_149),
.C(n_150),
.Y(n_175)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_139),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_161),
.B(n_140),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_143),
.A2(n_123),
.B1(n_119),
.B2(n_126),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_162),
.A2(n_165),
.B1(n_169),
.B2(n_134),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_151),
.A2(n_113),
.B(n_6),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_163),
.B(n_133),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_132),
.A2(n_113),
.B(n_66),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_145),
.A2(n_113),
.B1(n_73),
.B2(n_69),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_146),
.A2(n_73),
.B1(n_69),
.B2(n_8),
.Y(n_169)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_170),
.Y(n_196)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_166),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_172),
.B(n_173),
.Y(n_187)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_155),
.Y(n_173)
);

CKINVDCx14_ASAP7_75t_R g190 ( 
.A(n_174),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_175),
.B(n_184),
.C(n_167),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_157),
.B(n_132),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_177),
.B(n_180),
.Y(n_186)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_155),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_178),
.B(n_179),
.Y(n_188)
);

BUFx12_ASAP7_75t_L g179 ( 
.A(n_161),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_156),
.B(n_148),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_L g181 ( 
.A1(n_163),
.A2(n_142),
.B1(n_135),
.B2(n_138),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_181),
.A2(n_162),
.B(n_169),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_156),
.B(n_135),
.C(n_137),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_182),
.B(n_164),
.C(n_159),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_183),
.B(n_168),
.Y(n_185)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_160),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_185),
.B(n_193),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_189),
.B(n_191),
.C(n_192),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_175),
.B(n_153),
.C(n_168),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_182),
.B(n_147),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_194),
.A2(n_177),
.B(n_179),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_SL g195 ( 
.A(n_171),
.B(n_165),
.Y(n_195)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_195),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_189),
.A2(n_176),
.B(n_158),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_199),
.B(n_200),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_196),
.B(n_183),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_191),
.A2(n_171),
.B(n_180),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_201),
.B(n_202),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_187),
.B(n_179),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_203),
.B(n_204),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_190),
.A2(n_195),
.B1(n_193),
.B2(n_188),
.Y(n_204)
);

AOI31xp67_ASAP7_75t_L g206 ( 
.A1(n_204),
.A2(n_186),
.A3(n_6),
.B(n_8),
.Y(n_206)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_206),
.Y(n_214)
);

AOI322xp5_ASAP7_75t_L g207 ( 
.A1(n_197),
.A2(n_186),
.A3(n_73),
.B1(n_69),
.B2(n_66),
.C1(n_11),
.C2(n_5),
.Y(n_207)
);

AOI21xp33_ASAP7_75t_L g215 ( 
.A1(n_207),
.A2(n_9),
.B(n_10),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_205),
.B(n_8),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_210),
.B(n_211),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_205),
.B(n_9),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_208),
.B(n_201),
.C(n_198),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_213),
.B(n_215),
.Y(n_221)
);

A2O1A1O1Ixp25_ASAP7_75t_L g217 ( 
.A1(n_209),
.A2(n_9),
.B(n_10),
.C(n_11),
.D(n_12),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_217),
.B(n_13),
.Y(n_220)
);

NOR3xp33_ASAP7_75t_SL g218 ( 
.A(n_206),
.B(n_11),
.C(n_12),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_218),
.B(n_216),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_214),
.A2(n_212),
.B1(n_12),
.B2(n_13),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_219),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_220),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_222),
.B(n_217),
.C(n_221),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g226 ( 
.A(n_223),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_225),
.A2(n_224),
.B(n_220),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_227),
.B(n_226),
.Y(n_228)
);


endmodule