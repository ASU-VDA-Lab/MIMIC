module fake_jpeg_29943_n_379 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_379);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_379;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_377;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

HB1xp67_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

INVx13_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

BUFx24_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_11),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_11),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_12),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx16f_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_0),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_40),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_24),
.B(n_8),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_41),
.B(n_62),
.Y(n_73)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

BUFx2_ASAP7_75t_L g83 ( 
.A(n_42),
.Y(n_83)
);

BUFx24_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

INVx5_ASAP7_75t_SL g76 ( 
.A(n_43),
.Y(n_76)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_44),
.Y(n_96)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_45),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_46),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_47),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g112 ( 
.A(n_48),
.Y(n_112)
);

INVx3_ASAP7_75t_SL g49 ( 
.A(n_33),
.Y(n_49)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_49),
.Y(n_71)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_27),
.Y(n_50)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_50),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_51),
.Y(n_79)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_23),
.Y(n_52)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_52),
.Y(n_72)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_23),
.Y(n_53)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_53),
.Y(n_92)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_27),
.Y(n_54)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_54),
.Y(n_93)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_22),
.Y(n_55)
);

INVx13_ASAP7_75t_L g105 ( 
.A(n_55),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_19),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g108 ( 
.A(n_56),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_57),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_58),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_19),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_59),
.A2(n_26),
.B1(n_32),
.B2(n_33),
.Y(n_85)
);

HB1xp67_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_60),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_19),
.Y(n_61)
);

CKINVDCx14_ASAP7_75t_R g84 ( 
.A(n_61),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_18),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_63),
.B(n_64),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_18),
.Y(n_64)
);

AOI21xp33_ASAP7_75t_L g65 ( 
.A1(n_31),
.A2(n_8),
.B(n_15),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_65),
.B(n_67),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_21),
.B(n_16),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_66),
.B(n_68),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_18),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_21),
.B(n_16),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_24),
.B(n_15),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_69),
.B(n_25),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_40),
.A2(n_21),
.B1(n_28),
.B2(n_17),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_70),
.A2(n_87),
.B1(n_90),
.B2(n_95),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_69),
.B(n_37),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_74),
.B(n_77),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_41),
.B(n_37),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_46),
.B(n_29),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_81),
.B(n_94),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_85),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_49),
.A2(n_17),
.B1(n_23),
.B2(n_22),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_86),
.A2(n_102),
.B1(n_20),
.B2(n_32),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_47),
.A2(n_31),
.B1(n_38),
.B2(n_28),
.Y(n_87)
);

BUFx12_ASAP7_75t_L g89 ( 
.A(n_43),
.Y(n_89)
);

INVx4_ASAP7_75t_SL g122 ( 
.A(n_89),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_48),
.A2(n_28),
.B1(n_31),
.B2(n_29),
.Y(n_90)
);

CKINVDCx12_ASAP7_75t_R g91 ( 
.A(n_62),
.Y(n_91)
);

CKINVDCx14_ASAP7_75t_R g152 ( 
.A(n_91),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_60),
.B(n_30),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_51),
.A2(n_36),
.B1(n_22),
.B2(n_30),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_100),
.B(n_106),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_57),
.B(n_25),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_101),
.B(n_104),
.Y(n_130)
);

OAI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_58),
.A2(n_33),
.B1(n_36),
.B2(n_34),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_63),
.A2(n_38),
.B1(n_34),
.B2(n_33),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_103),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_64),
.B(n_38),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_67),
.B(n_12),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_41),
.B(n_34),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_111),
.B(n_16),
.Y(n_138)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_104),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_113),
.Y(n_187)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_72),
.Y(n_114)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_114),
.Y(n_170)
);

INVxp33_ASAP7_75t_L g115 ( 
.A(n_76),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_115),
.Y(n_156)
);

OA22x2_ASAP7_75t_L g116 ( 
.A1(n_87),
.A2(n_20),
.B1(n_32),
.B2(n_26),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_116),
.A2(n_120),
.B1(n_143),
.B2(n_83),
.Y(n_154)
);

BUFx12f_ASAP7_75t_L g118 ( 
.A(n_89),
.Y(n_118)
);

BUFx8_ASAP7_75t_L g185 ( 
.A(n_118),
.Y(n_185)
);

AO22x1_ASAP7_75t_SL g120 ( 
.A1(n_80),
.A2(n_20),
.B1(n_32),
.B2(n_26),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_72),
.Y(n_121)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_121),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_76),
.A2(n_36),
.B1(n_32),
.B2(n_26),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_123),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_88),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_124),
.Y(n_184)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_92),
.Y(n_125)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_125),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_126),
.A2(n_79),
.B1(n_108),
.B2(n_5),
.Y(n_175)
);

INVx2_ASAP7_75t_SL g127 ( 
.A(n_97),
.Y(n_127)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_127),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_89),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_128),
.B(n_129),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_71),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_78),
.B(n_32),
.C(n_20),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_131),
.B(n_141),
.C(n_144),
.Y(n_157)
);

BUFx2_ASAP7_75t_L g132 ( 
.A(n_112),
.Y(n_132)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_132),
.Y(n_180)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_92),
.Y(n_136)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_136),
.Y(n_189)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_81),
.B(n_101),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_137),
.B(n_139),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_138),
.B(n_148),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_73),
.B(n_71),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_74),
.B(n_0),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_140),
.B(n_142),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_110),
.B(n_20),
.C(n_15),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_77),
.B(n_0),
.Y(n_142)
);

OA22x2_ASAP7_75t_L g143 ( 
.A1(n_95),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_110),
.B(n_14),
.C(n_13),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_145),
.A2(n_146),
.B1(n_4),
.B2(n_6),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_82),
.A2(n_14),
.B1(n_10),
.B2(n_9),
.Y(n_146)
);

BUFx3_ASAP7_75t_L g147 ( 
.A(n_96),
.Y(n_147)
);

INVx6_ASAP7_75t_L g166 ( 
.A(n_147),
.Y(n_166)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_112),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_75),
.B(n_2),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_149),
.B(n_3),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_105),
.B(n_9),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_150),
.B(n_151),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_83),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_93),
.A2(n_9),
.B1(n_4),
.B2(n_5),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_153),
.A2(n_98),
.B1(n_82),
.B2(n_93),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g201 ( 
.A(n_154),
.B(n_155),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_SL g155 ( 
.A(n_120),
.B(n_96),
.C(n_84),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_158),
.A2(n_145),
.B1(n_127),
.B2(n_148),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_130),
.B(n_105),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_159),
.B(n_160),
.C(n_165),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_130),
.B(n_131),
.C(n_137),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_134),
.A2(n_97),
.B(n_109),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_161),
.A2(n_155),
.B(n_186),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_147),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_163),
.B(n_176),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_137),
.A2(n_98),
.B1(n_88),
.B2(n_109),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_164),
.A2(n_182),
.B1(n_122),
.B2(n_127),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_139),
.B(n_107),
.C(n_99),
.Y(n_165)
);

AND2x2_ASAP7_75t_SL g168 ( 
.A(n_120),
.B(n_107),
.Y(n_168)
);

CKINVDCx14_ASAP7_75t_R g205 ( 
.A(n_168),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_117),
.A2(n_99),
.B1(n_79),
.B2(n_108),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_172),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_175),
.A2(n_190),
.B1(n_128),
.B2(n_122),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_139),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_177),
.B(n_144),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_140),
.B(n_142),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_179),
.B(n_167),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_117),
.A2(n_79),
.B1(n_108),
.B2(n_6),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_132),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_183),
.B(n_115),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_119),
.A2(n_4),
.B(n_5),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_186),
.A2(n_149),
.B(n_141),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_192),
.Y(n_246)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_162),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_193),
.B(n_195),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_194),
.B(n_196),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_167),
.B(n_133),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_179),
.B(n_119),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_197),
.B(n_200),
.Y(n_241)
);

AND2x2_ASAP7_75t_L g257 ( 
.A(n_198),
.B(n_212),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_173),
.B(n_135),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_199),
.B(n_203),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_159),
.B(n_143),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_202),
.B(n_211),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_171),
.B(n_152),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_170),
.Y(n_204)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_204),
.Y(n_228)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_181),
.Y(n_206)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_206),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_207),
.A2(n_209),
.B1(n_215),
.B2(n_175),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_160),
.B(n_143),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g212 ( 
.A(n_154),
.B(n_116),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g213 ( 
.A(n_171),
.B(n_116),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_213),
.B(n_223),
.Y(n_253)
);

BUFx12f_ASAP7_75t_L g214 ( 
.A(n_184),
.Y(n_214)
);

BUFx10_ASAP7_75t_L g231 ( 
.A(n_214),
.Y(n_231)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_181),
.Y(n_216)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_216),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_169),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_217),
.B(n_219),
.Y(n_259)
);

NAND3xp33_ASAP7_75t_L g218 ( 
.A(n_178),
.B(n_136),
.C(n_114),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_218),
.B(n_220),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_177),
.B(n_143),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_180),
.Y(n_220)
);

INVx8_ASAP7_75t_L g221 ( 
.A(n_166),
.Y(n_221)
);

INVx6_ASAP7_75t_L g255 ( 
.A(n_221),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_187),
.B(n_118),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_222),
.B(n_224),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_157),
.B(n_116),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_161),
.B(n_118),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_157),
.B(n_7),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_225),
.B(n_185),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_188),
.A2(n_79),
.B(n_108),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_226),
.B(n_227),
.C(n_168),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_SL g227 ( 
.A(n_165),
.B(n_7),
.Y(n_227)
);

INVx2_ASAP7_75t_SL g232 ( 
.A(n_214),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_232),
.B(n_249),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_234),
.A2(n_235),
.B1(n_240),
.B2(n_251),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_197),
.A2(n_207),
.B1(n_219),
.B2(n_212),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_237),
.B(n_239),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_208),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_212),
.A2(n_168),
.B1(n_190),
.B2(n_188),
.Y(n_240)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_206),
.Y(n_243)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_243),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_204),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_244),
.B(n_247),
.Y(n_281)
);

CKINVDCx12_ASAP7_75t_R g245 ( 
.A(n_193),
.Y(n_245)
);

CKINVDCx16_ASAP7_75t_R g282 ( 
.A(n_245),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_225),
.B(n_174),
.Y(n_247)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_216),
.Y(n_250)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_250),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_223),
.A2(n_182),
.B1(n_156),
.B2(n_174),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_195),
.B(n_169),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_254),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_210),
.B(n_189),
.C(n_156),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_256),
.B(n_227),
.C(n_203),
.Y(n_272)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_221),
.Y(n_258)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_258),
.Y(n_271)
);

BUFx10_ASAP7_75t_L g260 ( 
.A(n_214),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_260),
.B(n_231),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_251),
.A2(n_201),
.B1(n_215),
.B2(n_213),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_262),
.A2(n_267),
.B1(n_246),
.B2(n_241),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_239),
.A2(n_201),
.B1(n_191),
.B2(n_200),
.Y(n_263)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_263),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_253),
.B(n_210),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_266),
.B(n_269),
.C(n_272),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_257),
.A2(n_201),
.B1(n_213),
.B2(n_205),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_257),
.A2(n_191),
.B1(n_198),
.B2(n_226),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_268),
.A2(n_275),
.B1(n_249),
.B2(n_246),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_253),
.B(n_211),
.Y(n_269)
);

INVx1_ASAP7_75t_SL g294 ( 
.A(n_274),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_236),
.A2(n_209),
.B1(n_196),
.B2(n_194),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_238),
.Y(n_276)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_276),
.Y(n_293)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_238),
.Y(n_277)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_277),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_252),
.B(n_202),
.Y(n_278)
);

XOR2x2_ASAP7_75t_L g289 ( 
.A(n_278),
.B(n_279),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_252),
.B(n_217),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_241),
.A2(n_220),
.B1(n_166),
.B2(n_184),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_280),
.A2(n_255),
.B1(n_242),
.B2(n_250),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_230),
.B(n_189),
.Y(n_283)
);

FAx1_ASAP7_75t_SL g296 ( 
.A(n_283),
.B(n_230),
.CI(n_248),
.CON(n_296),
.SN(n_296)
);

OAI21xp5_ASAP7_75t_L g285 ( 
.A1(n_257),
.A2(n_185),
.B(n_180),
.Y(n_285)
);

A2O1A1O1Ixp25_ASAP7_75t_L g287 ( 
.A1(n_285),
.A2(n_233),
.B(n_229),
.C(n_258),
.D(n_259),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_256),
.B(n_170),
.C(n_124),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_286),
.B(n_232),
.Y(n_302)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_287),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_274),
.Y(n_288)
);

OR2x2_ASAP7_75t_L g326 ( 
.A(n_288),
.B(n_305),
.Y(n_326)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_282),
.Y(n_290)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_290),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_291),
.A2(n_299),
.B1(n_277),
.B2(n_265),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_SL g310 ( 
.A(n_292),
.B(n_261),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_295),
.A2(n_303),
.B1(n_271),
.B2(n_276),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_296),
.B(n_269),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_284),
.A2(n_242),
.B1(n_243),
.B2(n_255),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_281),
.B(n_244),
.Y(n_301)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_301),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_302),
.B(n_286),
.C(n_301),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_280),
.A2(n_232),
.B1(n_228),
.B2(n_231),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_264),
.Y(n_304)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_304),
.Y(n_322)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_264),
.Y(n_305)
);

XOR2x1_ASAP7_75t_SL g306 ( 
.A(n_268),
.B(n_231),
.Y(n_306)
);

XNOR2x1_ASAP7_75t_SL g316 ( 
.A(n_306),
.B(n_285),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_273),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g325 ( 
.A1(n_307),
.A2(n_308),
.B1(n_271),
.B2(n_228),
.Y(n_325)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_265),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_SL g332 ( 
.A(n_309),
.B(n_323),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_310),
.B(n_313),
.C(n_314),
.Y(n_328)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_311),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_298),
.B(n_266),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_298),
.B(n_270),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_300),
.A2(n_261),
.B1(n_283),
.B2(n_279),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_315),
.A2(n_320),
.B1(n_306),
.B2(n_310),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_SL g331 ( 
.A1(n_316),
.A2(n_294),
.B(n_287),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_292),
.B(n_270),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_317),
.B(n_319),
.C(n_321),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_289),
.B(n_278),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_289),
.B(n_267),
.Y(n_321)
);

FAx1_ASAP7_75t_SL g323 ( 
.A(n_296),
.B(n_272),
.CI(n_262),
.CON(n_323),
.SN(n_323)
);

OAI22xp5_ASAP7_75t_L g335 ( 
.A1(n_324),
.A2(n_295),
.B1(n_303),
.B2(n_294),
.Y(n_335)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_325),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_327),
.B(n_296),
.C(n_308),
.Y(n_336)
);

XOR2xp5_ASAP7_75t_L g353 ( 
.A(n_329),
.B(n_315),
.Y(n_353)
);

AOI21xp5_ASAP7_75t_L g347 ( 
.A1(n_331),
.A2(n_342),
.B(n_316),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_326),
.Y(n_334)
);

NOR3xp33_ASAP7_75t_L g343 ( 
.A(n_334),
.B(n_340),
.C(n_297),
.Y(n_343)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_335),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_336),
.B(n_339),
.C(n_317),
.Y(n_344)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_326),
.Y(n_338)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_338),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_314),
.B(n_305),
.C(n_304),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_318),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_322),
.Y(n_341)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_341),
.Y(n_351)
);

OAI21xp5_ASAP7_75t_SL g342 ( 
.A1(n_312),
.A2(n_293),
.B(n_297),
.Y(n_342)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_343),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_SL g355 ( 
.A(n_344),
.B(n_349),
.Y(n_355)
);

BUFx24_ASAP7_75t_SL g346 ( 
.A(n_332),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_346),
.B(n_328),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_347),
.B(n_342),
.Y(n_358)
);

AOI21xp5_ASAP7_75t_L g349 ( 
.A1(n_331),
.A2(n_327),
.B(n_309),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_328),
.B(n_313),
.C(n_323),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g361 ( 
.A(n_350),
.B(n_352),
.Y(n_361)
);

NOR2xp67_ASAP7_75t_SL g352 ( 
.A(n_336),
.B(n_321),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_353),
.A2(n_329),
.B1(n_337),
.B2(n_333),
.Y(n_354)
);

INVxp67_ASAP7_75t_L g363 ( 
.A(n_354),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_348),
.A2(n_337),
.B1(n_333),
.B2(n_338),
.Y(n_356)
);

INVxp67_ASAP7_75t_L g368 ( 
.A(n_356),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_357),
.B(n_358),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_345),
.B(n_339),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_360),
.B(n_362),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_348),
.B(n_290),
.Y(n_362)
);

OAI221xp5_ASAP7_75t_L g364 ( 
.A1(n_359),
.A2(n_355),
.B1(n_361),
.B2(n_356),
.C(n_351),
.Y(n_364)
);

CKINVDCx16_ASAP7_75t_R g370 ( 
.A(n_364),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_354),
.B(n_353),
.C(n_330),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_366),
.B(n_369),
.Y(n_371)
);

NAND3xp33_ASAP7_75t_L g369 ( 
.A(n_359),
.B(n_341),
.C(n_293),
.Y(n_369)
);

AND2x2_ASAP7_75t_L g372 ( 
.A(n_367),
.B(n_330),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_SL g374 ( 
.A(n_372),
.B(n_373),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_365),
.B(n_214),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_371),
.B(n_363),
.C(n_368),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_375),
.B(n_370),
.C(n_319),
.Y(n_376)
);

HB1xp67_ASAP7_75t_L g377 ( 
.A(n_376),
.Y(n_377)
);

AOI21xp5_ASAP7_75t_L g378 ( 
.A1(n_377),
.A2(n_374),
.B(n_231),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_378),
.B(n_260),
.C(n_185),
.Y(n_379)
);


endmodule