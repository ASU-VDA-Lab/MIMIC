module fake_netlist_1_12371_n_520 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_73, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_71, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_74, n_72, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_520);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_73;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_71;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_74;
input n_72;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_520;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_206;
wire n_288;
wire n_383;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_211;
wire n_334;
wire n_389;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_476;
wire n_105;
wire n_227;
wire n_384;
wire n_434;
wire n_231;
wire n_452;
wire n_518;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_119;
wire n_141;
wire n_517;
wire n_479;
wire n_97;
wire n_167;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_502;
wire n_312;
wire n_455;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_482;
wire n_394;
wire n_415;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_133;
wire n_149;
wire n_81;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_516;
wire n_254;
wire n_262;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_98;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_420;
wire n_342;
wire n_423;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_245;
wire n_357;
wire n_90;
wire n_260;
wire n_78;
wire n_201;
wire n_197;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_265;
wire n_264;
wire n_208;
wire n_200;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_75;
wire n_376;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_121;
wire n_497;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_335;
wire n_272;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_418;
wire n_493;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_494;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_99;
wire n_109;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g75 ( .A(n_30), .Y(n_75) );
INVx1_ASAP7_75t_L g76 ( .A(n_1), .Y(n_76) );
CKINVDCx20_ASAP7_75t_R g77 ( .A(n_11), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_25), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_9), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_43), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_6), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_7), .Y(n_82) );
CKINVDCx16_ASAP7_75t_R g83 ( .A(n_19), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_0), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_12), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_22), .Y(n_86) );
BUFx2_ASAP7_75t_L g87 ( .A(n_31), .Y(n_87) );
INVxp33_ASAP7_75t_SL g88 ( .A(n_72), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_26), .Y(n_89) );
CKINVDCx5p33_ASAP7_75t_R g90 ( .A(n_18), .Y(n_90) );
CKINVDCx5p33_ASAP7_75t_R g91 ( .A(n_38), .Y(n_91) );
CKINVDCx20_ASAP7_75t_R g92 ( .A(n_14), .Y(n_92) );
CKINVDCx14_ASAP7_75t_R g93 ( .A(n_9), .Y(n_93) );
CKINVDCx20_ASAP7_75t_R g94 ( .A(n_46), .Y(n_94) );
CKINVDCx20_ASAP7_75t_R g95 ( .A(n_52), .Y(n_95) );
INVxp67_ASAP7_75t_SL g96 ( .A(n_34), .Y(n_96) );
INVxp67_ASAP7_75t_L g97 ( .A(n_2), .Y(n_97) );
INVxp33_ASAP7_75t_SL g98 ( .A(n_18), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_67), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_59), .Y(n_100) );
INVxp33_ASAP7_75t_L g101 ( .A(n_41), .Y(n_101) );
CKINVDCx16_ASAP7_75t_R g102 ( .A(n_24), .Y(n_102) );
CKINVDCx14_ASAP7_75t_R g103 ( .A(n_56), .Y(n_103) );
BUFx6f_ASAP7_75t_L g104 ( .A(n_3), .Y(n_104) );
INVxp33_ASAP7_75t_L g105 ( .A(n_57), .Y(n_105) );
CKINVDCx20_ASAP7_75t_R g106 ( .A(n_48), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_29), .Y(n_107) );
INVxp33_ASAP7_75t_L g108 ( .A(n_47), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_10), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_7), .Y(n_110) );
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_23), .Y(n_111) );
CKINVDCx20_ASAP7_75t_R g112 ( .A(n_1), .Y(n_112) );
INVxp33_ASAP7_75t_L g113 ( .A(n_16), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_44), .Y(n_114) );
INVx3_ASAP7_75t_L g115 ( .A(n_104), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_75), .Y(n_116) );
INVx2_ASAP7_75t_L g117 ( .A(n_75), .Y(n_117) );
OAI22xp5_ASAP7_75t_SL g118 ( .A1(n_77), .A2(n_0), .B1(n_2), .B2(n_3), .Y(n_118) );
INVx2_ASAP7_75t_L g119 ( .A(n_80), .Y(n_119) );
INVxp67_ASAP7_75t_L g120 ( .A(n_87), .Y(n_120) );
BUFx2_ASAP7_75t_L g121 ( .A(n_87), .Y(n_121) );
INVx3_ASAP7_75t_L g122 ( .A(n_104), .Y(n_122) );
BUFx6f_ASAP7_75t_L g123 ( .A(n_104), .Y(n_123) );
BUFx6f_ASAP7_75t_L g124 ( .A(n_104), .Y(n_124) );
INVx2_ASAP7_75t_L g125 ( .A(n_80), .Y(n_125) );
BUFx6f_ASAP7_75t_L g126 ( .A(n_104), .Y(n_126) );
AND2x2_ASAP7_75t_L g127 ( .A(n_113), .B(n_4), .Y(n_127) );
NAND2xp5_ASAP7_75t_L g128 ( .A(n_81), .B(n_4), .Y(n_128) );
INVx2_ASAP7_75t_L g129 ( .A(n_86), .Y(n_129) );
BUFx6f_ASAP7_75t_L g130 ( .A(n_86), .Y(n_130) );
NOR2xp33_ASAP7_75t_L g131 ( .A(n_101), .B(n_5), .Y(n_131) );
AND2x4_ASAP7_75t_L g132 ( .A(n_81), .B(n_5), .Y(n_132) );
BUFx6f_ASAP7_75t_L g133 ( .A(n_78), .Y(n_133) );
NAND2xp5_ASAP7_75t_SL g134 ( .A(n_105), .B(n_6), .Y(n_134) );
INVx3_ASAP7_75t_L g135 ( .A(n_89), .Y(n_135) );
BUFx6f_ASAP7_75t_L g136 ( .A(n_124), .Y(n_136) );
INVx1_ASAP7_75t_SL g137 ( .A(n_121), .Y(n_137) );
NAND2xp33_ASAP7_75t_L g138 ( .A(n_116), .B(n_91), .Y(n_138) );
NAND2xp5_ASAP7_75t_SL g139 ( .A(n_121), .B(n_102), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_120), .B(n_93), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_130), .Y(n_141) );
BUFx3_ASAP7_75t_L g142 ( .A(n_132), .Y(n_142) );
INVx2_ASAP7_75t_L g143 ( .A(n_124), .Y(n_143) );
NOR2xp33_ASAP7_75t_L g144 ( .A(n_120), .B(n_108), .Y(n_144) );
AND2x4_ASAP7_75t_L g145 ( .A(n_121), .B(n_82), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_130), .Y(n_146) );
BUFx6f_ASAP7_75t_L g147 ( .A(n_124), .Y(n_147) );
INVx2_ASAP7_75t_L g148 ( .A(n_124), .Y(n_148) );
INVx2_ASAP7_75t_L g149 ( .A(n_124), .Y(n_149) );
AND2x4_ASAP7_75t_L g150 ( .A(n_132), .B(n_82), .Y(n_150) );
INVxp67_ASAP7_75t_L g151 ( .A(n_127), .Y(n_151) );
AND2x6_ASAP7_75t_L g152 ( .A(n_132), .B(n_99), .Y(n_152) );
AOI22xp5_ASAP7_75t_L g153 ( .A1(n_127), .A2(n_98), .B1(n_83), .B2(n_90), .Y(n_153) );
NOR2xp33_ASAP7_75t_L g154 ( .A(n_116), .B(n_88), .Y(n_154) );
INVx2_ASAP7_75t_L g155 ( .A(n_124), .Y(n_155) );
NOR2xp33_ASAP7_75t_L g156 ( .A(n_135), .B(n_88), .Y(n_156) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_124), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_130), .Y(n_158) );
BUFx3_ASAP7_75t_L g159 ( .A(n_132), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_142), .Y(n_160) );
NOR2x1_ASAP7_75t_R g161 ( .A(n_145), .B(n_90), .Y(n_161) );
AOI22xp33_ASAP7_75t_SL g162 ( .A1(n_137), .A2(n_118), .B1(n_127), .B2(n_92), .Y(n_162) );
BUFx6f_ASAP7_75t_L g163 ( .A(n_142), .Y(n_163) );
INVx1_ASAP7_75t_L g164 ( .A(n_142), .Y(n_164) );
OAI22xp5_ASAP7_75t_L g165 ( .A1(n_151), .A2(n_106), .B1(n_94), .B2(n_95), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_159), .Y(n_166) );
NAND2xp33_ASAP7_75t_L g167 ( .A(n_152), .B(n_130), .Y(n_167) );
INVx4_ASAP7_75t_L g168 ( .A(n_152), .Y(n_168) );
BUFx3_ASAP7_75t_L g169 ( .A(n_152), .Y(n_169) );
INVx2_ASAP7_75t_L g170 ( .A(n_159), .Y(n_170) );
BUFx6f_ASAP7_75t_L g171 ( .A(n_159), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_150), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_150), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_154), .B(n_131), .Y(n_174) );
AO22x1_ASAP7_75t_L g175 ( .A1(n_152), .A2(n_132), .B1(n_98), .B2(n_96), .Y(n_175) );
CKINVDCx11_ASAP7_75t_R g176 ( .A(n_145), .Y(n_176) );
INVx1_ASAP7_75t_SL g177 ( .A(n_145), .Y(n_177) );
NAND2xp5_ASAP7_75t_SL g178 ( .A(n_145), .B(n_91), .Y(n_178) );
NOR2xp33_ASAP7_75t_L g179 ( .A(n_144), .B(n_131), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_150), .Y(n_180) );
INVx3_ASAP7_75t_L g181 ( .A(n_152), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_150), .Y(n_182) );
AOI22xp5_ASAP7_75t_L g183 ( .A1(n_152), .A2(n_118), .B1(n_135), .B2(n_128), .Y(n_183) );
INVx8_ASAP7_75t_L g184 ( .A(n_152), .Y(n_184) );
INVx2_ASAP7_75t_L g185 ( .A(n_141), .Y(n_185) );
NOR2xp33_ASAP7_75t_L g186 ( .A(n_140), .B(n_135), .Y(n_186) );
INVx3_ASAP7_75t_L g187 ( .A(n_152), .Y(n_187) );
INVx2_ASAP7_75t_L g188 ( .A(n_141), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_156), .B(n_135), .Y(n_189) );
INVxp67_ASAP7_75t_L g190 ( .A(n_139), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_177), .B(n_153), .Y(n_191) );
AOI22xp5_ASAP7_75t_L g192 ( .A1(n_179), .A2(n_153), .B1(n_138), .B2(n_134), .Y(n_192) );
BUFx6f_ASAP7_75t_L g193 ( .A(n_184), .Y(n_193) );
BUFx6f_ASAP7_75t_L g194 ( .A(n_184), .Y(n_194) );
NAND2xp5_ASAP7_75t_SL g195 ( .A(n_168), .B(n_111), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_175), .B(n_128), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_175), .B(n_134), .Y(n_197) );
BUFx6f_ASAP7_75t_L g198 ( .A(n_184), .Y(n_198) );
AOI21xp5_ASAP7_75t_L g199 ( .A1(n_189), .A2(n_158), .B(n_146), .Y(n_199) );
BUFx2_ASAP7_75t_SL g200 ( .A(n_168), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_172), .Y(n_201) );
CKINVDCx5p33_ASAP7_75t_R g202 ( .A(n_176), .Y(n_202) );
NOR2xp67_ASAP7_75t_L g203 ( .A(n_183), .B(n_111), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_172), .Y(n_204) );
INVx2_ASAP7_75t_SL g205 ( .A(n_184), .Y(n_205) );
BUFx6f_ASAP7_75t_L g206 ( .A(n_184), .Y(n_206) );
HB1xp67_ASAP7_75t_L g207 ( .A(n_165), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_173), .Y(n_208) );
A2O1A1Ixp33_ASAP7_75t_L g209 ( .A1(n_186), .A2(n_135), .B(n_119), .C(n_125), .Y(n_209) );
AO21x1_ASAP7_75t_L g210 ( .A1(n_174), .A2(n_125), .B(n_119), .Y(n_210) );
INVx3_ASAP7_75t_L g211 ( .A(n_163), .Y(n_211) );
INVx1_ASAP7_75t_L g212 ( .A(n_173), .Y(n_212) );
INVxp67_ASAP7_75t_L g213 ( .A(n_161), .Y(n_213) );
BUFx2_ASAP7_75t_L g214 ( .A(n_168), .Y(n_214) );
AOI22xp5_ASAP7_75t_L g215 ( .A1(n_183), .A2(n_112), .B1(n_97), .B2(n_103), .Y(n_215) );
O2A1O1Ixp33_ASAP7_75t_SL g216 ( .A1(n_160), .A2(n_158), .B(n_146), .C(n_107), .Y(n_216) );
NOR2xp33_ASAP7_75t_L g217 ( .A(n_190), .B(n_76), .Y(n_217) );
OAI22xp5_ASAP7_75t_L g218 ( .A1(n_168), .A2(n_129), .B1(n_125), .B2(n_119), .Y(n_218) );
INVx2_ASAP7_75t_L g219 ( .A(n_163), .Y(n_219) );
HB1xp67_ASAP7_75t_L g220 ( .A(n_169), .Y(n_220) );
INVx5_ASAP7_75t_L g221 ( .A(n_163), .Y(n_221) );
OAI22xp5_ASAP7_75t_L g222 ( .A1(n_203), .A2(n_180), .B1(n_182), .B2(n_169), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_201), .Y(n_223) );
NOR2xp33_ASAP7_75t_L g224 ( .A(n_207), .B(n_161), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_191), .B(n_180), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_192), .B(n_182), .Y(n_226) );
CKINVDCx5p33_ASAP7_75t_R g227 ( .A(n_202), .Y(n_227) );
INVx2_ASAP7_75t_L g228 ( .A(n_219), .Y(n_228) );
OAI22xp5_ASAP7_75t_SL g229 ( .A1(n_213), .A2(n_162), .B1(n_215), .B2(n_202), .Y(n_229) );
AOI222xp33_ASAP7_75t_L g230 ( .A1(n_217), .A2(n_178), .B1(n_84), .B2(n_85), .C1(n_109), .C2(n_79), .Y(n_230) );
AOI22xp33_ASAP7_75t_L g231 ( .A1(n_197), .A2(n_164), .B1(n_166), .B2(n_160), .Y(n_231) );
INVx2_ASAP7_75t_L g232 ( .A(n_219), .Y(n_232) );
HB1xp67_ASAP7_75t_L g233 ( .A(n_221), .Y(n_233) );
NAND2x1_ASAP7_75t_L g234 ( .A(n_211), .B(n_163), .Y(n_234) );
AOI21xp33_ASAP7_75t_L g235 ( .A1(n_196), .A2(n_166), .B(n_164), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_204), .Y(n_236) );
O2A1O1Ixp33_ASAP7_75t_SL g237 ( .A1(n_209), .A2(n_170), .B(n_114), .C(n_100), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_208), .B(n_170), .Y(n_238) );
NAND2xp5_ASAP7_75t_SL g239 ( .A(n_193), .B(n_169), .Y(n_239) );
INVx2_ASAP7_75t_L g240 ( .A(n_211), .Y(n_240) );
OR2x2_ASAP7_75t_L g241 ( .A(n_212), .B(n_163), .Y(n_241) );
BUFx6f_ASAP7_75t_L g242 ( .A(n_193), .Y(n_242) );
NAND2xp5_ASAP7_75t_SL g243 ( .A(n_193), .B(n_181), .Y(n_243) );
OAI22xp5_ASAP7_75t_L g244 ( .A1(n_200), .A2(n_129), .B1(n_117), .B2(n_163), .Y(n_244) );
OAI22xp5_ASAP7_75t_L g245 ( .A1(n_200), .A2(n_171), .B1(n_187), .B2(n_181), .Y(n_245) );
BUFx3_ASAP7_75t_L g246 ( .A(n_193), .Y(n_246) );
AOI22xp33_ASAP7_75t_L g247 ( .A1(n_214), .A2(n_171), .B1(n_187), .B2(n_181), .Y(n_247) );
AOI22xp33_ASAP7_75t_SL g248 ( .A1(n_214), .A2(n_181), .B1(n_187), .B2(n_171), .Y(n_248) );
BUFx4f_ASAP7_75t_SL g249 ( .A(n_246), .Y(n_249) );
AND2x4_ASAP7_75t_SL g250 ( .A(n_233), .B(n_193), .Y(n_250) );
BUFx5_ASAP7_75t_L g251 ( .A(n_246), .Y(n_251) );
AO21x1_ASAP7_75t_L g252 ( .A1(n_235), .A2(n_218), .B(n_199), .Y(n_252) );
OR2x2_ASAP7_75t_L g253 ( .A(n_226), .B(n_210), .Y(n_253) );
OAI22xp5_ASAP7_75t_L g254 ( .A1(n_224), .A2(n_221), .B1(n_220), .B2(n_205), .Y(n_254) );
OAI22xp5_ASAP7_75t_L g255 ( .A1(n_225), .A2(n_221), .B1(n_205), .B2(n_198), .Y(n_255) );
AOI22xp33_ASAP7_75t_L g256 ( .A1(n_229), .A2(n_210), .B1(n_171), .B2(n_195), .Y(n_256) );
AOI22xp33_ASAP7_75t_L g257 ( .A1(n_229), .A2(n_171), .B1(n_211), .B2(n_221), .Y(n_257) );
AO21x2_ASAP7_75t_L g258 ( .A1(n_237), .A2(n_216), .B(n_117), .Y(n_258) );
AOI22xp33_ASAP7_75t_L g259 ( .A1(n_230), .A2(n_171), .B1(n_221), .B2(n_167), .Y(n_259) );
AND2x4_ASAP7_75t_L g260 ( .A(n_223), .B(n_194), .Y(n_260) );
AOI221xp5_ASAP7_75t_L g261 ( .A1(n_223), .A2(n_110), .B1(n_84), .B2(n_85), .C(n_117), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_236), .Y(n_262) );
AOI22xp33_ASAP7_75t_L g263 ( .A1(n_230), .A2(n_206), .B1(n_198), .B2(n_194), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_236), .Y(n_264) );
AND2x2_ASAP7_75t_L g265 ( .A(n_241), .B(n_129), .Y(n_265) );
AOI22xp33_ASAP7_75t_L g266 ( .A1(n_222), .A2(n_206), .B1(n_198), .B2(n_194), .Y(n_266) );
BUFx3_ASAP7_75t_L g267 ( .A(n_246), .Y(n_267) );
OAI211xp5_ASAP7_75t_SL g268 ( .A1(n_231), .A2(n_115), .B(n_122), .C(n_143), .Y(n_268) );
AOI22xp33_ASAP7_75t_L g269 ( .A1(n_244), .A2(n_206), .B1(n_198), .B2(n_194), .Y(n_269) );
AOI22xp33_ASAP7_75t_L g270 ( .A1(n_244), .A2(n_206), .B1(n_198), .B2(n_194), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_238), .B(n_187), .Y(n_271) );
BUFx3_ASAP7_75t_L g272 ( .A(n_249), .Y(n_272) );
AOI221xp5_ASAP7_75t_L g273 ( .A1(n_261), .A2(n_227), .B1(n_133), .B2(n_130), .C(n_241), .Y(n_273) );
OAI221xp5_ASAP7_75t_SL g274 ( .A1(n_257), .A2(n_247), .B1(n_122), .B2(n_115), .C(n_240), .Y(n_274) );
NAND4xp25_ASAP7_75t_L g275 ( .A(n_256), .B(n_122), .C(n_115), .D(n_248), .Y(n_275) );
OAI221xp5_ASAP7_75t_L g276 ( .A1(n_263), .A2(n_234), .B1(n_133), .B2(n_130), .C(n_240), .Y(n_276) );
AOI22xp33_ASAP7_75t_L g277 ( .A1(n_260), .A2(n_240), .B1(n_133), .B2(n_242), .Y(n_277) );
AOI22xp5_ASAP7_75t_L g278 ( .A1(n_262), .A2(n_232), .B1(n_228), .B2(n_245), .Y(n_278) );
AOI221xp5_ASAP7_75t_L g279 ( .A1(n_262), .A2(n_133), .B1(n_130), .B2(n_115), .C(n_122), .Y(n_279) );
OAI221xp5_ASAP7_75t_L g280 ( .A1(n_259), .A2(n_234), .B1(n_133), .B2(n_130), .C(n_243), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_264), .Y(n_281) );
BUFx3_ASAP7_75t_L g282 ( .A(n_267), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_264), .Y(n_283) );
HB1xp67_ASAP7_75t_L g284 ( .A(n_265), .Y(n_284) );
AOI221xp5_ASAP7_75t_L g285 ( .A1(n_254), .A2(n_133), .B1(n_115), .B2(n_122), .C(n_228), .Y(n_285) );
OAI31xp33_ASAP7_75t_L g286 ( .A1(n_253), .A2(n_239), .A3(n_228), .B(n_232), .Y(n_286) );
OAI221xp5_ASAP7_75t_L g287 ( .A1(n_253), .A2(n_133), .B1(n_232), .B2(n_242), .C(n_123), .Y(n_287) );
AOI211xp5_ASAP7_75t_L g288 ( .A1(n_252), .A2(n_124), .B(n_126), .C(n_123), .Y(n_288) );
BUFx3_ASAP7_75t_L g289 ( .A(n_267), .Y(n_289) );
OR2x2_ASAP7_75t_L g290 ( .A(n_265), .B(n_242), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_260), .B(n_8), .Y(n_291) );
OAI21xp5_ASAP7_75t_SL g292 ( .A1(n_250), .A2(n_206), .B(n_242), .Y(n_292) );
OR2x2_ASAP7_75t_L g293 ( .A(n_260), .B(n_242), .Y(n_293) );
AND2x2_ASAP7_75t_L g294 ( .A(n_281), .B(n_252), .Y(n_294) );
AND2x2_ASAP7_75t_L g295 ( .A(n_281), .B(n_251), .Y(n_295) );
INVx2_ASAP7_75t_L g296 ( .A(n_283), .Y(n_296) );
AND2x2_ASAP7_75t_L g297 ( .A(n_283), .B(n_251), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_278), .Y(n_298) );
INVx1_ASAP7_75t_SL g299 ( .A(n_282), .Y(n_299) );
AOI22xp33_ASAP7_75t_L g300 ( .A1(n_284), .A2(n_260), .B1(n_258), .B2(n_268), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_278), .Y(n_301) );
AOI221x1_ASAP7_75t_L g302 ( .A1(n_275), .A2(n_255), .B1(n_123), .B2(n_126), .C(n_271), .Y(n_302) );
AND2x2_ASAP7_75t_L g303 ( .A(n_290), .B(n_251), .Y(n_303) );
AOI22xp33_ASAP7_75t_L g304 ( .A1(n_273), .A2(n_258), .B1(n_251), .B2(n_270), .Y(n_304) );
AND2x2_ASAP7_75t_L g305 ( .A(n_290), .B(n_293), .Y(n_305) );
AND2x2_ASAP7_75t_L g306 ( .A(n_293), .B(n_251), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_291), .Y(n_307) );
BUFx3_ASAP7_75t_L g308 ( .A(n_282), .Y(n_308) );
NAND3xp33_ASAP7_75t_L g309 ( .A(n_288), .B(n_123), .C(n_126), .Y(n_309) );
AND2x2_ASAP7_75t_L g310 ( .A(n_289), .B(n_251), .Y(n_310) );
AND2x2_ASAP7_75t_L g311 ( .A(n_289), .B(n_251), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_287), .Y(n_312) );
AO21x2_ASAP7_75t_L g313 ( .A1(n_276), .A2(n_258), .B(n_149), .Y(n_313) );
BUFx2_ASAP7_75t_L g314 ( .A(n_272), .Y(n_314) );
AOI22xp33_ASAP7_75t_L g315 ( .A1(n_280), .A2(n_251), .B1(n_269), .B2(n_250), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_292), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_279), .Y(n_317) );
INVx2_ASAP7_75t_L g318 ( .A(n_286), .Y(n_318) );
AND2x2_ASAP7_75t_L g319 ( .A(n_277), .B(n_126), .Y(n_319) );
AND2x2_ASAP7_75t_L g320 ( .A(n_272), .B(n_126), .Y(n_320) );
INVx3_ASAP7_75t_L g321 ( .A(n_274), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_305), .B(n_8), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_296), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_296), .Y(n_324) );
AND2x2_ASAP7_75t_L g325 ( .A(n_305), .B(n_123), .Y(n_325) );
O2A1O1Ixp33_ASAP7_75t_L g326 ( .A1(n_321), .A2(n_285), .B(n_266), .C(n_155), .Y(n_326) );
OAI21xp5_ASAP7_75t_L g327 ( .A1(n_302), .A2(n_155), .B(n_149), .Y(n_327) );
OAI31xp33_ASAP7_75t_L g328 ( .A1(n_321), .A2(n_10), .A3(n_11), .B(n_12), .Y(n_328) );
AND2x2_ASAP7_75t_L g329 ( .A(n_305), .B(n_123), .Y(n_329) );
AND2x4_ASAP7_75t_L g330 ( .A(n_294), .B(n_126), .Y(n_330) );
AND2x2_ASAP7_75t_L g331 ( .A(n_294), .B(n_123), .Y(n_331) );
OAI21xp5_ASAP7_75t_SL g332 ( .A1(n_314), .A2(n_321), .B(n_302), .Y(n_332) );
INVx1_ASAP7_75t_SL g333 ( .A(n_299), .Y(n_333) );
OR2x2_ASAP7_75t_L g334 ( .A(n_296), .B(n_126), .Y(n_334) );
NAND3xp33_ASAP7_75t_SL g335 ( .A(n_314), .B(n_13), .C(n_14), .Y(n_335) );
OR2x2_ASAP7_75t_L g336 ( .A(n_298), .B(n_126), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_307), .B(n_13), .Y(n_337) );
INVx2_ASAP7_75t_L g338 ( .A(n_295), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_294), .Y(n_339) );
HB1xp67_ASAP7_75t_L g340 ( .A(n_299), .Y(n_340) );
AND2x2_ASAP7_75t_L g341 ( .A(n_295), .B(n_15), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_295), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_297), .Y(n_343) );
OR2x2_ASAP7_75t_L g344 ( .A(n_298), .B(n_15), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_297), .Y(n_345) );
AND2x2_ASAP7_75t_L g346 ( .A(n_297), .B(n_16), .Y(n_346) );
AND2x2_ASAP7_75t_L g347 ( .A(n_303), .B(n_17), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_298), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_307), .B(n_17), .Y(n_349) );
O2A1O1Ixp33_ASAP7_75t_SL g350 ( .A1(n_316), .A2(n_19), .B(n_20), .C(n_21), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_301), .Y(n_351) );
AND2x2_ASAP7_75t_L g352 ( .A(n_303), .B(n_20), .Y(n_352) );
AND2x2_ASAP7_75t_L g353 ( .A(n_303), .B(n_21), .Y(n_353) );
BUFx3_ASAP7_75t_L g354 ( .A(n_308), .Y(n_354) );
AND2x2_ASAP7_75t_L g355 ( .A(n_306), .B(n_27), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_301), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_301), .Y(n_357) );
INVx2_ASAP7_75t_SL g358 ( .A(n_308), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_316), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_316), .Y(n_360) );
INVx2_ASAP7_75t_L g361 ( .A(n_307), .Y(n_361) );
AND2x4_ASAP7_75t_L g362 ( .A(n_306), .B(n_28), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_361), .Y(n_363) );
OR2x6_ASAP7_75t_L g364 ( .A(n_354), .B(n_308), .Y(n_364) );
INVx1_ASAP7_75t_SL g365 ( .A(n_333), .Y(n_365) );
NOR2xp67_ASAP7_75t_SL g366 ( .A(n_332), .B(n_314), .Y(n_366) );
AND2x2_ASAP7_75t_L g367 ( .A(n_340), .B(n_306), .Y(n_367) );
NOR2xp33_ASAP7_75t_L g368 ( .A(n_359), .B(n_320), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_325), .B(n_308), .Y(n_369) );
AOI21xp33_ASAP7_75t_L g370 ( .A1(n_328), .A2(n_320), .B(n_318), .Y(n_370) );
AND2x2_ASAP7_75t_L g371 ( .A(n_339), .B(n_310), .Y(n_371) );
INVxp33_ASAP7_75t_L g372 ( .A(n_347), .Y(n_372) );
OR2x2_ASAP7_75t_L g373 ( .A(n_342), .B(n_310), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_325), .B(n_310), .Y(n_374) );
OR2x2_ASAP7_75t_L g375 ( .A(n_342), .B(n_311), .Y(n_375) );
BUFx2_ASAP7_75t_L g376 ( .A(n_354), .Y(n_376) );
INVx1_ASAP7_75t_SL g377 ( .A(n_354), .Y(n_377) );
INVx1_ASAP7_75t_SL g378 ( .A(n_347), .Y(n_378) );
AND2x2_ASAP7_75t_L g379 ( .A(n_343), .B(n_311), .Y(n_379) );
AND2x2_ASAP7_75t_L g380 ( .A(n_343), .B(n_311), .Y(n_380) );
OAI22xp33_ASAP7_75t_L g381 ( .A1(n_344), .A2(n_321), .B1(n_302), .B2(n_318), .Y(n_381) );
INVxp67_ASAP7_75t_L g382 ( .A(n_329), .Y(n_382) );
HB1xp67_ASAP7_75t_L g383 ( .A(n_329), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_339), .B(n_318), .Y(n_384) );
AND2x2_ASAP7_75t_L g385 ( .A(n_338), .B(n_318), .Y(n_385) );
OAI21xp33_ASAP7_75t_L g386 ( .A1(n_359), .A2(n_320), .B(n_304), .Y(n_386) );
NAND4xp75_ASAP7_75t_L g387 ( .A(n_328), .B(n_312), .C(n_319), .D(n_317), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_345), .B(n_312), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_345), .B(n_312), .Y(n_389) );
INVxp67_ASAP7_75t_SL g390 ( .A(n_334), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_360), .Y(n_391) );
AND2x4_ASAP7_75t_L g392 ( .A(n_338), .B(n_313), .Y(n_392) );
AND2x2_ASAP7_75t_L g393 ( .A(n_360), .B(n_313), .Y(n_393) );
AO21x1_ASAP7_75t_L g394 ( .A1(n_352), .A2(n_319), .B(n_317), .Y(n_394) );
AND2x4_ASAP7_75t_L g395 ( .A(n_358), .B(n_313), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_341), .B(n_321), .Y(n_396) );
INVx2_ASAP7_75t_L g397 ( .A(n_323), .Y(n_397) );
AND2x2_ASAP7_75t_L g398 ( .A(n_331), .B(n_313), .Y(n_398) );
XNOR2x2_ASAP7_75t_L g399 ( .A(n_352), .B(n_309), .Y(n_399) );
NOR2x1p5_ASAP7_75t_L g400 ( .A(n_335), .B(n_321), .Y(n_400) );
NOR2xp33_ASAP7_75t_L g401 ( .A(n_322), .B(n_300), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_341), .B(n_300), .Y(n_402) );
AND2x4_ASAP7_75t_L g403 ( .A(n_358), .B(n_313), .Y(n_403) );
OAI31xp33_ASAP7_75t_L g404 ( .A1(n_353), .A2(n_309), .A3(n_315), .B(n_317), .Y(n_404) );
NOR2xp33_ASAP7_75t_L g405 ( .A(n_337), .B(n_319), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_323), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_324), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_324), .Y(n_408) );
INVxp67_ASAP7_75t_L g409 ( .A(n_353), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_346), .B(n_304), .Y(n_410) );
XOR2x2_ASAP7_75t_L g411 ( .A(n_378), .B(n_346), .Y(n_411) );
NAND2x1p5_ASAP7_75t_L g412 ( .A(n_376), .B(n_362), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_384), .B(n_357), .Y(n_413) );
XOR2xp5_ASAP7_75t_L g414 ( .A(n_372), .B(n_362), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_391), .B(n_357), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_371), .Y(n_416) );
AOI21xp33_ASAP7_75t_SL g417 ( .A1(n_372), .A2(n_344), .B(n_362), .Y(n_417) );
XOR2xp5_ASAP7_75t_L g418 ( .A(n_383), .B(n_362), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_371), .B(n_331), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_373), .Y(n_420) );
OAI21xp5_ASAP7_75t_L g421 ( .A1(n_387), .A2(n_350), .B(n_355), .Y(n_421) );
OR2x2_ASAP7_75t_L g422 ( .A(n_375), .B(n_356), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_406), .Y(n_423) );
NOR2xp33_ASAP7_75t_L g424 ( .A(n_365), .B(n_349), .Y(n_424) );
INVxp67_ASAP7_75t_L g425 ( .A(n_367), .Y(n_425) );
AND2x2_ASAP7_75t_L g426 ( .A(n_379), .B(n_330), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_388), .B(n_356), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_407), .Y(n_428) );
AOI22xp33_ASAP7_75t_L g429 ( .A1(n_400), .A2(n_351), .B1(n_348), .B2(n_330), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_408), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_389), .B(n_351), .Y(n_431) );
OR4x1_ASAP7_75t_L g432 ( .A(n_363), .B(n_348), .C(n_330), .D(n_355), .Y(n_432) );
NOR2xp33_ASAP7_75t_L g433 ( .A(n_409), .B(n_330), .Y(n_433) );
AOI321xp33_ASAP7_75t_L g434 ( .A1(n_401), .A2(n_315), .A3(n_336), .B1(n_326), .B2(n_334), .C(n_155), .Y(n_434) );
NOR2xp33_ASAP7_75t_L g435 ( .A(n_396), .B(n_336), .Y(n_435) );
OAI211xp5_ASAP7_75t_L g436 ( .A1(n_404), .A2(n_327), .B(n_149), .C(n_148), .Y(n_436) );
NOR2x1_ASAP7_75t_L g437 ( .A(n_364), .B(n_148), .Y(n_437) );
BUFx2_ASAP7_75t_L g438 ( .A(n_364), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_380), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_385), .B(n_32), .Y(n_440) );
XNOR2x2_ASAP7_75t_L g441 ( .A(n_399), .B(n_33), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_393), .B(n_35), .Y(n_442) );
NAND2xp5_ASAP7_75t_SL g443 ( .A(n_394), .B(n_157), .Y(n_443) );
OAI22xp5_ASAP7_75t_L g444 ( .A1(n_364), .A2(n_143), .B1(n_147), .B2(n_157), .Y(n_444) );
OR2x2_ASAP7_75t_L g445 ( .A(n_374), .B(n_36), .Y(n_445) );
INVxp67_ASAP7_75t_SL g446 ( .A(n_390), .Y(n_446) );
OR2x2_ASAP7_75t_L g447 ( .A(n_369), .B(n_37), .Y(n_447) );
AND2x2_ASAP7_75t_L g448 ( .A(n_382), .B(n_39), .Y(n_448) );
AOI221xp5_ASAP7_75t_L g449 ( .A1(n_370), .A2(n_157), .B1(n_147), .B2(n_136), .C(n_185), .Y(n_449) );
NAND4xp25_ASAP7_75t_L g450 ( .A(n_405), .B(n_40), .C(n_42), .D(n_45), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_397), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_368), .B(n_49), .Y(n_452) );
AOI22xp33_ASAP7_75t_L g453 ( .A1(n_405), .A2(n_157), .B1(n_147), .B2(n_136), .Y(n_453) );
OAI21xp5_ASAP7_75t_SL g454 ( .A1(n_381), .A2(n_50), .B(n_51), .Y(n_454) );
OAI22xp33_ASAP7_75t_SL g455 ( .A1(n_364), .A2(n_53), .B1(n_54), .B2(n_55), .Y(n_455) );
XOR2x2_ASAP7_75t_L g456 ( .A(n_399), .B(n_58), .Y(n_456) );
OAI22xp5_ASAP7_75t_L g457 ( .A1(n_402), .A2(n_157), .B1(n_147), .B2(n_136), .Y(n_457) );
INVxp67_ASAP7_75t_L g458 ( .A(n_368), .Y(n_458) );
AND2x2_ASAP7_75t_L g459 ( .A(n_377), .B(n_60), .Y(n_459) );
OR2x2_ASAP7_75t_L g460 ( .A(n_397), .B(n_61), .Y(n_460) );
AOI21xp5_ASAP7_75t_L g461 ( .A1(n_381), .A2(n_188), .B(n_185), .Y(n_461) );
OAI22xp5_ASAP7_75t_L g462 ( .A1(n_410), .A2(n_147), .B1(n_136), .B2(n_64), .Y(n_462) );
INVx2_ASAP7_75t_L g463 ( .A(n_392), .Y(n_463) );
XNOR2xp5_ASAP7_75t_L g464 ( .A(n_398), .B(n_62), .Y(n_464) );
AOI21xp5_ASAP7_75t_L g465 ( .A1(n_395), .A2(n_188), .B(n_136), .Y(n_465) );
INVxp67_ASAP7_75t_L g466 ( .A(n_366), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_393), .B(n_63), .Y(n_467) );
OAI211xp5_ASAP7_75t_L g468 ( .A1(n_386), .A2(n_65), .B(n_66), .C(n_68), .Y(n_468) );
OAI21xp33_ASAP7_75t_SL g469 ( .A1(n_398), .A2(n_69), .B(n_70), .Y(n_469) );
NOR2xp33_ASAP7_75t_L g470 ( .A(n_395), .B(n_71), .Y(n_470) );
NOR3xp33_ASAP7_75t_L g471 ( .A(n_395), .B(n_73), .C(n_74), .Y(n_471) );
AOI31xp33_ASAP7_75t_L g472 ( .A1(n_403), .A2(n_136), .A3(n_394), .B(n_372), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_403), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_403), .Y(n_474) );
OR2x2_ASAP7_75t_L g475 ( .A(n_392), .B(n_383), .Y(n_475) );
A2O1A1Ixp33_ASAP7_75t_L g476 ( .A1(n_392), .A2(n_366), .B(n_404), .C(n_372), .Y(n_476) );
AND2x2_ASAP7_75t_L g477 ( .A(n_367), .B(n_378), .Y(n_477) );
NOR2x1_ASAP7_75t_L g478 ( .A(n_400), .B(n_332), .Y(n_478) );
INVx2_ASAP7_75t_L g479 ( .A(n_475), .Y(n_479) );
NOR4xp75_ASAP7_75t_L g480 ( .A(n_421), .B(n_443), .C(n_456), .D(n_441), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_446), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_416), .Y(n_482) );
AND3x4_ASAP7_75t_L g483 ( .A(n_478), .B(n_471), .C(n_437), .Y(n_483) );
NOR3xp33_ASAP7_75t_L g484 ( .A(n_476), .B(n_454), .C(n_450), .Y(n_484) );
INVxp67_ASAP7_75t_SL g485 ( .A(n_465), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_458), .B(n_420), .Y(n_486) );
OAI21xp5_ASAP7_75t_L g487 ( .A1(n_469), .A2(n_472), .B(n_461), .Y(n_487) );
AOI221xp5_ASAP7_75t_L g488 ( .A1(n_424), .A2(n_425), .B1(n_417), .B2(n_432), .C(n_438), .Y(n_488) );
XNOR2xp5_ASAP7_75t_L g489 ( .A(n_411), .B(n_414), .Y(n_489) );
INVxp67_ASAP7_75t_L g490 ( .A(n_477), .Y(n_490) );
OA22x2_ASAP7_75t_L g491 ( .A1(n_466), .A2(n_464), .B1(n_418), .B2(n_474), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_428), .Y(n_492) );
OR2x2_ASAP7_75t_L g493 ( .A(n_422), .B(n_439), .Y(n_493) );
AOI31xp33_ASAP7_75t_L g494 ( .A1(n_412), .A2(n_429), .A3(n_461), .B(n_465), .Y(n_494) );
OAI211xp5_ASAP7_75t_L g495 ( .A1(n_434), .A2(n_436), .B(n_433), .C(n_449), .Y(n_495) );
OR2x2_ASAP7_75t_L g496 ( .A(n_473), .B(n_419), .Y(n_496) );
INVxp67_ASAP7_75t_L g497 ( .A(n_481), .Y(n_497) );
OAI22xp5_ASAP7_75t_L g498 ( .A1(n_491), .A2(n_412), .B1(n_426), .B2(n_463), .Y(n_498) );
OAI221xp5_ASAP7_75t_L g499 ( .A1(n_491), .A2(n_449), .B1(n_470), .B2(n_468), .C(n_427), .Y(n_499) );
AOI21xp33_ASAP7_75t_L g500 ( .A1(n_494), .A2(n_455), .B(n_445), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_492), .Y(n_501) );
AOI22xp5_ASAP7_75t_L g502 ( .A1(n_484), .A2(n_435), .B1(n_423), .B2(n_430), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_488), .B(n_431), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_482), .B(n_431), .Y(n_504) );
AOI221xp5_ASAP7_75t_L g505 ( .A1(n_494), .A2(n_427), .B1(n_413), .B2(n_415), .C(n_451), .Y(n_505) );
HB1xp67_ASAP7_75t_L g506 ( .A(n_479), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_497), .Y(n_507) );
NAND5xp2_ASAP7_75t_L g508 ( .A(n_505), .B(n_487), .C(n_495), .D(n_468), .E(n_480), .Y(n_508) );
AOI21xp5_ASAP7_75t_L g509 ( .A1(n_499), .A2(n_487), .B(n_483), .Y(n_509) );
NOR3xp33_ASAP7_75t_L g510 ( .A(n_500), .B(n_485), .C(n_462), .Y(n_510) );
OA22x2_ASAP7_75t_L g511 ( .A1(n_502), .A2(n_489), .B1(n_490), .B2(n_486), .Y(n_511) );
AND3x1_ASAP7_75t_L g512 ( .A(n_508), .B(n_503), .C(n_506), .Y(n_512) );
NAND3xp33_ASAP7_75t_SL g513 ( .A(n_509), .B(n_498), .C(n_501), .Y(n_513) );
OAI22xp5_ASAP7_75t_SL g514 ( .A1(n_511), .A2(n_452), .B1(n_453), .B2(n_447), .Y(n_514) );
AOI21xp5_ASAP7_75t_L g515 ( .A1(n_512), .A2(n_507), .B(n_510), .Y(n_515) );
OR2x2_ASAP7_75t_L g516 ( .A(n_513), .B(n_504), .Y(n_516) );
NOR2x1p5_ASAP7_75t_L g517 ( .A(n_516), .B(n_514), .Y(n_517) );
AOI222xp33_ASAP7_75t_L g518 ( .A1(n_517), .A2(n_515), .B1(n_448), .B2(n_442), .C1(n_459), .C2(n_467), .Y(n_518) );
AOI22x1_ASAP7_75t_L g519 ( .A1(n_518), .A2(n_496), .B1(n_493), .B2(n_460), .Y(n_519) );
AOI221xp5_ASAP7_75t_L g520 ( .A1(n_519), .A2(n_457), .B1(n_444), .B2(n_442), .C(n_440), .Y(n_520) );
endmodule