module fake_jpeg_12993_n_76 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_76);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_76;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_10;
wire n_23;
wire n_69;
wire n_27;
wire n_64;
wire n_55;
wire n_47;
wire n_22;
wire n_51;
wire n_14;
wire n_40;
wire n_73;
wire n_19;
wire n_20;
wire n_18;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_71;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_72;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_74;
wire n_11;
wire n_62;
wire n_25;
wire n_17;
wire n_56;
wire n_31;
wire n_67;
wire n_75;
wire n_29;
wire n_43;
wire n_50;
wire n_37;
wire n_12;
wire n_32;
wire n_70;
wire n_15;
wire n_66;

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_5),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_9),
.Y(n_12)
);

INVx3_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

BUFx3_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_2),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_0),
.B(n_8),
.Y(n_18)
);

CKINVDCx14_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

INVx5_ASAP7_75t_L g22 ( 
.A(n_20),
.Y(n_22)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_11),
.B(n_2),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_23),
.B(n_25),
.Y(n_32)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_11),
.B(n_3),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_18),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_26),
.B(n_27),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g27 ( 
.A(n_15),
.B(n_0),
.Y(n_27)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_19),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_28),
.B(n_15),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_27),
.B(n_17),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_30),
.B(n_42),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_26),
.B(n_12),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_39),
.B(n_41),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_22),
.A2(n_20),
.B1(n_13),
.B2(n_10),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_40),
.B(n_43),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_27),
.B(n_12),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

OR2x2_ASAP7_75t_L g43 ( 
.A(n_28),
.B(n_17),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_32),
.B(n_16),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_49),
.B(n_50),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_33),
.B(n_16),
.Y(n_50)
);

CKINVDCx5p33_ASAP7_75t_R g51 ( 
.A(n_43),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_51),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_30),
.B(n_13),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_52),
.B(n_47),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_14),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_53),
.B(n_54),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_37),
.B(n_29),
.Y(n_54)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

AOI21xp5_ASAP7_75t_L g63 ( 
.A1(n_56),
.A2(n_54),
.B(n_59),
.Y(n_63)
);

XOR2x1_ASAP7_75t_L g57 ( 
.A(n_51),
.B(n_37),
.Y(n_57)
);

XNOR2xp5_ASAP7_75t_L g65 ( 
.A(n_57),
.B(n_61),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_46),
.A2(n_21),
.B1(n_34),
.B2(n_31),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_58),
.A2(n_34),
.B1(n_31),
.B2(n_42),
.Y(n_62)
);

A2O1A1Ixp33_ASAP7_75t_SL g67 ( 
.A1(n_62),
.A2(n_64),
.B(n_29),
.C(n_60),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_63),
.B(n_36),
.Y(n_68)
);

AO22x1_ASAP7_75t_L g64 ( 
.A1(n_59),
.A2(n_57),
.B1(n_45),
.B2(n_44),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_55),
.B(n_44),
.C(n_54),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_66),
.B(n_36),
.C(n_6),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_67),
.B(n_68),
.C(n_69),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_69),
.B(n_66),
.C(n_65),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_71),
.B(n_65),
.C(n_64),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_72),
.B(n_73),
.C(n_4),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_70),
.B(n_4),
.Y(n_73)
);

NOR3xp33_ASAP7_75t_L g75 ( 
.A(n_74),
.B(n_6),
.C(n_7),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_L g76 ( 
.A(n_75),
.B(n_7),
.Y(n_76)
);


endmodule