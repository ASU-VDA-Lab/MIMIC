module fake_jpeg_1071_n_184 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_184);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_184;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_140;
wire n_128;
wire n_82;
wire n_96;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

INVx2_ASAP7_75t_SL g17 ( 
.A(n_0),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_13),
.B(n_8),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_11),
.B(n_14),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_10),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_9),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_34),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g35 ( 
.A(n_30),
.B(n_1),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_35),
.B(n_44),
.Y(n_51)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_36),
.Y(n_68)
);

BUFx10_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

BUFx2_ASAP7_75t_L g71 ( 
.A(n_37),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_50),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_17),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_40),
.A2(n_33),
.B1(n_24),
.B2(n_29),
.Y(n_54)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_26),
.B(n_32),
.Y(n_44)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_21),
.Y(n_46)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_46),
.Y(n_72)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_25),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_47),
.B(n_48),
.Y(n_62)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_21),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_20),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_49),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_27),
.Y(n_50)
);

OR2x4_ASAP7_75t_L g52 ( 
.A(n_35),
.B(n_17),
.Y(n_52)
);

AOI21xp33_ASAP7_75t_L g81 ( 
.A1(n_52),
.A2(n_54),
.B(n_22),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_34),
.B(n_25),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_53),
.B(n_67),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_46),
.B(n_18),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_59),
.B(n_61),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_48),
.B(n_18),
.Y(n_61)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_63),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_42),
.A2(n_29),
.B1(n_19),
.B2(n_28),
.Y(n_65)
);

OAI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_65),
.A2(n_76),
.B1(n_23),
.B2(n_37),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_38),
.B(n_28),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_49),
.B(n_19),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_69),
.B(n_5),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_36),
.A2(n_31),
.B1(n_23),
.B2(n_20),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_70),
.A2(n_23),
.B1(n_2),
.B2(n_5),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_45),
.B(n_16),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_74),
.B(n_8),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_41),
.B(n_32),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_75),
.B(n_6),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_40),
.A2(n_29),
.B1(n_33),
.B2(n_24),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_77),
.A2(n_64),
.B1(n_72),
.B2(n_68),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_51),
.B(n_12),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_78),
.Y(n_117)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_66),
.Y(n_80)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_80),
.Y(n_104)
);

OR2x2_ASAP7_75t_SL g109 ( 
.A(n_81),
.B(n_63),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_52),
.B(n_29),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_84),
.B(n_85),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_71),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_53),
.A2(n_43),
.B(n_31),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_86),
.A2(n_58),
.B(n_60),
.Y(n_111)
);

INVxp33_ASAP7_75t_L g87 ( 
.A(n_62),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_87),
.B(n_90),
.Y(n_108)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_66),
.Y(n_88)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_88),
.Y(n_116)
);

A2O1A1Ixp33_ASAP7_75t_L g89 ( 
.A1(n_51),
.A2(n_22),
.B(n_10),
.C(n_4),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_89),
.B(n_93),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_71),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_67),
.Y(n_91)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_91),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_92),
.A2(n_58),
.B1(n_68),
.B2(n_73),
.Y(n_112)
);

A2O1A1Ixp33_ASAP7_75t_L g93 ( 
.A1(n_74),
.A2(n_1),
.B(n_5),
.C(n_6),
.Y(n_93)
);

INVx13_ASAP7_75t_L g94 ( 
.A(n_57),
.Y(n_94)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_94),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_95),
.B(n_96),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_62),
.B(n_9),
.C(n_7),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_97),
.B(n_98),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_71),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_57),
.B(n_7),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_99),
.B(n_100),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_69),
.B(n_7),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_101),
.B(n_56),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_86),
.A2(n_70),
.B1(n_60),
.B2(n_73),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_103),
.A2(n_84),
.B1(n_100),
.B2(n_99),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_106),
.B(n_121),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_109),
.B(n_96),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_111),
.B(n_119),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_112),
.A2(n_115),
.B1(n_85),
.B2(n_90),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_91),
.A2(n_68),
.B1(n_55),
.B2(n_72),
.Y(n_115)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_88),
.Y(n_118)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_118),
.Y(n_130)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_80),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_122),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_111),
.A2(n_79),
.B1(n_92),
.B2(n_84),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_123),
.B(n_129),
.Y(n_143)
);

OR2x2_ASAP7_75t_L g125 ( 
.A(n_107),
.B(n_105),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_125),
.B(n_135),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_108),
.A2(n_79),
.B1(n_95),
.B2(n_83),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_126),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_SL g127 ( 
.A(n_105),
.B(n_83),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_127),
.B(n_113),
.C(n_114),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_108),
.A2(n_93),
.B(n_89),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_128),
.A2(n_138),
.B(n_110),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_119),
.A2(n_100),
.B1(n_99),
.B2(n_55),
.Y(n_129)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_104),
.Y(n_131)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_131),
.Y(n_140)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_132),
.Y(n_151)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_104),
.Y(n_133)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_133),
.Y(n_149)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_116),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_112),
.A2(n_101),
.B1(n_55),
.B2(n_97),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_136),
.A2(n_120),
.B(n_114),
.Y(n_148)
);

NOR3xp33_ASAP7_75t_L g141 ( 
.A(n_137),
.B(n_120),
.C(n_117),
.Y(n_141)
);

AOI22x1_ASAP7_75t_L g138 ( 
.A1(n_109),
.A2(n_113),
.B1(n_115),
.B2(n_107),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_125),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_139),
.B(n_146),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_141),
.B(n_144),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_124),
.B(n_102),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_147),
.B(n_110),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_148),
.A2(n_150),
.B1(n_138),
.B2(n_128),
.Y(n_153)
);

HB1xp67_ASAP7_75t_L g165 ( 
.A(n_153),
.Y(n_165)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_154),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_145),
.A2(n_136),
.B1(n_134),
.B2(n_132),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_155),
.B(n_156),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_140),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_157),
.A2(n_158),
.B(n_161),
.Y(n_163)
);

OA21x2_ASAP7_75t_L g158 ( 
.A1(n_150),
.A2(n_134),
.B(n_151),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_144),
.B(n_127),
.C(n_123),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_159),
.B(n_160),
.C(n_143),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_148),
.B(n_143),
.C(n_145),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_151),
.B(n_134),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_162),
.B(n_158),
.C(n_64),
.Y(n_173)
);

AOI322xp5_ASAP7_75t_L g167 ( 
.A1(n_152),
.A2(n_142),
.A3(n_149),
.B1(n_129),
.B2(n_94),
.C1(n_130),
.C2(n_121),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_167),
.A2(n_158),
.B(n_161),
.Y(n_170)
);

MAJx2_ASAP7_75t_L g168 ( 
.A(n_159),
.B(n_142),
.C(n_116),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_168),
.B(n_160),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_169),
.B(n_173),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_170),
.A2(n_166),
.B1(n_82),
.B2(n_98),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_164),
.B(n_130),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_171),
.B(n_172),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_166),
.B(n_118),
.Y(n_172)
);

NOR3xp33_ASAP7_75t_SL g174 ( 
.A(n_173),
.B(n_163),
.C(n_165),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_174),
.B(n_82),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_177),
.B(n_175),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_178),
.B(n_179),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_176),
.A2(n_94),
.B(n_174),
.Y(n_179)
);

HB1xp67_ASAP7_75t_L g182 ( 
.A(n_180),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_182),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_183),
.B(n_181),
.Y(n_184)
);


endmodule