module real_aes_8861_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_503;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_578;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_725;
wire n_119;
wire n_310;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_363;
wire n_182;
wire n_449;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_552;
wire n_617;
wire n_602;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_741;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_175;
wire n_168;
wire n_241;
wire n_687;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g509 ( .A1(n_0), .A2(n_152), .B(n_510), .C(n_511), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_1), .B(n_171), .Y(n_513) );
NAND3xp33_ASAP7_75t_SL g106 ( .A(n_2), .B(n_107), .C(n_108), .Y(n_106) );
INVx1_ASAP7_75t_L g119 ( .A(n_2), .Y(n_119) );
A2O1A1Ixp33_ASAP7_75t_L g180 ( .A1(n_3), .A2(n_138), .B(n_143), .C(n_181), .Y(n_180) );
AOI21xp5_ASAP7_75t_L g229 ( .A1(n_4), .A2(n_133), .B(n_230), .Y(n_229) );
NAND2xp5_ASAP7_75t_SL g500 ( .A(n_5), .B(n_208), .Y(n_500) );
AOI21xp5_ASAP7_75t_L g454 ( .A1(n_6), .A2(n_133), .B(n_455), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_7), .B(n_171), .Y(n_237) );
AO21x2_ASAP7_75t_L g463 ( .A1(n_8), .A2(n_156), .B(n_464), .Y(n_463) );
AND2x6_ASAP7_75t_L g138 ( .A(n_9), .B(n_139), .Y(n_138) );
A2O1A1Ixp33_ASAP7_75t_L g520 ( .A1(n_10), .A2(n_138), .B(n_143), .C(n_521), .Y(n_520) );
INVx1_ASAP7_75t_L g150 ( .A(n_11), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g105 ( .A(n_12), .B(n_41), .Y(n_105) );
NOR2xp33_ASAP7_75t_L g120 ( .A(n_12), .B(n_41), .Y(n_120) );
NAND2xp5_ASAP7_75t_SL g185 ( .A(n_13), .B(n_148), .Y(n_185) );
INVx1_ASAP7_75t_L g131 ( .A(n_14), .Y(n_131) );
NAND2xp5_ASAP7_75t_SL g470 ( .A(n_15), .B(n_208), .Y(n_470) );
A2O1A1Ixp33_ASAP7_75t_L g164 ( .A1(n_16), .A2(n_151), .B(n_165), .C(n_169), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_17), .B(n_171), .Y(n_170) );
CKINVDCx20_ASAP7_75t_R g732 ( .A(n_18), .Y(n_732) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_19), .B(n_277), .Y(n_276) );
A2O1A1Ixp33_ASAP7_75t_L g194 ( .A1(n_20), .A2(n_195), .B(n_196), .C(n_198), .Y(n_194) );
A2O1A1Ixp33_ASAP7_75t_L g488 ( .A1(n_21), .A2(n_143), .B(n_212), .C(n_489), .Y(n_488) );
NAND2xp5_ASAP7_75t_SL g223 ( .A(n_22), .B(n_148), .Y(n_223) );
NAND2xp5_ASAP7_75t_SL g209 ( .A(n_23), .B(n_148), .Y(n_209) );
CKINVDCx16_ASAP7_75t_R g219 ( .A(n_24), .Y(n_219) );
INVx1_ASAP7_75t_L g207 ( .A(n_25), .Y(n_207) );
A2O1A1Ixp33_ASAP7_75t_L g466 ( .A1(n_26), .A2(n_143), .B(n_212), .C(n_467), .Y(n_466) );
BUFx6f_ASAP7_75t_L g137 ( .A(n_27), .Y(n_137) );
CKINVDCx20_ASAP7_75t_R g178 ( .A(n_28), .Y(n_178) );
INVx1_ASAP7_75t_L g273 ( .A(n_29), .Y(n_273) );
AOI21xp5_ASAP7_75t_L g506 ( .A1(n_30), .A2(n_133), .B(n_507), .Y(n_506) );
INVx2_ASAP7_75t_L g136 ( .A(n_31), .Y(n_136) );
A2O1A1Ixp33_ASAP7_75t_L g478 ( .A1(n_32), .A2(n_224), .B(n_445), .C(n_479), .Y(n_478) );
CKINVDCx20_ASAP7_75t_R g188 ( .A(n_33), .Y(n_188) );
A2O1A1Ixp33_ASAP7_75t_L g232 ( .A1(n_34), .A2(n_195), .B(n_233), .C(n_235), .Y(n_232) );
INVxp67_ASAP7_75t_L g274 ( .A(n_35), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_36), .B(n_469), .Y(n_468) );
A2O1A1Ixp33_ASAP7_75t_L g205 ( .A1(n_37), .A2(n_143), .B(n_206), .C(n_212), .Y(n_205) );
CKINVDCx14_ASAP7_75t_R g231 ( .A(n_38), .Y(n_231) );
OAI22xp5_ASAP7_75t_SL g739 ( .A1(n_39), .A2(n_46), .B1(n_740), .B2(n_741), .Y(n_739) );
INVx1_ASAP7_75t_L g740 ( .A(n_39), .Y(n_740) );
OAI22xp5_ASAP7_75t_L g723 ( .A1(n_40), .A2(n_45), .B1(n_724), .B2(n_725), .Y(n_723) );
INVx1_ASAP7_75t_L g725 ( .A(n_40), .Y(n_725) );
A2O1A1Ixp33_ASAP7_75t_L g146 ( .A1(n_42), .A2(n_147), .B(n_149), .C(n_152), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_43), .B(n_268), .Y(n_487) );
CKINVDCx20_ASAP7_75t_R g525 ( .A(n_44), .Y(n_525) );
CKINVDCx20_ASAP7_75t_R g724 ( .A(n_45), .Y(n_724) );
INVx1_ASAP7_75t_L g741 ( .A(n_46), .Y(n_741) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_47), .B(n_208), .Y(n_448) );
CKINVDCx20_ASAP7_75t_R g747 ( .A(n_48), .Y(n_747) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_49), .B(n_133), .Y(n_465) );
CKINVDCx20_ASAP7_75t_R g214 ( .A(n_50), .Y(n_214) );
CKINVDCx20_ASAP7_75t_R g270 ( .A(n_51), .Y(n_270) );
A2O1A1Ixp33_ASAP7_75t_L g444 ( .A1(n_52), .A2(n_224), .B(n_445), .C(n_446), .Y(n_444) );
INVx1_ASAP7_75t_L g512 ( .A(n_53), .Y(n_512) );
INVx1_ASAP7_75t_L g447 ( .A(n_54), .Y(n_447) );
INVx1_ASAP7_75t_L g193 ( .A(n_55), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_56), .B(n_133), .Y(n_443) );
CKINVDCx20_ASAP7_75t_R g493 ( .A(n_57), .Y(n_493) );
CKINVDCx14_ASAP7_75t_R g141 ( .A(n_58), .Y(n_141) );
AOI22xp33_ASAP7_75t_L g101 ( .A1(n_59), .A2(n_102), .B1(n_111), .B2(n_750), .Y(n_101) );
INVx1_ASAP7_75t_L g139 ( .A(n_60), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_61), .B(n_133), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_62), .B(n_171), .Y(n_461) );
A2O1A1Ixp33_ASAP7_75t_L g457 ( .A1(n_63), .A2(n_211), .B(n_458), .C(n_459), .Y(n_457) );
INVx1_ASAP7_75t_L g130 ( .A(n_64), .Y(n_130) );
INVx1_ASAP7_75t_SL g234 ( .A(n_65), .Y(n_234) );
CKINVDCx20_ASAP7_75t_R g735 ( .A(n_66), .Y(n_735) );
NAND2xp5_ASAP7_75t_SL g481 ( .A(n_67), .B(n_208), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_68), .B(n_171), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_69), .B(n_151), .Y(n_522) );
INVx1_ASAP7_75t_L g222 ( .A(n_70), .Y(n_222) );
CKINVDCx16_ASAP7_75t_R g508 ( .A(n_71), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_72), .B(n_184), .Y(n_490) );
A2O1A1Ixp33_ASAP7_75t_L g497 ( .A1(n_73), .A2(n_143), .B(n_224), .C(n_498), .Y(n_497) );
CKINVDCx16_ASAP7_75t_R g456 ( .A(n_74), .Y(n_456) );
INVx1_ASAP7_75t_L g110 ( .A(n_75), .Y(n_110) );
AOI21xp5_ASAP7_75t_L g132 ( .A1(n_76), .A2(n_133), .B(n_140), .Y(n_132) );
CKINVDCx20_ASAP7_75t_R g226 ( .A(n_77), .Y(n_226) );
AOI21xp5_ASAP7_75t_L g161 ( .A1(n_78), .A2(n_133), .B(n_162), .Y(n_161) );
AOI21xp5_ASAP7_75t_L g267 ( .A1(n_79), .A2(n_268), .B(n_269), .Y(n_267) );
INVx1_ASAP7_75t_L g163 ( .A(n_80), .Y(n_163) );
CKINVDCx16_ASAP7_75t_R g204 ( .A(n_81), .Y(n_204) );
NAND2xp5_ASAP7_75t_SL g491 ( .A(n_82), .B(n_183), .Y(n_491) );
CKINVDCx20_ASAP7_75t_R g483 ( .A(n_83), .Y(n_483) );
AOI21xp5_ASAP7_75t_L g191 ( .A1(n_84), .A2(n_133), .B(n_192), .Y(n_191) );
INVx1_ASAP7_75t_L g166 ( .A(n_85), .Y(n_166) );
INVx2_ASAP7_75t_L g128 ( .A(n_86), .Y(n_128) );
INVx1_ASAP7_75t_L g182 ( .A(n_87), .Y(n_182) );
CKINVDCx20_ASAP7_75t_R g504 ( .A(n_88), .Y(n_504) );
NAND2xp5_ASAP7_75t_SL g523 ( .A(n_89), .B(n_148), .Y(n_523) );
INVx2_ASAP7_75t_L g107 ( .A(n_90), .Y(n_107) );
OR2x2_ASAP7_75t_L g436 ( .A(n_90), .B(n_118), .Y(n_436) );
OR2x2_ASAP7_75t_L g743 ( .A(n_90), .B(n_731), .Y(n_743) );
A2O1A1Ixp33_ASAP7_75t_L g220 ( .A1(n_91), .A2(n_143), .B(n_221), .C(n_224), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_92), .B(n_133), .Y(n_477) );
INVx1_ASAP7_75t_L g480 ( .A(n_93), .Y(n_480) );
INVxp67_ASAP7_75t_L g460 ( .A(n_94), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_95), .B(n_156), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_96), .B(n_110), .Y(n_109) );
INVx2_ASAP7_75t_L g197 ( .A(n_97), .Y(n_197) );
INVx1_ASAP7_75t_L g499 ( .A(n_98), .Y(n_499) );
INVx1_ASAP7_75t_L g519 ( .A(n_99), .Y(n_519) );
AND2x2_ASAP7_75t_L g450 ( .A(n_100), .B(n_127), .Y(n_450) );
INVx1_ASAP7_75t_SL g102 ( .A(n_103), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
INVx1_ASAP7_75t_SL g750 ( .A(n_104), .Y(n_750) );
NOR2xp33_ASAP7_75t_L g104 ( .A(n_105), .B(n_106), .Y(n_104) );
OR2x2_ASAP7_75t_L g117 ( .A(n_107), .B(n_118), .Y(n_117) );
NOR2x2_ASAP7_75t_L g730 ( .A(n_107), .B(n_731), .Y(n_730) );
INVx1_ASAP7_75t_SL g108 ( .A(n_109), .Y(n_108) );
AO221x1_ASAP7_75t_L g111 ( .A1(n_112), .A2(n_733), .B1(n_736), .B2(n_744), .C(n_746), .Y(n_111) );
OAI222xp33_ASAP7_75t_L g112 ( .A1(n_113), .A2(n_722), .B1(n_723), .B2(n_726), .C1(n_729), .C2(n_732), .Y(n_112) );
AOI22xp5_ASAP7_75t_L g113 ( .A1(n_114), .A2(n_121), .B1(n_433), .B2(n_437), .Y(n_113) );
AOI22x1_ASAP7_75t_SL g726 ( .A1(n_114), .A2(n_433), .B1(n_727), .B2(n_728), .Y(n_726) );
INVx1_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
INVx2_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
INVx2_ASAP7_75t_L g731 ( .A(n_118), .Y(n_731) );
AND2x2_ASAP7_75t_L g118 ( .A(n_119), .B(n_120), .Y(n_118) );
INVx2_ASAP7_75t_L g727 ( .A(n_121), .Y(n_727) );
OR2x2_ASAP7_75t_L g121 ( .A(n_122), .B(n_363), .Y(n_121) );
NAND5xp2_ASAP7_75t_L g122 ( .A(n_123), .B(n_278), .C(n_310), .D(n_327), .E(n_350), .Y(n_122) );
AOI221xp5_ASAP7_75t_L g123 ( .A1(n_124), .A2(n_201), .B1(n_238), .B2(n_242), .C(n_246), .Y(n_123) );
INVx1_ASAP7_75t_L g390 ( .A(n_124), .Y(n_390) );
AND2x2_ASAP7_75t_L g124 ( .A(n_125), .B(n_173), .Y(n_124) );
AND3x2_ASAP7_75t_L g365 ( .A(n_125), .B(n_175), .C(n_366), .Y(n_365) );
AND2x2_ASAP7_75t_L g125 ( .A(n_126), .B(n_158), .Y(n_125) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_126), .B(n_244), .Y(n_243) );
BUFx3_ASAP7_75t_L g253 ( .A(n_126), .Y(n_253) );
AND2x2_ASAP7_75t_L g257 ( .A(n_126), .B(n_189), .Y(n_257) );
INVx2_ASAP7_75t_L g287 ( .A(n_126), .Y(n_287) );
OR2x2_ASAP7_75t_L g298 ( .A(n_126), .B(n_190), .Y(n_298) );
NOR2xp33_ASAP7_75t_L g317 ( .A(n_126), .B(n_174), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_126), .B(n_336), .Y(n_335) );
AND2x2_ASAP7_75t_L g377 ( .A(n_126), .B(n_190), .Y(n_377) );
OA21x2_ASAP7_75t_L g126 ( .A1(n_127), .A2(n_132), .B(n_155), .Y(n_126) );
INVx1_ASAP7_75t_L g176 ( .A(n_127), .Y(n_176) );
O2A1O1Ixp33_ASAP7_75t_L g203 ( .A1(n_127), .A2(n_179), .B(n_204), .C(n_205), .Y(n_203) );
INVx2_ASAP7_75t_L g227 ( .A(n_127), .Y(n_227) );
AOI21xp5_ASAP7_75t_L g442 ( .A1(n_127), .A2(n_443), .B(n_444), .Y(n_442) );
AOI21xp5_ASAP7_75t_L g476 ( .A1(n_127), .A2(n_477), .B(n_478), .Y(n_476) );
AND2x2_ASAP7_75t_SL g127 ( .A(n_128), .B(n_129), .Y(n_127) );
AND2x2_ASAP7_75t_L g157 ( .A(n_128), .B(n_129), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g129 ( .A(n_130), .B(n_131), .Y(n_129) );
BUFx2_ASAP7_75t_L g268 ( .A(n_133), .Y(n_268) );
AND2x4_ASAP7_75t_L g133 ( .A(n_134), .B(n_138), .Y(n_133) );
NAND2x1p5_ASAP7_75t_L g179 ( .A(n_134), .B(n_138), .Y(n_179) );
AND2x2_ASAP7_75t_L g134 ( .A(n_135), .B(n_137), .Y(n_134) );
INVx1_ASAP7_75t_L g211 ( .A(n_135), .Y(n_211) );
INVx1_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
INVx2_ASAP7_75t_L g144 ( .A(n_136), .Y(n_144) );
INVx1_ASAP7_75t_L g199 ( .A(n_136), .Y(n_199) );
INVx1_ASAP7_75t_L g145 ( .A(n_137), .Y(n_145) );
BUFx6f_ASAP7_75t_L g148 ( .A(n_137), .Y(n_148) );
INVx3_ASAP7_75t_L g151 ( .A(n_137), .Y(n_151) );
BUFx6f_ASAP7_75t_L g168 ( .A(n_137), .Y(n_168) );
INVx1_ASAP7_75t_L g469 ( .A(n_137), .Y(n_469) );
INVx4_ASAP7_75t_SL g154 ( .A(n_138), .Y(n_154) );
BUFx3_ASAP7_75t_L g212 ( .A(n_138), .Y(n_212) );
O2A1O1Ixp33_ASAP7_75t_SL g140 ( .A1(n_141), .A2(n_142), .B(n_146), .C(n_154), .Y(n_140) );
O2A1O1Ixp33_ASAP7_75t_SL g162 ( .A1(n_142), .A2(n_154), .B(n_163), .C(n_164), .Y(n_162) );
O2A1O1Ixp33_ASAP7_75t_SL g192 ( .A1(n_142), .A2(n_154), .B(n_193), .C(n_194), .Y(n_192) );
O2A1O1Ixp33_ASAP7_75t_L g230 ( .A1(n_142), .A2(n_154), .B(n_231), .C(n_232), .Y(n_230) );
O2A1O1Ixp33_ASAP7_75t_SL g269 ( .A1(n_142), .A2(n_154), .B(n_270), .C(n_271), .Y(n_269) );
INVx2_ASAP7_75t_L g445 ( .A(n_142), .Y(n_445) );
O2A1O1Ixp33_ASAP7_75t_L g455 ( .A1(n_142), .A2(n_154), .B(n_456), .C(n_457), .Y(n_455) );
O2A1O1Ixp33_ASAP7_75t_SL g507 ( .A1(n_142), .A2(n_154), .B(n_508), .C(n_509), .Y(n_507) );
INVx5_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
AND2x6_ASAP7_75t_L g143 ( .A(n_144), .B(n_145), .Y(n_143) );
BUFx3_ASAP7_75t_L g153 ( .A(n_144), .Y(n_153) );
BUFx6f_ASAP7_75t_L g236 ( .A(n_144), .Y(n_236) );
INVx2_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx4_ASAP7_75t_L g195 ( .A(n_148), .Y(n_195) );
NOR2xp33_ASAP7_75t_L g149 ( .A(n_150), .B(n_151), .Y(n_149) );
INVx5_ASAP7_75t_L g208 ( .A(n_151), .Y(n_208) );
INVx2_ASAP7_75t_L g186 ( .A(n_152), .Y(n_186) );
INVx2_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx1_ASAP7_75t_L g169 ( .A(n_153), .Y(n_169) );
HB1xp67_ASAP7_75t_L g449 ( .A(n_153), .Y(n_449) );
INVx1_ASAP7_75t_L g224 ( .A(n_154), .Y(n_224) );
HB1xp67_ASAP7_75t_L g160 ( .A(n_156), .Y(n_160) );
INVx4_ASAP7_75t_L g172 ( .A(n_156), .Y(n_172) );
AOI21xp5_ASAP7_75t_L g464 ( .A1(n_156), .A2(n_465), .B(n_466), .Y(n_464) );
BUFx6f_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVx1_ASAP7_75t_L g265 ( .A(n_157), .Y(n_265) );
HB1xp67_ASAP7_75t_L g256 ( .A(n_158), .Y(n_256) );
AND2x2_ASAP7_75t_L g318 ( .A(n_158), .B(n_319), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_158), .B(n_174), .Y(n_337) );
INVx1_ASAP7_75t_SL g158 ( .A(n_159), .Y(n_158) );
OR2x2_ASAP7_75t_L g245 ( .A(n_159), .B(n_174), .Y(n_245) );
HB1xp67_ASAP7_75t_L g252 ( .A(n_159), .Y(n_252) );
AND2x2_ASAP7_75t_L g304 ( .A(n_159), .B(n_190), .Y(n_304) );
NAND3xp33_ASAP7_75t_L g329 ( .A(n_159), .B(n_173), .C(n_287), .Y(n_329) );
AND2x2_ASAP7_75t_L g394 ( .A(n_159), .B(n_175), .Y(n_394) );
AND2x2_ASAP7_75t_L g428 ( .A(n_159), .B(n_174), .Y(n_428) );
OA21x2_ASAP7_75t_L g159 ( .A1(n_160), .A2(n_161), .B(n_170), .Y(n_159) );
OA21x2_ASAP7_75t_L g190 ( .A1(n_160), .A2(n_191), .B(n_200), .Y(n_190) );
OA21x2_ASAP7_75t_L g228 ( .A1(n_160), .A2(n_229), .B(n_237), .Y(n_228) );
OA21x2_ASAP7_75t_L g453 ( .A1(n_160), .A2(n_454), .B(n_461), .Y(n_453) );
NOR2xp33_ASAP7_75t_L g165 ( .A(n_166), .B(n_167), .Y(n_165) );
NOR2xp33_ASAP7_75t_L g196 ( .A(n_167), .B(n_197), .Y(n_196) );
OAI22xp33_ASAP7_75t_L g272 ( .A1(n_167), .A2(n_208), .B1(n_273), .B2(n_274), .Y(n_272) );
INVx1_ASAP7_75t_L g458 ( .A(n_167), .Y(n_458) );
INVx4_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
INVx2_ASAP7_75t_L g184 ( .A(n_168), .Y(n_184) );
OA21x2_ASAP7_75t_L g505 ( .A1(n_171), .A2(n_506), .B(n_513), .Y(n_505) );
INVx3_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
NOR2xp33_ASAP7_75t_L g187 ( .A(n_172), .B(n_188), .Y(n_187) );
NOR2xp33_ASAP7_75t_L g213 ( .A(n_172), .B(n_214), .Y(n_213) );
AO21x2_ASAP7_75t_L g217 ( .A1(n_172), .A2(n_218), .B(n_225), .Y(n_217) );
NOR2xp33_ASAP7_75t_L g482 ( .A(n_172), .B(n_483), .Y(n_482) );
AO21x2_ASAP7_75t_L g495 ( .A1(n_172), .A2(n_496), .B(n_503), .Y(n_495) );
NOR2xp33_ASAP7_75t_L g503 ( .A(n_172), .B(n_504), .Y(n_503) );
AO21x2_ASAP7_75t_L g517 ( .A1(n_172), .A2(n_518), .B(n_524), .Y(n_517) );
INVxp67_ASAP7_75t_L g254 ( .A(n_173), .Y(n_254) );
AND2x2_ASAP7_75t_L g173 ( .A(n_174), .B(n_189), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_174), .B(n_287), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_174), .B(n_318), .Y(n_326) );
AND2x2_ASAP7_75t_L g376 ( .A(n_174), .B(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g404 ( .A(n_174), .Y(n_404) );
INVx4_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
AND2x2_ASAP7_75t_L g311 ( .A(n_175), .B(n_304), .Y(n_311) );
BUFx3_ASAP7_75t_L g343 ( .A(n_175), .Y(n_343) );
AO21x2_ASAP7_75t_L g175 ( .A1(n_176), .A2(n_177), .B(n_187), .Y(n_175) );
NOR2xp33_ASAP7_75t_L g492 ( .A(n_176), .B(n_493), .Y(n_492) );
OAI21xp5_ASAP7_75t_L g177 ( .A1(n_178), .A2(n_179), .B(n_180), .Y(n_177) );
OAI21xp5_ASAP7_75t_L g218 ( .A1(n_179), .A2(n_219), .B(n_220), .Y(n_218) );
OAI21xp5_ASAP7_75t_L g518 ( .A1(n_179), .A2(n_519), .B(n_520), .Y(n_518) );
O2A1O1Ixp5_ASAP7_75t_L g181 ( .A1(n_182), .A2(n_183), .B(n_185), .C(n_186), .Y(n_181) );
O2A1O1Ixp33_ASAP7_75t_L g221 ( .A1(n_183), .A2(n_186), .B(n_222), .C(n_223), .Y(n_221) );
O2A1O1Ixp33_ASAP7_75t_L g446 ( .A1(n_183), .A2(n_447), .B(n_448), .C(n_449), .Y(n_446) );
O2A1O1Ixp33_ASAP7_75t_L g479 ( .A1(n_183), .A2(n_449), .B(n_480), .C(n_481), .Y(n_479) );
INVx2_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
INVx2_ASAP7_75t_L g319 ( .A(n_189), .Y(n_319) );
INVx2_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
HB1xp67_ASAP7_75t_L g288 ( .A(n_190), .Y(n_288) );
NOR2xp33_ASAP7_75t_L g233 ( .A(n_195), .B(n_234), .Y(n_233) );
NOR2xp33_ASAP7_75t_L g511 ( .A(n_195), .B(n_512), .Y(n_511) );
INVx2_ASAP7_75t_L g471 ( .A(n_198), .Y(n_471) );
INVx3_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
AOI22xp33_ASAP7_75t_L g378 ( .A1(n_201), .A2(n_379), .B1(n_381), .B2(n_382), .Y(n_378) );
AND2x2_ASAP7_75t_L g201 ( .A(n_202), .B(n_215), .Y(n_201) );
AND2x2_ASAP7_75t_L g238 ( .A(n_202), .B(n_239), .Y(n_238) );
INVx3_ASAP7_75t_SL g249 ( .A(n_202), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_202), .B(n_282), .Y(n_314) );
OR2x2_ASAP7_75t_L g333 ( .A(n_202), .B(n_216), .Y(n_333) );
AND2x2_ASAP7_75t_L g338 ( .A(n_202), .B(n_290), .Y(n_338) );
AND2x2_ASAP7_75t_L g341 ( .A(n_202), .B(n_283), .Y(n_341) );
AND2x2_ASAP7_75t_L g353 ( .A(n_202), .B(n_228), .Y(n_353) );
AND2x2_ASAP7_75t_L g369 ( .A(n_202), .B(n_217), .Y(n_369) );
AND2x4_ASAP7_75t_L g372 ( .A(n_202), .B(n_240), .Y(n_372) );
OR2x2_ASAP7_75t_L g389 ( .A(n_202), .B(n_325), .Y(n_389) );
OR2x2_ASAP7_75t_L g420 ( .A(n_202), .B(n_262), .Y(n_420) );
NAND2xp5_ASAP7_75t_SL g422 ( .A(n_202), .B(n_348), .Y(n_422) );
OR2x6_ASAP7_75t_L g202 ( .A(n_203), .B(n_213), .Y(n_202) );
O2A1O1Ixp33_ASAP7_75t_L g206 ( .A1(n_207), .A2(n_208), .B(n_209), .C(n_210), .Y(n_206) );
NOR2xp33_ASAP7_75t_L g459 ( .A(n_208), .B(n_460), .Y(n_459) );
INVx2_ASAP7_75t_L g510 ( .A(n_208), .Y(n_510) );
AOI21xp5_ASAP7_75t_L g489 ( .A1(n_210), .A2(n_490), .B(n_491), .Y(n_489) );
INVx2_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
NAND2xp5_ASAP7_75t_SL g271 ( .A(n_211), .B(n_272), .Y(n_271) );
AND2x2_ASAP7_75t_L g296 ( .A(n_215), .B(n_260), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_215), .B(n_283), .Y(n_415) );
AND2x2_ASAP7_75t_L g215 ( .A(n_216), .B(n_228), .Y(n_215) );
AND2x2_ASAP7_75t_L g248 ( .A(n_216), .B(n_249), .Y(n_248) );
AND2x2_ASAP7_75t_L g282 ( .A(n_216), .B(n_283), .Y(n_282) );
AND2x2_ASAP7_75t_L g290 ( .A(n_216), .B(n_262), .Y(n_290) );
AND2x2_ASAP7_75t_L g308 ( .A(n_216), .B(n_240), .Y(n_308) );
OR2x2_ASAP7_75t_L g325 ( .A(n_216), .B(n_283), .Y(n_325) );
INVx2_ASAP7_75t_SL g216 ( .A(n_217), .Y(n_216) );
BUFx2_ASAP7_75t_L g241 ( .A(n_217), .Y(n_241) );
AND2x2_ASAP7_75t_L g348 ( .A(n_217), .B(n_228), .Y(n_348) );
NOR2xp33_ASAP7_75t_L g225 ( .A(n_226), .B(n_227), .Y(n_225) );
INVx1_ASAP7_75t_L g277 ( .A(n_227), .Y(n_277) );
INVx2_ASAP7_75t_L g240 ( .A(n_228), .Y(n_240) );
INVx1_ASAP7_75t_L g360 ( .A(n_228), .Y(n_360) );
AND2x2_ASAP7_75t_L g410 ( .A(n_228), .B(n_249), .Y(n_410) );
INVx3_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
HB1xp67_ASAP7_75t_L g501 ( .A(n_236), .Y(n_501) );
AND2x2_ASAP7_75t_L g259 ( .A(n_239), .B(n_260), .Y(n_259) );
AND2x2_ASAP7_75t_L g294 ( .A(n_239), .B(n_249), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_239), .B(n_341), .Y(n_340) );
AND2x2_ASAP7_75t_L g239 ( .A(n_240), .B(n_241), .Y(n_239) );
AND2x2_ASAP7_75t_L g281 ( .A(n_240), .B(n_249), .Y(n_281) );
OR2x2_ASAP7_75t_L g397 ( .A(n_241), .B(n_371), .Y(n_397) );
INVx1_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_244), .B(n_377), .Y(n_383) );
INVx2_ASAP7_75t_SL g244 ( .A(n_245), .Y(n_244) );
OAI32xp33_ASAP7_75t_L g339 ( .A1(n_245), .A2(n_340), .A3(n_342), .B1(n_344), .B2(n_345), .Y(n_339) );
OR2x2_ASAP7_75t_L g356 ( .A(n_245), .B(n_298), .Y(n_356) );
OAI21xp33_ASAP7_75t_SL g381 ( .A1(n_245), .A2(n_255), .B(n_286), .Y(n_381) );
OAI22xp33_ASAP7_75t_L g246 ( .A1(n_247), .A2(n_250), .B1(n_255), .B2(n_258), .Y(n_246) );
INVxp33_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_248), .B(n_322), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_249), .B(n_290), .Y(n_289) );
AND2x2_ASAP7_75t_L g307 ( .A(n_249), .B(n_308), .Y(n_307) );
AND2x2_ASAP7_75t_L g407 ( .A(n_249), .B(n_348), .Y(n_407) );
OR2x2_ASAP7_75t_L g431 ( .A(n_249), .B(n_325), .Y(n_431) );
AOI21xp33_ASAP7_75t_L g414 ( .A1(n_250), .A2(n_313), .B(n_415), .Y(n_414) );
OR2x2_ASAP7_75t_L g250 ( .A(n_251), .B(n_254), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_252), .B(n_253), .Y(n_251) );
INVx1_ASAP7_75t_L g291 ( .A(n_252), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_252), .B(n_257), .Y(n_309) );
AND2x2_ASAP7_75t_L g331 ( .A(n_253), .B(n_304), .Y(n_331) );
INVx1_ASAP7_75t_L g344 ( .A(n_253), .Y(n_344) );
OR2x2_ASAP7_75t_L g349 ( .A(n_253), .B(n_283), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_256), .B(n_257), .Y(n_255) );
NOR2xp33_ASAP7_75t_L g297 ( .A(n_256), .B(n_298), .Y(n_297) );
OAI22xp33_ASAP7_75t_L g279 ( .A1(n_257), .A2(n_280), .B1(n_285), .B2(n_289), .Y(n_279) );
INVx1_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
OAI22xp5_ASAP7_75t_L g328 ( .A1(n_260), .A2(n_322), .B1(n_329), .B2(n_330), .Y(n_328) );
AND2x2_ASAP7_75t_L g406 ( .A(n_260), .B(n_407), .Y(n_406) );
INVx2_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
INVx1_ASAP7_75t_SL g261 ( .A(n_262), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_262), .B(n_360), .Y(n_359) );
AND2x2_ASAP7_75t_L g425 ( .A(n_262), .B(n_308), .Y(n_425) );
AO21x2_ASAP7_75t_L g262 ( .A1(n_263), .A2(n_266), .B(n_275), .Y(n_262) );
INVx1_ASAP7_75t_L g284 ( .A(n_263), .Y(n_284) );
INVx1_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
INVx2_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
NOR2xp33_ASAP7_75t_L g524 ( .A(n_265), .B(n_525), .Y(n_524) );
INVx1_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
OA21x2_ASAP7_75t_L g283 ( .A1(n_267), .A2(n_276), .B(n_284), .Y(n_283) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
AOI21xp5_ASAP7_75t_SL g486 ( .A1(n_277), .A2(n_487), .B(n_488), .Y(n_486) );
AOI221xp5_ASAP7_75t_L g278 ( .A1(n_279), .A2(n_291), .B1(n_292), .B2(n_297), .C(n_299), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_281), .B(n_282), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_281), .B(n_283), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_281), .B(n_324), .Y(n_323) );
INVx1_ASAP7_75t_L g300 ( .A(n_282), .Y(n_300) );
O2A1O1Ixp33_ASAP7_75t_L g387 ( .A1(n_282), .A2(n_388), .B(n_389), .C(n_390), .Y(n_387) );
AND2x2_ASAP7_75t_L g392 ( .A(n_282), .B(n_372), .Y(n_392) );
O2A1O1Ixp33_ASAP7_75t_SL g430 ( .A1(n_282), .A2(n_371), .B(n_431), .C(n_432), .Y(n_430) );
BUFx3_ASAP7_75t_L g322 ( .A(n_283), .Y(n_322) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_286), .B(n_343), .Y(n_386) );
AOI211xp5_ASAP7_75t_L g405 ( .A1(n_286), .A2(n_406), .B(n_408), .C(n_414), .Y(n_405) );
AND2x2_ASAP7_75t_L g286 ( .A(n_287), .B(n_288), .Y(n_286) );
INVxp67_ASAP7_75t_L g366 ( .A(n_288), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_290), .B(n_410), .Y(n_409) );
NAND2xp5_ASAP7_75t_SL g292 ( .A(n_293), .B(n_295), .Y(n_292) );
INVx1_ASAP7_75t_SL g293 ( .A(n_294), .Y(n_293) );
AOI211xp5_ASAP7_75t_L g310 ( .A1(n_294), .A2(n_311), .B(n_312), .C(n_320), .Y(n_310) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
INVx1_ASAP7_75t_L g395 ( .A(n_298), .Y(n_395) );
OR2x2_ASAP7_75t_L g412 ( .A(n_298), .B(n_342), .Y(n_412) );
OAI22xp5_ASAP7_75t_L g299 ( .A1(n_300), .A2(n_301), .B1(n_306), .B2(n_309), .Y(n_299) );
OAI22xp33_ASAP7_75t_L g312 ( .A1(n_301), .A2(n_313), .B1(n_314), .B2(n_315), .Y(n_312) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
NOR2xp33_ASAP7_75t_L g302 ( .A(n_303), .B(n_305), .Y(n_302) );
OR2x2_ASAP7_75t_L g399 ( .A(n_303), .B(n_343), .Y(n_399) );
INVx1_ASAP7_75t_SL g303 ( .A(n_304), .Y(n_303) );
AND2x2_ASAP7_75t_L g354 ( .A(n_304), .B(n_344), .Y(n_354) );
INVx1_ASAP7_75t_L g362 ( .A(n_305), .Y(n_362) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_308), .B(n_322), .Y(n_370) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
AND2x2_ASAP7_75t_L g316 ( .A(n_317), .B(n_318), .Y(n_316) );
NAND2xp5_ASAP7_75t_SL g361 ( .A(n_318), .B(n_362), .Y(n_361) );
INVx2_ASAP7_75t_L g427 ( .A(n_319), .Y(n_427) );
AOI21xp33_ASAP7_75t_L g320 ( .A1(n_321), .A2(n_323), .B(n_326), .Y(n_320) );
INVx1_ASAP7_75t_L g357 ( .A(n_321), .Y(n_357) );
NAND2xp5_ASAP7_75t_SL g332 ( .A(n_322), .B(n_333), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_322), .B(n_353), .Y(n_352) );
NAND2x1p5_ASAP7_75t_L g373 ( .A(n_322), .B(n_348), .Y(n_373) );
NAND2xp5_ASAP7_75t_SL g380 ( .A(n_322), .B(n_369), .Y(n_380) );
OAI211xp5_ASAP7_75t_L g384 ( .A1(n_322), .A2(n_332), .B(n_372), .C(n_385), .Y(n_384) );
INVx1_ASAP7_75t_SL g324 ( .A(n_325), .Y(n_324) );
AOI221xp5_ASAP7_75t_SL g327 ( .A1(n_328), .A2(n_332), .B1(n_334), .B2(n_338), .C(n_339), .Y(n_327) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
INVxp67_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_336), .B(n_344), .Y(n_418) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
O2A1O1Ixp33_ASAP7_75t_L g429 ( .A1(n_338), .A2(n_353), .B(n_355), .C(n_430), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_341), .B(n_348), .Y(n_413) );
NAND2xp5_ASAP7_75t_SL g432 ( .A(n_342), .B(n_395), .Y(n_432) );
CKINVDCx16_ASAP7_75t_R g342 ( .A(n_343), .Y(n_342) );
INVxp33_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
NOR2xp33_ASAP7_75t_L g346 ( .A(n_347), .B(n_349), .Y(n_346) );
AOI21xp33_ASAP7_75t_SL g358 ( .A1(n_347), .A2(n_359), .B(n_361), .Y(n_358) );
NOR2xp33_ASAP7_75t_L g419 ( .A(n_347), .B(n_420), .Y(n_419) );
INVx2_ASAP7_75t_SL g347 ( .A(n_348), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_348), .B(n_402), .Y(n_401) );
AOI221xp5_ASAP7_75t_L g350 ( .A1(n_351), .A2(n_354), .B1(n_355), .B2(n_357), .C(n_358), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_354), .B(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
INVx1_ASAP7_75t_L g388 ( .A(n_360), .Y(n_388) );
NAND5xp2_ASAP7_75t_L g363 ( .A(n_364), .B(n_391), .C(n_405), .D(n_416), .E(n_429), .Y(n_363) );
AOI211xp5_ASAP7_75t_L g364 ( .A1(n_365), .A2(n_367), .B(n_374), .C(n_387), .Y(n_364) );
INVx2_ASAP7_75t_SL g411 ( .A(n_365), .Y(n_411) );
NAND4xp25_ASAP7_75t_SL g367 ( .A(n_368), .B(n_370), .C(n_371), .D(n_373), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVx3_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
OAI211xp5_ASAP7_75t_SL g374 ( .A1(n_373), .A2(n_375), .B(n_378), .C(n_384), .Y(n_374) );
CKINVDCx20_ASAP7_75t_R g375 ( .A(n_376), .Y(n_375) );
AOI221xp5_ASAP7_75t_L g416 ( .A1(n_376), .A2(n_417), .B1(n_419), .B2(n_421), .C(n_423), .Y(n_416) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
AOI221xp5_ASAP7_75t_SL g391 ( .A1(n_392), .A2(n_393), .B1(n_396), .B2(n_398), .C(n_400), .Y(n_391) );
AND2x2_ASAP7_75t_L g393 ( .A(n_394), .B(n_395), .Y(n_393) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
OAI22xp5_ASAP7_75t_L g423 ( .A1(n_399), .A2(n_422), .B1(n_424), .B2(n_426), .Y(n_423) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx1_ASAP7_75t_SL g402 ( .A(n_403), .Y(n_402) );
OAI22xp5_ASAP7_75t_L g408 ( .A1(n_409), .A2(n_411), .B1(n_412), .B2(n_413), .Y(n_408) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx1_ASAP7_75t_SL g424 ( .A(n_425), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_427), .B(n_428), .Y(n_426) );
INVx1_ASAP7_75t_SL g433 ( .A(n_434), .Y(n_433) );
INVx2_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx4_ASAP7_75t_L g728 ( .A(n_437), .Y(n_728) );
XOR2xp5_ASAP7_75t_L g738 ( .A(n_437), .B(n_739), .Y(n_738) );
BUFx6f_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
OR5x1_ASAP7_75t_L g438 ( .A(n_439), .B(n_595), .C(n_673), .D(n_697), .E(n_714), .Y(n_438) );
OAI211xp5_ASAP7_75t_SL g439 ( .A1(n_440), .A2(n_472), .B(n_514), .C(n_572), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_441), .B(n_451), .Y(n_440) );
AND2x2_ASAP7_75t_L g526 ( .A(n_441), .B(n_453), .Y(n_526) );
INVx5_ASAP7_75t_SL g554 ( .A(n_441), .Y(n_554) );
AND2x2_ASAP7_75t_L g590 ( .A(n_441), .B(n_575), .Y(n_590) );
OR2x2_ASAP7_75t_L g629 ( .A(n_441), .B(n_452), .Y(n_629) );
OR2x2_ASAP7_75t_L g660 ( .A(n_441), .B(n_551), .Y(n_660) );
NOR2xp33_ASAP7_75t_L g696 ( .A(n_441), .B(n_564), .Y(n_696) );
AND2x2_ASAP7_75t_L g708 ( .A(n_441), .B(n_551), .Y(n_708) );
OR2x6_ASAP7_75t_L g441 ( .A(n_442), .B(n_450), .Y(n_441) );
AND2x2_ASAP7_75t_L g707 ( .A(n_451), .B(n_708), .Y(n_707) );
INVx1_ASAP7_75t_SL g451 ( .A(n_452), .Y(n_451) );
OR2x2_ASAP7_75t_L g570 ( .A(n_452), .B(n_571), .Y(n_570) );
OR2x2_ASAP7_75t_L g452 ( .A(n_453), .B(n_462), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_453), .B(n_551), .Y(n_550) );
HB1xp67_ASAP7_75t_L g563 ( .A(n_453), .Y(n_563) );
INVx3_ASAP7_75t_L g578 ( .A(n_453), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_453), .B(n_462), .Y(n_602) );
OR2x2_ASAP7_75t_L g611 ( .A(n_453), .B(n_554), .Y(n_611) );
AND2x2_ASAP7_75t_L g615 ( .A(n_453), .B(n_575), .Y(n_615) );
AND2x2_ASAP7_75t_L g621 ( .A(n_453), .B(n_622), .Y(n_621) );
INVxp67_ASAP7_75t_L g658 ( .A(n_453), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_453), .B(n_517), .Y(n_672) );
O2A1O1Ixp33_ASAP7_75t_L g498 ( .A1(n_458), .A2(n_499), .B(n_500), .C(n_501), .Y(n_498) );
OR2x2_ASAP7_75t_L g564 ( .A(n_462), .B(n_517), .Y(n_564) );
AND2x2_ASAP7_75t_L g575 ( .A(n_462), .B(n_551), .Y(n_575) );
AND2x2_ASAP7_75t_L g587 ( .A(n_462), .B(n_578), .Y(n_587) );
NAND2xp5_ASAP7_75t_SL g610 ( .A(n_462), .B(n_517), .Y(n_610) );
INVx1_ASAP7_75t_SL g622 ( .A(n_462), .Y(n_622) );
INVx2_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
AND2x2_ASAP7_75t_L g516 ( .A(n_463), .B(n_517), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_463), .B(n_554), .Y(n_553) );
AOI21xp5_ASAP7_75t_L g467 ( .A1(n_468), .A2(n_470), .B(n_471), .Y(n_467) );
AOI21xp5_ASAP7_75t_L g521 ( .A1(n_471), .A2(n_522), .B(n_523), .Y(n_521) );
INVx1_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
AND2x2_ASAP7_75t_L g473 ( .A(n_474), .B(n_484), .Y(n_473) );
AND2x2_ASAP7_75t_L g535 ( .A(n_474), .B(n_536), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_474), .B(n_494), .Y(n_539) );
AND2x2_ASAP7_75t_L g542 ( .A(n_474), .B(n_543), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_474), .B(n_545), .Y(n_544) );
OR2x2_ASAP7_75t_L g567 ( .A(n_474), .B(n_558), .Y(n_567) );
HB1xp67_ASAP7_75t_L g586 ( .A(n_474), .Y(n_586) );
AND2x2_ASAP7_75t_L g607 ( .A(n_474), .B(n_608), .Y(n_607) );
OR2x2_ASAP7_75t_L g617 ( .A(n_474), .B(n_618), .Y(n_617) );
AND2x2_ASAP7_75t_L g663 ( .A(n_474), .B(n_546), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_474), .B(n_569), .Y(n_690) );
INVx5_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
BUFx2_ASAP7_75t_L g560 ( .A(n_475), .Y(n_560) );
AND2x2_ASAP7_75t_L g626 ( .A(n_475), .B(n_558), .Y(n_626) );
AND2x2_ASAP7_75t_L g710 ( .A(n_475), .B(n_578), .Y(n_710) );
OR2x6_ASAP7_75t_L g475 ( .A(n_476), .B(n_482), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_484), .B(n_696), .Y(n_695) );
INVx1_ASAP7_75t_L g699 ( .A(n_484), .Y(n_699) );
AND2x2_ASAP7_75t_L g484 ( .A(n_485), .B(n_494), .Y(n_484) );
AND2x2_ASAP7_75t_L g529 ( .A(n_485), .B(n_530), .Y(n_529) );
AND2x4_ASAP7_75t_L g538 ( .A(n_485), .B(n_536), .Y(n_538) );
INVx5_ASAP7_75t_L g546 ( .A(n_485), .Y(n_546) );
AND2x2_ASAP7_75t_L g569 ( .A(n_485), .B(n_505), .Y(n_569) );
HB1xp67_ASAP7_75t_L g606 ( .A(n_485), .Y(n_606) );
OR2x6_ASAP7_75t_L g485 ( .A(n_486), .B(n_492), .Y(n_485) );
INVx1_ASAP7_75t_L g647 ( .A(n_494), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_494), .B(n_663), .Y(n_662) );
AND2x2_ASAP7_75t_L g680 ( .A(n_494), .B(n_546), .Y(n_680) );
A2O1A1Ixp33_ASAP7_75t_L g709 ( .A1(n_494), .A2(n_603), .B(n_710), .C(n_711), .Y(n_709) );
AND2x2_ASAP7_75t_L g494 ( .A(n_495), .B(n_505), .Y(n_494) );
BUFx2_ASAP7_75t_L g530 ( .A(n_495), .Y(n_530) );
INVx2_ASAP7_75t_L g534 ( .A(n_495), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_497), .B(n_502), .Y(n_496) );
INVx2_ASAP7_75t_L g536 ( .A(n_505), .Y(n_536) );
AND2x2_ASAP7_75t_L g543 ( .A(n_505), .B(n_534), .Y(n_543) );
AND2x2_ASAP7_75t_L g634 ( .A(n_505), .B(n_546), .Y(n_634) );
AOI211x1_ASAP7_75t_SL g514 ( .A1(n_515), .A2(n_527), .B(n_540), .C(n_565), .Y(n_514) );
INVx1_ASAP7_75t_L g631 ( .A(n_515), .Y(n_631) );
AND2x2_ASAP7_75t_L g515 ( .A(n_516), .B(n_526), .Y(n_515) );
INVx5_ASAP7_75t_SL g551 ( .A(n_517), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_517), .B(n_621), .Y(n_620) );
AOI311xp33_ASAP7_75t_L g639 ( .A1(n_517), .A2(n_640), .A3(n_642), .B(n_643), .C(n_649), .Y(n_639) );
A2O1A1Ixp33_ASAP7_75t_L g674 ( .A1(n_517), .A2(n_587), .B(n_675), .C(n_678), .Y(n_674) );
INVxp67_ASAP7_75t_L g594 ( .A(n_526), .Y(n_594) );
NAND4xp25_ASAP7_75t_SL g527 ( .A(n_528), .B(n_531), .C(n_537), .D(n_539), .Y(n_527) );
NOR2xp33_ASAP7_75t_L g592 ( .A(n_528), .B(n_593), .Y(n_592) );
INVx2_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
AND2x2_ASAP7_75t_L g585 ( .A(n_529), .B(n_586), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_532), .B(n_535), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_532), .B(n_538), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_532), .B(n_545), .Y(n_665) );
BUFx2_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_533), .B(n_546), .Y(n_683) );
HB1xp67_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
INVx2_ASAP7_75t_L g558 ( .A(n_534), .Y(n_558) );
INVxp67_ASAP7_75t_L g593 ( .A(n_535), .Y(n_593) );
AND2x4_ASAP7_75t_L g545 ( .A(n_536), .B(n_546), .Y(n_545) );
AND2x2_ASAP7_75t_L g619 ( .A(n_536), .B(n_558), .Y(n_619) );
INVx1_ASAP7_75t_L g646 ( .A(n_536), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_536), .B(n_633), .Y(n_693) );
NOR2xp33_ASAP7_75t_L g627 ( .A(n_537), .B(n_607), .Y(n_627) );
INVx1_ASAP7_75t_SL g537 ( .A(n_538), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_538), .B(n_560), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_538), .B(n_607), .Y(n_706) );
INVx1_ASAP7_75t_L g717 ( .A(n_539), .Y(n_717) );
A2O1A1Ixp33_ASAP7_75t_L g540 ( .A1(n_541), .A2(n_544), .B(n_547), .C(n_555), .Y(n_540) );
INVx1_ASAP7_75t_SL g541 ( .A(n_542), .Y(n_541) );
AND2x2_ASAP7_75t_L g559 ( .A(n_543), .B(n_560), .Y(n_559) );
AND2x2_ASAP7_75t_L g597 ( .A(n_543), .B(n_598), .Y(n_597) );
INVx1_ASAP7_75t_L g579 ( .A(n_544), .Y(n_579) );
AND2x2_ASAP7_75t_L g556 ( .A(n_545), .B(n_557), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_545), .B(n_607), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_545), .B(n_626), .Y(n_650) );
OR2x2_ASAP7_75t_L g566 ( .A(n_546), .B(n_567), .Y(n_566) );
INVx2_ASAP7_75t_L g598 ( .A(n_546), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_546), .B(n_558), .Y(n_613) );
AND2x2_ASAP7_75t_L g670 ( .A(n_546), .B(n_626), .Y(n_670) );
HB1xp67_ASAP7_75t_L g677 ( .A(n_546), .Y(n_677) );
INVx1_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
AOI221xp5_ASAP7_75t_L g681 ( .A1(n_548), .A2(n_560), .B1(n_682), .B2(n_684), .C(n_687), .Y(n_681) );
AND2x2_ASAP7_75t_L g548 ( .A(n_549), .B(n_552), .Y(n_548) );
INVx1_ASAP7_75t_SL g549 ( .A(n_550), .Y(n_549) );
OR2x2_ASAP7_75t_L g571 ( .A(n_551), .B(n_554), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_551), .B(n_621), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_551), .B(n_578), .Y(n_686) );
INVx1_ASAP7_75t_SL g552 ( .A(n_553), .Y(n_552) );
OR2x2_ASAP7_75t_L g671 ( .A(n_553), .B(n_672), .Y(n_671) );
OR2x2_ASAP7_75t_L g685 ( .A(n_553), .B(n_686), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_554), .B(n_578), .Y(n_577) );
AND2x2_ASAP7_75t_L g582 ( .A(n_554), .B(n_575), .Y(n_582) );
AND2x2_ASAP7_75t_L g652 ( .A(n_554), .B(n_653), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_554), .B(n_601), .Y(n_698) );
NOR2xp33_ASAP7_75t_L g701 ( .A(n_554), .B(n_702), .Y(n_701) );
OAI21xp5_ASAP7_75t_SL g555 ( .A1(n_556), .A2(n_559), .B(n_561), .Y(n_555) );
INVx2_ASAP7_75t_L g588 ( .A(n_556), .Y(n_588) );
HB1xp67_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
INVx1_ASAP7_75t_L g608 ( .A(n_558), .Y(n_608) );
OR2x2_ASAP7_75t_L g612 ( .A(n_560), .B(n_613), .Y(n_612) );
OR2x2_ASAP7_75t_L g715 ( .A(n_560), .B(n_683), .Y(n_715) );
INVx1_ASAP7_75t_SL g561 ( .A(n_562), .Y(n_561) );
OR2x2_ASAP7_75t_L g562 ( .A(n_563), .B(n_564), .Y(n_562) );
AOI21xp33_ASAP7_75t_SL g565 ( .A1(n_566), .A2(n_568), .B(n_570), .Y(n_565) );
INVx1_ASAP7_75t_L g719 ( .A(n_566), .Y(n_719) );
INVx2_ASAP7_75t_SL g633 ( .A(n_567), .Y(n_633) );
INVx1_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
A2O1A1Ixp33_ASAP7_75t_L g714 ( .A1(n_570), .A2(n_651), .B(n_715), .C(n_716), .Y(n_714) );
OAI322xp33_ASAP7_75t_SL g583 ( .A1(n_571), .A2(n_584), .A3(n_587), .B1(n_588), .B2(n_589), .C1(n_591), .C2(n_594), .Y(n_583) );
INVx2_ASAP7_75t_L g603 ( .A(n_571), .Y(n_603) );
AOI221xp5_ASAP7_75t_L g572 ( .A1(n_573), .A2(n_579), .B1(n_580), .B2(n_582), .C(n_583), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
OAI22xp33_ASAP7_75t_SL g649 ( .A1(n_574), .A2(n_650), .B1(n_651), .B2(n_654), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_575), .B(n_576), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_575), .B(n_578), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_575), .B(n_713), .Y(n_712) );
INVx2_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
OR2x2_ASAP7_75t_L g648 ( .A(n_577), .B(n_610), .Y(n_648) );
INVx1_ASAP7_75t_L g638 ( .A(n_578), .Y(n_638) );
INVx1_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
AOI21xp5_ASAP7_75t_L g691 ( .A1(n_582), .A2(n_692), .B(n_694), .Y(n_691) );
AOI21xp33_ASAP7_75t_L g616 ( .A1(n_584), .A2(n_617), .B(n_620), .Y(n_616) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
NOR2xp67_ASAP7_75t_SL g645 ( .A(n_586), .B(n_646), .Y(n_645) );
NOR2xp33_ASAP7_75t_L g678 ( .A(n_586), .B(n_679), .Y(n_678) );
INVx1_ASAP7_75t_SL g702 ( .A(n_587), .Y(n_702) );
INVx1_ASAP7_75t_SL g589 ( .A(n_590), .Y(n_589) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
NAND4xp25_ASAP7_75t_L g595 ( .A(n_596), .B(n_623), .C(n_639), .D(n_655), .Y(n_595) );
AOI211xp5_ASAP7_75t_L g596 ( .A1(n_597), .A2(n_599), .B(n_604), .C(n_616), .Y(n_596) );
INVx1_ASAP7_75t_L g688 ( .A(n_597), .Y(n_688) );
AND2x2_ASAP7_75t_L g636 ( .A(n_598), .B(n_619), .Y(n_636) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_601), .B(n_603), .Y(n_600) );
INVx1_ASAP7_75t_SL g601 ( .A(n_602), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_603), .B(n_638), .Y(n_637) );
OAI22xp33_ASAP7_75t_L g604 ( .A1(n_605), .A2(n_609), .B1(n_612), .B2(n_614), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_606), .B(n_607), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_606), .B(n_626), .Y(n_625) );
INVx1_ASAP7_75t_L g654 ( .A(n_607), .Y(n_654) );
O2A1O1Ixp33_ASAP7_75t_L g668 ( .A1(n_607), .A2(n_646), .B(n_669), .C(n_671), .Y(n_668) );
OR2x2_ASAP7_75t_L g609 ( .A(n_610), .B(n_611), .Y(n_609) );
INVx1_ASAP7_75t_L g653 ( .A(n_610), .Y(n_653) );
INVx1_ASAP7_75t_L g713 ( .A(n_611), .Y(n_713) );
NAND2xp33_ASAP7_75t_SL g703 ( .A(n_612), .B(n_704), .Y(n_703) );
INVx1_ASAP7_75t_SL g614 ( .A(n_615), .Y(n_614) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
INVx2_ASAP7_75t_L g642 ( .A(n_621), .Y(n_642) );
O2A1O1Ixp33_ASAP7_75t_L g623 ( .A1(n_624), .A2(n_627), .B(n_628), .C(n_630), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
OAI22xp5_ASAP7_75t_L g630 ( .A1(n_631), .A2(n_632), .B1(n_635), .B2(n_637), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_633), .B(n_634), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_633), .B(n_677), .Y(n_676) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_638), .B(n_659), .Y(n_721) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
AOI21xp33_ASAP7_75t_SL g643 ( .A1(n_644), .A2(n_647), .B(n_648), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
INVx1_ASAP7_75t_SL g651 ( .A(n_652), .Y(n_651) );
AOI221xp5_ASAP7_75t_L g655 ( .A1(n_656), .A2(n_661), .B1(n_664), .B2(n_666), .C(n_668), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_658), .B(n_659), .Y(n_657) );
INVx1_ASAP7_75t_SL g659 ( .A(n_660), .Y(n_659) );
INVx1_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
INVxp67_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
OAI22xp5_ASAP7_75t_L g687 ( .A1(n_671), .A2(n_688), .B1(n_689), .B2(n_690), .Y(n_687) );
NAND3xp33_ASAP7_75t_SL g673 ( .A(n_674), .B(n_681), .C(n_691), .Y(n_673) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
INVx1_ASAP7_75t_SL g679 ( .A(n_680), .Y(n_679) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
CKINVDCx16_ASAP7_75t_R g684 ( .A(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
INVxp67_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
OAI211xp5_ASAP7_75t_L g697 ( .A1(n_698), .A2(n_699), .B(n_700), .C(n_709), .Y(n_697) );
INVx1_ASAP7_75t_L g718 ( .A(n_698), .Y(n_718) );
AOI22xp33_ASAP7_75t_L g700 ( .A1(n_701), .A2(n_703), .B1(n_705), .B2(n_707), .Y(n_700) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVx1_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
AOI22xp5_ASAP7_75t_L g716 ( .A1(n_717), .A2(n_718), .B1(n_719), .B2(n_720), .Y(n_716) );
INVx1_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
CKINVDCx16_ASAP7_75t_R g722 ( .A(n_723), .Y(n_722) );
INVx2_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
BUFx2_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
INVx2_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
INVx1_ASAP7_75t_L g745 ( .A(n_735), .Y(n_745) );
INVxp67_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
NAND2xp5_ASAP7_75t_L g737 ( .A(n_738), .B(n_742), .Y(n_737) );
BUFx2_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
INVx2_ASAP7_75t_L g749 ( .A(n_743), .Y(n_749) );
INVx1_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
NOR2xp33_ASAP7_75t_L g746 ( .A(n_747), .B(n_748), .Y(n_746) );
INVx1_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
endmodule