module fake_jpeg_21685_n_208 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_208);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_208;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

BUFx3_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_3),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx16_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx14_ASAP7_75t_R g23 ( 
.A(n_12),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_19),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_19),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

INVx13_ASAP7_75t_L g29 ( 
.A(n_25),
.Y(n_29)
);

INVx5_ASAP7_75t_SL g46 ( 
.A(n_29),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_19),
.Y(n_30)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

AND2x2_ASAP7_75t_SL g31 ( 
.A(n_25),
.B(n_0),
.Y(n_31)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_31),
.B(n_24),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_19),
.Y(n_32)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_13),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_33),
.B(n_35),
.Y(n_38)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_34),
.A2(n_24),
.B1(n_18),
.B2(n_17),
.Y(n_41)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_37),
.B(n_30),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_41),
.A2(n_44),
.B1(n_49),
.B2(n_26),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_31),
.A2(n_18),
.B1(n_22),
.B2(n_15),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_43),
.A2(n_45),
.B1(n_48),
.B2(n_35),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_34),
.A2(n_20),
.B1(n_15),
.B2(n_22),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_31),
.A2(n_23),
.B1(n_17),
.B2(n_16),
.Y(n_45)
);

AO22x1_ASAP7_75t_SL g48 ( 
.A1(n_31),
.A2(n_23),
.B1(n_14),
.B2(n_21),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_34),
.A2(n_20),
.B1(n_16),
.B2(n_14),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_50),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_51),
.A2(n_57),
.B1(n_59),
.B2(n_43),
.Y(n_69)
);

AND2x4_ASAP7_75t_L g52 ( 
.A(n_37),
.B(n_31),
.Y(n_52)
);

OR2x2_ASAP7_75t_L g83 ( 
.A(n_52),
.B(n_47),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_37),
.B(n_33),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_53),
.B(n_65),
.Y(n_71)
);

HAxp5_ASAP7_75t_SL g54 ( 
.A(n_48),
.B(n_21),
.CON(n_54),
.SN(n_54)
);

OR2x2_ASAP7_75t_SL g74 ( 
.A(n_54),
.B(n_63),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_38),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_55),
.B(n_58),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_56),
.Y(n_67)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_38),
.A2(n_26),
.B1(n_27),
.B2(n_28),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_38),
.B(n_29),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_60),
.B(n_48),
.Y(n_73)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_61),
.Y(n_70)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_62),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_37),
.A2(n_14),
.B1(n_29),
.B2(n_27),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g64 ( 
.A(n_44),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_64),
.B(n_46),
.Y(n_78)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_66),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_69),
.A2(n_63),
.B1(n_52),
.B2(n_41),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_60),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_72),
.B(n_73),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_53),
.B(n_52),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_75),
.B(n_79),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_55),
.B(n_45),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_76),
.B(n_84),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g85 ( 
.A1(n_78),
.A2(n_64),
.B(n_63),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_57),
.B(n_48),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_65),
.B(n_48),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_80),
.B(n_83),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_59),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_85),
.A2(n_78),
.B1(n_49),
.B2(n_46),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g86 ( 
.A(n_75),
.B(n_52),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_86),
.B(n_89),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_79),
.A2(n_65),
.B1(n_52),
.B2(n_51),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_88),
.A2(n_83),
.B1(n_69),
.B2(n_101),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g89 ( 
.A(n_71),
.B(n_52),
.Y(n_89)
);

BUFx2_ASAP7_75t_L g90 ( 
.A(n_68),
.Y(n_90)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_90),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_81),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_92),
.B(n_96),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_94),
.A2(n_84),
.B1(n_74),
.B2(n_71),
.Y(n_106)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_81),
.Y(n_95)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_95),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_70),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_77),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_97),
.Y(n_102)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_77),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_99),
.B(n_100),
.Y(n_107)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_68),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_83),
.B(n_65),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_101),
.A2(n_74),
.B1(n_76),
.B2(n_72),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_87),
.A2(n_73),
.B(n_80),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_103),
.A2(n_113),
.B1(n_116),
.B2(n_117),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_98),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_104),
.B(n_108),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_105),
.A2(n_46),
.B1(n_36),
.B2(n_100),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_106),
.A2(n_110),
.B1(n_112),
.B2(n_93),
.Y(n_120)
);

OA22x2_ASAP7_75t_L g111 ( 
.A1(n_97),
.A2(n_62),
.B1(n_36),
.B2(n_47),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_111),
.A2(n_114),
.B1(n_67),
.B2(n_36),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_94),
.A2(n_58),
.B1(n_50),
.B2(n_47),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_99),
.B(n_82),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_88),
.A2(n_62),
.B1(n_67),
.B2(n_61),
.Y(n_114)
);

NAND2xp33_ASAP7_75t_SL g116 ( 
.A(n_85),
.B(n_30),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_120),
.B(n_114),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_118),
.B(n_86),
.C(n_89),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_121),
.B(n_131),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_102),
.B(n_91),
.Y(n_122)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_122),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_118),
.B(n_91),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_123),
.B(n_127),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_104),
.A2(n_93),
.B1(n_92),
.B2(n_95),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_124),
.A2(n_126),
.B1(n_132),
.B2(n_109),
.Y(n_146)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_107),
.Y(n_125)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_125),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_103),
.B(n_70),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_115),
.B(n_82),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_128),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_129),
.A2(n_113),
.B(n_116),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_111),
.B(n_90),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_130),
.B(n_134),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_106),
.B(n_66),
.Y(n_131)
);

HB1xp67_ASAP7_75t_L g133 ( 
.A(n_110),
.Y(n_133)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_133),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_117),
.B(n_113),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_111),
.B(n_66),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_135),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_105),
.B(n_112),
.Y(n_136)
);

MAJx2_ASAP7_75t_L g148 ( 
.A(n_136),
.B(n_111),
.C(n_28),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_137),
.A2(n_140),
.B1(n_121),
.B2(n_109),
.Y(n_154)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_132),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_139),
.B(n_150),
.Y(n_153)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_129),
.Y(n_145)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_145),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_146),
.A2(n_149),
.B1(n_39),
.B2(n_67),
.Y(n_160)
);

MAJx2_ASAP7_75t_L g163 ( 
.A(n_148),
.B(n_32),
.C(n_46),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_119),
.A2(n_136),
.B1(n_131),
.B2(n_127),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_123),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_154),
.B(n_155),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_144),
.B(n_68),
.C(n_28),
.Y(n_155)
);

BUFx12_ASAP7_75t_L g156 ( 
.A(n_151),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_156),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_144),
.B(n_30),
.C(n_32),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_157),
.B(n_160),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_138),
.B(n_10),
.Y(n_159)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_159),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_143),
.B(n_8),
.Y(n_161)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_161),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_152),
.B(n_32),
.C(n_40),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_162),
.B(n_163),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_152),
.B(n_40),
.C(n_56),
.Y(n_164)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_164),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_147),
.B(n_7),
.Y(n_165)
);

INVxp67_ASAP7_75t_SL g170 ( 
.A(n_165),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_153),
.A2(n_139),
.B1(n_140),
.B2(n_145),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_166),
.B(n_167),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_158),
.A2(n_141),
.B1(n_137),
.B2(n_142),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_164),
.A2(n_142),
.B1(n_148),
.B2(n_56),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_169),
.B(n_162),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_167),
.B(n_157),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_177),
.B(n_181),
.Y(n_193)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_179),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_174),
.A2(n_155),
.B1(n_163),
.B2(n_156),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_180),
.A2(n_169),
.B1(n_172),
.B2(n_166),
.Y(n_186)
);

BUFx2_ASAP7_75t_L g181 ( 
.A(n_170),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_171),
.B(n_156),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_182),
.A2(n_183),
.B(n_184),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_168),
.A2(n_7),
.B(n_12),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_171),
.A2(n_6),
.B(n_12),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_176),
.B(n_40),
.C(n_61),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_185),
.B(n_176),
.C(n_40),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_186),
.B(n_188),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_178),
.A2(n_182),
.B1(n_173),
.B2(n_175),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_189),
.B(n_0),
.C(n_1),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_185),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_190),
.B(n_0),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_181),
.B(n_5),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_191),
.B(n_4),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_195),
.B(n_196),
.Y(n_202)
);

AOI322xp5_ASAP7_75t_L g200 ( 
.A1(n_197),
.A2(n_198),
.A3(n_190),
.B1(n_11),
.B2(n_8),
.C1(n_10),
.C2(n_1),
.Y(n_200)
);

OAI21x1_ASAP7_75t_L g198 ( 
.A1(n_187),
.A2(n_3),
.B(n_6),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_192),
.B(n_3),
.C(n_6),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_199),
.A2(n_11),
.B(n_1),
.Y(n_203)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_200),
.Y(n_205)
);

AOI322xp5_ASAP7_75t_L g201 ( 
.A1(n_194),
.A2(n_193),
.A3(n_189),
.B1(n_8),
.B2(n_10),
.C1(n_11),
.C2(n_2),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_201),
.B(n_203),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_205),
.A2(n_202),
.B(n_2),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_206),
.B(n_204),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_207),
.B(n_2),
.Y(n_208)
);


endmodule