module fake_jpeg_603_n_132 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_132);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_132;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_30),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_22),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

CKINVDCx5p33_ASAP7_75t_R g42 ( 
.A(n_33),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_3),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_11),
.Y(n_47)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_49),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_50),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

CKINVDCx6p67_ASAP7_75t_R g64 ( 
.A(n_51),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_52),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_42),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_53),
.B(n_42),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_54),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_55),
.B(n_57),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_50),
.B(n_40),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_52),
.B(n_35),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_58),
.B(n_60),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_52),
.B(n_47),
.Y(n_60)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_56),
.Y(n_65)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_65),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_61),
.A2(n_54),
.B1(n_46),
.B2(n_38),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_66),
.B(n_68),
.Y(n_83)
);

OA21x2_ASAP7_75t_L g67 ( 
.A1(n_57),
.A2(n_43),
.B(n_44),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_67),
.Y(n_77)
);

INVx1_ASAP7_75t_SL g68 ( 
.A(n_62),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_64),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_69),
.B(n_71),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_64),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_61),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_72),
.B(n_75),
.Y(n_80)
);

INVx13_ASAP7_75t_L g74 ( 
.A(n_64),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_74),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_59),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_63),
.B(n_45),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_76),
.B(n_63),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_72),
.B(n_34),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_82),
.B(n_84),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_73),
.B(n_39),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_70),
.B(n_37),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_L g90 ( 
.A(n_85),
.B(n_87),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_86),
.B(n_89),
.Y(n_103)
);

A2O1A1Ixp33_ASAP7_75t_L g87 ( 
.A1(n_69),
.A2(n_37),
.B(n_40),
.C(n_2),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_71),
.B(n_59),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_SL g100 ( 
.A(n_88),
.B(n_5),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_67),
.B(n_46),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_77),
.A2(n_67),
.B1(n_75),
.B2(n_68),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_91),
.A2(n_94),
.B1(n_96),
.B2(n_99),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_81),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_92),
.B(n_93),
.Y(n_114)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_82),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_83),
.A2(n_74),
.B1(n_62),
.B2(n_3),
.Y(n_94)
);

OA22x2_ASAP7_75t_L g95 ( 
.A1(n_83),
.A2(n_62),
.B1(n_14),
.B2(n_15),
.Y(n_95)
);

AO21x1_ASAP7_75t_L g109 ( 
.A1(n_95),
.A2(n_16),
.B(n_28),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_88),
.A2(n_0),
.B1(n_1),
.B2(n_4),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_87),
.B(n_80),
.C(n_78),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_97),
.B(n_102),
.C(n_31),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_79),
.Y(n_98)
);

CKINVDCx14_ASAP7_75t_R g105 ( 
.A(n_98),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_77),
.A2(n_0),
.B1(n_4),
.B2(n_5),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_100),
.B(n_6),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_85),
.B(n_20),
.C(n_29),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_101),
.B(n_6),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_104),
.B(n_106),
.Y(n_117)
);

NAND3xp33_ASAP7_75t_L g106 ( 
.A(n_103),
.B(n_90),
.C(n_98),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_92),
.Y(n_107)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_107),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_108),
.B(n_115),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_109),
.A2(n_111),
.B1(n_113),
.B2(n_7),
.Y(n_118)
);

NAND3xp33_ASAP7_75t_L g110 ( 
.A(n_103),
.B(n_13),
.C(n_27),
.Y(n_110)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_110),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_95),
.B(n_7),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_97),
.A2(n_12),
.B(n_26),
.Y(n_113)
);

O2A1O1Ixp33_ASAP7_75t_L g116 ( 
.A1(n_112),
.A2(n_25),
.B(n_24),
.C(n_23),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_116),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_118),
.B(n_8),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_117),
.A2(n_106),
.B1(n_114),
.B2(n_105),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_122),
.A2(n_120),
.B1(n_116),
.B2(n_119),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_121),
.B(n_110),
.C(n_109),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_124),
.B(n_125),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_126),
.A2(n_127),
.B(n_123),
.Y(n_128)
);

FAx1_ASAP7_75t_SL g129 ( 
.A(n_128),
.B(n_124),
.CI(n_121),
.CON(n_129),
.SN(n_129)
);

BUFx24_ASAP7_75t_SL g130 ( 
.A(n_129),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_130),
.B(n_129),
.C(n_10),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_131),
.A2(n_8),
.B(n_10),
.Y(n_132)
);


endmodule