module fake_jpeg_31157_n_137 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_137);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_137;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_57;
wire n_21;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_11),
.Y(n_12)
);

INVx4_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

INVxp67_ASAP7_75t_L g14 ( 
.A(n_11),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_8),
.Y(n_15)
);

INVx6_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx14_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g28 ( 
.A(n_19),
.B(n_7),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_28),
.B(n_30),
.Y(n_37)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_25),
.Y(n_29)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_14),
.B(n_0),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_19),
.B(n_1),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_32),
.B(n_34),
.Y(n_44)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_27),
.B(n_0),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

INVx6_ASAP7_75t_SL g36 ( 
.A(n_14),
.Y(n_36)
);

INVx1_ASAP7_75t_SL g43 ( 
.A(n_36),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

BUFx2_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

NOR2x1_ASAP7_75t_L g45 ( 
.A(n_28),
.B(n_24),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_45),
.B(n_32),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_34),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_46),
.B(n_36),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_46),
.B(n_39),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_48),
.B(n_49),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_39),
.B(n_42),
.C(n_30),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_44),
.A2(n_31),
.B1(n_16),
.B2(n_13),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_50),
.B(n_52),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_51),
.B(n_57),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_L g52 ( 
.A(n_37),
.B(n_45),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_45),
.B(n_21),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_53),
.B(n_54),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_38),
.A2(n_13),
.B1(n_22),
.B2(n_21),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_55),
.B(n_58),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_43),
.B(n_18),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_38),
.A2(n_29),
.B1(n_25),
.B2(n_17),
.Y(n_58)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_60),
.Y(n_75)
);

HAxp5_ASAP7_75t_SL g82 ( 
.A(n_61),
.B(n_53),
.CON(n_82),
.SN(n_82)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_62),
.Y(n_77)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_63),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_41),
.B(n_20),
.Y(n_64)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_64),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_38),
.A2(n_29),
.B1(n_25),
.B2(n_22),
.Y(n_65)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_65),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_40),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_66),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g73 ( 
.A1(n_48),
.A2(n_56),
.B(n_49),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_73),
.B(n_54),
.Y(n_86)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_60),
.Y(n_74)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_74),
.Y(n_84)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_63),
.Y(n_80)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_80),
.Y(n_87)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_62),
.Y(n_81)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_81),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_82),
.B(n_35),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_78),
.B(n_52),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_83),
.B(n_85),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_70),
.B(n_23),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_86),
.B(n_91),
.C(n_93),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_88),
.A2(n_95),
.B(n_86),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_72),
.B(n_26),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_89),
.B(n_94),
.Y(n_105)
);

MAJx2_ASAP7_75t_L g91 ( 
.A(n_67),
.B(n_26),
.C(n_23),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_74),
.Y(n_92)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_92),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_73),
.B(n_35),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_69),
.B(n_12),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_82),
.B(n_40),
.C(n_15),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_95),
.Y(n_97)
);

AO22x1_ASAP7_75t_SL g96 ( 
.A1(n_88),
.A2(n_68),
.B1(n_76),
.B2(n_71),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_96),
.B(n_100),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_93),
.A2(n_68),
.B1(n_79),
.B2(n_80),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_98),
.A2(n_106),
.B1(n_75),
.B2(n_77),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_99),
.B(n_103),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_84),
.Y(n_100)
);

OR2x2_ASAP7_75t_L g103 ( 
.A(n_91),
.B(n_71),
.Y(n_103)
);

A2O1A1Ixp33_ASAP7_75t_SL g106 ( 
.A1(n_87),
.A2(n_59),
.B(n_81),
.C(n_75),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_101),
.B(n_90),
.C(n_77),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_108),
.B(n_110),
.Y(n_117)
);

INVx1_ASAP7_75t_SL g118 ( 
.A(n_109),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_97),
.B(n_59),
.C(n_25),
.Y(n_110)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_104),
.Y(n_112)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_112),
.Y(n_115)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_96),
.Y(n_113)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_113),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_105),
.B(n_2),
.Y(n_114)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_114),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_111),
.A2(n_103),
.B(n_97),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_116),
.A2(n_102),
.B(n_108),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_117),
.A2(n_107),
.B(n_110),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_121),
.A2(n_124),
.B(n_125),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_122),
.B(n_123),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_120),
.B(n_3),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_115),
.B(n_8),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_119),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_121),
.B(n_118),
.C(n_106),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_126),
.B(n_106),
.C(n_10),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_121),
.B(n_118),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_128),
.B(n_106),
.Y(n_131)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_129),
.Y(n_130)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_130),
.Y(n_133)
);

OR2x2_ASAP7_75t_L g134 ( 
.A(n_131),
.B(n_132),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_133),
.B(n_127),
.Y(n_135)
);

MAJx2_ASAP7_75t_L g136 ( 
.A(n_135),
.B(n_134),
.C(n_128),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_136),
.B(n_10),
.Y(n_137)
);


endmodule