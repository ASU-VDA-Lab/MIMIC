module fake_jpeg_30673_n_47 (n_3, n_2, n_1, n_0, n_4, n_5, n_47);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_47;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_44;
wire n_26;
wire n_38;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

BUFx2_ASAP7_75t_L g6 ( 
.A(n_3),
.Y(n_6)
);

INVx1_ASAP7_75t_L g7 ( 
.A(n_5),
.Y(n_7)
);

INVx8_ASAP7_75t_L g8 ( 
.A(n_5),
.Y(n_8)
);

BUFx3_ASAP7_75t_L g9 ( 
.A(n_0),
.Y(n_9)
);

INVx3_ASAP7_75t_L g10 ( 
.A(n_5),
.Y(n_10)
);

INVx4_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

INVx8_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_12),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_14),
.B(n_16),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_L g15 ( 
.A1(n_12),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_15)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_15),
.A2(n_17),
.B1(n_7),
.B2(n_21),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_11),
.B(n_0),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_L g17 ( 
.A1(n_10),
.A2(n_3),
.B1(n_4),
.B2(n_0),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_18),
.B(n_20),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_11),
.B(n_0),
.C(n_1),
.Y(n_19)
);

AOI21xp5_ASAP7_75t_L g23 ( 
.A1(n_19),
.A2(n_1),
.B(n_9),
.Y(n_23)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_6),
.B(n_1),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_SL g26 ( 
.A(n_21),
.B(n_6),
.Y(n_26)
);

OAI21xp5_ASAP7_75t_L g30 ( 
.A1(n_23),
.A2(n_9),
.B(n_14),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_24),
.A2(n_15),
.B1(n_19),
.B2(n_17),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_16),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_25),
.Y(n_33)
);

XOR2xp5_ASAP7_75t_L g31 ( 
.A(n_26),
.B(n_27),
.Y(n_31)
);

OAI21xp5_ASAP7_75t_SL g27 ( 
.A1(n_19),
.A2(n_10),
.B(n_7),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_29),
.A2(n_23),
.B1(n_18),
.B2(n_20),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_30),
.B(n_32),
.Y(n_36)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_28),
.Y(n_32)
);

AOI21xp33_ASAP7_75t_SL g34 ( 
.A1(n_31),
.A2(n_26),
.B(n_27),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_34),
.B(n_31),
.C(n_36),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_30),
.A2(n_24),
.B1(n_22),
.B2(n_14),
.Y(n_35)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_35),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_37),
.B(n_18),
.C(n_20),
.Y(n_41)
);

XOR2xp5_ASAP7_75t_L g42 ( 
.A(n_39),
.B(n_40),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_37),
.B(n_32),
.C(n_33),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_41),
.B(n_35),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_43),
.A2(n_44),
.B1(n_13),
.B2(n_8),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_38),
.B(n_8),
.Y(n_44)
);

AOI21xp5_ASAP7_75t_L g46 ( 
.A1(n_45),
.A2(n_42),
.B(n_1),
.Y(n_46)
);

AO21x1_ASAP7_75t_L g47 ( 
.A1(n_46),
.A2(n_42),
.B(n_13),
.Y(n_47)
);


endmodule