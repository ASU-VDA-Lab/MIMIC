module real_aes_2443_n_100 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_100);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_100;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_659;
wire n_547;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_754;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_769;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_733;
wire n_602;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_768;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_288;
wire n_150;
wire n_147;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_749;
wire n_162;
wire n_358;
wire n_275;
wire n_214;
wire n_385;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_420;
wire n_336;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_762;
wire n_210;
wire n_212;
wire n_325;
wire n_575;
wire n_338;
wire n_479;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_SL g515 ( .A(n_0), .B(n_144), .Y(n_515) );
AOI21xp5_ASAP7_75t_L g462 ( .A1(n_1), .A2(n_152), .B(n_463), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g105 ( .A(n_2), .B(n_106), .Y(n_105) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_3), .B(n_144), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_4), .B(n_171), .Y(n_183) );
NAND2xp5_ASAP7_75t_SL g497 ( .A(n_5), .B(n_171), .Y(n_497) );
INVx1_ASAP7_75t_L g140 ( .A(n_6), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_7), .B(n_171), .Y(n_546) );
CKINVDCx16_ASAP7_75t_R g106 ( .A(n_8), .Y(n_106) );
OAI22xp5_ASAP7_75t_L g767 ( .A1(n_9), .A2(n_13), .B1(n_768), .B2(n_769), .Y(n_767) );
CKINVDCx20_ASAP7_75t_R g768 ( .A(n_9), .Y(n_768) );
NAND2xp33_ASAP7_75t_L g538 ( .A(n_10), .B(n_169), .Y(n_538) );
AND2x2_ASAP7_75t_L g174 ( .A(n_11), .B(n_175), .Y(n_174) );
AND2x2_ASAP7_75t_L g185 ( .A(n_12), .B(n_186), .Y(n_185) );
AOI222xp33_ASAP7_75t_SL g100 ( .A1(n_13), .A2(n_101), .B1(n_116), .B2(n_760), .C1(n_762), .C2(n_773), .Y(n_100) );
CKINVDCx20_ASAP7_75t_R g769 ( .A(n_13), .Y(n_769) );
INVx2_ASAP7_75t_L g131 ( .A(n_14), .Y(n_131) );
AOI221x1_ASAP7_75t_L g482 ( .A1(n_15), .A2(n_26), .B1(n_144), .B2(n_152), .C(n_483), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_16), .B(n_171), .Y(n_211) );
CKINVDCx16_ASAP7_75t_R g110 ( .A(n_17), .Y(n_110) );
NAND2xp5_ASAP7_75t_SL g534 ( .A(n_18), .B(n_144), .Y(n_534) );
AO21x2_ASAP7_75t_L g532 ( .A1(n_19), .A2(n_186), .B(n_533), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_20), .B(n_129), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_21), .B(n_171), .Y(n_471) );
AO21x1_ASAP7_75t_L g492 ( .A1(n_22), .A2(n_144), .B(n_493), .Y(n_492) );
NAND2xp5_ASAP7_75t_SL g227 ( .A(n_23), .B(n_144), .Y(n_227) );
INVx1_ASAP7_75t_L g114 ( .A(n_24), .Y(n_114) );
AOI22xp33_ASAP7_75t_L g134 ( .A1(n_25), .A2(n_88), .B1(n_135), .B2(n_144), .Y(n_134) );
NAND2x1_ASAP7_75t_L g513 ( .A(n_27), .B(n_171), .Y(n_513) );
NAND2x1_ASAP7_75t_L g545 ( .A(n_28), .B(n_169), .Y(n_545) );
OR2x2_ASAP7_75t_L g132 ( .A(n_29), .B(n_85), .Y(n_132) );
OA21x2_ASAP7_75t_L g164 ( .A1(n_29), .A2(n_85), .B(n_131), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_30), .B(n_169), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_31), .B(n_171), .Y(n_537) );
AO21x2_ASAP7_75t_L g206 ( .A1(n_32), .A2(n_175), .B(n_207), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_33), .B(n_169), .Y(n_496) );
AOI21xp5_ASAP7_75t_L g180 ( .A1(n_34), .A2(n_152), .B(n_181), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_35), .B(n_171), .Y(n_241) );
AOI21xp5_ASAP7_75t_L g502 ( .A1(n_36), .A2(n_152), .B(n_503), .Y(n_502) );
AND2x2_ASAP7_75t_L g142 ( .A(n_37), .B(n_143), .Y(n_142) );
AND2x2_ASAP7_75t_L g150 ( .A(n_37), .B(n_140), .Y(n_150) );
INVx1_ASAP7_75t_L g156 ( .A(n_37), .Y(n_156) );
OR2x6_ASAP7_75t_L g112 ( .A(n_38), .B(n_113), .Y(n_112) );
NAND2xp5_ASAP7_75t_SL g506 ( .A(n_39), .B(n_144), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_40), .B(n_144), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_41), .B(n_171), .Y(n_222) );
CKINVDCx20_ASAP7_75t_R g475 ( .A(n_42), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_43), .B(n_169), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_44), .B(n_144), .Y(n_193) );
AOI21xp5_ASAP7_75t_L g166 ( .A1(n_45), .A2(n_152), .B(n_167), .Y(n_166) );
AOI21xp5_ASAP7_75t_L g543 ( .A1(n_46), .A2(n_152), .B(n_544), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_47), .B(n_169), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_48), .B(n_169), .Y(n_514) );
NAND2xp5_ASAP7_75t_SL g208 ( .A(n_49), .B(n_144), .Y(n_208) );
INVx1_ASAP7_75t_L g138 ( .A(n_50), .Y(n_138) );
INVx1_ASAP7_75t_L g147 ( .A(n_50), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_51), .B(n_171), .Y(n_170) );
AND2x2_ASAP7_75t_L g217 ( .A(n_52), .B(n_129), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_53), .B(n_169), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_54), .B(n_171), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_55), .B(n_169), .Y(n_240) );
AOI21xp5_ASAP7_75t_L g511 ( .A1(n_56), .A2(n_152), .B(n_512), .Y(n_511) );
NAND2xp5_ASAP7_75t_SL g173 ( .A(n_57), .B(n_144), .Y(n_173) );
NAND2xp5_ASAP7_75t_SL g219 ( .A(n_58), .B(n_144), .Y(n_219) );
AOI21xp5_ASAP7_75t_L g238 ( .A1(n_59), .A2(n_152), .B(n_239), .Y(n_238) );
AND2x2_ASAP7_75t_L g233 ( .A(n_60), .B(n_130), .Y(n_233) );
AO21x1_ASAP7_75t_L g494 ( .A1(n_61), .A2(n_152), .B(n_495), .Y(n_494) );
NAND2xp5_ASAP7_75t_SL g461 ( .A(n_62), .B(n_144), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_63), .B(n_169), .Y(n_223) );
NAND2xp5_ASAP7_75t_SL g547 ( .A(n_64), .B(n_144), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_65), .B(n_169), .Y(n_212) );
AOI22xp5_ASAP7_75t_L g151 ( .A1(n_66), .A2(n_92), .B1(n_152), .B2(n_154), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_67), .B(n_171), .Y(n_230) );
AND2x2_ASAP7_75t_L g507 ( .A(n_68), .B(n_130), .Y(n_507) );
INVx1_ASAP7_75t_L g143 ( .A(n_69), .Y(n_143) );
INVx1_ASAP7_75t_L g149 ( .A(n_69), .Y(n_149) );
AND2x2_ASAP7_75t_L g548 ( .A(n_70), .B(n_175), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_71), .B(n_169), .Y(n_182) );
AOI21xp5_ASAP7_75t_L g220 ( .A1(n_72), .A2(n_152), .B(n_221), .Y(n_220) );
AOI22xp5_ASAP7_75t_SL g748 ( .A1(n_73), .A2(n_79), .B1(n_749), .B2(n_750), .Y(n_748) );
CKINVDCx20_ASAP7_75t_R g750 ( .A(n_73), .Y(n_750) );
AOI21xp5_ASAP7_75t_L g194 ( .A1(n_74), .A2(n_152), .B(n_195), .Y(n_194) );
AOI21xp5_ASAP7_75t_L g209 ( .A1(n_75), .A2(n_152), .B(n_210), .Y(n_209) );
CKINVDCx20_ASAP7_75t_R g756 ( .A(n_76), .Y(n_756) );
AND2x2_ASAP7_75t_L g243 ( .A(n_77), .B(n_130), .Y(n_243) );
NAND2xp5_ASAP7_75t_SL g128 ( .A(n_78), .B(n_129), .Y(n_128) );
INVx1_ASAP7_75t_L g749 ( .A(n_79), .Y(n_749) );
INVx1_ASAP7_75t_L g115 ( .A(n_80), .Y(n_115) );
AND2x2_ASAP7_75t_L g459 ( .A(n_81), .B(n_175), .Y(n_459) );
NAND2xp5_ASAP7_75t_SL g473 ( .A(n_82), .B(n_144), .Y(n_473) );
AND2x2_ASAP7_75t_L g198 ( .A(n_83), .B(n_186), .Y(n_198) );
AND2x2_ASAP7_75t_L g493 ( .A(n_84), .B(n_213), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_86), .B(n_169), .Y(n_472) );
AND2x2_ASAP7_75t_L g516 ( .A(n_87), .B(n_175), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_89), .B(n_171), .Y(n_505) );
AOI21xp5_ASAP7_75t_L g469 ( .A1(n_90), .A2(n_152), .B(n_470), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_91), .B(n_169), .Y(n_484) );
AOI21xp5_ASAP7_75t_L g228 ( .A1(n_93), .A2(n_152), .B(n_229), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_94), .B(n_171), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_95), .B(n_171), .Y(n_464) );
BUFx2_ASAP7_75t_L g232 ( .A(n_96), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g771 ( .A(n_97), .B(n_772), .Y(n_771) );
BUFx2_ASAP7_75t_L g107 ( .A(n_98), .Y(n_107) );
BUFx2_ASAP7_75t_SL g777 ( .A(n_98), .Y(n_777) );
AOI21xp5_ASAP7_75t_L g535 ( .A1(n_99), .A2(n_152), .B(n_536), .Y(n_535) );
AND2x2_ASAP7_75t_L g101 ( .A(n_102), .B(n_108), .Y(n_101) );
INVxp67_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
NAND2xp5_ASAP7_75t_SL g103 ( .A(n_104), .B(n_107), .Y(n_103) );
INVx2_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
OR2x2_ASAP7_75t_SL g761 ( .A(n_105), .B(n_107), .Y(n_761) );
AOI21xp5_ASAP7_75t_L g774 ( .A1(n_105), .A2(n_775), .B(n_778), .Y(n_774) );
INVx1_ASAP7_75t_SL g765 ( .A(n_108), .Y(n_765) );
INVx2_ASAP7_75t_L g772 ( .A(n_108), .Y(n_772) );
BUFx2_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
BUFx2_ASAP7_75t_L g779 ( .A(n_109), .Y(n_779) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_110), .B(n_111), .Y(n_109) );
AND2x6_ASAP7_75t_SL g451 ( .A(n_110), .B(n_112), .Y(n_451) );
OR2x6_ASAP7_75t_SL g746 ( .A(n_110), .B(n_111), .Y(n_746) );
OR2x2_ASAP7_75t_L g759 ( .A(n_110), .B(n_112), .Y(n_759) );
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_112), .Y(n_111) );
NAND2xp5_ASAP7_75t_L g113 ( .A(n_114), .B(n_115), .Y(n_113) );
INVxp33_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
AOI221xp5_ASAP7_75t_L g117 ( .A1(n_118), .A2(n_747), .B1(n_748), .B2(n_751), .C(n_755), .Y(n_117) );
OAI22xp5_ASAP7_75t_L g118 ( .A1(n_119), .A2(n_448), .B1(n_452), .B2(n_744), .Y(n_118) );
INVx3_ASAP7_75t_L g752 ( .A(n_119), .Y(n_752) );
OAI22xp5_ASAP7_75t_L g766 ( .A1(n_119), .A2(n_752), .B1(n_767), .B2(n_770), .Y(n_766) );
AND2x4_ASAP7_75t_L g119 ( .A(n_120), .B(n_373), .Y(n_119) );
NOR3xp33_ASAP7_75t_L g120 ( .A(n_121), .B(n_309), .C(n_356), .Y(n_120) );
NAND4xp25_ASAP7_75t_SL g121 ( .A(n_122), .B(n_244), .C(n_262), .D(n_288), .Y(n_121) );
OAI21xp33_ASAP7_75t_SL g122 ( .A1(n_123), .A2(n_202), .B(n_203), .Y(n_122) );
NAND2xp5_ASAP7_75t_SL g123 ( .A(n_124), .B(n_187), .Y(n_123) );
INVx1_ASAP7_75t_L g424 ( .A(n_124), .Y(n_424) );
OR2x2_ASAP7_75t_L g124 ( .A(n_125), .B(n_159), .Y(n_124) );
INVx2_ASAP7_75t_L g248 ( .A(n_125), .Y(n_248) );
AND2x2_ASAP7_75t_L g268 ( .A(n_125), .B(n_269), .Y(n_268) );
OR2x2_ASAP7_75t_L g370 ( .A(n_125), .B(n_189), .Y(n_370) );
AND2x2_ASAP7_75t_L g430 ( .A(n_125), .B(n_249), .Y(n_430) );
INVx2_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_126), .B(n_283), .Y(n_282) );
INVx2_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
OR2x2_ASAP7_75t_L g314 ( .A(n_127), .B(n_162), .Y(n_314) );
BUFx3_ASAP7_75t_L g324 ( .A(n_127), .Y(n_324) );
AND2x2_ASAP7_75t_L g387 ( .A(n_127), .B(n_388), .Y(n_387) );
AND2x4_ASAP7_75t_L g127 ( .A(n_128), .B(n_133), .Y(n_127) );
AND2x4_ASAP7_75t_L g201 ( .A(n_128), .B(n_133), .Y(n_201) );
AO21x2_ASAP7_75t_L g133 ( .A1(n_129), .A2(n_134), .B(n_151), .Y(n_133) );
CKINVDCx5p33_ASAP7_75t_R g178 ( .A(n_129), .Y(n_178) );
AOI21xp5_ASAP7_75t_L g192 ( .A1(n_129), .A2(n_193), .B(n_194), .Y(n_192) );
AOI21xp5_ASAP7_75t_L g460 ( .A1(n_129), .A2(n_461), .B(n_462), .Y(n_460) );
OA21x2_ASAP7_75t_L g481 ( .A1(n_129), .A2(n_482), .B(n_486), .Y(n_481) );
OA21x2_ASAP7_75t_L g552 ( .A1(n_129), .A2(n_482), .B(n_486), .Y(n_552) );
BUFx6f_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
AND2x2_ASAP7_75t_SL g130 ( .A(n_131), .B(n_132), .Y(n_130) );
AND2x4_ASAP7_75t_L g213 ( .A(n_131), .B(n_132), .Y(n_213) );
AND2x4_ASAP7_75t_L g135 ( .A(n_136), .B(n_141), .Y(n_135) );
AND2x2_ASAP7_75t_L g136 ( .A(n_137), .B(n_139), .Y(n_136) );
INVx2_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
AND2x2_ASAP7_75t_L g153 ( .A(n_138), .B(n_140), .Y(n_153) );
AND2x4_ASAP7_75t_L g171 ( .A(n_138), .B(n_148), .Y(n_171) );
HB1xp67_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
BUFx3_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
AND2x6_ASAP7_75t_L g152 ( .A(n_142), .B(n_153), .Y(n_152) );
INVx2_ASAP7_75t_L g158 ( .A(n_143), .Y(n_158) );
AND2x6_ASAP7_75t_L g169 ( .A(n_143), .B(n_146), .Y(n_169) );
AND2x4_ASAP7_75t_L g144 ( .A(n_145), .B(n_150), .Y(n_144) );
AND2x4_ASAP7_75t_L g145 ( .A(n_146), .B(n_148), .Y(n_145) );
INVx2_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx2_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx5_ASAP7_75t_L g172 ( .A(n_150), .Y(n_172) );
AND2x4_ASAP7_75t_L g154 ( .A(n_153), .B(n_155), .Y(n_154) );
NOR2x1p5_ASAP7_75t_L g155 ( .A(n_156), .B(n_157), .Y(n_155) );
INVx3_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx1_ASAP7_75t_SL g159 ( .A(n_160), .Y(n_159) );
INVx1_ASAP7_75t_L g433 ( .A(n_160), .Y(n_433) );
AND2x2_ASAP7_75t_L g160 ( .A(n_161), .B(n_176), .Y(n_160) );
AND2x2_ASAP7_75t_L g200 ( .A(n_161), .B(n_201), .Y(n_200) );
INVx1_ASAP7_75t_L g388 ( .A(n_161), .Y(n_388) );
INVx2_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
AND2x2_ASAP7_75t_L g202 ( .A(n_162), .B(n_191), .Y(n_202) );
AND2x2_ASAP7_75t_L g265 ( .A(n_162), .B(n_176), .Y(n_265) );
INVx2_ASAP7_75t_L g270 ( .A(n_162), .Y(n_270) );
AND2x2_ASAP7_75t_L g272 ( .A(n_162), .B(n_177), .Y(n_272) );
AO21x2_ASAP7_75t_L g162 ( .A1(n_163), .A2(n_165), .B(n_174), .Y(n_162) );
INVx4_ASAP7_75t_L g175 ( .A(n_163), .Y(n_175) );
INVx3_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
BUFx4f_ASAP7_75t_L g186 ( .A(n_164), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_166), .B(n_173), .Y(n_165) );
AOI21xp5_ASAP7_75t_L g167 ( .A1(n_168), .A2(n_170), .B(n_172), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_169), .B(n_232), .Y(n_231) );
AOI21xp5_ASAP7_75t_L g181 ( .A1(n_172), .A2(n_182), .B(n_183), .Y(n_181) );
AOI21xp5_ASAP7_75t_L g195 ( .A1(n_172), .A2(n_196), .B(n_197), .Y(n_195) );
AOI21xp5_ASAP7_75t_L g210 ( .A1(n_172), .A2(n_211), .B(n_212), .Y(n_210) );
AOI21xp5_ASAP7_75t_L g221 ( .A1(n_172), .A2(n_222), .B(n_223), .Y(n_221) );
AOI21xp5_ASAP7_75t_L g229 ( .A1(n_172), .A2(n_230), .B(n_231), .Y(n_229) );
AOI21xp5_ASAP7_75t_L g239 ( .A1(n_172), .A2(n_240), .B(n_241), .Y(n_239) );
AOI21xp5_ASAP7_75t_L g463 ( .A1(n_172), .A2(n_464), .B(n_465), .Y(n_463) );
AOI21xp5_ASAP7_75t_L g470 ( .A1(n_172), .A2(n_471), .B(n_472), .Y(n_470) );
AOI21xp5_ASAP7_75t_L g483 ( .A1(n_172), .A2(n_484), .B(n_485), .Y(n_483) );
AOI21xp5_ASAP7_75t_L g495 ( .A1(n_172), .A2(n_496), .B(n_497), .Y(n_495) );
AOI21xp5_ASAP7_75t_L g503 ( .A1(n_172), .A2(n_504), .B(n_505), .Y(n_503) );
AOI21xp5_ASAP7_75t_L g512 ( .A1(n_172), .A2(n_513), .B(n_514), .Y(n_512) );
AOI21xp5_ASAP7_75t_L g536 ( .A1(n_172), .A2(n_537), .B(n_538), .Y(n_536) );
AOI21xp5_ASAP7_75t_L g544 ( .A1(n_172), .A2(n_545), .B(n_546), .Y(n_544) );
INVx3_ASAP7_75t_L g236 ( .A(n_175), .Y(n_236) );
INVx1_ASAP7_75t_L g250 ( .A(n_176), .Y(n_250) );
INVx2_ASAP7_75t_L g254 ( .A(n_176), .Y(n_254) );
AND2x4_ASAP7_75t_SL g285 ( .A(n_176), .B(n_191), .Y(n_285) );
HB1xp67_ASAP7_75t_L g317 ( .A(n_176), .Y(n_317) );
INVx3_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
HB1xp67_ASAP7_75t_L g199 ( .A(n_177), .Y(n_199) );
AOI21x1_ASAP7_75t_L g177 ( .A1(n_178), .A2(n_179), .B(n_185), .Y(n_177) );
AO21x2_ASAP7_75t_L g541 ( .A1(n_178), .A2(n_542), .B(n_548), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_180), .B(n_184), .Y(n_179) );
AOI21xp5_ASAP7_75t_L g226 ( .A1(n_186), .A2(n_227), .B(n_228), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_188), .B(n_200), .Y(n_187) );
AND2x2_ASAP7_75t_L g351 ( .A(n_188), .B(n_296), .Y(n_351) );
INVx2_ASAP7_75t_SL g439 ( .A(n_188), .Y(n_439) );
INVx1_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_190), .B(n_199), .Y(n_189) );
NAND2x1p5_ASAP7_75t_L g252 ( .A(n_190), .B(n_253), .Y(n_252) );
AND2x2_ASAP7_75t_L g359 ( .A(n_190), .B(n_272), .Y(n_359) );
INVx4_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
BUFx2_ASAP7_75t_L g247 ( .A(n_191), .Y(n_247) );
AND2x4_ASAP7_75t_L g249 ( .A(n_191), .B(n_250), .Y(n_249) );
NOR2x1_ASAP7_75t_L g269 ( .A(n_191), .B(n_270), .Y(n_269) );
INVx1_ASAP7_75t_L g342 ( .A(n_191), .Y(n_342) );
AND2x2_ASAP7_75t_L g361 ( .A(n_191), .B(n_300), .Y(n_361) );
AND2x2_ASAP7_75t_L g392 ( .A(n_191), .B(n_301), .Y(n_392) );
OR2x6_ASAP7_75t_L g191 ( .A(n_192), .B(n_198), .Y(n_191) );
AND2x2_ASAP7_75t_L g331 ( .A(n_200), .B(n_285), .Y(n_331) );
NAND2xp5_ASAP7_75t_SL g367 ( .A(n_200), .B(n_342), .Y(n_367) );
AOI22xp5_ASAP7_75t_L g441 ( .A1(n_200), .A2(n_442), .B1(n_444), .B2(n_445), .Y(n_441) );
AND2x2_ASAP7_75t_L g444 ( .A(n_200), .B(n_251), .Y(n_444) );
INVx3_ASAP7_75t_L g297 ( .A(n_201), .Y(n_297) );
AND2x2_ASAP7_75t_L g300 ( .A(n_201), .B(n_301), .Y(n_300) );
AND2x2_ASAP7_75t_L g316 ( .A(n_202), .B(n_317), .Y(n_316) );
INVx1_ASAP7_75t_L g325 ( .A(n_202), .Y(n_325) );
AND2x4_ASAP7_75t_SL g203 ( .A(n_204), .B(n_214), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_204), .B(n_337), .Y(n_336) );
AND2x2_ASAP7_75t_L g376 ( .A(n_204), .B(n_377), .Y(n_376) );
NOR3xp33_ASAP7_75t_L g428 ( .A(n_204), .B(n_338), .C(n_429), .Y(n_428) );
OR2x2_ASAP7_75t_L g446 ( .A(n_204), .B(n_340), .Y(n_446) );
INVx3_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
OR2x2_ASAP7_75t_L g261 ( .A(n_206), .B(n_225), .Y(n_261) );
INVx1_ASAP7_75t_L g278 ( .A(n_206), .Y(n_278) );
INVx2_ASAP7_75t_L g291 ( .A(n_206), .Y(n_291) );
HB1xp67_ASAP7_75t_L g306 ( .A(n_206), .Y(n_306) );
AND2x2_ASAP7_75t_L g320 ( .A(n_206), .B(n_293), .Y(n_320) );
AND2x2_ASAP7_75t_L g399 ( .A(n_206), .B(n_216), .Y(n_399) );
AOI21xp5_ASAP7_75t_L g207 ( .A1(n_208), .A2(n_209), .B(n_213), .Y(n_207) );
AOI21xp5_ASAP7_75t_L g218 ( .A1(n_213), .A2(n_219), .B(n_220), .Y(n_218) );
INVx1_ASAP7_75t_SL g467 ( .A(n_213), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_213), .B(n_499), .Y(n_498) );
AOI21xp5_ASAP7_75t_L g533 ( .A1(n_213), .A2(n_534), .B(n_535), .Y(n_533) );
AOI221xp5_ASAP7_75t_L g262 ( .A1(n_214), .A2(n_263), .B1(n_266), .B2(n_273), .C(n_279), .Y(n_262) );
AOI221xp5_ASAP7_75t_L g391 ( .A1(n_214), .A2(n_392), .B1(n_393), .B2(n_394), .C(n_395), .Y(n_391) );
AND2x2_ASAP7_75t_L g214 ( .A(n_215), .B(n_224), .Y(n_214) );
INVx2_ASAP7_75t_L g333 ( .A(n_215), .Y(n_333) );
AND2x2_ASAP7_75t_L g393 ( .A(n_215), .B(n_277), .Y(n_393) );
AND2x2_ASAP7_75t_L g403 ( .A(n_215), .B(n_289), .Y(n_403) );
OR2x2_ASAP7_75t_L g443 ( .A(n_215), .B(n_327), .Y(n_443) );
INVx2_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
OR2x2_ASAP7_75t_SL g260 ( .A(n_216), .B(n_261), .Y(n_260) );
NAND2x1_ASAP7_75t_L g276 ( .A(n_216), .B(n_225), .Y(n_276) );
INVx4_ASAP7_75t_L g305 ( .A(n_216), .Y(n_305) );
OR2x2_ASAP7_75t_L g347 ( .A(n_216), .B(n_234), .Y(n_347) );
OR2x6_ASAP7_75t_L g216 ( .A(n_217), .B(n_218), .Y(n_216) );
AND2x2_ASAP7_75t_L g398 ( .A(n_224), .B(n_399), .Y(n_398) );
AND2x2_ASAP7_75t_L g224 ( .A(n_225), .B(n_234), .Y(n_224) );
INVx2_ASAP7_75t_SL g286 ( .A(n_225), .Y(n_286) );
NOR2x1_ASAP7_75t_SL g292 ( .A(n_225), .B(n_293), .Y(n_292) );
AND2x2_ASAP7_75t_L g307 ( .A(n_225), .B(n_308), .Y(n_307) );
OR2x2_ASAP7_75t_L g338 ( .A(n_225), .B(n_305), .Y(n_338) );
AND2x2_ASAP7_75t_L g345 ( .A(n_225), .B(n_291), .Y(n_345) );
BUFx2_ASAP7_75t_L g379 ( .A(n_225), .Y(n_379) );
AND2x2_ASAP7_75t_L g390 ( .A(n_225), .B(n_305), .Y(n_390) );
OR2x6_ASAP7_75t_L g225 ( .A(n_226), .B(n_233), .Y(n_225) );
HB1xp67_ASAP7_75t_L g258 ( .A(n_234), .Y(n_258) );
AND2x2_ASAP7_75t_L g277 ( .A(n_234), .B(n_278), .Y(n_277) );
INVx2_ASAP7_75t_L g308 ( .A(n_234), .Y(n_308) );
AND2x2_ASAP7_75t_L g334 ( .A(n_234), .B(n_290), .Y(n_334) );
INVx3_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
AO21x2_ASAP7_75t_L g235 ( .A1(n_236), .A2(n_237), .B(n_243), .Y(n_235) );
AO21x1_ASAP7_75t_SL g293 ( .A1(n_236), .A2(n_237), .B(n_243), .Y(n_293) );
AO21x2_ASAP7_75t_L g500 ( .A1(n_236), .A2(n_501), .B(n_507), .Y(n_500) );
AO21x2_ASAP7_75t_L g509 ( .A1(n_236), .A2(n_510), .B(n_516), .Y(n_509) );
AO21x2_ASAP7_75t_L g522 ( .A1(n_236), .A2(n_510), .B(n_516), .Y(n_522) );
AO21x2_ASAP7_75t_L g525 ( .A1(n_236), .A2(n_501), .B(n_507), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_238), .B(n_242), .Y(n_237) );
OAI31xp33_ASAP7_75t_L g244 ( .A1(n_245), .A2(n_249), .A3(n_251), .B(n_255), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_247), .B(n_248), .Y(n_246) );
INVx2_ASAP7_75t_L g353 ( .A(n_247), .Y(n_353) );
NOR2xp67_ASAP7_75t_L g263 ( .A(n_248), .B(n_264), .Y(n_263) );
AOI322xp5_ASAP7_75t_L g343 ( .A1(n_248), .A2(n_337), .A3(n_344), .B1(n_348), .B2(n_349), .C1(n_351), .C2(n_352), .Y(n_343) );
AND2x2_ASAP7_75t_L g415 ( .A(n_248), .B(n_392), .Y(n_415) );
AOI221xp5_ASAP7_75t_SL g328 ( .A1(n_249), .A2(n_329), .B1(n_331), .B2(n_332), .C(n_335), .Y(n_328) );
INVx2_ASAP7_75t_L g348 ( .A(n_249), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_251), .B(n_313), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_251), .B(n_344), .Y(n_447) );
INVx1_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
OR2x2_ASAP7_75t_L g322 ( .A(n_252), .B(n_297), .Y(n_322) );
INVx1_ASAP7_75t_SL g253 ( .A(n_254), .Y(n_253) );
AND2x2_ASAP7_75t_L g301 ( .A(n_254), .B(n_270), .Y(n_301) );
AND2x4_ASAP7_75t_L g255 ( .A(n_256), .B(n_259), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
INVx1_ASAP7_75t_L g372 ( .A(n_258), .Y(n_372) );
O2A1O1Ixp5_ASAP7_75t_L g363 ( .A1(n_259), .A2(n_364), .B(n_366), .C(n_368), .Y(n_363) );
INVx2_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
OAI22xp5_ASAP7_75t_L g395 ( .A1(n_260), .A2(n_396), .B1(n_397), .B2(n_400), .Y(n_395) );
OR2x2_ASAP7_75t_L g350 ( .A(n_261), .B(n_347), .Y(n_350) );
INVx1_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
NAND2xp5_ASAP7_75t_SL g266 ( .A(n_267), .B(n_271), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
INVx1_ASAP7_75t_L g283 ( .A(n_270), .Y(n_283) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_272), .B(n_296), .Y(n_295) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_275), .B(n_277), .Y(n_274) );
INVx3_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
OR2x2_ASAP7_75t_L g326 ( .A(n_276), .B(n_327), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_276), .B(n_277), .Y(n_369) );
OR2x2_ASAP7_75t_L g371 ( .A(n_276), .B(n_372), .Y(n_371) );
NOR2xp33_ASAP7_75t_L g419 ( .A(n_276), .B(n_420), .Y(n_419) );
BUFx2_ASAP7_75t_L g287 ( .A(n_278), .Y(n_287) );
NOR4xp25_ASAP7_75t_L g279 ( .A(n_280), .B(n_284), .C(n_286), .D(n_287), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
AND2x2_ASAP7_75t_L g407 ( .A(n_281), .B(n_408), .Y(n_407) );
AND2x2_ASAP7_75t_L g435 ( .A(n_281), .B(n_284), .Y(n_435) );
INVx2_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
INVx1_ASAP7_75t_L g365 ( .A(n_283), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_284), .B(n_313), .Y(n_400) );
AOI321xp33_ASAP7_75t_L g402 ( .A1(n_284), .A2(n_403), .A3(n_404), .B1(n_405), .B2(n_407), .C(n_410), .Y(n_402) );
INVx2_ASAP7_75t_SL g284 ( .A(n_285), .Y(n_284) );
AND2x2_ASAP7_75t_SL g364 ( .A(n_285), .B(n_365), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_285), .B(n_324), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_286), .B(n_308), .Y(n_413) );
OR2x2_ASAP7_75t_L g440 ( .A(n_287), .B(n_324), .Y(n_440) );
AOI21xp5_ASAP7_75t_L g288 ( .A1(n_289), .A2(n_294), .B(n_298), .Y(n_288) );
AND2x2_ASAP7_75t_L g329 ( .A(n_289), .B(n_330), .Y(n_329) );
AND2x2_ASAP7_75t_L g289 ( .A(n_290), .B(n_292), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
AND2x2_ASAP7_75t_L g355 ( .A(n_291), .B(n_293), .Y(n_355) );
INVx2_ASAP7_75t_L g340 ( .A(n_292), .Y(n_340) );
INVx1_ASAP7_75t_SL g294 ( .A(n_295), .Y(n_294) );
NOR2xp33_ASAP7_75t_L g410 ( .A(n_295), .B(n_411), .Y(n_410) );
OR2x2_ASAP7_75t_L g396 ( .A(n_296), .B(n_348), .Y(n_396) );
INVx2_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
AND2x2_ASAP7_75t_L g354 ( .A(n_297), .B(n_355), .Y(n_354) );
NOR2x1_ASAP7_75t_L g432 ( .A(n_297), .B(n_433), .Y(n_432) );
NOR2xp67_ASAP7_75t_L g298 ( .A(n_299), .B(n_302), .Y(n_298) );
INVx2_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
INVx1_ASAP7_75t_L g383 ( .A(n_301), .Y(n_383) );
INVx2_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
AND2x2_ASAP7_75t_L g303 ( .A(n_304), .B(n_307), .Y(n_303) );
NOR2xp67_ASAP7_75t_L g304 ( .A(n_305), .B(n_306), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_305), .B(n_320), .Y(n_319) );
INVx1_ASAP7_75t_L g330 ( .A(n_305), .Y(n_330) );
BUFx2_ASAP7_75t_L g412 ( .A(n_305), .Y(n_412) );
INVxp67_ASAP7_75t_L g420 ( .A(n_308), .Y(n_420) );
NAND3xp33_ASAP7_75t_L g309 ( .A(n_310), .B(n_328), .C(n_343), .Y(n_309) );
AOI21xp5_ASAP7_75t_L g310 ( .A1(n_311), .A2(n_318), .B(n_321), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_312), .B(n_315), .Y(n_311) );
INVx2_ASAP7_75t_SL g313 ( .A(n_314), .Y(n_313) );
OR2x2_ASAP7_75t_L g341 ( .A(n_314), .B(n_342), .Y(n_341) );
INVx2_ASAP7_75t_L g394 ( .A(n_315), .Y(n_394) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
INVx2_ASAP7_75t_L g409 ( .A(n_317), .Y(n_409) );
AOI21xp5_ASAP7_75t_L g414 ( .A1(n_318), .A2(n_415), .B(n_416), .Y(n_414) );
INVx1_ASAP7_75t_SL g318 ( .A(n_319), .Y(n_318) );
INVx2_ASAP7_75t_SL g327 ( .A(n_320), .Y(n_327) );
AND2x2_ASAP7_75t_L g389 ( .A(n_320), .B(n_390), .Y(n_389) );
AOI21xp33_ASAP7_75t_L g321 ( .A1(n_322), .A2(n_323), .B(n_326), .Y(n_321) );
OAI22xp5_ASAP7_75t_L g368 ( .A1(n_322), .A2(n_369), .B1(n_370), .B2(n_371), .Y(n_368) );
OR2x2_ASAP7_75t_L g323 ( .A(n_324), .B(n_325), .Y(n_323) );
INVx1_ASAP7_75t_L g358 ( .A(n_324), .Y(n_358) );
OR2x2_ASAP7_75t_L g406 ( .A(n_327), .B(n_338), .Y(n_406) );
NOR4xp25_ASAP7_75t_L g438 ( .A(n_330), .B(n_379), .C(n_439), .D(n_440), .Y(n_438) );
AND2x2_ASAP7_75t_L g332 ( .A(n_333), .B(n_334), .Y(n_332) );
OR2x2_ASAP7_75t_L g339 ( .A(n_333), .B(n_340), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_333), .B(n_355), .Y(n_437) );
AOI21xp33_ASAP7_75t_SL g335 ( .A1(n_336), .A2(n_339), .B(n_341), .Y(n_335) );
INVx2_ASAP7_75t_SL g337 ( .A(n_338), .Y(n_337) );
OR2x2_ASAP7_75t_L g426 ( .A(n_338), .B(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g434 ( .A(n_340), .Y(n_434) );
AND2x4_ASAP7_75t_L g344 ( .A(n_345), .B(n_346), .Y(n_344) );
INVxp67_ASAP7_75t_L g362 ( .A(n_345), .Y(n_362) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
OR2x2_ASAP7_75t_L g378 ( .A(n_347), .B(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
AND2x2_ASAP7_75t_L g352 ( .A(n_353), .B(n_354), .Y(n_352) );
AND2x2_ASAP7_75t_L g381 ( .A(n_353), .B(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g427 ( .A(n_355), .Y(n_427) );
A2O1A1Ixp33_ASAP7_75t_L g356 ( .A1(n_357), .A2(n_360), .B(n_362), .C(n_363), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_358), .B(n_359), .Y(n_357) );
INVx1_ASAP7_75t_L g417 ( .A(n_359), .Y(n_417) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
INVxp67_ASAP7_75t_L g421 ( .A(n_364), .Y(n_421) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
NOR3xp33_ASAP7_75t_L g373 ( .A(n_374), .B(n_401), .C(n_422), .Y(n_373) );
OAI211xp5_ASAP7_75t_SL g374 ( .A1(n_375), .A2(n_380), .B(n_384), .C(n_391), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx1_ASAP7_75t_SL g377 ( .A(n_378), .Y(n_377) );
INVxp67_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx2_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
OAI21xp5_ASAP7_75t_SL g384 ( .A1(n_385), .A2(n_387), .B(n_389), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
O2A1O1Ixp33_ASAP7_75t_L g423 ( .A1(n_387), .A2(n_424), .B(n_425), .C(n_428), .Y(n_423) );
BUFx2_ASAP7_75t_L g404 ( .A(n_388), .Y(n_404) );
INVx2_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_402), .B(n_414), .Y(n_401) );
INVx2_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx2_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
OAI22xp5_ASAP7_75t_L g416 ( .A1(n_411), .A2(n_417), .B1(n_418), .B2(n_421), .Y(n_416) );
OR2x2_ASAP7_75t_L g411 ( .A(n_412), .B(n_413), .Y(n_411) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
NAND4xp25_ASAP7_75t_L g422 ( .A(n_423), .B(n_431), .C(n_441), .D(n_447), .Y(n_422) );
INVx2_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
AOI221xp5_ASAP7_75t_L g431 ( .A1(n_432), .A2(n_434), .B1(n_435), .B2(n_436), .C(n_438), .Y(n_431) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
CKINVDCx6p67_ASAP7_75t_R g448 ( .A(n_449), .Y(n_448) );
INVx3_ASAP7_75t_SL g449 ( .A(n_450), .Y(n_449) );
OAI22xp5_ASAP7_75t_L g751 ( .A1(n_450), .A2(n_752), .B1(n_753), .B2(n_754), .Y(n_751) );
CKINVDCx5p33_ASAP7_75t_R g450 ( .A(n_451), .Y(n_450) );
INVx3_ASAP7_75t_SL g754 ( .A(n_452), .Y(n_754) );
NOR2x2_ASAP7_75t_L g452 ( .A(n_453), .B(n_631), .Y(n_452) );
AO211x2_ASAP7_75t_L g453 ( .A1(n_454), .A2(n_476), .B(n_526), .C(n_599), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVxp67_ASAP7_75t_SL g455 ( .A(n_456), .Y(n_455) );
AND3x2_ASAP7_75t_L g680 ( .A(n_456), .B(n_561), .C(n_577), .Y(n_680) );
AND2x4_ASAP7_75t_L g683 ( .A(n_456), .B(n_684), .Y(n_683) );
AND2x2_ASAP7_75t_L g456 ( .A(n_457), .B(n_466), .Y(n_456) );
NAND2x1p5_ASAP7_75t_L g539 ( .A(n_457), .B(n_540), .Y(n_539) );
INVx4_ASAP7_75t_L g592 ( .A(n_457), .Y(n_592) );
AND2x2_ASAP7_75t_SL g677 ( .A(n_457), .B(n_586), .Y(n_677) );
AND2x2_ASAP7_75t_L g720 ( .A(n_457), .B(n_541), .Y(n_720) );
INVx5_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
BUFx2_ASAP7_75t_L g569 ( .A(n_458), .Y(n_569) );
AND2x2_ASAP7_75t_L g588 ( .A(n_458), .B(n_532), .Y(n_588) );
AND2x2_ASAP7_75t_L g606 ( .A(n_458), .B(n_541), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_458), .B(n_540), .Y(n_666) );
NOR2x1_ASAP7_75t_SL g693 ( .A(n_458), .B(n_466), .Y(n_693) );
OR2x6_ASAP7_75t_L g458 ( .A(n_459), .B(n_460), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_466), .B(n_532), .Y(n_531) );
AO21x2_ASAP7_75t_L g466 ( .A1(n_467), .A2(n_468), .B(n_474), .Y(n_466) );
NOR2xp33_ASAP7_75t_L g474 ( .A(n_467), .B(n_475), .Y(n_474) );
AO21x2_ASAP7_75t_L g565 ( .A1(n_467), .A2(n_468), .B(n_474), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_469), .B(n_473), .Y(n_468) );
AO21x1_ASAP7_75t_L g476 ( .A1(n_477), .A2(n_508), .B(n_517), .Y(n_476) );
INVx2_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
OAI22xp33_ASAP7_75t_L g574 ( .A1(n_478), .A2(n_575), .B1(n_579), .B2(n_580), .Y(n_574) );
OR2x2_ASAP7_75t_L g478 ( .A(n_479), .B(n_487), .Y(n_478) );
AND2x2_ASAP7_75t_L g635 ( .A(n_479), .B(n_523), .Y(n_635) );
BUFx2_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
AND2x4_ASAP7_75t_L g568 ( .A(n_480), .B(n_551), .Y(n_568) );
AND2x2_ASAP7_75t_L g640 ( .A(n_480), .B(n_525), .Y(n_640) );
AND2x2_ASAP7_75t_L g659 ( .A(n_480), .B(n_625), .Y(n_659) );
INVx2_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
INVx2_ASAP7_75t_L g518 ( .A(n_481), .Y(n_518) );
HB1xp67_ASAP7_75t_L g646 ( .A(n_481), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_487), .B(n_629), .Y(n_628) );
INVx2_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
AND2x2_ASAP7_75t_L g619 ( .A(n_488), .B(n_520), .Y(n_619) );
AND2x4_ASAP7_75t_L g488 ( .A(n_489), .B(n_500), .Y(n_488) );
AND2x2_ASAP7_75t_L g523 ( .A(n_489), .B(n_524), .Y(n_523) );
OR2x2_ASAP7_75t_L g556 ( .A(n_489), .B(n_557), .Y(n_556) );
AND2x2_ASAP7_75t_SL g616 ( .A(n_489), .B(n_552), .Y(n_616) );
INVx2_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
BUFx2_ASAP7_75t_L g709 ( .A(n_490), .Y(n_709) );
INVx2_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
INVx2_ASAP7_75t_L g551 ( .A(n_491), .Y(n_551) );
OAI21x1_ASAP7_75t_SL g491 ( .A1(n_492), .A2(n_494), .B(n_498), .Y(n_491) );
INVx1_ASAP7_75t_L g499 ( .A(n_493), .Y(n_499) );
INVx2_ASAP7_75t_L g557 ( .A(n_500), .Y(n_557) );
HB1xp67_ASAP7_75t_L g657 ( .A(n_500), .Y(n_657) );
NAND2xp5_ASAP7_75t_SL g501 ( .A(n_502), .B(n_506), .Y(n_501) );
INVx2_ASAP7_75t_L g553 ( .A(n_508), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_508), .B(n_685), .Y(n_711) );
AND2x2_ASAP7_75t_L g730 ( .A(n_508), .B(n_720), .Y(n_730) );
BUFx2_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
AND2x4_ASAP7_75t_SL g598 ( .A(n_509), .B(n_557), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_511), .B(n_515), .Y(n_510) );
AND2x2_ASAP7_75t_SL g517 ( .A(n_518), .B(n_519), .Y(n_517) );
AND2x2_ASAP7_75t_L g597 ( .A(n_518), .B(n_598), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_518), .B(n_567), .Y(n_602) );
INVx1_ASAP7_75t_SL g729 ( .A(n_518), .Y(n_729) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_519), .B(n_680), .Y(n_679) );
AND2x2_ASAP7_75t_L g519 ( .A(n_520), .B(n_523), .Y(n_519) );
INVx1_ASAP7_75t_L g555 ( .A(n_520), .Y(n_555) );
AND2x2_ASAP7_75t_L g741 ( .A(n_520), .B(n_742), .Y(n_741) );
BUFx2_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
AND2x2_ASAP7_75t_L g617 ( .A(n_521), .B(n_524), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_521), .B(n_630), .Y(n_629) );
AND2x2_ASAP7_75t_L g671 ( .A(n_521), .B(n_525), .Y(n_671) );
AND2x2_ASAP7_75t_L g702 ( .A(n_521), .B(n_703), .Y(n_702) );
INVx2_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
AND2x2_ASAP7_75t_L g567 ( .A(n_522), .B(n_525), .Y(n_567) );
INVxp67_ASAP7_75t_L g584 ( .A(n_522), .Y(n_584) );
BUFx3_ASAP7_75t_L g625 ( .A(n_522), .Y(n_625) );
AND2x2_ASAP7_75t_L g645 ( .A(n_523), .B(n_646), .Y(n_645) );
NAND2xp33_ASAP7_75t_L g658 ( .A(n_523), .B(n_659), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_524), .B(n_551), .Y(n_614) );
AND2x2_ASAP7_75t_L g703 ( .A(n_524), .B(n_552), .Y(n_703) );
INVx2_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
AND2x2_ASAP7_75t_L g630 ( .A(n_525), .B(n_552), .Y(n_630) );
OR3x1_ASAP7_75t_L g526 ( .A(n_527), .B(n_574), .C(n_589), .Y(n_526) );
OAI321xp33_ASAP7_75t_L g527 ( .A1(n_528), .A2(n_539), .A3(n_549), .B1(n_554), .B2(n_558), .C(n_566), .Y(n_527) );
INVx1_ASAP7_75t_SL g528 ( .A(n_529), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
INVxp67_ASAP7_75t_SL g605 ( .A(n_531), .Y(n_605) );
INVxp67_ASAP7_75t_SL g623 ( .A(n_531), .Y(n_623) );
OR2x2_ASAP7_75t_L g627 ( .A(n_531), .B(n_539), .Y(n_627) );
BUFx3_ASAP7_75t_L g561 ( .A(n_532), .Y(n_561) );
AND2x2_ASAP7_75t_L g578 ( .A(n_532), .B(n_564), .Y(n_578) );
INVx1_ASAP7_75t_L g595 ( .A(n_532), .Y(n_595) );
INVx2_ASAP7_75t_L g611 ( .A(n_532), .Y(n_611) );
OR2x2_ASAP7_75t_L g650 ( .A(n_532), .B(n_540), .Y(n_650) );
INVx2_ASAP7_75t_L g638 ( .A(n_539), .Y(n_638) );
AND2x2_ASAP7_75t_L g562 ( .A(n_540), .B(n_563), .Y(n_562) );
INVx2_ASAP7_75t_L g577 ( .A(n_540), .Y(n_577) );
AND2x4_ASAP7_75t_L g586 ( .A(n_540), .B(n_587), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_540), .B(n_563), .Y(n_609) );
AND2x2_ASAP7_75t_L g716 ( .A(n_540), .B(n_611), .Y(n_716) );
INVx4_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
HB1xp67_ASAP7_75t_L g675 ( .A(n_541), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_543), .B(n_547), .Y(n_542) );
INVx1_ASAP7_75t_L g603 ( .A(n_549), .Y(n_603) );
NAND2xp5_ASAP7_75t_SL g549 ( .A(n_550), .B(n_553), .Y(n_549) );
AND2x2_ASAP7_75t_L g690 ( .A(n_550), .B(n_617), .Y(n_690) );
INVx1_ASAP7_75t_SL g707 ( .A(n_550), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g736 ( .A(n_550), .B(n_683), .Y(n_736) );
AND2x4_ASAP7_75t_L g550 ( .A(n_551), .B(n_552), .Y(n_550) );
OR2x2_ASAP7_75t_L g579 ( .A(n_551), .B(n_552), .Y(n_579) );
AND2x2_ASAP7_75t_L g672 ( .A(n_553), .B(n_568), .Y(n_672) );
OR2x2_ASAP7_75t_L g554 ( .A(n_555), .B(n_556), .Y(n_554) );
NAND2xp5_ASAP7_75t_SL g695 ( .A(n_557), .B(n_568), .Y(n_695) );
INVx2_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
AOI22xp33_ASAP7_75t_L g712 ( .A1(n_559), .A2(n_708), .B1(n_713), .B2(n_715), .Y(n_712) );
AND2x4_ASAP7_75t_L g559 ( .A(n_560), .B(n_562), .Y(n_559) );
AND2x2_ASAP7_75t_L g637 ( .A(n_560), .B(n_638), .Y(n_637) );
OR2x2_ASAP7_75t_L g732 ( .A(n_560), .B(n_733), .Y(n_732) );
INVx2_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
AND2x2_ASAP7_75t_L g688 ( .A(n_561), .B(n_606), .Y(n_688) );
AND2x4_ASAP7_75t_L g642 ( .A(n_562), .B(n_588), .Y(n_642) );
INVx1_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
HB1xp67_ASAP7_75t_L g740 ( .A(n_564), .Y(n_740) );
INVx2_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
INVx1_ASAP7_75t_L g573 ( .A(n_565), .Y(n_573) );
INVx1_ASAP7_75t_L g587 ( .A(n_565), .Y(n_587) );
NAND4xp25_ASAP7_75t_L g566 ( .A(n_567), .B(n_568), .C(n_569), .D(n_570), .Y(n_566) );
AND2x2_ASAP7_75t_L g724 ( .A(n_567), .B(n_709), .Y(n_724) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_567), .B(n_735), .Y(n_734) );
NOR2xp33_ASAP7_75t_L g643 ( .A(n_568), .B(n_644), .Y(n_643) );
OAI322xp33_ASAP7_75t_L g651 ( .A1(n_568), .A2(n_652), .A3(n_656), .B1(n_658), .B2(n_660), .C1(n_662), .C2(n_667), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_568), .B(n_617), .Y(n_667) );
INVx1_ASAP7_75t_L g735 ( .A(n_568), .Y(n_735) );
INVx2_ASAP7_75t_L g581 ( .A(n_569), .Y(n_581) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
INVx2_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_572), .B(n_675), .Y(n_674) );
INVx2_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_573), .B(n_592), .Y(n_649) );
INVx1_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_576), .B(n_619), .Y(n_618) );
AND2x2_ASAP7_75t_L g576 ( .A(n_577), .B(n_578), .Y(n_576) );
INVx1_ASAP7_75t_L g622 ( .A(n_577), .Y(n_622) );
AND2x2_ASAP7_75t_L g694 ( .A(n_577), .B(n_605), .Y(n_694) );
AOI31xp33_ASAP7_75t_L g580 ( .A1(n_578), .A2(n_581), .A3(n_582), .B(n_585), .Y(n_580) );
AND2x2_ASAP7_75t_L g591 ( .A(n_578), .B(n_592), .Y(n_591) );
AND2x2_ASAP7_75t_L g719 ( .A(n_578), .B(n_720), .Y(n_719) );
AND2x2_ASAP7_75t_SL g726 ( .A(n_578), .B(n_606), .Y(n_726) );
INVx1_ASAP7_75t_L g727 ( .A(n_578), .Y(n_727) );
INVx1_ASAP7_75t_SL g685 ( .A(n_579), .Y(n_685) );
NAND3xp33_ASAP7_75t_SL g713 ( .A(n_579), .B(n_707), .C(n_714), .Y(n_713) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
OR2x2_ASAP7_75t_L g613 ( .A(n_584), .B(n_614), .Y(n_613) );
AND2x2_ASAP7_75t_L g585 ( .A(n_586), .B(n_588), .Y(n_585) );
AND2x2_ASAP7_75t_L g594 ( .A(n_586), .B(n_595), .Y(n_594) );
INVx2_ASAP7_75t_L g655 ( .A(n_586), .Y(n_655) );
AOI322xp5_ASAP7_75t_L g737 ( .A1(n_586), .A2(n_616), .A3(n_619), .B1(n_738), .B2(n_739), .C1(n_741), .C2(n_743), .Y(n_737) );
AND2x2_ASAP7_75t_L g743 ( .A(n_586), .B(n_592), .Y(n_743) );
AOI21xp5_ASAP7_75t_L g589 ( .A1(n_590), .A2(n_593), .B(n_596), .Y(n_589) );
INVx1_ASAP7_75t_SL g590 ( .A(n_591), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_592), .B(n_611), .Y(n_610) );
AND2x4_ASAP7_75t_L g738 ( .A(n_592), .B(n_625), .Y(n_738) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
INVx1_ASAP7_75t_L g664 ( .A(n_595), .Y(n_664) );
AND2x2_ASAP7_75t_L g692 ( .A(n_595), .B(n_693), .Y(n_692) );
AND2x2_ASAP7_75t_L g739 ( .A(n_595), .B(n_740), .Y(n_739) );
INVx1_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
INVx1_ASAP7_75t_L g644 ( .A(n_598), .Y(n_644) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
O2A1O1Ixp5_ASAP7_75t_L g600 ( .A1(n_601), .A2(n_603), .B(n_604), .C(n_607), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
AND2x2_ASAP7_75t_L g604 ( .A(n_605), .B(n_606), .Y(n_604) );
AND2x2_ASAP7_75t_L g661 ( .A(n_606), .B(n_611), .Y(n_661) );
OAI211xp5_ASAP7_75t_L g607 ( .A1(n_608), .A2(n_612), .B(n_618), .C(n_620), .Y(n_607) );
OAI221xp5_ASAP7_75t_L g633 ( .A1(n_608), .A2(n_634), .B1(n_636), .B2(n_639), .C(n_641), .Y(n_633) );
OR2x2_ASAP7_75t_L g608 ( .A(n_609), .B(n_610), .Y(n_608) );
INVx1_ASAP7_75t_L g653 ( .A(n_610), .Y(n_653) );
OR2x2_ASAP7_75t_L g673 ( .A(n_610), .B(n_674), .Y(n_673) );
AND2x2_ASAP7_75t_L g612 ( .A(n_613), .B(n_615), .Y(n_612) );
INVx1_ASAP7_75t_L g718 ( .A(n_613), .Y(n_718) );
INVx1_ASAP7_75t_L g742 ( .A(n_614), .Y(n_742) );
NAND2xp5_ASAP7_75t_SL g615 ( .A(n_616), .B(n_617), .Y(n_615) );
AND2x2_ASAP7_75t_L g624 ( .A(n_616), .B(n_625), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_616), .B(n_686), .Y(n_698) );
INVx1_ASAP7_75t_L g678 ( .A(n_617), .Y(n_678) );
AOI22xp5_ASAP7_75t_L g620 ( .A1(n_621), .A2(n_624), .B1(n_626), .B2(n_628), .Y(n_620) );
AND2x2_ASAP7_75t_L g621 ( .A(n_622), .B(n_623), .Y(n_621) );
INVx1_ASAP7_75t_SL g686 ( .A(n_625), .Y(n_686) );
INVx2_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
NAND4xp75_ASAP7_75t_L g631 ( .A(n_632), .B(n_668), .C(n_696), .D(n_721), .Y(n_631) );
NOR2xp67_ASAP7_75t_L g632 ( .A(n_633), .B(n_651), .Y(n_632) );
INVx1_ASAP7_75t_SL g634 ( .A(n_635), .Y(n_634) );
INVx2_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
AND2x2_ASAP7_75t_SL g708 ( .A(n_640), .B(n_709), .Y(n_708) );
AOI22xp5_ASAP7_75t_L g641 ( .A1(n_642), .A2(n_643), .B1(n_645), .B2(n_647), .Y(n_641) );
NOR2xp33_ASAP7_75t_L g706 ( .A(n_644), .B(n_707), .Y(n_706) );
INVx2_ASAP7_75t_SL g647 ( .A(n_648), .Y(n_647) );
OR2x2_ASAP7_75t_L g648 ( .A(n_649), .B(n_650), .Y(n_648) );
INVx2_ASAP7_75t_L g684 ( .A(n_650), .Y(n_684) );
OR2x2_ASAP7_75t_L g699 ( .A(n_650), .B(n_700), .Y(n_699) );
NAND2xp5_ASAP7_75t_SL g652 ( .A(n_653), .B(n_654), .Y(n_652) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
INVx1_ASAP7_75t_L g714 ( .A(n_659), .Y(n_714) );
INVx1_ASAP7_75t_SL g660 ( .A(n_661), .Y(n_660) );
OAI21xp5_ASAP7_75t_SL g705 ( .A1(n_661), .A2(n_706), .B(n_708), .Y(n_705) );
INVxp67_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
AND2x2_ASAP7_75t_L g663 ( .A(n_664), .B(n_665), .Y(n_663) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
NOR2x1_ASAP7_75t_L g668 ( .A(n_669), .B(n_681), .Y(n_668) );
OAI221xp5_ASAP7_75t_L g669 ( .A1(n_670), .A2(n_673), .B1(n_676), .B2(n_678), .C(n_679), .Y(n_669) );
NOR2xp33_ASAP7_75t_L g670 ( .A(n_671), .B(n_672), .Y(n_670) );
OAI21xp33_ASAP7_75t_L g717 ( .A1(n_671), .A2(n_718), .B(n_719), .Y(n_717) );
INVx3_ASAP7_75t_SL g676 ( .A(n_677), .Y(n_676) );
OAI322xp33_ASAP7_75t_L g681 ( .A1(n_682), .A2(n_685), .A3(n_686), .B1(n_687), .B2(n_689), .C1(n_691), .C2(n_695), .Y(n_681) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
INVx1_ASAP7_75t_SL g689 ( .A(n_690), .Y(n_689) );
NOR2x1_ASAP7_75t_L g691 ( .A(n_692), .B(n_694), .Y(n_691) );
INVx1_ASAP7_75t_L g704 ( .A(n_692), .Y(n_704) );
INVx1_ASAP7_75t_L g700 ( .A(n_693), .Y(n_700) );
AND2x2_ASAP7_75t_L g715 ( .A(n_693), .B(n_716), .Y(n_715) );
NOR2x1_ASAP7_75t_L g696 ( .A(n_697), .B(n_710), .Y(n_696) );
OAI221xp5_ASAP7_75t_L g697 ( .A1(n_698), .A2(n_699), .B1(n_701), .B2(n_704), .C(n_705), .Y(n_697) );
INVx1_ASAP7_75t_SL g701 ( .A(n_702), .Y(n_701) );
OAI211xp5_ASAP7_75t_SL g710 ( .A1(n_704), .A2(n_711), .B(n_712), .C(n_717), .Y(n_710) );
INVx2_ASAP7_75t_SL g733 ( .A(n_720), .Y(n_733) );
NOR2x1_ASAP7_75t_L g721 ( .A(n_722), .B(n_731), .Y(n_721) );
OAI22xp33_ASAP7_75t_L g722 ( .A1(n_723), .A2(n_725), .B1(n_727), .B2(n_728), .Y(n_722) );
INVx1_ASAP7_75t_SL g723 ( .A(n_724), .Y(n_723) );
INVx2_ASAP7_75t_SL g725 ( .A(n_726), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_729), .B(n_730), .Y(n_728) );
OAI211xp5_ASAP7_75t_SL g731 ( .A1(n_732), .A2(n_734), .B(n_736), .C(n_737), .Y(n_731) );
CKINVDCx20_ASAP7_75t_R g744 ( .A(n_745), .Y(n_744) );
INVx1_ASAP7_75t_SL g753 ( .A(n_745), .Y(n_753) );
CKINVDCx11_ASAP7_75t_R g745 ( .A(n_746), .Y(n_745) );
CKINVDCx12_ASAP7_75t_R g747 ( .A(n_748), .Y(n_747) );
NOR2xp33_ASAP7_75t_L g755 ( .A(n_756), .B(n_757), .Y(n_755) );
INVx1_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
INVx3_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
INVx1_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
OAI21xp33_ASAP7_75t_L g762 ( .A1(n_763), .A2(n_766), .B(n_771), .Y(n_762) );
CKINVDCx11_ASAP7_75t_R g763 ( .A(n_764), .Y(n_763) );
INVx1_ASAP7_75t_SL g764 ( .A(n_765), .Y(n_764) );
INVx1_ASAP7_75t_L g770 ( .A(n_767), .Y(n_770) );
INVx1_ASAP7_75t_SL g773 ( .A(n_774), .Y(n_773) );
CKINVDCx11_ASAP7_75t_R g775 ( .A(n_776), .Y(n_775) );
CKINVDCx8_ASAP7_75t_R g776 ( .A(n_777), .Y(n_776) );
INVx2_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
endmodule