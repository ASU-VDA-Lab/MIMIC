module fake_jpeg_30513_n_319 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_319);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_319;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx6_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_13),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_16),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx24_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_7),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_9),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_13),
.B(n_11),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

BUFx16f_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

BUFx12_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_12),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

INVx1_ASAP7_75t_SL g41 ( 
.A(n_6),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_14),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_43),
.Y(n_83)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_44),
.Y(n_104)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_45),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_32),
.B(n_7),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_46),
.B(n_52),
.Y(n_87)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_19),
.Y(n_47)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_47),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_20),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_20),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_49),
.Y(n_89)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_19),
.Y(n_50)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_50),
.Y(n_85)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_51),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_35),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_53),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_32),
.B(n_16),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_54),
.B(n_63),
.Y(n_94)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_27),
.Y(n_55)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_55),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_26),
.Y(n_56)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_56),
.Y(n_96)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_26),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_57),
.Y(n_90)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_26),
.Y(n_58)
);

INVx1_ASAP7_75t_SL g81 ( 
.A(n_58),
.Y(n_81)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g105 ( 
.A(n_59),
.Y(n_105)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_60),
.Y(n_108)
);

INVx4_ASAP7_75t_SL g61 ( 
.A(n_35),
.Y(n_61)
);

INVx4_ASAP7_75t_SL g75 ( 
.A(n_61),
.Y(n_75)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_20),
.Y(n_62)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_62),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_34),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_34),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_64),
.B(n_65),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_42),
.B(n_6),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_22),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_66),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_22),
.Y(n_67)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_67),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_22),
.A2(n_6),
.B1(n_14),
.B2(n_2),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_68),
.A2(n_30),
.B1(n_31),
.B2(n_28),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_44),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_69),
.B(n_97),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_53),
.B(n_42),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_70),
.B(n_78),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_51),
.B(n_41),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_72),
.B(n_93),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_43),
.A2(n_41),
.B1(n_39),
.B2(n_36),
.Y(n_74)
);

AO21x1_ASAP7_75t_L g116 ( 
.A1(n_74),
.A2(n_95),
.B(n_102),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

INVx5_ASAP7_75t_SL g139 ( 
.A(n_76),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_52),
.B(n_21),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_61),
.B(n_21),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_79),
.B(n_55),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_82),
.A2(n_37),
.B1(n_29),
.B2(n_24),
.Y(n_127)
);

BUFx12_ASAP7_75t_L g88 ( 
.A(n_60),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_88),
.B(n_75),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_62),
.A2(n_41),
.B1(n_17),
.B2(n_40),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_91),
.A2(n_98),
.B1(n_106),
.B2(n_1),
.Y(n_144)
);

NAND2xp33_ASAP7_75t_SL g93 ( 
.A(n_45),
.B(n_17),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_43),
.A2(n_39),
.B1(n_36),
.B2(n_19),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_59),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_48),
.A2(n_17),
.B1(n_25),
.B2(n_36),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_49),
.A2(n_18),
.B1(n_31),
.B2(n_30),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g132 ( 
.A1(n_99),
.A2(n_24),
.B1(n_23),
.B2(n_4),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_59),
.B(n_38),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_100),
.B(n_101),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_56),
.B(n_28),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_56),
.A2(n_19),
.B1(n_18),
.B2(n_38),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_67),
.A2(n_19),
.B1(n_25),
.B2(n_29),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_58),
.A2(n_37),
.B1(n_29),
.B2(n_24),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_107),
.A2(n_66),
.B1(n_57),
.B2(n_37),
.Y(n_117)
);

OA22x2_ASAP7_75t_L g111 ( 
.A1(n_50),
.A2(n_29),
.B1(n_24),
.B2(n_23),
.Y(n_111)
);

OA22x2_ASAP7_75t_L g135 ( 
.A1(n_111),
.A2(n_23),
.B1(n_1),
.B2(n_4),
.Y(n_135)
);

OR2x2_ASAP7_75t_SL g113 ( 
.A(n_72),
.B(n_58),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_R g183 ( 
.A(n_113),
.B(n_135),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_115),
.B(n_118),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_117),
.A2(n_127),
.B1(n_81),
.B2(n_96),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_71),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_104),
.B(n_66),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_119),
.B(n_123),
.Y(n_154)
);

OR2x2_ASAP7_75t_L g120 ( 
.A(n_103),
.B(n_37),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_120),
.B(n_125),
.Y(n_151)
);

BUFx5_ASAP7_75t_L g121 ( 
.A(n_105),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g161 ( 
.A(n_121),
.Y(n_161)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_90),
.Y(n_122)
);

INVx1_ASAP7_75t_SL g181 ( 
.A(n_122),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_110),
.B(n_0),
.Y(n_123)
);

BUFx2_ASAP7_75t_L g124 ( 
.A(n_90),
.Y(n_124)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_124),
.Y(n_170)
);

OAI32xp33_ASAP7_75t_L g125 ( 
.A1(n_93),
.A2(n_94),
.A3(n_87),
.B1(n_72),
.B2(n_86),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_75),
.B(n_0),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_126),
.B(n_138),
.Y(n_155)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_77),
.Y(n_128)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_128),
.Y(n_159)
);

NAND3xp33_ASAP7_75t_L g129 ( 
.A(n_83),
.B(n_10),
.C(n_2),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_129),
.B(n_133),
.Y(n_153)
);

INVx1_ASAP7_75t_SL g130 ( 
.A(n_83),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_130),
.B(n_135),
.Y(n_157)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_92),
.Y(n_131)
);

BUFx4f_ASAP7_75t_SL g179 ( 
.A(n_131),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_132),
.A2(n_142),
.B1(n_127),
.B2(n_138),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_111),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_134),
.B(n_136),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_71),
.Y(n_136)
);

BUFx12f_ASAP7_75t_L g137 ( 
.A(n_92),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_137),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_106),
.B(n_1),
.Y(n_138)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_84),
.Y(n_141)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_141),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_109),
.A2(n_23),
.B1(n_3),
.B2(n_5),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_77),
.Y(n_143)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_143),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_144),
.A2(n_147),
.B1(n_8),
.B2(n_12),
.Y(n_150)
);

INVx8_ASAP7_75t_L g145 ( 
.A(n_109),
.Y(n_145)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_145),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_76),
.B(n_5),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_146),
.B(n_14),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_73),
.A2(n_5),
.B1(n_8),
.B2(n_10),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_111),
.B(n_1),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_149),
.B(n_111),
.C(n_81),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_150),
.A2(n_184),
.B1(n_169),
.B2(n_158),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_152),
.B(n_158),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_123),
.B(n_89),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_156),
.B(n_165),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_162),
.B(n_176),
.Y(n_198)
);

NAND2x1p5_ASAP7_75t_L g163 ( 
.A(n_140),
.B(n_96),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_163),
.A2(n_128),
.B(n_141),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_126),
.B(n_140),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_140),
.B(n_73),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_166),
.B(n_169),
.Y(n_194)
);

AND2x2_ASAP7_75t_SL g167 ( 
.A(n_119),
.B(n_84),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_167),
.B(n_180),
.C(n_156),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_149),
.B(n_120),
.Y(n_169)
);

OAI21xp33_ASAP7_75t_SL g210 ( 
.A1(n_171),
.A2(n_183),
.B(n_157),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_125),
.A2(n_89),
.B1(n_85),
.B2(n_80),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_174),
.A2(n_178),
.B1(n_147),
.B2(n_131),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_112),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_116),
.A2(n_139),
.B1(n_80),
.B2(n_135),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_177),
.A2(n_137),
.B1(n_136),
.B2(n_121),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_149),
.A2(n_85),
.B1(n_108),
.B2(n_15),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_113),
.A2(n_105),
.B(n_108),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_180),
.A2(n_88),
.B(n_166),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_114),
.B(n_105),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_182),
.B(n_118),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_L g184 ( 
.A1(n_144),
.A2(n_88),
.B1(n_135),
.B2(n_116),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_176),
.B(n_148),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_186),
.B(n_188),
.Y(n_231)
);

OA21x2_ASAP7_75t_L g187 ( 
.A1(n_151),
.A2(n_139),
.B(n_143),
.Y(n_187)
);

A2O1A1Ixp33_ASAP7_75t_SL g225 ( 
.A1(n_187),
.A2(n_213),
.B(n_179),
.C(n_181),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_182),
.B(n_130),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_189),
.A2(n_197),
.B1(n_203),
.B2(n_210),
.Y(n_239)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_159),
.Y(n_190)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_190),
.Y(n_217)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_172),
.Y(n_192)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_192),
.Y(n_233)
);

BUFx12f_ASAP7_75t_L g193 ( 
.A(n_161),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_193),
.B(n_201),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_195),
.B(n_204),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_196),
.B(n_205),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_150),
.A2(n_145),
.B1(n_122),
.B2(n_124),
.Y(n_197)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_172),
.Y(n_199)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_199),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_200),
.A2(n_181),
.B1(n_168),
.B2(n_175),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_160),
.B(n_137),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_202),
.A2(n_173),
.B(n_179),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_157),
.A2(n_164),
.B(n_183),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_154),
.B(n_155),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_206),
.B(n_208),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_154),
.B(n_155),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_207),
.B(n_211),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_165),
.B(n_167),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_161),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_209),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_168),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_159),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_212),
.B(n_190),
.Y(n_229)
);

OA22x2_ASAP7_75t_L g213 ( 
.A1(n_174),
.A2(n_163),
.B1(n_157),
.B2(n_167),
.Y(n_213)
);

AND2x6_ASAP7_75t_L g214 ( 
.A(n_163),
.B(n_153),
.Y(n_214)
);

A2O1A1O1Ixp25_ASAP7_75t_L g227 ( 
.A1(n_214),
.A2(n_170),
.B(n_202),
.C(n_191),
.D(n_196),
.Y(n_227)
);

INVx13_ASAP7_75t_L g215 ( 
.A(n_179),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_215),
.B(n_216),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_173),
.B(n_152),
.C(n_175),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_220),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_222),
.A2(n_225),
.B(n_220),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_211),
.B(n_162),
.Y(n_224)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_224),
.Y(n_242)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_227),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_216),
.A2(n_170),
.B1(n_205),
.B2(n_194),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_228),
.B(n_234),
.Y(n_256)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_229),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_187),
.B(n_209),
.Y(n_230)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_230),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_206),
.B(n_185),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_185),
.B(n_194),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_235),
.B(n_240),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_187),
.B(n_198),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_237),
.B(n_241),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_208),
.B(n_203),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_192),
.Y(n_241)
);

OAI322xp33_ASAP7_75t_L g243 ( 
.A1(n_223),
.A2(n_214),
.A3(n_204),
.B1(n_213),
.B2(n_195),
.C1(n_189),
.C2(n_212),
.Y(n_243)
);

OAI322xp33_ASAP7_75t_L g277 ( 
.A1(n_243),
.A2(n_255),
.A3(n_225),
.B1(n_221),
.B2(n_236),
.C1(n_232),
.C2(n_241),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_228),
.B(n_213),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_246),
.B(n_247),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_219),
.B(n_231),
.Y(n_247)
);

OR2x2_ASAP7_75t_L g273 ( 
.A(n_248),
.B(n_225),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_223),
.B(n_213),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_250),
.B(n_253),
.Y(n_270)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_229),
.Y(n_252)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_252),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_218),
.B(n_199),
.C(n_197),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_218),
.B(n_193),
.C(n_215),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_254),
.B(n_261),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_SL g255 ( 
.A(n_240),
.B(n_193),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_239),
.A2(n_193),
.B1(n_225),
.B2(n_235),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_259),
.B(n_239),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_234),
.B(n_226),
.Y(n_260)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_260),
.Y(n_266)
);

CKINVDCx16_ASAP7_75t_R g261 ( 
.A(n_217),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_217),
.Y(n_262)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_262),
.Y(n_267)
);

A2O1A1Ixp33_ASAP7_75t_L g263 ( 
.A1(n_244),
.A2(n_226),
.B(n_222),
.C(n_227),
.Y(n_263)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_263),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_265),
.A2(n_253),
.B1(n_249),
.B2(n_252),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_242),
.B(n_231),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_268),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_245),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_271),
.B(n_276),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_273),
.A2(n_248),
.B(n_225),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_260),
.B(n_236),
.Y(n_274)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_274),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_257),
.B(n_251),
.Y(n_275)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_275),
.Y(n_284)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_262),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_277),
.B(n_271),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_270),
.B(n_250),
.C(n_246),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_279),
.B(n_287),
.C(n_288),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_281),
.B(n_265),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_264),
.A2(n_259),
.B1(n_249),
.B2(n_275),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_283),
.B(n_258),
.Y(n_300)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_286),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_272),
.B(n_254),
.C(n_255),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_269),
.B(n_256),
.C(n_251),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_273),
.A2(n_232),
.B(n_256),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_SL g298 ( 
.A1(n_289),
.A2(n_290),
.B(n_284),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_291),
.B(n_293),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_287),
.B(n_263),
.C(n_274),
.Y(n_293)
);

AOI31xp67_ASAP7_75t_SL g294 ( 
.A1(n_278),
.A2(n_268),
.A3(n_264),
.B(n_266),
.Y(n_294)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_294),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_SL g295 ( 
.A(n_282),
.B(n_266),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_295),
.A2(n_297),
.B(n_298),
.Y(n_303)
);

NOR2xp67_ASAP7_75t_SL g297 ( 
.A(n_285),
.B(n_273),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_279),
.B(n_267),
.C(n_276),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_299),
.B(n_288),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_300),
.B(n_283),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_301),
.B(n_305),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_293),
.A2(n_282),
.B(n_286),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_306),
.B(n_307),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_292),
.B(n_281),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_303),
.B(n_302),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_308),
.B(n_311),
.Y(n_315)
);

AOI21x1_ASAP7_75t_L g311 ( 
.A1(n_304),
.A2(n_296),
.B(n_289),
.Y(n_311)
);

NOR4xp25_ASAP7_75t_L g312 ( 
.A(n_307),
.B(n_292),
.C(n_258),
.D(n_280),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_312),
.B(n_301),
.C(n_267),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_313),
.B(n_314),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_309),
.B(n_233),
.C(n_238),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_315),
.A2(n_310),
.B1(n_233),
.B2(n_238),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_316),
.B(n_317),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_318),
.B(n_316),
.Y(n_319)
);


endmodule