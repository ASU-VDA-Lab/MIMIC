module fake_jpeg_16967_n_347 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_347);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_347;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_11),
.B(n_4),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_8),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_13),
.Y(n_24)
);

BUFx24_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx16f_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

HB1xp67_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_16),
.B(n_15),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_43),
.Y(n_51)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_35),
.Y(n_38)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_41),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_16),
.B(n_18),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_44),
.B(n_32),
.Y(n_55)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_23),
.Y(n_47)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_23),
.Y(n_49)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_L g50 ( 
.A1(n_44),
.A2(n_31),
.B(n_19),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_50),
.A2(n_53),
.B(n_25),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g53 ( 
.A1(n_37),
.A2(n_31),
.B(n_19),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_55),
.B(n_59),
.Y(n_112)
);

BUFx2_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_58),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_39),
.B(n_23),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_39),
.A2(n_20),
.B1(n_29),
.B2(n_22),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_60),
.A2(n_62),
.B1(n_75),
.B2(n_26),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_40),
.A2(n_20),
.B1(n_29),
.B2(n_22),
.Y(n_62)
);

OR2x2_ASAP7_75t_L g63 ( 
.A(n_40),
.B(n_19),
.Y(n_63)
);

A2O1A1Ixp33_ASAP7_75t_L g113 ( 
.A1(n_63),
.A2(n_48),
.B(n_42),
.C(n_46),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_45),
.B(n_32),
.Y(n_65)
);

OR2x2_ASAP7_75t_L g96 ( 
.A(n_65),
.B(n_73),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_45),
.A2(n_20),
.B1(n_22),
.B2(n_31),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_66),
.A2(n_70),
.B1(n_72),
.B2(n_25),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_42),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_69),
.B(n_43),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_49),
.A2(n_31),
.B1(n_33),
.B2(n_18),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_49),
.A2(n_31),
.B1(n_32),
.B2(n_33),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_43),
.B(n_26),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_38),
.A2(n_26),
.B1(n_33),
.B2(n_18),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_L g76 ( 
.A(n_50),
.B(n_36),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_76),
.B(n_100),
.C(n_112),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_71),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g114 ( 
.A(n_77),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_79),
.A2(n_98),
.B(n_51),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_80),
.Y(n_118)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_57),
.Y(n_81)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_81),
.Y(n_125)
);

OAI22xp33_ASAP7_75t_L g82 ( 
.A1(n_59),
.A2(n_41),
.B1(n_48),
.B2(n_42),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_82),
.A2(n_90),
.B1(n_100),
.B2(n_103),
.Y(n_123)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_74),
.Y(n_83)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_83),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_50),
.B(n_46),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_84),
.B(n_89),
.Y(n_126)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_61),
.Y(n_85)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_85),
.Y(n_134)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_71),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_86),
.A2(n_88),
.B1(n_97),
.B2(n_108),
.Y(n_129)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_61),
.Y(n_87)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_87),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_57),
.A2(n_21),
.B1(n_30),
.B2(n_24),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_63),
.B(n_46),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_53),
.A2(n_38),
.B1(n_21),
.B2(n_24),
.Y(n_90)
);

O2A1O1Ixp33_ASAP7_75t_L g91 ( 
.A1(n_75),
.A2(n_30),
.B(n_27),
.C(n_28),
.Y(n_91)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_91),
.Y(n_139)
);

BUFx2_ASAP7_75t_L g92 ( 
.A(n_52),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_92),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_63),
.B(n_46),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_93),
.B(n_113),
.Y(n_140)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_71),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_94),
.B(n_95),
.Y(n_127)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_56),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_57),
.A2(n_28),
.B1(n_27),
.B2(n_14),
.Y(n_97)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_99),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_53),
.A2(n_36),
.B1(n_34),
.B2(n_25),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_74),
.A2(n_15),
.B1(n_14),
.B2(n_2),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_101),
.A2(n_106),
.B1(n_55),
.B2(n_1),
.Y(n_120)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_52),
.Y(n_102)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_102),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_65),
.A2(n_34),
.B1(n_35),
.B2(n_25),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_60),
.A2(n_34),
.B1(n_25),
.B2(n_15),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_104),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_51),
.B(n_48),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_105),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_74),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_68),
.Y(n_107)
);

INVx1_ASAP7_75t_SL g122 ( 
.A(n_107),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_62),
.A2(n_69),
.B1(n_56),
.B2(n_67),
.Y(n_108)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_58),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_109),
.Y(n_133)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_68),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_110),
.Y(n_143)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_70),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_111),
.B(n_70),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_115),
.B(n_119),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_111),
.A2(n_64),
.B1(n_67),
.B2(n_73),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_116),
.A2(n_121),
.B1(n_128),
.B2(n_86),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_117),
.A2(n_89),
.B1(n_104),
.B2(n_101),
.Y(n_151)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_76),
.B(n_64),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_120),
.A2(n_124),
.B1(n_3),
.B2(n_5),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_84),
.A2(n_66),
.B1(n_72),
.B2(n_58),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_98),
.A2(n_3),
.B(n_4),
.Y(n_128)
);

A2O1A1Ixp33_ASAP7_75t_L g131 ( 
.A1(n_96),
.A2(n_3),
.B(n_4),
.C(n_5),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_131),
.B(n_91),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_SL g148 ( 
.A(n_137),
.B(n_117),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_112),
.B(n_41),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_138),
.B(n_106),
.Y(n_157)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_130),
.Y(n_144)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_144),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_118),
.B(n_96),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_145),
.B(n_149),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_118),
.B(n_81),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_146),
.B(n_172),
.Y(n_182)
);

OR2x2_ASAP7_75t_SL g147 ( 
.A(n_138),
.B(n_93),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_147),
.A2(n_174),
.B(n_176),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_148),
.B(n_161),
.C(n_171),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_132),
.B(n_95),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_130),
.Y(n_150)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_150),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_151),
.B(n_122),
.Y(n_188)
);

BUFx2_ASAP7_75t_L g152 ( 
.A(n_114),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_152),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_116),
.B(n_83),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_153),
.B(n_162),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_154),
.A2(n_128),
.B(n_139),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_141),
.A2(n_99),
.B1(n_82),
.B2(n_113),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_155),
.A2(n_166),
.B1(n_122),
.B2(n_136),
.Y(n_190)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_127),
.Y(n_156)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_156),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_157),
.B(n_163),
.Y(n_210)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_127),
.Y(n_158)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_158),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_159),
.A2(n_175),
.B1(n_129),
.B2(n_125),
.Y(n_180)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_142),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_160),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_126),
.B(n_78),
.C(n_54),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_126),
.B(n_87),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_142),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_134),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_164),
.B(n_165),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_119),
.B(n_85),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_141),
.A2(n_78),
.B1(n_109),
.B2(n_110),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_134),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_167),
.B(n_169),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_168),
.A2(n_136),
.B1(n_143),
.B2(n_7),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_140),
.B(n_92),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_119),
.B(n_107),
.Y(n_170)
);

OR2x2_ASAP7_75t_L g205 ( 
.A(n_170),
.B(n_6),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_137),
.B(n_54),
.C(n_77),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_125),
.B(n_92),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_135),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_139),
.A2(n_94),
.B1(n_102),
.B2(n_7),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_135),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_114),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_177),
.A2(n_143),
.B(n_54),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_178),
.B(n_183),
.Y(n_217)
);

NOR3xp33_ASAP7_75t_L g179 ( 
.A(n_154),
.B(n_140),
.C(n_120),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_179),
.B(n_192),
.Y(n_214)
);

OAI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_180),
.A2(n_202),
.B1(n_174),
.B2(n_150),
.Y(n_224)
);

A2O1A1O1Ixp25_ASAP7_75t_L g183 ( 
.A1(n_148),
.A2(n_123),
.B(n_121),
.C(n_131),
.D(n_115),
.Y(n_183)
);

NOR3xp33_ASAP7_75t_SL g184 ( 
.A(n_170),
.B(n_131),
.C(n_124),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_184),
.B(n_185),
.Y(n_225)
);

AOI31xp33_ASAP7_75t_L g185 ( 
.A1(n_151),
.A2(n_123),
.A3(n_133),
.B(n_122),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_188),
.B(n_163),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_190),
.A2(n_155),
.B1(n_158),
.B2(n_156),
.Y(n_223)
);

INVx1_ASAP7_75t_SL g192 ( 
.A(n_152),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_194),
.A2(n_175),
.B1(n_159),
.B2(n_169),
.Y(n_216)
);

INVx8_ASAP7_75t_L g197 ( 
.A(n_152),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_197),
.B(n_198),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_149),
.Y(n_198)
);

XOR2x1_ASAP7_75t_SL g199 ( 
.A(n_147),
.B(n_5),
.Y(n_199)
);

OAI32xp33_ASAP7_75t_L g218 ( 
.A1(n_199),
.A2(n_145),
.A3(n_153),
.B1(n_157),
.B2(n_165),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_166),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_203),
.A2(n_206),
.B(n_211),
.Y(n_226)
);

AND2x6_ASAP7_75t_L g204 ( 
.A(n_173),
.B(n_5),
.Y(n_204)
);

BUFx3_ASAP7_75t_L g219 ( 
.A(n_204),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_205),
.B(n_6),
.Y(n_227)
);

A2O1A1Ixp33_ASAP7_75t_SL g206 ( 
.A1(n_168),
.A2(n_114),
.B(n_7),
.C(n_8),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_177),
.Y(n_207)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_207),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_173),
.A2(n_6),
.B(n_8),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_181),
.Y(n_212)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_212),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_203),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_213),
.B(n_221),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_195),
.B(n_171),
.C(n_161),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_215),
.B(n_220),
.C(n_230),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g252 ( 
.A(n_216),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_218),
.A2(n_199),
.B(n_205),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_195),
.B(n_162),
.C(n_173),
.Y(n_220)
);

CKINVDCx14_ASAP7_75t_R g221 ( 
.A(n_209),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_223),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_224),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_227),
.B(n_209),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_207),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g257 ( 
.A(n_228),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_202),
.A2(n_144),
.B1(n_176),
.B2(n_160),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_229),
.A2(n_236),
.B1(n_184),
.B2(n_198),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_188),
.B(n_167),
.C(n_164),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_231),
.B(n_240),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_181),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_232),
.B(n_233),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_187),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_210),
.B(n_6),
.Y(n_234)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_234),
.Y(n_249)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_187),
.Y(n_235)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_235),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_183),
.A2(n_9),
.B1(n_10),
.B2(n_12),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_189),
.Y(n_237)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_237),
.Y(n_256)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_201),
.Y(n_238)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_238),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_200),
.B(n_114),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_242),
.A2(n_253),
.B1(n_263),
.B2(n_236),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_232),
.B(n_191),
.Y(n_245)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_245),
.Y(n_266)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_246),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_248),
.B(n_262),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_L g253 ( 
.A1(n_226),
.A2(n_178),
.B(n_191),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_233),
.B(n_208),
.Y(n_254)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_254),
.Y(n_276)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_212),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_260),
.B(n_261),
.Y(n_278)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_235),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_239),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_L g263 ( 
.A1(n_226),
.A2(n_193),
.B(n_211),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_234),
.B(n_189),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_264),
.B(n_265),
.Y(n_279)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_222),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_244),
.B(n_231),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_267),
.B(n_271),
.C(n_274),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_SL g288 ( 
.A(n_268),
.B(n_246),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_252),
.A2(n_223),
.B1(n_213),
.B2(n_214),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_269),
.A2(n_281),
.B1(n_263),
.B2(n_206),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_259),
.B(n_215),
.C(n_220),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_241),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_272),
.B(n_275),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_259),
.B(n_230),
.Y(n_274)
);

INVx1_ASAP7_75t_SL g275 ( 
.A(n_241),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_244),
.B(n_217),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_277),
.B(n_280),
.C(n_282),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_244),
.B(n_217),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_252),
.A2(n_194),
.B1(n_219),
.B2(n_229),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_259),
.B(n_240),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_253),
.B(n_245),
.C(n_255),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_283),
.B(n_285),
.C(n_219),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_254),
.B(n_208),
.Y(n_284)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_284),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_255),
.B(n_200),
.C(n_238),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_248),
.B(n_258),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_286),
.B(n_264),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_L g287 ( 
.A1(n_273),
.A2(n_251),
.B(n_243),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_SL g312 ( 
.A(n_287),
.B(n_288),
.Y(n_312)
);

INVxp67_ASAP7_75t_SL g304 ( 
.A(n_289),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_291),
.B(n_302),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_275),
.A2(n_265),
.B1(n_258),
.B2(n_256),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_292),
.A2(n_279),
.B1(n_278),
.B2(n_270),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_L g293 ( 
.A1(n_283),
.A2(n_242),
.B(n_225),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_293),
.B(n_297),
.C(n_303),
.Y(n_305)
);

HB1xp67_ASAP7_75t_L g296 ( 
.A(n_285),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_296),
.B(n_269),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_274),
.B(n_218),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_276),
.A2(n_256),
.B1(n_261),
.B2(n_260),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_299),
.A2(n_300),
.B1(n_301),
.B2(n_196),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_L g300 ( 
.A1(n_266),
.A2(n_247),
.B1(n_250),
.B2(n_249),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_284),
.A2(n_247),
.B1(n_250),
.B2(n_249),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_278),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_290),
.B(n_297),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_306),
.B(n_309),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_308),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_303),
.A2(n_279),
.B1(n_281),
.B2(n_268),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_310),
.B(n_311),
.Y(n_320)
);

HB1xp67_ASAP7_75t_L g313 ( 
.A(n_298),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_313),
.B(n_314),
.Y(n_327)
);

NOR3xp33_ASAP7_75t_SL g314 ( 
.A(n_293),
.B(n_204),
.C(n_206),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_290),
.B(n_271),
.C(n_282),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_315),
.B(n_295),
.C(n_267),
.Y(n_318)
);

BUFx24_ASAP7_75t_SL g316 ( 
.A(n_292),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_316),
.A2(n_182),
.B(n_206),
.Y(n_325)
);

OR2x2_ASAP7_75t_L g317 ( 
.A(n_294),
.B(n_196),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_317),
.A2(n_206),
.B(n_227),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_318),
.B(n_319),
.C(n_277),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_305),
.B(n_295),
.C(n_288),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_SL g321 ( 
.A1(n_307),
.A2(n_257),
.B(n_186),
.Y(n_321)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_321),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_304),
.A2(n_287),
.B1(n_289),
.B2(n_257),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_322),
.B(n_325),
.Y(n_336)
);

AND2x2_ASAP7_75t_L g324 ( 
.A(n_312),
.B(n_280),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_324),
.B(n_314),
.Y(n_330)
);

AOI221xp5_ASAP7_75t_L g333 ( 
.A1(n_328),
.A2(n_216),
.B1(n_190),
.B2(n_192),
.C(n_186),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_329),
.B(n_332),
.C(n_319),
.Y(n_337)
);

AO21x1_ASAP7_75t_L g340 ( 
.A1(n_330),
.A2(n_334),
.B(n_324),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_320),
.A2(n_304),
.B1(n_312),
.B2(n_317),
.Y(n_332)
);

AO21x2_ASAP7_75t_L g339 ( 
.A1(n_333),
.A2(n_335),
.B(n_328),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_323),
.B(n_239),
.Y(n_334)
);

NOR3xp33_ASAP7_75t_SL g335 ( 
.A(n_327),
.B(n_262),
.C(n_197),
.Y(n_335)
);

INVxp67_ASAP7_75t_L g343 ( 
.A(n_337),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_331),
.B(n_326),
.C(n_318),
.Y(n_338)
);

AOI21xp5_ASAP7_75t_L g342 ( 
.A1(n_338),
.A2(n_339),
.B(n_340),
.Y(n_342)
);

AOI31xp67_ASAP7_75t_L g341 ( 
.A1(n_335),
.A2(n_322),
.A3(n_10),
.B(n_12),
.Y(n_341)
);

OAI21xp5_ASAP7_75t_L g344 ( 
.A1(n_343),
.A2(n_341),
.B(n_336),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_344),
.B(n_342),
.C(n_333),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_345),
.B(n_9),
.C(n_10),
.Y(n_346)
);

AOI21xp5_ASAP7_75t_L g347 ( 
.A1(n_346),
.A2(n_9),
.B(n_10),
.Y(n_347)
);


endmodule