module fake_jpeg_23523_n_73 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_73);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_73;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_10;
wire n_23;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_59;
wire n_20;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_71;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_72;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_11;
wire n_62;
wire n_17;
wire n_25;
wire n_56;
wire n_31;
wire n_67;
wire n_37;
wire n_43;
wire n_29;
wire n_50;
wire n_12;
wire n_32;
wire n_70;
wire n_15;
wire n_66;

INVx6_ASAP7_75t_L g10 ( 
.A(n_9),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_3),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_SL g12 ( 
.A(n_0),
.B(n_9),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_7),
.Y(n_14)
);

CKINVDCx16_ASAP7_75t_R g15 ( 
.A(n_5),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx16f_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

HB1xp67_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx4f_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_18),
.Y(n_22)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

AOI21xp33_ASAP7_75t_L g23 ( 
.A1(n_14),
.A2(n_1),
.B(n_2),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_23),
.A2(n_28),
.B1(n_24),
.B2(n_17),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_14),
.B(n_1),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_24),
.B(n_28),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_19),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_25),
.B(n_15),
.Y(n_39)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_26),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_27),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_19),
.B(n_3),
.Y(n_28)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_32),
.B(n_4),
.Y(n_42)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_35),
.Y(n_45)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_26),
.A2(n_13),
.B1(n_17),
.B2(n_12),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_36),
.A2(n_37),
.B1(n_11),
.B2(n_16),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_26),
.A2(n_13),
.B1(n_12),
.B2(n_11),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_38),
.B(n_41),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_39),
.B(n_6),
.Y(n_49)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_42),
.B(n_48),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_43),
.B(n_47),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_33),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_44),
.Y(n_56)
);

AOI21xp5_ASAP7_75t_L g46 ( 
.A1(n_33),
.A2(n_27),
.B(n_22),
.Y(n_46)
);

XOR2xp5_ASAP7_75t_L g55 ( 
.A(n_46),
.B(n_27),
.Y(n_55)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_49),
.Y(n_52)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

BUFx2_ASAP7_75t_L g58 ( 
.A(n_50),
.Y(n_58)
);

XOR2xp5_ASAP7_75t_L g63 ( 
.A(n_55),
.B(n_42),
.Y(n_63)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_57),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_55),
.B(n_51),
.C(n_48),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_59),
.B(n_60),
.C(n_63),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_54),
.B(n_32),
.C(n_46),
.Y(n_60)
);

NAND3xp33_ASAP7_75t_L g62 ( 
.A(n_52),
.B(n_42),
.C(n_40),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_62),
.A2(n_53),
.B1(n_57),
.B2(n_30),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_62),
.A2(n_43),
.B1(n_56),
.B2(n_30),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_64),
.B(n_61),
.C(n_31),
.Y(n_67)
);

XNOR2xp5_ASAP7_75t_L g68 ( 
.A(n_65),
.B(n_20),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_67),
.B(n_66),
.C(n_58),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_68),
.B(n_20),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_69),
.B(n_70),
.C(n_58),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_71),
.A2(n_20),
.B1(n_16),
.B2(n_7),
.Y(n_72)
);

XOR2xp5_ASAP7_75t_L g73 ( 
.A(n_72),
.B(n_6),
.Y(n_73)
);


endmodule