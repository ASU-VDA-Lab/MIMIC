module real_jpeg_16925_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_553;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_214;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_559;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_323;
wire n_215;
wire n_176;
wire n_166;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_548;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_546;
wire n_531;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_450;
wire n_333;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_534;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_568;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx2_ASAP7_75t_SL g21 ( 
.A(n_0),
.Y(n_21)
);

AND2x2_ASAP7_75t_L g22 ( 
.A(n_0),
.B(n_23),
.Y(n_22)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_1),
.B(n_64),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_1),
.B(n_80),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_1),
.B(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_1),
.B(n_144),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_1),
.B(n_158),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g250 ( 
.A(n_1),
.B(n_251),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_1),
.B(n_254),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_1),
.A2(n_7),
.B1(n_287),
.B2(n_291),
.Y(n_286)
);

CKINVDCx16_ASAP7_75t_R g404 ( 
.A(n_1),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_2),
.B(n_307),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_2),
.B(n_392),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_SL g418 ( 
.A(n_2),
.B(n_419),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_2),
.B(n_450),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_2),
.B(n_492),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g503 ( 
.A(n_2),
.B(n_504),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_SL g512 ( 
.A(n_2),
.B(n_513),
.Y(n_512)
);

BUFx3_ASAP7_75t_L g170 ( 
.A(n_3),
.Y(n_170)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_3),
.Y(n_290)
);

BUFx5_ASAP7_75t_L g389 ( 
.A(n_3),
.Y(n_389)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_4),
.Y(n_172)
);

NAND2x1_ASAP7_75t_L g175 ( 
.A(n_4),
.B(n_176),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g241 ( 
.A(n_4),
.B(n_242),
.Y(n_241)
);

AND2x2_ASAP7_75t_SL g256 ( 
.A(n_4),
.B(n_31),
.Y(n_256)
);

AND2x2_ASAP7_75t_L g302 ( 
.A(n_4),
.B(n_303),
.Y(n_302)
);

AND2x2_ASAP7_75t_L g360 ( 
.A(n_4),
.B(n_113),
.Y(n_360)
);

AND2x2_ASAP7_75t_L g384 ( 
.A(n_4),
.B(n_385),
.Y(n_384)
);

AND2x2_ASAP7_75t_L g468 ( 
.A(n_4),
.B(n_248),
.Y(n_468)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_5),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_5),
.Y(n_83)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_5),
.Y(n_110)
);

BUFx5_ASAP7_75t_L g394 ( 
.A(n_5),
.Y(n_394)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_6),
.A2(n_20),
.B(n_22),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_7),
.B(n_103),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_7),
.B(n_235),
.Y(n_234)
);

AND2x2_ASAP7_75t_L g357 ( 
.A(n_7),
.B(n_358),
.Y(n_357)
);

AND2x2_ASAP7_75t_L g397 ( 
.A(n_7),
.B(n_398),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_SL g421 ( 
.A(n_7),
.B(n_238),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_SL g453 ( 
.A(n_7),
.B(n_454),
.Y(n_453)
);

AND2x2_ASAP7_75t_L g460 ( 
.A(n_7),
.B(n_461),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_7),
.B(n_168),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_8),
.B(n_103),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_8),
.B(n_154),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_8),
.B(n_178),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_8),
.B(n_200),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_8),
.B(n_238),
.Y(n_237)
);

AND2x2_ASAP7_75t_L g308 ( 
.A(n_8),
.B(n_309),
.Y(n_308)
);

CKINVDCx16_ASAP7_75t_R g351 ( 
.A(n_8),
.Y(n_351)
);

AND2x2_ASAP7_75t_L g387 ( 
.A(n_8),
.B(n_388),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_9),
.B(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_9),
.B(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_9),
.B(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_9),
.B(n_99),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_9),
.B(n_148),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_9),
.B(n_144),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g218 ( 
.A(n_9),
.B(n_219),
.Y(n_218)
);

AND2x2_ASAP7_75t_L g247 ( 
.A(n_9),
.B(n_248),
.Y(n_247)
);

BUFx5_ASAP7_75t_L g113 ( 
.A(n_10),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_10),
.Y(n_149)
);

BUFx5_ASAP7_75t_L g254 ( 
.A(n_10),
.Y(n_254)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_10),
.Y(n_311)
);

BUFx6f_ASAP7_75t_L g457 ( 
.A(n_10),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_11),
.B(n_68),
.Y(n_67)
);

INVxp33_ASAP7_75t_L g107 ( 
.A(n_11),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_11),
.B(n_130),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_11),
.B(n_151),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_11),
.B(n_204),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_11),
.B(n_298),
.Y(n_297)
);

AND2x2_ASAP7_75t_L g313 ( 
.A(n_11),
.B(n_314),
.Y(n_313)
);

AND2x2_ASAP7_75t_SL g352 ( 
.A(n_11),
.B(n_353),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_12),
.B(n_208),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_12),
.B(n_210),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g295 ( 
.A(n_12),
.B(n_296),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_12),
.B(n_317),
.Y(n_316)
);

AND2x2_ASAP7_75t_L g361 ( 
.A(n_12),
.B(n_362),
.Y(n_361)
);

AND2x2_ASAP7_75t_L g462 ( 
.A(n_12),
.B(n_463),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_12),
.B(n_467),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_SL g481 ( 
.A(n_12),
.B(n_482),
.Y(n_481)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_13),
.Y(n_141)
);

BUFx4f_ASAP7_75t_L g220 ( 
.A(n_13),
.Y(n_220)
);

BUFx12f_ASAP7_75t_L g252 ( 
.A(n_13),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_14),
.B(n_31),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_14),
.B(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_SL g49 ( 
.A(n_14),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_14),
.B(n_72),
.Y(n_71)
);

AND2x4_ASAP7_75t_SL g167 ( 
.A(n_14),
.B(n_168),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_14),
.B(n_564),
.Y(n_563)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g160 ( 
.A(n_15),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_15),
.Y(n_202)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_16),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g146 ( 
.A(n_16),
.Y(n_146)
);

BUFx3_ASAP7_75t_L g206 ( 
.A(n_16),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_16),
.Y(n_239)
);

INVx3_ASAP7_75t_L g305 ( 
.A(n_16),
.Y(n_305)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_16),
.Y(n_495)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_17),
.Y(n_89)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_18),
.Y(n_57)
);

BUFx8_ASAP7_75t_L g65 ( 
.A(n_18),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

O2A1O1Ixp33_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_559),
.B(n_566),
.C(n_568),
.Y(n_23)
);

OAI21x1_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_121),
.B(n_558),
.Y(n_24)
);

CKINVDCx16_ASAP7_75t_R g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_75),
.Y(n_26)
);

OR2x2_ASAP7_75t_L g558 ( 
.A(n_27),
.B(n_75),
.Y(n_558)
);

XOR2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_58),
.Y(n_27)
);

XNOR2xp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_44),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g567 ( 
.A(n_29),
.B(n_44),
.C(n_58),
.Y(n_567)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_33),
.C(n_37),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_30),
.A2(n_46),
.B1(n_50),
.B2(n_51),
.Y(n_45)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_30),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_30),
.A2(n_33),
.B1(n_50),
.B2(n_62),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_SL g561 ( 
.A(n_30),
.B(n_46),
.C(n_52),
.Y(n_561)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_32),
.Y(n_96)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_32),
.Y(n_179)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_32),
.Y(n_293)
);

INVx1_ASAP7_75t_SL g62 ( 
.A(n_33),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_33),
.B(n_67),
.C(n_70),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_33),
.A2(n_62),
.B1(n_70),
.B2(n_71),
.Y(n_116)
);

BUFx2_ASAP7_75t_L g151 ( 
.A(n_34),
.Y(n_151)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_35),
.Y(n_101)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_35),
.Y(n_452)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

XOR2xp5_ASAP7_75t_L g60 ( 
.A(n_37),
.B(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

XNOR2xp5_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_52),
.Y(n_44)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_46),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g562 ( 
.A1(n_46),
.A2(n_51),
.B1(n_563),
.B2(n_566),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_47),
.B(n_49),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_48),
.Y(n_155)
);

OR2x2_ASAP7_75t_L g111 ( 
.A(n_49),
.B(n_112),
.Y(n_111)
);

OR2x2_ASAP7_75t_L g138 ( 
.A(n_49),
.B(n_139),
.Y(n_138)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_56),
.Y(n_69)
);

INVx8_ASAP7_75t_L g176 ( 
.A(n_56),
.Y(n_176)
);

INVx4_ASAP7_75t_L g565 ( 
.A(n_56),
.Y(n_565)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_57),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_63),
.C(n_66),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_59),
.A2(n_60),
.B1(n_119),
.B2(n_120),
.Y(n_118)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

XNOR2xp5_ASAP7_75t_SL g120 ( 
.A(n_63),
.B(n_66),
.Y(n_120)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_65),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_67),
.B(n_116),
.Y(n_115)
);

INVx3_ASAP7_75t_SL g68 ( 
.A(n_69),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_70),
.A2(n_71),
.B1(n_111),
.B2(n_136),
.Y(n_182)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_SL g105 ( 
.A(n_71),
.B(n_106),
.C(n_111),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_117),
.C(n_118),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_76),
.B(n_189),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_105),
.C(n_114),
.Y(n_76)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_77),
.B(n_187),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_90),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_84),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_79),
.B(n_84),
.C(n_90),
.Y(n_117)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

HB1xp67_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

OR2x2_ASAP7_75t_L g171 ( 
.A(n_82),
.B(n_172),
.Y(n_171)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_89),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g318 ( 
.A(n_89),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g402 ( 
.A(n_89),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_97),
.C(n_102),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_91),
.A2(n_92),
.B1(n_97),
.B2(n_98),
.Y(n_163)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

XNOR2x1_ASAP7_75t_L g162 ( 
.A(n_102),
.B(n_163),
.Y(n_162)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_105),
.B(n_115),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_SL g181 ( 
.A(n_106),
.B(n_182),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_108),
.Y(n_106)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_110),
.Y(n_208)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_110),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_111),
.A2(n_136),
.B1(n_137),
.B2(n_138),
.Y(n_135)
);

INVx1_ASAP7_75t_SL g136 ( 
.A(n_111),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_111),
.B(n_129),
.C(n_137),
.Y(n_183)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

HB1xp67_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_117),
.B(n_118),
.Y(n_189)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

AOI21x1_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_276),
.B(n_553),
.Y(n_121)
);

NOR3xp33_ASAP7_75t_SL g122 ( 
.A(n_123),
.B(n_190),
.C(n_270),
.Y(n_122)
);

OAI21x1_ASAP7_75t_SL g553 ( 
.A1(n_123),
.A2(n_554),
.B(n_557),
.Y(n_553)
);

NOR2x1_ASAP7_75t_R g123 ( 
.A(n_124),
.B(n_188),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_124),
.B(n_188),
.Y(n_557)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_180),
.C(n_185),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_125),
.B(n_273),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_162),
.C(n_164),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_127),
.B(n_267),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_142),
.C(n_152),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_128),
.B(n_227),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_135),
.Y(n_128)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_137),
.A2(n_138),
.B1(n_167),
.B2(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_SL g137 ( 
.A(n_138),
.Y(n_137)
);

MAJx2_ASAP7_75t_L g166 ( 
.A(n_138),
.B(n_167),
.C(n_171),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_140),
.Y(n_516)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g386 ( 
.A(n_141),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_142),
.B(n_152),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_147),
.C(n_150),
.Y(n_142)
);

XNOR2x1_ASAP7_75t_L g215 ( 
.A(n_143),
.B(n_150),
.Y(n_215)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

XNOR2x1_ASAP7_75t_L g214 ( 
.A(n_147),
.B(n_215),
.Y(n_214)
);

BUFx2_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx6_ASAP7_75t_L g483 ( 
.A(n_149),
.Y(n_483)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_156),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_153),
.B(n_157),
.C(n_161),
.Y(n_184)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_161),
.Y(n_156)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

BUFx3_ASAP7_75t_L g296 ( 
.A(n_160),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_162),
.B(n_164),
.Y(n_267)
);

MAJx2_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_173),
.C(n_177),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_165),
.A2(n_166),
.B1(n_195),
.B2(n_196),
.Y(n_194)
);

INVx1_ASAP7_75t_SL g165 ( 
.A(n_166),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_167),
.B(n_217),
.C(n_218),
.Y(n_216)
);

INVx1_ASAP7_75t_SL g225 ( 
.A(n_167),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_167),
.A2(n_218),
.B1(n_225),
.B2(n_232),
.Y(n_231)
);

INVx5_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_170),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_171),
.A2(n_222),
.B1(n_223),
.B2(n_224),
.Y(n_221)
);

INVx1_ASAP7_75t_SL g222 ( 
.A(n_171),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_171),
.A2(n_222),
.B1(n_297),
.B2(n_345),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_173),
.B(n_284),
.Y(n_283)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_SL g195 ( 
.A(n_175),
.B(n_177),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_175),
.B(n_247),
.C(n_250),
.Y(n_246)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_177),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_177),
.A2(n_209),
.B1(n_212),
.B2(n_259),
.Y(n_258)
);

INVx6_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_180),
.A2(n_185),
.B1(n_186),
.B2(n_274),
.Y(n_273)
);

INVxp67_ASAP7_75t_SL g274 ( 
.A(n_180),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_183),
.C(n_184),
.Y(n_180)
);

XNOR2x2_ASAP7_75t_L g264 ( 
.A(n_181),
.B(n_265),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_183),
.B(n_184),
.Y(n_265)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_260),
.Y(n_190)
);

NOR2x1_ASAP7_75t_L g555 ( 
.A(n_191),
.B(n_260),
.Y(n_555)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_226),
.C(n_228),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_192),
.B(n_226),
.Y(n_374)
);

XNOR2x1_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_213),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_197),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_194),
.B(n_197),
.C(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_195),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_209),
.C(n_212),
.Y(n_197)
);

XNOR2x1_ASAP7_75t_L g257 ( 
.A(n_198),
.B(n_258),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_203),
.C(n_207),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_199),
.B(n_207),
.Y(n_244)
);

HB1xp67_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx6_ASAP7_75t_L g359 ( 
.A(n_201),
.Y(n_359)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

BUFx5_ASAP7_75t_L g242 ( 
.A(n_202),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_203),
.B(n_244),
.Y(n_243)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_209),
.Y(n_259)
);

INVx6_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx4_ASAP7_75t_L g307 ( 
.A(n_211),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_213),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_216),
.C(n_221),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_214),
.B(n_216),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_217),
.B(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_218),
.Y(n_232)
);

BUFx2_ASAP7_75t_L g461 ( 
.A(n_219),
.Y(n_461)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_220),
.Y(n_350)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_221),
.B(n_325),
.Y(n_324)
);

MAJx2_ASAP7_75t_L g294 ( 
.A(n_222),
.B(n_295),
.C(n_297),
.Y(n_294)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g373 ( 
.A(n_228),
.B(n_374),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_245),
.C(n_257),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_SL g326 ( 
.A(n_229),
.B(n_327),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_233),
.C(n_243),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_230),
.B(n_233),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_237),
.C(n_240),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_234),
.A2(n_240),
.B1(n_241),
.B2(n_371),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_234),
.Y(n_371)
);

HB1xp67_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g369 ( 
.A(n_237),
.B(n_370),
.Y(n_369)
);

BUFx12f_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_240),
.B(n_418),
.C(n_421),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_L g475 ( 
.A1(n_240),
.A2(n_241),
.B1(n_418),
.B2(n_476),
.Y(n_475)
);

INVx2_ASAP7_75t_SL g240 ( 
.A(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_243),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_245),
.B(n_257),
.Y(n_327)
);

MAJx2_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_253),
.C(n_255),
.Y(n_245)
);

XNOR2x1_ASAP7_75t_SL g320 ( 
.A(n_246),
.B(n_321),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_247),
.B(n_250),
.Y(n_284)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx3_ASAP7_75t_L g299 ( 
.A(n_252),
.Y(n_299)
);

BUFx3_ASAP7_75t_L g467 ( 
.A(n_252),
.Y(n_467)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_253),
.A2(n_255),
.B1(n_256),
.B2(n_322),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_253),
.Y(n_322)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_254),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g535 ( 
.A1(n_255),
.A2(n_256),
.B1(n_390),
.B2(n_391),
.Y(n_535)
);

INVx2_ASAP7_75t_SL g255 ( 
.A(n_256),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_256),
.B(n_383),
.C(n_390),
.Y(n_382)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_263),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_261),
.B(n_264),
.C(n_268),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_264),
.A2(n_266),
.B1(n_268),
.B2(n_269),
.Y(n_263)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_264),
.Y(n_269)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_266),
.Y(n_268)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

AOI21x1_ASAP7_75t_L g554 ( 
.A1(n_271),
.A2(n_555),
.B(n_556),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_275),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g556 ( 
.A(n_272),
.B(n_275),
.Y(n_556)
);

AO21x2_ASAP7_75t_L g276 ( 
.A1(n_277),
.A2(n_377),
.B(n_550),
.Y(n_276)
);

NOR2xp67_ASAP7_75t_SL g277 ( 
.A(n_278),
.B(n_372),
.Y(n_277)
);

AND2x2_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_330),
.Y(n_278)
);

OR2x2_ASAP7_75t_L g551 ( 
.A(n_279),
.B(n_330),
.Y(n_551)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_323),
.Y(n_279)
);

INVxp67_ASAP7_75t_SL g376 ( 
.A(n_280),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_300),
.C(n_319),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_282),
.B(n_334),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_285),
.C(n_294),
.Y(n_282)
);

XNOR2x2_ASAP7_75t_L g429 ( 
.A(n_283),
.B(n_430),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_SL g430 ( 
.A1(n_285),
.A2(n_286),
.B1(n_294),
.B2(n_431),
.Y(n_430)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g396 ( 
.A1(n_286),
.A2(n_397),
.B(n_403),
.Y(n_396)
);

INVx6_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx6_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx3_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_290),
.Y(n_355)
);

BUFx3_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx2_ASAP7_75t_SL g292 ( 
.A(n_293),
.Y(n_292)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_294),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_295),
.B(n_344),
.Y(n_343)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_297),
.Y(n_345)
);

INVx4_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_300),
.A2(n_319),
.B1(n_320),
.B2(n_335),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_300),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_312),
.C(n_316),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_306),
.C(n_308),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_302),
.B(n_306),
.C(n_308),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g409 ( 
.A(n_302),
.B(n_308),
.Y(n_409)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_302),
.Y(n_447)
);

HB1xp67_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_305),
.Y(n_364)
);

XOR2xp5_ASAP7_75t_L g408 ( 
.A(n_306),
.B(n_409),
.Y(n_408)
);

INVx8_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

BUFx6f_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_311),
.Y(n_508)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_312),
.A2(n_313),
.B1(n_316),
.B2(n_367),
.Y(n_366)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_316),
.Y(n_367)
);

BUFx6f_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx4_ASAP7_75t_L g420 ( 
.A(n_318),
.Y(n_420)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_324),
.A2(n_326),
.B1(n_328),
.B2(n_329),
.Y(n_323)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_324),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_324),
.B(n_329),
.C(n_376),
.Y(n_375)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_326),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_331),
.B(n_336),
.C(n_339),
.Y(n_330)
);

HB1xp67_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_SL g437 ( 
.A1(n_332),
.A2(n_333),
.B1(n_336),
.B2(n_438),
.Y(n_437)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_336),
.Y(n_438)
);

XOR2x2_ASAP7_75t_L g336 ( 
.A(n_337),
.B(n_338),
.Y(n_336)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g436 ( 
.A(n_340),
.B(n_437),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_341),
.B(n_365),
.C(n_369),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_SL g432 ( 
.A(n_341),
.B(n_433),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_342),
.B(n_346),
.C(n_356),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

XNOR2x1_ASAP7_75t_L g424 ( 
.A(n_343),
.B(n_425),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_346),
.B(n_356),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_347),
.B(n_352),
.Y(n_346)
);

XOR2xp5_ASAP7_75t_L g423 ( 
.A(n_347),
.B(n_352),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_348),
.B(n_351),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

BUFx6f_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_354),
.Y(n_464)
);

BUFx6f_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_357),
.B(n_360),
.C(n_361),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_SL g413 ( 
.A1(n_357),
.A2(n_360),
.B1(n_414),
.B2(n_415),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_357),
.Y(n_414)
);

INVx8_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_360),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_SL g489 ( 
.A1(n_360),
.A2(n_415),
.B1(n_490),
.B2(n_491),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_360),
.B(n_490),
.C(n_496),
.Y(n_523)
);

XOR2xp5_ASAP7_75t_L g412 ( 
.A(n_361),
.B(n_413),
.Y(n_412)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

INVx5_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g433 ( 
.A(n_365),
.B(n_369),
.Y(n_433)
);

XOR2xp5_ASAP7_75t_L g365 ( 
.A(n_366),
.B(n_368),
.Y(n_365)
);

OAI21xp5_ASAP7_75t_L g550 ( 
.A1(n_372),
.A2(n_551),
.B(n_552),
.Y(n_550)
);

AND2x2_ASAP7_75t_L g372 ( 
.A(n_373),
.B(n_375),
.Y(n_372)
);

OR2x2_ASAP7_75t_L g552 ( 
.A(n_373),
.B(n_375),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_378),
.B(n_546),
.Y(n_377)
);

NAND3xp33_ASAP7_75t_SL g378 ( 
.A(n_379),
.B(n_434),
.C(n_439),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_380),
.B(n_426),
.Y(n_379)
);

NOR2xp67_ASAP7_75t_SL g549 ( 
.A(n_380),
.B(n_426),
.Y(n_549)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_381),
.B(n_410),
.C(n_424),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g543 ( 
.A(n_381),
.B(n_544),
.Y(n_543)
);

XOR2xp5_ASAP7_75t_L g381 ( 
.A(n_382),
.B(n_395),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_382),
.B(n_396),
.C(n_408),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_SL g534 ( 
.A(n_383),
.B(n_535),
.Y(n_534)
);

AND2x2_ASAP7_75t_L g383 ( 
.A(n_384),
.B(n_387),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_L g480 ( 
.A(n_384),
.B(n_387),
.Y(n_480)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_384),
.Y(n_499)
);

AOI22xp5_ASAP7_75t_L g509 ( 
.A1(n_384),
.A2(n_499),
.B1(n_500),
.B2(n_510),
.Y(n_509)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

BUFx3_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

INVx3_ASAP7_75t_L g407 ( 
.A(n_389),
.Y(n_407)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

INVx3_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g395 ( 
.A(n_396),
.B(n_408),
.Y(n_395)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

INVx3_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_404),
.B(n_405),
.Y(n_403)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

HB1xp67_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_L g544 ( 
.A(n_411),
.B(n_424),
.Y(n_544)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_412),
.B(n_416),
.C(n_422),
.Y(n_411)
);

XOR2xp5_ASAP7_75t_L g529 ( 
.A(n_412),
.B(n_530),
.Y(n_529)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_L g530 ( 
.A(n_417),
.B(n_423),
.Y(n_530)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_418),
.Y(n_476)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

XOR2xp5_ASAP7_75t_L g474 ( 
.A(n_421),
.B(n_475),
.Y(n_474)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

XOR2xp5_ASAP7_75t_L g426 ( 
.A(n_427),
.B(n_432),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_428),
.B(n_429),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_428),
.B(n_429),
.C(n_432),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_435),
.B(n_436),
.Y(n_434)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_435),
.Y(n_548)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_436),
.Y(n_547)
);

OAI21xp5_ASAP7_75t_SL g439 ( 
.A1(n_440),
.A2(n_541),
.B(n_545),
.Y(n_439)
);

AOI21xp5_ASAP7_75t_L g440 ( 
.A1(n_441),
.A2(n_526),
.B(n_540),
.Y(n_440)
);

OAI21xp5_ASAP7_75t_SL g441 ( 
.A1(n_442),
.A2(n_484),
.B(n_525),
.Y(n_441)
);

AND2x2_ASAP7_75t_L g442 ( 
.A(n_443),
.B(n_471),
.Y(n_442)
);

OR2x2_ASAP7_75t_L g525 ( 
.A(n_443),
.B(n_471),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_444),
.B(n_458),
.C(n_465),
.Y(n_443)
);

HB1xp67_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);

XOR2xp5_ASAP7_75t_L g520 ( 
.A(n_445),
.B(n_521),
.Y(n_520)
);

XNOR2xp5_ASAP7_75t_L g445 ( 
.A(n_446),
.B(n_448),
.Y(n_445)
);

INVx1_ASAP7_75t_SL g446 ( 
.A(n_447),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_447),
.B(n_449),
.C(n_453),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_449),
.B(n_453),
.Y(n_448)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_451),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_452),
.Y(n_451)
);

HB1xp67_ASAP7_75t_L g454 ( 
.A(n_455),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_456),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_457),
.Y(n_456)
);

AOI22xp5_ASAP7_75t_L g521 ( 
.A1(n_458),
.A2(n_459),
.B1(n_465),
.B2(n_522),
.Y(n_521)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_459),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_460),
.B(n_462),
.Y(n_459)
);

XNOR2xp5_ASAP7_75t_SL g497 ( 
.A(n_460),
.B(n_462),
.Y(n_497)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_464),
.Y(n_463)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_465),
.Y(n_522)
);

AO22x1_ASAP7_75t_SL g465 ( 
.A1(n_466),
.A2(n_468),
.B1(n_469),
.B2(n_470),
.Y(n_465)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_466),
.Y(n_469)
);

INVx1_ASAP7_75t_SL g470 ( 
.A(n_468),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_468),
.B(n_469),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_470),
.B(n_512),
.Y(n_511)
);

XOR2xp5_ASAP7_75t_L g471 ( 
.A(n_472),
.B(n_477),
.Y(n_471)
);

XNOR2xp5_ASAP7_75t_L g472 ( 
.A(n_473),
.B(n_474),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g538 ( 
.A(n_473),
.B(n_477),
.C(n_539),
.Y(n_538)
);

HB1xp67_ASAP7_75t_L g539 ( 
.A(n_474),
.Y(n_539)
);

XOR2xp5_ASAP7_75t_L g477 ( 
.A(n_478),
.B(n_479),
.Y(n_477)
);

MAJx2_ASAP7_75t_L g537 ( 
.A(n_478),
.B(n_480),
.C(n_481),
.Y(n_537)
);

XNOR2xp5_ASAP7_75t_L g479 ( 
.A(n_480),
.B(n_481),
.Y(n_479)
);

INVx4_ASAP7_75t_L g482 ( 
.A(n_483),
.Y(n_482)
);

AOI21xp5_ASAP7_75t_L g484 ( 
.A1(n_485),
.A2(n_519),
.B(n_524),
.Y(n_484)
);

OAI21xp5_ASAP7_75t_SL g485 ( 
.A1(n_486),
.A2(n_501),
.B(n_518),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_487),
.B(n_498),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_487),
.B(n_498),
.Y(n_518)
);

OAI22xp5_ASAP7_75t_SL g487 ( 
.A1(n_488),
.A2(n_489),
.B1(n_496),
.B2(n_497),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_489),
.Y(n_488)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_491),
.Y(n_490)
);

INVx3_ASAP7_75t_L g492 ( 
.A(n_493),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_494),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_495),
.Y(n_494)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_497),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_SL g498 ( 
.A(n_499),
.B(n_500),
.Y(n_498)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_500),
.Y(n_510)
);

AOI21x1_ASAP7_75t_SL g501 ( 
.A1(n_502),
.A2(n_511),
.B(n_517),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_503),
.B(n_509),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_503),
.B(n_509),
.Y(n_517)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_505),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_506),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_507),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_508),
.Y(n_507)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_514),
.Y(n_513)
);

HB1xp67_ASAP7_75t_L g514 ( 
.A(n_515),
.Y(n_514)
);

INVx3_ASAP7_75t_L g515 ( 
.A(n_516),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_SL g519 ( 
.A(n_520),
.B(n_523),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_520),
.B(n_523),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_SL g526 ( 
.A(n_527),
.B(n_538),
.Y(n_526)
);

NOR2xp67_ASAP7_75t_L g540 ( 
.A(n_527),
.B(n_538),
.Y(n_540)
);

AOI22xp5_ASAP7_75t_L g527 ( 
.A1(n_528),
.A2(n_529),
.B1(n_531),
.B2(n_532),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g542 ( 
.A(n_528),
.B(n_533),
.C(n_537),
.Y(n_542)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_529),
.Y(n_528)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_532),
.Y(n_531)
);

AOI22xp5_ASAP7_75t_L g532 ( 
.A1(n_533),
.A2(n_534),
.B1(n_536),
.B2(n_537),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_534),
.Y(n_533)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_537),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_542),
.B(n_543),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_542),
.B(n_543),
.Y(n_545)
);

MAJIxp5_ASAP7_75t_L g546 ( 
.A(n_547),
.B(n_548),
.C(n_549),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_L g559 ( 
.A(n_560),
.B(n_567),
.Y(n_559)
);

AND2x2_ASAP7_75t_L g569 ( 
.A(n_560),
.B(n_567),
.Y(n_569)
);

XNOR2xp5_ASAP7_75t_L g560 ( 
.A(n_561),
.B(n_562),
.Y(n_560)
);

CKINVDCx16_ASAP7_75t_R g566 ( 
.A(n_563),
.Y(n_566)
);

BUFx6f_ASAP7_75t_L g564 ( 
.A(n_565),
.Y(n_564)
);

CKINVDCx20_ASAP7_75t_R g568 ( 
.A(n_569),
.Y(n_568)
);


endmodule