module fake_netlist_1_8692_n_23 (n_1, n_2, n_6, n_4, n_3, n_5, n_0, n_23);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_5;
input n_0;
output n_23;
wire n_20;
wire n_8;
wire n_22;
wire n_11;
wire n_16;
wire n_13;
wire n_18;
wire n_12;
wire n_9;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_19;
wire n_21;
wire n_7;
INVx2_ASAP7_75t_L g7 ( .A(n_3), .Y(n_7) );
CKINVDCx20_ASAP7_75t_R g8 ( .A(n_4), .Y(n_8) );
INVx2_ASAP7_75t_L g9 ( .A(n_4), .Y(n_9) );
INVx1_ASAP7_75t_L g10 ( .A(n_3), .Y(n_10) );
INVx1_ASAP7_75t_L g11 ( .A(n_5), .Y(n_11) );
OAI21x1_ASAP7_75t_L g12 ( .A1(n_11), .A2(n_6), .B(n_1), .Y(n_12) );
NOR2xp33_ASAP7_75t_L g13 ( .A(n_11), .B(n_0), .Y(n_13) );
AND2x4_ASAP7_75t_L g14 ( .A(n_13), .B(n_7), .Y(n_14) );
AND2x2_ASAP7_75t_L g15 ( .A(n_14), .B(n_10), .Y(n_15) );
INVxp67_ASAP7_75t_SL g16 ( .A(n_15), .Y(n_16) );
INVx2_ASAP7_75t_L g17 ( .A(n_15), .Y(n_17) );
AOI221xp5_ASAP7_75t_L g18 ( .A1(n_16), .A2(n_17), .B1(n_14), .B2(n_8), .C(n_10), .Y(n_18) );
O2A1O1Ixp33_ASAP7_75t_L g19 ( .A1(n_17), .A2(n_14), .B(n_9), .C(n_7), .Y(n_19) );
HB1xp67_ASAP7_75t_L g20 ( .A(n_18), .Y(n_20) );
INVx1_ASAP7_75t_L g21 ( .A(n_19), .Y(n_21) );
INVx1_ASAP7_75t_L g22 ( .A(n_20), .Y(n_22) );
AOI22xp5_ASAP7_75t_L g23 ( .A1(n_22), .A2(n_21), .B1(n_12), .B2(n_2), .Y(n_23) );
endmodule