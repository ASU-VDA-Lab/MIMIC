module fake_jpeg_11656_n_510 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_510);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_510;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_6),
.B(n_10),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_5),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_17),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx16f_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_6),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

CKINVDCx14_ASAP7_75t_R g33 ( 
.A(n_10),
.Y(n_33)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

BUFx2_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_8),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

INVx1_ASAP7_75t_SL g43 ( 
.A(n_17),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_1),
.Y(n_44)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_13),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_2),
.Y(n_48)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_49),
.Y(n_111)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_23),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_50),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_18),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_51),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_18),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_52),
.Y(n_151)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_53),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_18),
.Y(n_54)
);

INVx6_ASAP7_75t_L g143 ( 
.A(n_54),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_43),
.B(n_15),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_55),
.B(n_60),
.Y(n_116)
);

INVx6_ASAP7_75t_SL g56 ( 
.A(n_29),
.Y(n_56)
);

CKINVDCx14_ASAP7_75t_R g103 ( 
.A(n_56),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

INVx6_ASAP7_75t_L g147 ( 
.A(n_57),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_58),
.Y(n_148)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_29),
.Y(n_59)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_59),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_43),
.B(n_0),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g146 ( 
.A(n_61),
.Y(n_146)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_28),
.Y(n_62)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_62),
.Y(n_97)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_25),
.Y(n_63)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_63),
.Y(n_106)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_28),
.Y(n_64)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_64),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

INVx6_ASAP7_75t_L g152 ( 
.A(n_65),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

BUFx2_ASAP7_75t_L g100 ( 
.A(n_66),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g145 ( 
.A(n_67),
.Y(n_145)
);

INVx13_ASAP7_75t_L g68 ( 
.A(n_33),
.Y(n_68)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_68),
.Y(n_101)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_29),
.Y(n_69)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_69),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_70),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_71),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_72),
.Y(n_139)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_36),
.Y(n_73)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_73),
.Y(n_117)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_29),
.Y(n_74)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_74),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_47),
.Y(n_75)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_75),
.Y(n_144)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_36),
.Y(n_76)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_76),
.Y(n_118)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_24),
.Y(n_77)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_77),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_47),
.Y(n_78)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_78),
.Y(n_155)
);

OR2x2_ASAP7_75t_L g79 ( 
.A(n_25),
.B(n_32),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_79),
.B(n_27),
.Y(n_105)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_24),
.Y(n_80)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_80),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_43),
.B(n_0),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_81),
.B(n_92),
.Y(n_99)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_24),
.Y(n_82)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_82),
.Y(n_134)
);

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_46),
.Y(n_83)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_83),
.Y(n_154)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_32),
.Y(n_84)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_84),
.Y(n_126)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_42),
.Y(n_85)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_85),
.Y(n_120)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_42),
.Y(n_86)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_86),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_23),
.Y(n_87)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_87),
.Y(n_135)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_42),
.Y(n_88)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_88),
.Y(n_141)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_42),
.Y(n_89)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_89),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_23),
.Y(n_90)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_90),
.Y(n_156)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_20),
.Y(n_91)
);

HB1xp67_ASAP7_75t_L g98 ( 
.A(n_91),
.Y(n_98)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_34),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_34),
.Y(n_93)
);

NOR3xp33_ASAP7_75t_L g130 ( 
.A(n_93),
.B(n_94),
.C(n_95),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_34),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_46),
.Y(n_95)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_20),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_96),
.B(n_41),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_61),
.A2(n_35),
.B1(n_46),
.B2(n_41),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_102),
.A2(n_107),
.B1(n_110),
.B2(n_114),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_105),
.B(n_124),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_66),
.A2(n_35),
.B1(n_41),
.B2(n_20),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_67),
.A2(n_35),
.B1(n_41),
.B2(n_20),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_55),
.A2(n_21),
.B1(n_60),
.B2(n_81),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_113),
.A2(n_137),
.B1(n_11),
.B2(n_12),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_71),
.A2(n_41),
.B1(n_20),
.B2(n_83),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g205 ( 
.A(n_121),
.B(n_129),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_79),
.B(n_21),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_123),
.B(n_125),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_96),
.B(n_27),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_95),
.B(n_48),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_93),
.B(n_48),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_127),
.B(n_133),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_68),
.B(n_30),
.Y(n_129)
);

NAND2x1p5_ASAP7_75t_L g131 ( 
.A(n_72),
.B(n_44),
.Y(n_131)
);

AO22x1_ASAP7_75t_L g192 ( 
.A1(n_131),
.A2(n_140),
.B1(n_3),
.B2(n_4),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_94),
.B(n_44),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_87),
.A2(n_40),
.B1(n_31),
.B2(n_26),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_90),
.A2(n_38),
.B1(n_30),
.B2(n_31),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_75),
.B(n_40),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_149),
.B(n_153),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_78),
.B(n_26),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_L g157 ( 
.A1(n_51),
.A2(n_38),
.B1(n_22),
.B2(n_19),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_157),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_98),
.Y(n_158)
);

HB1xp67_ASAP7_75t_L g222 ( 
.A(n_158),
.Y(n_222)
);

INVx4_ASAP7_75t_SL g160 ( 
.A(n_103),
.Y(n_160)
);

INVx5_ASAP7_75t_SL g233 ( 
.A(n_160),
.Y(n_233)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_106),
.Y(n_161)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_161),
.Y(n_226)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_145),
.Y(n_163)
);

INVx4_ASAP7_75t_L g234 ( 
.A(n_163),
.Y(n_234)
);

INVx8_ASAP7_75t_L g164 ( 
.A(n_142),
.Y(n_164)
);

INVx5_ASAP7_75t_L g239 ( 
.A(n_164),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_116),
.B(n_22),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_165),
.B(n_179),
.Y(n_256)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_156),
.Y(n_166)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_166),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_142),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_167),
.Y(n_261)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_126),
.Y(n_169)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_169),
.Y(n_241)
);

INVx1_ASAP7_75t_SL g170 ( 
.A(n_129),
.Y(n_170)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_170),
.B(n_186),
.Y(n_220)
);

INVx8_ASAP7_75t_L g171 ( 
.A(n_151),
.Y(n_171)
);

INVx3_ASAP7_75t_L g244 ( 
.A(n_171),
.Y(n_244)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_119),
.Y(n_172)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_172),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_100),
.A2(n_19),
.B1(n_58),
.B2(n_57),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_173),
.Y(n_228)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_97),
.Y(n_174)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_174),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_100),
.A2(n_65),
.B1(n_54),
.B2(n_52),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g246 ( 
.A(n_175),
.Y(n_246)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_115),
.Y(n_176)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_176),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_177),
.A2(n_208),
.B1(n_152),
.B2(n_148),
.Y(n_224)
);

BUFx3_ASAP7_75t_L g178 ( 
.A(n_146),
.Y(n_178)
);

BUFx3_ASAP7_75t_L g262 ( 
.A(n_178),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_99),
.B(n_101),
.Y(n_179)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_117),
.Y(n_180)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_180),
.Y(n_217)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_145),
.Y(n_181)
);

BUFx2_ASAP7_75t_SL g221 ( 
.A(n_181),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_151),
.Y(n_182)
);

INVx6_ASAP7_75t_L g240 ( 
.A(n_182),
.Y(n_240)
);

INVx5_ASAP7_75t_L g183 ( 
.A(n_145),
.Y(n_183)
);

INVx6_ASAP7_75t_L g257 ( 
.A(n_183),
.Y(n_257)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_118),
.Y(n_184)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_184),
.Y(n_219)
);

OA22x2_ASAP7_75t_L g185 ( 
.A1(n_131),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_185)
);

OA22x2_ASAP7_75t_L g247 ( 
.A1(n_185),
.A2(n_197),
.B1(n_14),
.B2(n_192),
.Y(n_247)
);

INVx1_ASAP7_75t_SL g186 ( 
.A(n_146),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_122),
.Y(n_187)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_187),
.Y(n_236)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_136),
.Y(n_188)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_188),
.Y(n_254)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_150),
.Y(n_189)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_189),
.Y(n_259)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_134),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_190),
.B(n_193),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_192),
.A2(n_203),
.B1(n_204),
.B2(n_186),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_98),
.Y(n_193)
);

INVx13_ASAP7_75t_L g195 ( 
.A(n_104),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g249 ( 
.A(n_195),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_112),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_196),
.A2(n_210),
.B1(n_214),
.B2(n_102),
.Y(n_227)
);

OA22x2_ASAP7_75t_L g197 ( 
.A1(n_157),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_108),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_198),
.B(n_199),
.Y(n_231)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_109),
.Y(n_199)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_128),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_200),
.B(n_202),
.Y(n_251)
);

INVx3_ASAP7_75t_SL g201 ( 
.A(n_143),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_201),
.Y(n_253)
);

BUFx3_ASAP7_75t_L g202 ( 
.A(n_112),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_143),
.Y(n_203)
);

BUFx2_ASAP7_75t_L g204 ( 
.A(n_128),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_99),
.B(n_7),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_206),
.B(n_207),
.Y(n_223)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_120),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_107),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_121),
.B(n_9),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_209),
.B(n_211),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_130),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_111),
.B(n_10),
.Y(n_211)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_138),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_212),
.B(n_213),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_139),
.B(n_11),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_139),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_215),
.B(n_216),
.Y(n_260)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_141),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_224),
.A2(n_232),
.B1(n_237),
.B2(n_242),
.Y(n_273)
);

OAI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_214),
.A2(n_114),
.B1(n_110),
.B2(n_130),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_225),
.A2(n_227),
.B1(n_182),
.B2(n_167),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_168),
.A2(n_144),
.B1(n_155),
.B2(n_132),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_229),
.A2(n_250),
.B1(n_252),
.B2(n_201),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_162),
.A2(n_152),
.B1(n_148),
.B2(n_147),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_205),
.A2(n_154),
.B(n_155),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_235),
.A2(n_251),
.B(n_219),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_168),
.A2(n_147),
.B1(n_144),
.B2(n_135),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_L g242 ( 
.A1(n_170),
.A2(n_132),
.B1(n_12),
.B2(n_13),
.Y(n_242)
);

AND2x2_ASAP7_75t_SL g243 ( 
.A(n_185),
.B(n_11),
.Y(n_243)
);

AND2x2_ASAP7_75t_L g293 ( 
.A(n_243),
.B(n_247),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_205),
.B(n_13),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_245),
.B(n_189),
.C(n_188),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_159),
.A2(n_14),
.B1(n_213),
.B2(n_185),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_185),
.A2(n_14),
.B1(n_194),
.B2(n_197),
.Y(n_252)
);

A2O1A1Ixp33_ASAP7_75t_L g263 ( 
.A1(n_205),
.A2(n_14),
.B(n_209),
.C(n_197),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_263),
.B(n_264),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_197),
.B(n_176),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_174),
.B(n_184),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_265),
.B(n_166),
.Y(n_279)
);

CKINVDCx16_ASAP7_75t_R g297 ( 
.A(n_266),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_260),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_268),
.B(n_271),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_243),
.A2(n_191),
.B(n_160),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g316 ( 
.A(n_269),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_256),
.B(n_180),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_270),
.B(n_282),
.Y(n_317)
);

INVxp33_ASAP7_75t_L g271 ( 
.A(n_233),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_SL g349 ( 
.A(n_272),
.B(n_307),
.Y(n_349)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_265),
.Y(n_274)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_274),
.Y(n_315)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_260),
.Y(n_275)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_275),
.Y(n_350)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_236),
.Y(n_277)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_277),
.Y(n_328)
);

BUFx24_ASAP7_75t_SL g278 ( 
.A(n_226),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_278),
.B(n_283),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_279),
.B(n_280),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_255),
.B(n_200),
.Y(n_280)
);

BUFx3_ASAP7_75t_L g281 ( 
.A(n_262),
.Y(n_281)
);

HB1xp67_ASAP7_75t_L g324 ( 
.A(n_281),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_255),
.B(n_158),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_SL g283 ( 
.A(n_230),
.B(n_212),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_220),
.Y(n_284)
);

HB1xp67_ASAP7_75t_L g346 ( 
.A(n_284),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_264),
.A2(n_232),
.B1(n_224),
.B2(n_246),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_285),
.A2(n_294),
.B1(n_300),
.B2(n_306),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_L g327 ( 
.A1(n_286),
.A2(n_292),
.B1(n_303),
.B2(n_310),
.Y(n_327)
);

AOI22xp33_ASAP7_75t_SL g287 ( 
.A1(n_228),
.A2(n_202),
.B1(n_204),
.B2(n_178),
.Y(n_287)
);

AOI22xp33_ASAP7_75t_SL g318 ( 
.A1(n_287),
.A2(n_262),
.B1(n_257),
.B2(n_261),
.Y(n_318)
);

OR2x2_ASAP7_75t_L g288 ( 
.A(n_233),
.B(n_163),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_SL g326 ( 
.A1(n_288),
.A2(n_289),
.B(n_296),
.Y(n_326)
);

HB1xp67_ASAP7_75t_L g290 ( 
.A(n_239),
.Y(n_290)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_290),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_231),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_291),
.B(n_295),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_229),
.A2(n_203),
.B1(n_171),
.B2(n_164),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g294 ( 
.A1(n_228),
.A2(n_181),
.B1(n_183),
.B2(n_195),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_218),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_223),
.B(n_230),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_263),
.B(n_245),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_298),
.B(n_309),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_223),
.B(n_220),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_299),
.B(n_272),
.C(n_268),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_237),
.A2(n_266),
.B1(n_247),
.B2(n_235),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_243),
.A2(n_220),
.B1(n_247),
.B2(n_253),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_SL g341 ( 
.A1(n_301),
.A2(n_304),
.B(n_297),
.Y(n_341)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_236),
.Y(n_302)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_302),
.Y(n_331)
);

AOI22xp33_ASAP7_75t_L g303 ( 
.A1(n_244),
.A2(n_247),
.B1(n_219),
.B2(n_259),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_222),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_305),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_241),
.A2(n_248),
.B1(n_244),
.B2(n_254),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_217),
.A2(n_254),
.B1(n_259),
.B2(n_267),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_307),
.A2(n_261),
.B1(n_273),
.B2(n_285),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_217),
.Y(n_308)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_308),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_258),
.B(n_238),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_239),
.A2(n_240),
.B1(n_258),
.B2(n_238),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g311 ( 
.A(n_249),
.Y(n_311)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_311),
.Y(n_345)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_240),
.Y(n_312)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_312),
.Y(n_352)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_221),
.Y(n_313)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_313),
.Y(n_353)
);

OA21x2_ASAP7_75t_L g314 ( 
.A1(n_300),
.A2(n_257),
.B(n_234),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_314),
.B(n_321),
.Y(n_354)
);

INVxp67_ASAP7_75t_L g357 ( 
.A(n_318),
.Y(n_357)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_299),
.B(n_234),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_320),
.B(n_325),
.C(n_329),
.Y(n_361)
);

INVxp33_ASAP7_75t_L g321 ( 
.A(n_288),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_323),
.B(n_310),
.Y(n_355)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_275),
.B(n_282),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_274),
.B(n_280),
.C(n_296),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_332),
.B(n_333),
.C(n_344),
.Y(n_368)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_276),
.B(n_298),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_L g335 ( 
.A1(n_286),
.A2(n_289),
.B1(n_303),
.B2(n_301),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_335),
.A2(n_314),
.B1(n_327),
.B2(n_321),
.Y(n_372)
);

AOI21xp5_ASAP7_75t_L g336 ( 
.A1(n_288),
.A2(n_304),
.B(n_293),
.Y(n_336)
);

AOI21xp5_ASAP7_75t_SL g381 ( 
.A1(n_336),
.A2(n_344),
.B(n_333),
.Y(n_381)
);

OAI21xp5_ASAP7_75t_L g360 ( 
.A1(n_341),
.A2(n_351),
.B(n_309),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_273),
.A2(n_297),
.B1(n_293),
.B2(n_276),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_342),
.A2(n_347),
.B1(n_281),
.B2(n_319),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_293),
.A2(n_283),
.B1(n_295),
.B2(n_294),
.Y(n_343)
);

OAI211xp5_ASAP7_75t_L g387 ( 
.A1(n_343),
.A2(n_336),
.B(n_316),
.C(n_301),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_269),
.B(n_293),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_279),
.A2(n_305),
.B1(n_292),
.B2(n_306),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_349),
.B(n_329),
.C(n_320),
.Y(n_374)
);

OAI21xp5_ASAP7_75t_SL g351 ( 
.A1(n_270),
.A2(n_291),
.B(n_302),
.Y(n_351)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_355),
.Y(n_392)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_328),
.Y(n_356)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_356),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_340),
.B(n_277),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_SL g403 ( 
.A(n_358),
.B(n_380),
.Y(n_403)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_328),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_359),
.B(n_363),
.Y(n_394)
);

OAI21xp5_ASAP7_75t_SL g388 ( 
.A1(n_360),
.A2(n_375),
.B(n_381),
.Y(n_388)
);

OAI21xp5_ASAP7_75t_L g362 ( 
.A1(n_316),
.A2(n_313),
.B(n_290),
.Y(n_362)
);

AOI21xp5_ASAP7_75t_L g396 ( 
.A1(n_362),
.A2(n_367),
.B(n_360),
.Y(n_396)
);

AO22x1_ASAP7_75t_SL g363 ( 
.A1(n_315),
.A2(n_281),
.B1(n_312),
.B2(n_350),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_337),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_364),
.B(n_366),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_SL g402 ( 
.A1(n_365),
.A2(n_377),
.B1(n_382),
.B2(n_387),
.Y(n_402)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_331),
.Y(n_366)
);

OAI21xp5_ASAP7_75t_L g367 ( 
.A1(n_316),
.A2(n_336),
.B(n_341),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_338),
.B(n_351),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_369),
.B(n_370),
.Y(n_416)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_331),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_338),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_371),
.B(n_373),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_SL g407 ( 
.A1(n_372),
.A2(n_385),
.B1(n_355),
.B2(n_354),
.Y(n_407)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_352),
.Y(n_373)
);

MAJx2_ASAP7_75t_L g391 ( 
.A(n_374),
.B(n_361),
.C(n_368),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_346),
.A2(n_314),
.B1(n_326),
.B2(n_348),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_332),
.B(n_317),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_376),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_L g377 ( 
.A1(n_323),
.A2(n_342),
.B1(n_319),
.B2(n_343),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_325),
.B(n_347),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_378),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_326),
.B(n_322),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_379),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_322),
.B(n_334),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_L g382 ( 
.A1(n_352),
.A2(n_334),
.B1(n_330),
.B2(n_349),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_330),
.B(n_339),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_383),
.B(n_384),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_353),
.B(n_345),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_353),
.A2(n_335),
.B1(n_314),
.B2(n_327),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_345),
.B(n_324),
.Y(n_386)
);

XOR2xp5_ASAP7_75t_L g389 ( 
.A(n_386),
.B(n_378),
.Y(n_389)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_389),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_391),
.B(n_397),
.C(n_399),
.Y(n_421)
);

OAI21xp5_ASAP7_75t_SL g432 ( 
.A1(n_396),
.A2(n_400),
.B(n_411),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_374),
.B(n_361),
.C(n_368),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_374),
.B(n_361),
.C(n_368),
.Y(n_399)
);

OA21x2_ASAP7_75t_L g400 ( 
.A1(n_354),
.A2(n_375),
.B(n_372),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_382),
.B(n_376),
.C(n_381),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_401),
.B(n_414),
.C(n_410),
.Y(n_428)
);

XOR2xp5_ASAP7_75t_L g406 ( 
.A(n_379),
.B(n_381),
.Y(n_406)
);

XOR2xp5_ASAP7_75t_L g434 ( 
.A(n_406),
.B(n_410),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_407),
.A2(n_400),
.B1(n_404),
.B2(n_389),
.Y(n_436)
);

AOI22x1_ASAP7_75t_L g409 ( 
.A1(n_377),
.A2(n_365),
.B1(n_387),
.B2(n_369),
.Y(n_409)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_409),
.Y(n_423)
);

XOR2xp5_ASAP7_75t_L g410 ( 
.A(n_380),
.B(n_367),
.Y(n_410)
);

AOI21xp5_ASAP7_75t_L g411 ( 
.A1(n_362),
.A2(n_357),
.B(n_385),
.Y(n_411)
);

OA21x2_ASAP7_75t_L g412 ( 
.A1(n_384),
.A2(n_358),
.B(n_386),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_412),
.B(n_413),
.Y(n_417)
);

OA21x2_ASAP7_75t_L g413 ( 
.A1(n_363),
.A2(n_371),
.B(n_359),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_383),
.B(n_364),
.C(n_363),
.Y(n_414)
);

AOI21xp5_ASAP7_75t_L g415 ( 
.A1(n_356),
.A2(n_366),
.B(n_370),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_415),
.B(n_413),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_398),
.B(n_363),
.Y(n_418)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_418),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_402),
.A2(n_373),
.B1(n_411),
.B2(n_392),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_L g452 ( 
.A1(n_419),
.A2(n_431),
.B1(n_406),
.B2(n_391),
.Y(n_452)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_420),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_SL g424 ( 
.A(n_398),
.B(n_393),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_SL g453 ( 
.A(n_424),
.B(n_425),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_416),
.B(n_395),
.Y(n_425)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_425),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_395),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_426),
.B(n_435),
.Y(n_443)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_416),
.Y(n_427)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_427),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_428),
.B(n_397),
.C(n_399),
.Y(n_441)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_413),
.Y(n_429)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_429),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_412),
.B(n_394),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g450 ( 
.A(n_430),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_SL g431 ( 
.A1(n_402),
.A2(n_392),
.B1(n_414),
.B2(n_394),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_412),
.B(n_390),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g459 ( 
.A(n_433),
.Y(n_459)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_408),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_L g445 ( 
.A1(n_436),
.A2(n_401),
.B1(n_409),
.B2(n_407),
.Y(n_445)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_408),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_437),
.B(n_438),
.Y(n_448)
);

NOR3xp33_ASAP7_75t_SL g438 ( 
.A(n_388),
.B(n_403),
.C(n_396),
.Y(n_438)
);

CKINVDCx14_ASAP7_75t_R g439 ( 
.A(n_415),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_439),
.B(n_440),
.Y(n_458)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_409),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_441),
.B(n_453),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_426),
.B(n_405),
.Y(n_444)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_444),
.Y(n_471)
);

AND2x2_ASAP7_75t_L g466 ( 
.A(n_445),
.B(n_452),
.Y(n_466)
);

OAI21xp5_ASAP7_75t_SL g451 ( 
.A1(n_439),
.A2(n_400),
.B(n_388),
.Y(n_451)
);

AOI21xp5_ASAP7_75t_L g467 ( 
.A1(n_451),
.A2(n_432),
.B(n_420),
.Y(n_467)
);

XOR2xp5_ASAP7_75t_L g454 ( 
.A(n_428),
.B(n_434),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_454),
.B(n_421),
.C(n_422),
.Y(n_464)
);

CKINVDCx16_ASAP7_75t_R g456 ( 
.A(n_417),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_456),
.B(n_457),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_421),
.B(n_434),
.C(n_422),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_424),
.B(n_437),
.Y(n_460)
);

CKINVDCx16_ASAP7_75t_R g473 ( 
.A(n_460),
.Y(n_473)
);

BUFx24_ASAP7_75t_SL g461 ( 
.A(n_448),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_SL g483 ( 
.A(n_461),
.B(n_463),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_448),
.B(n_431),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_464),
.B(n_470),
.C(n_475),
.Y(n_487)
);

AOI21xp5_ASAP7_75t_SL g477 ( 
.A1(n_467),
.A2(n_451),
.B(n_446),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_SL g468 ( 
.A(n_441),
.B(n_453),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_SL g485 ( 
.A(n_468),
.B(n_469),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_SL g469 ( 
.A(n_441),
.B(n_433),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_454),
.B(n_436),
.C(n_432),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_SL g472 ( 
.A(n_444),
.B(n_427),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_472),
.B(n_474),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_SL g474 ( 
.A(n_457),
.B(n_438),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_454),
.B(n_419),
.C(n_418),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_464),
.B(n_445),
.C(n_452),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_476),
.B(n_478),
.Y(n_492)
);

AOI21xp5_ASAP7_75t_SL g491 ( 
.A1(n_477),
.A2(n_486),
.B(n_447),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_466),
.B(n_446),
.C(n_442),
.Y(n_478)
);

OAI21xp5_ASAP7_75t_SL g479 ( 
.A1(n_462),
.A2(n_456),
.B(n_458),
.Y(n_479)
);

AOI21xp5_ASAP7_75t_L g488 ( 
.A1(n_479),
.A2(n_480),
.B(n_482),
.Y(n_488)
);

AOI21xp5_ASAP7_75t_L g480 ( 
.A1(n_465),
.A2(n_458),
.B(n_460),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_475),
.B(n_459),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_470),
.B(n_459),
.Y(n_484)
);

AOI21xp5_ASAP7_75t_L g493 ( 
.A1(n_484),
.A2(n_447),
.B(n_443),
.Y(n_493)
);

OR2x2_ASAP7_75t_L g486 ( 
.A(n_471),
.B(n_449),
.Y(n_486)
);

XOR2xp5_ASAP7_75t_SL g489 ( 
.A(n_481),
.B(n_466),
.Y(n_489)
);

XOR2xp5_ASAP7_75t_L g499 ( 
.A(n_489),
.B(n_494),
.Y(n_499)
);

XOR2xp5_ASAP7_75t_L g490 ( 
.A(n_487),
.B(n_467),
.Y(n_490)
);

AND2x2_ASAP7_75t_L g500 ( 
.A(n_490),
.B(n_476),
.Y(n_500)
);

OAI21xp5_ASAP7_75t_L g497 ( 
.A1(n_491),
.A2(n_495),
.B(n_486),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_SL g496 ( 
.A(n_493),
.B(n_473),
.Y(n_496)
);

OAI21xp33_ASAP7_75t_L g494 ( 
.A1(n_477),
.A2(n_438),
.B(n_450),
.Y(n_494)
);

MAJx2_ASAP7_75t_L g495 ( 
.A(n_485),
.B(n_443),
.C(n_449),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_496),
.B(n_500),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_497),
.B(n_498),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_492),
.B(n_483),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_499),
.B(n_478),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_502),
.B(n_496),
.C(n_423),
.Y(n_505)
);

NOR2xp67_ASAP7_75t_L g504 ( 
.A(n_501),
.B(n_488),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_504),
.B(n_505),
.C(n_503),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_506),
.B(n_435),
.C(n_455),
.Y(n_507)
);

BUFx24_ASAP7_75t_SL g508 ( 
.A(n_507),
.Y(n_508)
);

XNOR2xp5_ASAP7_75t_L g509 ( 
.A(n_508),
.B(n_494),
.Y(n_509)
);

AOI21xp5_ASAP7_75t_L g510 ( 
.A1(n_509),
.A2(n_430),
.B(n_417),
.Y(n_510)
);


endmodule