module fake_jpeg_12698_n_37 (n_3, n_2, n_1, n_0, n_4, n_5, n_37);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_37;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx3_ASAP7_75t_L g6 ( 
.A(n_1),
.Y(n_6)
);

INVx2_ASAP7_75t_L g7 ( 
.A(n_3),
.Y(n_7)
);

BUFx5_ASAP7_75t_L g8 ( 
.A(n_2),
.Y(n_8)
);

BUFx12f_ASAP7_75t_L g9 ( 
.A(n_3),
.Y(n_9)
);

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_3),
.Y(n_10)
);

NOR2xp33_ASAP7_75t_L g11 ( 
.A(n_2),
.B(n_4),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_11),
.B(n_0),
.Y(n_12)
);

AND2x2_ASAP7_75t_L g18 ( 
.A(n_12),
.B(n_13),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_7),
.B(n_0),
.Y(n_13)
);

INVx6_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

BUFx2_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

CKINVDCx12_ASAP7_75t_R g15 ( 
.A(n_9),
.Y(n_15)
);

INVx13_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

AOI22xp33_ASAP7_75t_L g16 ( 
.A1(n_7),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_16)
);

AND2x2_ASAP7_75t_SL g22 ( 
.A(n_16),
.B(n_17),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g17 ( 
.A1(n_6),
.A2(n_1),
.B(n_4),
.Y(n_17)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_21),
.B(n_9),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_L g23 ( 
.A1(n_22),
.A2(n_17),
.B(n_13),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_SL g27 ( 
.A1(n_23),
.A2(n_24),
.B(n_25),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_22),
.A2(n_14),
.B1(n_16),
.B2(n_6),
.Y(n_25)
);

AOI221xp5_ASAP7_75t_L g26 ( 
.A1(n_22),
.A2(n_12),
.B1(n_5),
.B2(n_9),
.C(n_10),
.Y(n_26)
);

OAI21xp33_ASAP7_75t_L g29 ( 
.A1(n_26),
.A2(n_18),
.B(n_5),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_23),
.A2(n_18),
.B1(n_9),
.B2(n_20),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g30 ( 
.A(n_28),
.B(n_29),
.C(n_18),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_L g32 ( 
.A(n_30),
.B(n_31),
.C(n_19),
.Y(n_32)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_27),
.Y(n_31)
);

OAI21xp5_ASAP7_75t_L g34 ( 
.A1(n_32),
.A2(n_33),
.B(n_21),
.Y(n_34)
);

OAI21xp5_ASAP7_75t_L g33 ( 
.A1(n_31),
.A2(n_19),
.B(n_21),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_L g35 ( 
.A1(n_34),
.A2(n_21),
.B1(n_14),
.B2(n_20),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_35),
.B(n_20),
.C(n_8),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_36),
.B(n_8),
.Y(n_37)
);


endmodule