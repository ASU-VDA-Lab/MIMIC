module fake_jpeg_13862_n_32 (n_3, n_2, n_1, n_0, n_4, n_5, n_32);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_32;

wire n_13;
wire n_21;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_12;
wire n_8;
wire n_15;
wire n_7;

BUFx12f_ASAP7_75t_L g6 ( 
.A(n_5),
.Y(n_6)
);

INVx1_ASAP7_75t_L g7 ( 
.A(n_5),
.Y(n_7)
);

AOI21xp33_ASAP7_75t_L g8 ( 
.A1(n_0),
.A2(n_1),
.B(n_2),
.Y(n_8)
);

INVx8_ASAP7_75t_L g9 ( 
.A(n_1),
.Y(n_9)
);

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_3),
.Y(n_10)
);

BUFx12f_ASAP7_75t_L g11 ( 
.A(n_3),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

AOI22xp5_ASAP7_75t_L g13 ( 
.A1(n_10),
.A2(n_12),
.B1(n_8),
.B2(n_9),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_13),
.B(n_18),
.Y(n_23)
);

HB1xp67_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_6),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_15),
.B(n_16),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_SL g16 ( 
.A(n_6),
.B(n_4),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_SL g21 ( 
.A(n_17),
.B(n_19),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_L g18 ( 
.A1(n_10),
.A2(n_0),
.B1(n_4),
.B2(n_12),
.Y(n_18)
);

INVx5_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

MAJx2_ASAP7_75t_L g25 ( 
.A(n_23),
.B(n_13),
.C(n_20),
.Y(n_25)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_25),
.Y(n_27)
);

XNOR2xp5_ASAP7_75t_SL g26 ( 
.A(n_22),
.B(n_11),
.Y(n_26)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_26),
.Y(n_28)
);

AOI21xp5_ASAP7_75t_L g29 ( 
.A1(n_28),
.A2(n_23),
.B(n_21),
.Y(n_29)
);

AOI21xp5_ASAP7_75t_SL g30 ( 
.A1(n_29),
.A2(n_27),
.B(n_28),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_30),
.Y(n_31)
);

AOI221xp5_ASAP7_75t_L g32 ( 
.A1(n_31),
.A2(n_24),
.B1(n_0),
.B2(n_20),
.C(n_19),
.Y(n_32)
);


endmodule