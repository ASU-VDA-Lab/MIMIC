module fake_jpeg_31041_n_479 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_479);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_479;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_13),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_4),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx8_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

HB1xp67_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_6),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_11),
.Y(n_39)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_7),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_10),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_4),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_1),
.Y(n_45)
);

INVx11_ASAP7_75t_SL g46 ( 
.A(n_8),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_0),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_3),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_5),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_14),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_18),
.Y(n_51)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_51),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_21),
.B(n_8),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_52),
.B(n_84),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_18),
.Y(n_53)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_53),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_46),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_54),
.B(n_71),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_55),
.Y(n_108)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

INVx11_ASAP7_75t_L g115 ( 
.A(n_56),
.Y(n_115)
);

INVx6_ASAP7_75t_SL g57 ( 
.A(n_46),
.Y(n_57)
);

INVx1_ASAP7_75t_SL g118 ( 
.A(n_57),
.Y(n_118)
);

BUFx4f_ASAP7_75t_L g58 ( 
.A(n_29),
.Y(n_58)
);

INVx3_ASAP7_75t_SL g105 ( 
.A(n_58),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_18),
.Y(n_59)
);

INVx6_ASAP7_75t_L g145 ( 
.A(n_59),
.Y(n_145)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_18),
.Y(n_60)
);

INVx6_ASAP7_75t_L g147 ( 
.A(n_60),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_24),
.Y(n_61)
);

INVx8_ASAP7_75t_L g109 ( 
.A(n_61),
.Y(n_109)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

INVx8_ASAP7_75t_L g142 ( 
.A(n_62),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_24),
.Y(n_63)
);

INVx11_ASAP7_75t_L g128 ( 
.A(n_63),
.Y(n_128)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_64),
.Y(n_116)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_65),
.Y(n_126)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_26),
.Y(n_66)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_66),
.Y(n_101)
);

BUFx8_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

INVx2_ASAP7_75t_SL g106 ( 
.A(n_67),
.Y(n_106)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_34),
.Y(n_68)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_68),
.Y(n_100)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_34),
.Y(n_69)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_69),
.Y(n_102)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_70),
.Y(n_130)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_21),
.Y(n_71)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_38),
.Y(n_72)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_72),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_29),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_73),
.B(n_74),
.Y(n_112)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_21),
.Y(n_74)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_39),
.Y(n_75)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_75),
.Y(n_139)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_24),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_76),
.B(n_81),
.Y(n_120)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_26),
.Y(n_77)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_77),
.Y(n_132)
);

BUFx24_ASAP7_75t_L g78 ( 
.A(n_29),
.Y(n_78)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_78),
.Y(n_110)
);

INVx11_ASAP7_75t_L g79 ( 
.A(n_24),
.Y(n_79)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_79),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_31),
.Y(n_80)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_80),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_29),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_32),
.B(n_9),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_82),
.B(n_86),
.Y(n_123)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_39),
.Y(n_83)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_83),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_25),
.B(n_9),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_33),
.Y(n_85)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_85),
.Y(n_141)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_33),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_26),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_87),
.B(n_88),
.Y(n_140)
);

BUFx12f_ASAP7_75t_L g88 ( 
.A(n_31),
.Y(n_88)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_23),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_89),
.B(n_90),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_19),
.B(n_9),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_31),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_91),
.A2(n_94),
.B1(n_42),
.B2(n_35),
.Y(n_124)
);

AND2x2_ASAP7_75t_SL g92 ( 
.A(n_31),
.B(n_0),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_92),
.B(n_44),
.C(n_43),
.Y(n_127)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_35),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_93),
.B(n_95),
.Y(n_99)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_39),
.Y(n_94)
);

INVx2_ASAP7_75t_SL g95 ( 
.A(n_22),
.Y(n_95)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_29),
.Y(n_96)
);

OA22x2_ASAP7_75t_L g150 ( 
.A1(n_96),
.A2(n_78),
.B1(n_58),
.B2(n_72),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_19),
.B(n_7),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_97),
.B(n_98),
.Y(n_144)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_22),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_52),
.A2(n_92),
.B1(n_84),
.B2(n_95),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_113),
.A2(n_117),
.B1(n_133),
.B2(n_134),
.Y(n_154)
);

OAI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_60),
.A2(n_22),
.B1(n_40),
.B2(n_35),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_51),
.A2(n_50),
.B1(n_49),
.B2(n_41),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_119),
.A2(n_121),
.B1(n_122),
.B2(n_125),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_92),
.A2(n_40),
.B1(n_35),
.B2(n_17),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_68),
.A2(n_69),
.B1(n_80),
.B2(n_53),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_124),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_59),
.A2(n_40),
.B1(n_20),
.B2(n_27),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_127),
.B(n_43),
.C(n_44),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_85),
.A2(n_42),
.B1(n_20),
.B2(n_27),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_129),
.A2(n_136),
.B1(n_137),
.B2(n_78),
.Y(n_167)
);

OAI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_86),
.A2(n_93),
.B1(n_61),
.B2(n_63),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_79),
.A2(n_25),
.B1(n_45),
.B2(n_47),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_66),
.A2(n_42),
.B1(n_96),
.B2(n_57),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_77),
.A2(n_42),
.B1(n_20),
.B2(n_27),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_91),
.A2(n_17),
.B1(n_49),
.B2(n_41),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_138),
.A2(n_146),
.B1(n_149),
.B2(n_28),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_75),
.A2(n_17),
.B1(n_28),
.B2(n_30),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_83),
.B(n_45),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_148),
.B(n_153),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_55),
.A2(n_47),
.B1(n_23),
.B2(n_50),
.Y(n_149)
);

INVx2_ASAP7_75t_SL g186 ( 
.A(n_150),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_58),
.A2(n_14),
.B(n_16),
.Y(n_152)
);

A2O1A1Ixp33_ASAP7_75t_L g204 ( 
.A1(n_152),
.A2(n_12),
.B(n_13),
.C(n_2),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_94),
.B(n_37),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_111),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_156),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_107),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_157),
.B(n_159),
.Y(n_207)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_100),
.Y(n_158)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_158),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_123),
.B(n_30),
.Y(n_159)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_104),
.Y(n_160)
);

INVx13_ASAP7_75t_L g212 ( 
.A(n_160),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_135),
.B(n_48),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_161),
.B(n_166),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_135),
.B(n_37),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_162),
.B(n_174),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_111),
.Y(n_163)
);

INVx6_ASAP7_75t_L g205 ( 
.A(n_163),
.Y(n_205)
);

INVx1_ASAP7_75t_SL g164 ( 
.A(n_110),
.Y(n_164)
);

AND2x2_ASAP7_75t_L g242 ( 
.A(n_164),
.B(n_173),
.Y(n_242)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_104),
.Y(n_165)
);

INVx13_ASAP7_75t_L g232 ( 
.A(n_165),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_135),
.B(n_48),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_167),
.A2(n_187),
.B1(n_106),
.B2(n_118),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_168),
.A2(n_195),
.B1(n_118),
.B2(n_145),
.Y(n_236)
);

INVx4_ASAP7_75t_SL g170 ( 
.A(n_132),
.Y(n_170)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_170),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_114),
.Y(n_171)
);

INVx5_ASAP7_75t_L g214 ( 
.A(n_171),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_143),
.B(n_67),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_172),
.B(n_188),
.Y(n_219)
);

INVx1_ASAP7_75t_SL g173 ( 
.A(n_110),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_144),
.B(n_48),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_175),
.B(n_180),
.C(n_191),
.Y(n_238)
);

AO22x1_ASAP7_75t_SL g176 ( 
.A1(n_113),
.A2(n_65),
.B1(n_70),
.B2(n_64),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_176),
.A2(n_185),
.B1(n_193),
.B2(n_197),
.Y(n_240)
);

INVx8_ASAP7_75t_L g177 ( 
.A(n_126),
.Y(n_177)
);

INVx5_ASAP7_75t_L g230 ( 
.A(n_177),
.Y(n_230)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_100),
.Y(n_178)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_178),
.Y(n_237)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_139),
.Y(n_179)
);

HB1xp67_ASAP7_75t_L g228 ( 
.A(n_179),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_127),
.B(n_56),
.C(n_67),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_148),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_181),
.B(n_183),
.Y(n_217)
);

INVx6_ASAP7_75t_L g182 ( 
.A(n_109),
.Y(n_182)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_182),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_153),
.Y(n_183)
);

INVx5_ASAP7_75t_L g184 ( 
.A(n_115),
.Y(n_184)
);

BUFx12f_ASAP7_75t_L g210 ( 
.A(n_184),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_L g185 ( 
.A1(n_149),
.A2(n_88),
.B1(n_76),
.B2(n_44),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_102),
.A2(n_42),
.B1(n_76),
.B2(n_88),
.Y(n_187)
);

FAx1_ASAP7_75t_SL g188 ( 
.A(n_144),
.B(n_62),
.CI(n_43),
.CON(n_188),
.SN(n_188)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_112),
.B(n_7),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_190),
.B(n_199),
.Y(n_224)
);

NAND2x1_ASAP7_75t_L g191 ( 
.A(n_152),
.B(n_0),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_102),
.Y(n_192)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_192),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_L g193 ( 
.A1(n_147),
.A2(n_11),
.B1(n_15),
.B2(n_14),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_99),
.B(n_5),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_194),
.B(n_202),
.Y(n_216)
);

OAI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_147),
.A2(n_11),
.B1(n_15),
.B2(n_13),
.Y(n_195)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_139),
.Y(n_196)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_196),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_L g197 ( 
.A1(n_114),
.A2(n_16),
.B1(n_15),
.B2(n_13),
.Y(n_197)
);

BUFx3_ASAP7_75t_L g198 ( 
.A(n_142),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_198),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_146),
.B(n_16),
.Y(n_199)
);

HB1xp67_ASAP7_75t_L g200 ( 
.A(n_101),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_200),
.Y(n_221)
);

HB1xp67_ASAP7_75t_L g201 ( 
.A(n_101),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_201),
.B(n_203),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_99),
.B(n_12),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_134),
.Y(n_203)
);

OAI21xp33_ASAP7_75t_SL g234 ( 
.A1(n_204),
.A2(n_150),
.B(n_126),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_L g206 ( 
.A1(n_203),
.A2(n_168),
.B1(n_186),
.B2(n_189),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_206),
.A2(n_236),
.B1(n_249),
.B2(n_154),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_186),
.A2(n_122),
.B1(n_121),
.B2(n_125),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_208),
.A2(n_211),
.B1(n_227),
.B2(n_169),
.Y(n_252)
);

OAI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_188),
.A2(n_176),
.B1(n_181),
.B2(n_183),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_155),
.B(n_141),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_218),
.B(n_222),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_155),
.B(n_141),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_SL g259 ( 
.A1(n_223),
.A2(n_106),
.B(n_204),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_186),
.A2(n_138),
.B1(n_145),
.B2(n_103),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_157),
.B(n_120),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_229),
.B(n_235),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_198),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_233),
.B(n_247),
.Y(n_255)
);

OAI21xp33_ASAP7_75t_L g289 ( 
.A1(n_234),
.A2(n_116),
.B(n_106),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_194),
.B(n_140),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_202),
.B(n_103),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_241),
.B(n_243),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_172),
.B(n_105),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_188),
.B(n_105),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_245),
.B(n_246),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_161),
.B(n_105),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_158),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_169),
.A2(n_176),
.B1(n_154),
.B2(n_191),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_209),
.Y(n_250)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_250),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_251),
.A2(n_283),
.B1(n_227),
.B2(n_240),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_252),
.A2(n_278),
.B1(n_284),
.B2(n_220),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_226),
.A2(n_191),
.B(n_180),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_253),
.A2(n_259),
.B(n_261),
.Y(n_297)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_209),
.Y(n_254)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_254),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_207),
.B(n_178),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_256),
.B(n_260),
.Y(n_302)
);

AND2x2_ASAP7_75t_L g257 ( 
.A(n_226),
.B(n_150),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g311 ( 
.A(n_257),
.B(n_289),
.Y(n_311)
);

FAx1_ASAP7_75t_L g258 ( 
.A(n_249),
.B(n_175),
.CI(n_166),
.CON(n_258),
.SN(n_258)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_258),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_216),
.B(n_192),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_245),
.A2(n_164),
.B(n_173),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_217),
.B(n_177),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_SL g303 ( 
.A(n_262),
.B(n_274),
.Y(n_303)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_237),
.Y(n_263)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_263),
.Y(n_295)
);

CKINVDCx16_ASAP7_75t_R g264 ( 
.A(n_242),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_264),
.B(n_266),
.Y(n_294)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_228),
.Y(n_265)
);

INVx1_ASAP7_75t_SL g326 ( 
.A(n_265),
.Y(n_326)
);

CKINVDCx16_ASAP7_75t_R g266 ( 
.A(n_242),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_207),
.B(n_165),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_267),
.B(n_273),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_238),
.B(n_150),
.C(n_160),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_268),
.B(n_280),
.C(n_282),
.Y(n_308)
);

BUFx3_ASAP7_75t_L g269 ( 
.A(n_230),
.Y(n_269)
);

BUFx4f_ASAP7_75t_L g315 ( 
.A(n_269),
.Y(n_315)
);

INVx5_ASAP7_75t_L g270 ( 
.A(n_225),
.Y(n_270)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_270),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_238),
.A2(n_242),
.B(n_219),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_271),
.A2(n_253),
.B(n_261),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_217),
.B(n_196),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_224),
.B(n_179),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_224),
.B(n_170),
.Y(n_275)
);

CKINVDCx16_ASAP7_75t_R g313 ( 
.A(n_275),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_216),
.B(n_151),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_276),
.B(n_220),
.Y(n_319)
);

NAND3xp33_ASAP7_75t_L g277 ( 
.A(n_219),
.B(n_116),
.C(n_130),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_277),
.B(n_288),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_208),
.A2(n_151),
.B1(n_109),
.B2(n_171),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_237),
.Y(n_279)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_279),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_213),
.B(n_131),
.C(n_130),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_229),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_281),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_213),
.B(n_131),
.C(n_108),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_236),
.A2(n_128),
.B1(n_156),
.B2(n_163),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_240),
.A2(n_182),
.B1(n_128),
.B2(n_132),
.Y(n_284)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_243),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_247),
.B(n_170),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_290),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_296),
.A2(n_301),
.B1(n_272),
.B2(n_286),
.Y(n_337)
);

AOI21xp5_ASAP7_75t_L g351 ( 
.A1(n_299),
.A2(n_259),
.B(n_275),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_300),
.A2(n_309),
.B1(n_310),
.B2(n_316),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_251),
.A2(n_246),
.B1(n_218),
.B2(n_222),
.Y(n_301)
);

AND2x2_ASAP7_75t_SL g304 ( 
.A(n_287),
.B(n_244),
.Y(n_304)
);

CKINVDCx16_ASAP7_75t_R g338 ( 
.A(n_304),
.Y(n_338)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_290),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_306),
.B(n_321),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_252),
.A2(n_241),
.B1(n_235),
.B2(n_244),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_284),
.A2(n_215),
.B1(n_233),
.B2(n_231),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_278),
.A2(n_215),
.B1(n_231),
.B2(n_239),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_258),
.B(n_248),
.C(n_221),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_317),
.B(n_320),
.C(n_268),
.Y(n_332)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_250),
.Y(n_318)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_318),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_SL g344 ( 
.A(n_319),
.B(n_276),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_258),
.B(n_248),
.C(n_228),
.Y(n_320)
);

AOI32xp33_ASAP7_75t_L g321 ( 
.A1(n_258),
.A2(n_205),
.A3(n_230),
.B1(n_239),
.B2(n_212),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_254),
.Y(n_322)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_322),
.Y(n_339)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_263),
.Y(n_323)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_323),
.Y(n_350)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_255),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_324),
.B(n_262),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_255),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_327),
.Y(n_349)
);

BUFx12f_ASAP7_75t_SL g330 ( 
.A(n_312),
.Y(n_330)
);

INVxp67_ASAP7_75t_L g361 ( 
.A(n_330),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_SL g384 ( 
.A(n_332),
.B(n_341),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_327),
.B(n_292),
.Y(n_333)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_333),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_L g334 ( 
.A1(n_296),
.A2(n_257),
.B1(n_281),
.B2(n_268),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_334),
.A2(n_336),
.B1(n_337),
.B2(n_346),
.Y(n_366)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_335),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_L g336 ( 
.A1(n_298),
.A2(n_257),
.B1(n_286),
.B2(n_285),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_300),
.A2(n_257),
.B1(n_283),
.B2(n_260),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_340),
.A2(n_307),
.B1(n_294),
.B2(n_321),
.Y(n_369)
);

MAJx2_ASAP7_75t_L g341 ( 
.A(n_308),
.B(n_287),
.C(n_285),
.Y(n_341)
);

XNOR2x1_ASAP7_75t_L g342 ( 
.A(n_308),
.B(n_280),
.Y(n_342)
);

XOR2xp5_ASAP7_75t_L g362 ( 
.A(n_342),
.B(n_344),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_317),
.B(n_271),
.C(n_280),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_343),
.B(n_354),
.C(n_311),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_SL g345 ( 
.A(n_292),
.B(n_256),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_SL g363 ( 
.A(n_345),
.B(n_355),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_L g346 ( 
.A1(n_301),
.A2(n_272),
.B1(n_273),
.B2(n_282),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_309),
.B(n_274),
.Y(n_347)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_347),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_302),
.B(n_267),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_348),
.B(n_356),
.Y(n_377)
);

INVxp67_ASAP7_75t_L g381 ( 
.A(n_351),
.Y(n_381)
);

BUFx12f_ASAP7_75t_L g352 ( 
.A(n_315),
.Y(n_352)
);

BUFx6f_ASAP7_75t_L g374 ( 
.A(n_352),
.Y(n_374)
);

INVx13_ASAP7_75t_L g353 ( 
.A(n_315),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_353),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_299),
.B(n_277),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_303),
.B(n_265),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_302),
.B(n_279),
.Y(n_356)
);

OAI32xp33_ASAP7_75t_L g357 ( 
.A1(n_325),
.A2(n_266),
.A3(n_264),
.B1(n_210),
.B2(n_269),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_L g365 ( 
.A1(n_357),
.A2(n_360),
.B1(n_325),
.B2(n_313),
.Y(n_365)
);

AOI21xp5_ASAP7_75t_L g358 ( 
.A1(n_311),
.A2(n_269),
.B(n_184),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_358),
.A2(n_359),
.B1(n_313),
.B2(n_311),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_320),
.A2(n_205),
.B1(n_225),
.B2(n_214),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_291),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_365),
.B(n_369),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_367),
.A2(n_389),
.B1(n_338),
.B2(n_371),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_L g368 ( 
.A1(n_328),
.A2(n_297),
.B1(n_303),
.B2(n_304),
.Y(n_368)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_368),
.Y(n_404)
);

XOR2xp5_ASAP7_75t_L g370 ( 
.A(n_342),
.B(n_297),
.Y(n_370)
);

XOR2xp5_ASAP7_75t_L g402 ( 
.A(n_370),
.B(n_359),
.Y(n_402)
);

NOR2x1_ASAP7_75t_SL g371 ( 
.A(n_330),
.B(n_304),
.Y(n_371)
);

A2O1A1O1Ixp25_ASAP7_75t_L g400 ( 
.A1(n_371),
.A2(n_356),
.B(n_349),
.C(n_357),
.D(n_338),
.Y(n_400)
);

XNOR2x1_ASAP7_75t_L g412 ( 
.A(n_372),
.B(n_315),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_SL g373 ( 
.A1(n_329),
.A2(n_307),
.B1(n_304),
.B2(n_294),
.Y(n_373)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_373),
.Y(n_392)
);

BUFx24_ASAP7_75t_SL g375 ( 
.A(n_341),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_SL g407 ( 
.A(n_375),
.B(n_331),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_332),
.B(n_319),
.C(n_310),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_376),
.B(n_380),
.C(n_382),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_333),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_SL g409 ( 
.A(n_378),
.B(n_350),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_SL g379 ( 
.A1(n_329),
.A2(n_316),
.B1(n_323),
.B2(n_322),
.Y(n_379)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_379),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_343),
.B(n_293),
.C(n_318),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_346),
.B(n_291),
.C(n_314),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_334),
.B(n_293),
.C(n_295),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_383),
.B(n_387),
.C(n_349),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_340),
.A2(n_295),
.B1(n_314),
.B2(n_326),
.Y(n_385)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_385),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_344),
.B(n_336),
.C(n_351),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_SL g417 ( 
.A1(n_390),
.A2(n_369),
.B1(n_385),
.B2(n_379),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_363),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_393),
.B(n_394),
.Y(n_420)
);

NOR2x1_ASAP7_75t_L g394 ( 
.A(n_373),
.B(n_345),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_SL g395 ( 
.A(n_370),
.B(n_354),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_395),
.B(n_396),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_376),
.B(n_337),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_397),
.B(n_399),
.C(n_402),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g399 ( 
.A(n_387),
.B(n_348),
.Y(n_399)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_400),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_383),
.B(n_331),
.Y(n_401)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_401),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_384),
.B(n_358),
.C(n_360),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_405),
.B(n_411),
.C(n_412),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_407),
.B(n_410),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_388),
.B(n_350),
.Y(n_408)
);

INVxp67_ASAP7_75t_L g429 ( 
.A(n_408),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_409),
.B(n_377),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_386),
.B(n_339),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_L g411 ( 
.A(n_382),
.B(n_339),
.Y(n_411)
);

AOI22xp33_ASAP7_75t_SL g413 ( 
.A1(n_389),
.A2(n_352),
.B1(n_315),
.B2(n_305),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_L g419 ( 
.A1(n_413),
.A2(n_374),
.B1(n_367),
.B2(n_364),
.Y(n_419)
);

NOR2xp67_ASAP7_75t_L g414 ( 
.A(n_394),
.B(n_361),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_414),
.B(n_416),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_SL g434 ( 
.A1(n_417),
.A2(n_403),
.B1(n_398),
.B2(n_406),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_L g437 ( 
.A1(n_419),
.A2(n_398),
.B1(n_406),
.B2(n_402),
.Y(n_437)
);

A2O1A1Ixp33_ASAP7_75t_L g421 ( 
.A1(n_392),
.A2(n_377),
.B(n_381),
.C(n_361),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_SL g438 ( 
.A(n_421),
.B(n_426),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_391),
.B(n_380),
.C(n_396),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_422),
.B(n_428),
.C(n_430),
.Y(n_436)
);

OAI21xp5_ASAP7_75t_SL g426 ( 
.A1(n_404),
.A2(n_381),
.B(n_372),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_SL g427 ( 
.A(n_399),
.B(n_366),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_427),
.B(n_400),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_391),
.B(n_384),
.C(n_362),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_397),
.B(n_362),
.C(n_366),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_392),
.B(n_326),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_432),
.B(n_403),
.Y(n_433)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_433),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_SL g447 ( 
.A(n_434),
.B(n_439),
.Y(n_447)
);

XOR2xp5_ASAP7_75t_SL g435 ( 
.A(n_420),
.B(n_390),
.Y(n_435)
);

NAND2x1_ASAP7_75t_SL g458 ( 
.A(n_435),
.B(n_425),
.Y(n_458)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_437),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_422),
.B(n_412),
.C(n_411),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_429),
.B(n_374),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_440),
.B(n_443),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_441),
.B(n_444),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_L g443 ( 
.A1(n_423),
.A2(n_305),
.B1(n_270),
.B2(n_205),
.Y(n_443)
);

BUFx6f_ASAP7_75t_L g444 ( 
.A(n_424),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_431),
.B(n_352),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_445),
.B(n_416),
.Y(n_448)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_448),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g449 ( 
.A(n_439),
.B(n_436),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_449),
.B(n_454),
.Y(n_460)
);

NOR2xp67_ASAP7_75t_L g450 ( 
.A(n_442),
.B(n_435),
.Y(n_450)
);

INVxp67_ASAP7_75t_L g465 ( 
.A(n_450),
.Y(n_465)
);

OAI321xp33_ASAP7_75t_L g453 ( 
.A1(n_433),
.A2(n_421),
.A3(n_429),
.B1(n_417),
.B2(n_426),
.C(n_418),
.Y(n_453)
);

AOI22xp33_ASAP7_75t_L g464 ( 
.A1(n_453),
.A2(n_270),
.B1(n_353),
.B2(n_210),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_SL g454 ( 
.A(n_444),
.B(n_425),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_440),
.B(n_415),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_455),
.B(n_436),
.Y(n_462)
);

OAI21xp5_ASAP7_75t_L g456 ( 
.A1(n_438),
.A2(n_430),
.B(n_428),
.Y(n_456)
);

INVxp67_ASAP7_75t_L g466 ( 
.A(n_458),
.Y(n_466)
);

NAND2xp33_ASAP7_75t_SL g459 ( 
.A(n_451),
.B(n_434),
.Y(n_459)
);

AOI322xp5_ASAP7_75t_L g468 ( 
.A1(n_459),
.A2(n_465),
.A3(n_446),
.B1(n_466),
.B2(n_457),
.C1(n_461),
.C2(n_452),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_447),
.B(n_225),
.C(n_352),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_464),
.B(n_467),
.Y(n_472)
);

OAI21xp5_ASAP7_75t_SL g467 ( 
.A1(n_456),
.A2(n_210),
.B(n_212),
.Y(n_467)
);

AOI322xp5_ASAP7_75t_L g474 ( 
.A1(n_468),
.A2(n_470),
.A3(n_232),
.B1(n_115),
.B2(n_12),
.C1(n_3),
.C2(n_0),
.Y(n_474)
);

AND2x2_ASAP7_75t_L g469 ( 
.A(n_460),
.B(n_463),
.Y(n_469)
);

OAI22xp5_ASAP7_75t_L g470 ( 
.A1(n_465),
.A2(n_458),
.B1(n_214),
.B2(n_108),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_466),
.B(n_210),
.C(n_142),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_471),
.B(n_232),
.C(n_212),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_473),
.B(n_474),
.Y(n_477)
);

AOI322xp5_ASAP7_75t_L g475 ( 
.A1(n_472),
.A2(n_232),
.A3(n_12),
.B1(n_3),
.B2(n_4),
.C1(n_2),
.C2(n_1),
.Y(n_475)
);

AOI321xp33_ASAP7_75t_SL g476 ( 
.A1(n_475),
.A2(n_1),
.A3(n_2),
.B1(n_3),
.B2(n_4),
.C(n_469),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_477),
.B(n_2),
.C(n_462),
.Y(n_478)
);

FAx1_ASAP7_75t_SL g479 ( 
.A(n_478),
.B(n_333),
.CI(n_476),
.CON(n_479),
.SN(n_479)
);


endmodule