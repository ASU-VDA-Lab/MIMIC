module fake_netlist_1_9975_n_40 (n_11, n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_40);
input n_11;
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_40;
wire n_20;
wire n_38;
wire n_36;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
wire n_39;
INVx3_ASAP7_75t_L g12 ( .A(n_3), .Y(n_12) );
CKINVDCx5p33_ASAP7_75t_R g13 ( .A(n_2), .Y(n_13) );
AND2x2_ASAP7_75t_L g14 ( .A(n_0), .B(n_2), .Y(n_14) );
INVx2_ASAP7_75t_L g15 ( .A(n_4), .Y(n_15) );
INVx1_ASAP7_75t_L g16 ( .A(n_0), .Y(n_16) );
INVx2_ASAP7_75t_L g17 ( .A(n_9), .Y(n_17) );
BUFx3_ASAP7_75t_L g18 ( .A(n_12), .Y(n_18) );
BUFx2_ASAP7_75t_L g19 ( .A(n_13), .Y(n_19) );
O2A1O1Ixp33_ASAP7_75t_L g20 ( .A1(n_16), .A2(n_1), .B(n_5), .C(n_6), .Y(n_20) );
NAND2xp5_ASAP7_75t_L g21 ( .A(n_12), .B(n_1), .Y(n_21) );
O2A1O1Ixp33_ASAP7_75t_SL g22 ( .A1(n_21), .A2(n_15), .B(n_17), .C(n_14), .Y(n_22) );
AND2x2_ASAP7_75t_L g23 ( .A(n_19), .B(n_13), .Y(n_23) );
AND2x4_ASAP7_75t_L g24 ( .A(n_18), .B(n_15), .Y(n_24) );
AND2x2_ASAP7_75t_L g25 ( .A(n_23), .B(n_21), .Y(n_25) );
BUFx6f_ASAP7_75t_L g26 ( .A(n_24), .Y(n_26) );
BUFx2_ASAP7_75t_L g27 ( .A(n_25), .Y(n_27) );
CKINVDCx20_ASAP7_75t_R g28 ( .A(n_26), .Y(n_28) );
INVx1_ASAP7_75t_L g29 ( .A(n_27), .Y(n_29) );
AND2x2_ASAP7_75t_L g30 ( .A(n_28), .B(n_23), .Y(n_30) );
O2A1O1Ixp5_ASAP7_75t_L g31 ( .A1(n_29), .A2(n_24), .B(n_22), .C(n_26), .Y(n_31) );
NAND2xp33_ASAP7_75t_SL g32 ( .A(n_30), .B(n_26), .Y(n_32) );
INVx1_ASAP7_75t_L g33 ( .A(n_30), .Y(n_33) );
INVx1_ASAP7_75t_L g34 ( .A(n_33), .Y(n_34) );
NAND4xp75_ASAP7_75t_L g35 ( .A(n_31), .B(n_20), .C(n_8), .D(n_10), .Y(n_35) );
OAI21xp5_ASAP7_75t_L g36 ( .A1(n_33), .A2(n_24), .B(n_7), .Y(n_36) );
AND2x2_ASAP7_75t_L g37 ( .A(n_34), .B(n_36), .Y(n_37) );
INVx1_ASAP7_75t_L g38 ( .A(n_35), .Y(n_38) );
OAI22xp5_ASAP7_75t_L g39 ( .A1(n_37), .A2(n_35), .B1(n_32), .B2(n_11), .Y(n_39) );
NAND3xp33_ASAP7_75t_L g40 ( .A(n_39), .B(n_38), .C(n_37), .Y(n_40) );
endmodule