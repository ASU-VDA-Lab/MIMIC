module fake_jpeg_13002_n_175 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_175);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_175;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_93;
wire n_91;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx2_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_23),
.Y(n_47)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_18),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_34),
.Y(n_50)
);

CKINVDCx5p33_ASAP7_75t_R g51 ( 
.A(n_14),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_26),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_20),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_31),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

BUFx12_ASAP7_75t_L g56 ( 
.A(n_27),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_19),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_9),
.B(n_8),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_7),
.Y(n_59)
);

INVx6_ASAP7_75t_SL g60 ( 
.A(n_24),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_28),
.B(n_12),
.Y(n_61)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_8),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_6),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_5),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_43),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_38),
.Y(n_68)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_36),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_33),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_17),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_59),
.B(n_0),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_72),
.B(n_76),
.Y(n_88)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_60),
.Y(n_73)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_73),
.Y(n_84)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_53),
.Y(n_74)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_74),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_71),
.Y(n_75)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_75),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_58),
.B(n_0),
.Y(n_76)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_71),
.Y(n_77)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_77),
.Y(n_90)
);

INVx2_ASAP7_75t_SL g78 ( 
.A(n_57),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_78),
.B(n_79),
.Y(n_89)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_64),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_58),
.B(n_1),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_80),
.B(n_1),
.Y(n_92)
);

NOR2x1_ASAP7_75t_L g81 ( 
.A(n_74),
.B(n_65),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_81),
.B(n_83),
.Y(n_96)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_75),
.Y(n_82)
);

INVx1_ASAP7_75t_SL g102 ( 
.A(n_82),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_77),
.Y(n_83)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_78),
.Y(n_85)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_85),
.Y(n_116)
);

INVx4_ASAP7_75t_SL g86 ( 
.A(n_73),
.Y(n_86)
);

CKINVDCx14_ASAP7_75t_R g99 ( 
.A(n_86),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_73),
.B(n_50),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_87),
.B(n_93),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_92),
.B(n_95),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_80),
.B(n_50),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_80),
.B(n_67),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_88),
.B(n_89),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_97),
.B(n_107),
.Y(n_119)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_91),
.Y(n_98)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_98),
.Y(n_129)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_89),
.Y(n_100)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_100),
.Y(n_121)
);

AND2x6_ASAP7_75t_L g101 ( 
.A(n_88),
.B(n_37),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_101),
.B(n_110),
.Y(n_126)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_90),
.Y(n_103)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_103),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_92),
.Y(n_104)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_104),
.Y(n_134)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_94),
.Y(n_106)
);

BUFx2_ASAP7_75t_L g120 ( 
.A(n_106),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_84),
.B(n_54),
.Y(n_107)
);

INVxp67_ASAP7_75t_SL g109 ( 
.A(n_82),
.Y(n_109)
);

INVx13_ASAP7_75t_L g132 ( 
.A(n_109),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_93),
.B(n_61),
.Y(n_110)
);

INVx11_ASAP7_75t_L g111 ( 
.A(n_86),
.Y(n_111)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_111),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_89),
.A2(n_55),
.B(n_63),
.Y(n_112)
);

NOR3xp33_ASAP7_75t_L g118 ( 
.A(n_112),
.B(n_51),
.C(n_66),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_90),
.A2(n_62),
.B1(n_57),
.B2(n_70),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_113),
.A2(n_99),
.B1(n_48),
.B2(n_56),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_95),
.B(n_68),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_114),
.B(n_47),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_93),
.B(n_61),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_SL g135 ( 
.A(n_115),
.B(n_99),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_96),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_117),
.B(n_118),
.Y(n_141)
);

OAI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_113),
.A2(n_45),
.B1(n_46),
.B2(n_69),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_122),
.A2(n_128),
.B1(n_3),
.B2(n_4),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_123),
.B(n_119),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_105),
.B(n_52),
.Y(n_124)
);

NAND3xp33_ASAP7_75t_L g139 ( 
.A(n_124),
.B(n_130),
.C(n_3),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_108),
.B(n_62),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_125),
.A2(n_4),
.B(n_5),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_116),
.B(n_2),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_127),
.B(n_137),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_106),
.A2(n_109),
.B1(n_48),
.B2(n_102),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_101),
.B(n_49),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_131),
.B(n_25),
.Y(n_150)
);

NOR4xp25_ASAP7_75t_L g151 ( 
.A(n_135),
.B(n_29),
.C(n_40),
.D(n_10),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_104),
.B(n_2),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_98),
.Y(n_138)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_138),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_139),
.B(n_145),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_124),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_140),
.B(n_144),
.Y(n_156)
);

OR2x2_ASAP7_75t_L g143 ( 
.A(n_121),
.B(n_56),
.Y(n_143)
);

INVxp33_ASAP7_75t_L g162 ( 
.A(n_143),
.Y(n_162)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_133),
.Y(n_144)
);

INVxp33_ASAP7_75t_L g163 ( 
.A(n_146),
.Y(n_163)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_129),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_147),
.B(n_149),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_148),
.B(n_150),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_134),
.B(n_6),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_151),
.B(n_152),
.Y(n_160)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_136),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_120),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_153),
.A2(n_155),
.B(n_126),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_130),
.A2(n_7),
.B1(n_9),
.B2(n_11),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_161),
.B(n_125),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_SL g164 ( 
.A(n_156),
.B(n_157),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_164),
.B(n_166),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_163),
.A2(n_154),
.B1(n_143),
.B2(n_149),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_165),
.A2(n_167),
.B(n_139),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_162),
.A2(n_141),
.B(n_142),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_169),
.B(n_159),
.C(n_158),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_170),
.B(n_168),
.Y(n_171)
);

AOI322xp5_ASAP7_75t_L g172 ( 
.A1(n_171),
.A2(n_160),
.A3(n_132),
.B1(n_15),
.B2(n_16),
.C1(n_21),
.C2(n_22),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_172),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_173),
.A2(n_163),
.B(n_150),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_174),
.B(n_13),
.Y(n_175)
);


endmodule