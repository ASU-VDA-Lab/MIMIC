module real_aes_9126_n_77 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_77);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_77;
wire n_480;
wire n_113;
wire n_476;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_522;
wire n_485;
wire n_222;
wire n_503;
wire n_287;
wire n_357;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_540;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_341;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_260;
wire n_97;
wire n_186;
wire n_138;
wire n_379;
wire n_374;
wire n_453;
wire n_235;
wire n_399;
wire n_378;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_145;
wire n_415;
wire n_227;
wire n_92;
wire n_519;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_462;
wire n_289;
wire n_280;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_408;
wire n_184;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_506;
wire n_513;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_164;
wire n_231;
wire n_102;
wire n_454;
wire n_122;
wire n_443;
wire n_534;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_204;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_331;
wire n_93;
wire n_182;
wire n_417;
wire n_449;
wire n_363;
wire n_323;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_368;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_250;
wire n_85;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_402;
wire n_87;
wire n_171;
wire n_78;
wire n_531;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_501;
wire n_488;
wire n_251;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_158;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_109;
wire n_536;
wire n_203;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_526;
wire n_155;
wire n_243;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_446;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_266;
wire n_183;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_180;
wire n_212;
wire n_210;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_371;
wire n_103;
wire n_166;
wire n_224;
wire n_151;
wire n_130;
wire n_253;
wire n_459;
wire n_99;
wire n_440;
wire n_525;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_305;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_465;
wire n_473;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_340;
wire n_483;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_206;
wire n_307;
wire n_500;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_264;
wire n_237;
wire n_91;
A2O1A1Ixp33_ASAP7_75t_L g293 ( .A1(n_0), .A2(n_196), .B(n_199), .C(n_294), .Y(n_293) );
AOI21xp5_ASAP7_75t_L g320 ( .A1(n_1), .A2(n_231), .B(n_321), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_2), .B(n_271), .Y(n_328) );
AOI22xp33_ASAP7_75t_L g145 ( .A1(n_3), .A2(n_42), .B1(n_146), .B2(n_153), .Y(n_145) );
INVx1_ASAP7_75t_L g182 ( .A(n_4), .Y(n_182) );
AND2x6_ASAP7_75t_L g196 ( .A(n_4), .B(n_180), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_4), .B(n_534), .Y(n_533) );
INVx1_ASAP7_75t_L g254 ( .A(n_5), .Y(n_254) );
NAND2xp5_ASAP7_75t_SL g298 ( .A(n_6), .B(n_207), .Y(n_298) );
AO22x2_ASAP7_75t_L g99 ( .A1(n_7), .A2(n_24), .B1(n_91), .B2(n_96), .Y(n_99) );
INVx1_ASAP7_75t_L g215 ( .A(n_8), .Y(n_215) );
A2O1A1Ixp33_ASAP7_75t_L g278 ( .A1(n_9), .A2(n_205), .B(n_279), .C(n_281), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_10), .B(n_271), .Y(n_282) );
AO22x2_ASAP7_75t_L g101 ( .A1(n_11), .A2(n_26), .B1(n_91), .B2(n_92), .Y(n_101) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_12), .B(n_244), .Y(n_243) );
CKINVDCx20_ASAP7_75t_R g144 ( .A(n_13), .Y(n_144) );
A2O1A1Ixp33_ASAP7_75t_L g264 ( .A1(n_14), .A2(n_265), .B(n_266), .C(n_268), .Y(n_264) );
NAND2xp5_ASAP7_75t_SL g315 ( .A(n_15), .B(n_207), .Y(n_315) );
NAND2xp5_ASAP7_75t_SL g206 ( .A(n_16), .B(n_207), .Y(n_206) );
CKINVDCx16_ASAP7_75t_R g311 ( .A(n_17), .Y(n_311) );
INVx1_ASAP7_75t_L g203 ( .A(n_18), .Y(n_203) );
BUFx6f_ASAP7_75t_L g195 ( .A(n_19), .Y(n_195) );
CKINVDCx20_ASAP7_75t_R g292 ( .A(n_20), .Y(n_292) );
AOI22xp5_ASAP7_75t_L g514 ( .A1(n_20), .A2(n_292), .B1(n_515), .B2(n_516), .Y(n_514) );
CKINVDCx20_ASAP7_75t_R g126 ( .A(n_21), .Y(n_126) );
INVx1_ASAP7_75t_L g237 ( .A(n_22), .Y(n_237) );
INVx2_ASAP7_75t_L g194 ( .A(n_23), .Y(n_194) );
CKINVDCx20_ASAP7_75t_R g301 ( .A(n_25), .Y(n_301) );
OAI221xp5_ASAP7_75t_L g524 ( .A1(n_26), .A2(n_43), .B1(n_54), .B2(n_525), .C(n_526), .Y(n_524) );
INVxp67_ASAP7_75t_L g527 ( .A(n_26), .Y(n_527) );
A2O1A1Ixp33_ASAP7_75t_L g323 ( .A1(n_27), .A2(n_265), .B(n_324), .C(n_326), .Y(n_323) );
AOI22xp33_ASAP7_75t_L g106 ( .A1(n_28), .A2(n_56), .B1(n_107), .B2(n_114), .Y(n_106) );
INVxp67_ASAP7_75t_L g238 ( .A(n_29), .Y(n_238) );
A2O1A1Ixp33_ASAP7_75t_L g198 ( .A1(n_30), .A2(n_199), .B(n_202), .C(n_210), .Y(n_198) );
CKINVDCx14_ASAP7_75t_R g322 ( .A(n_31), .Y(n_322) );
A2O1A1Ixp33_ASAP7_75t_L g251 ( .A1(n_32), .A2(n_252), .B(n_253), .C(n_255), .Y(n_251) );
INVx1_ASAP7_75t_L g538 ( .A(n_32), .Y(n_538) );
CKINVDCx20_ASAP7_75t_R g132 ( .A(n_33), .Y(n_132) );
AOI22xp33_ASAP7_75t_L g84 ( .A1(n_34), .A2(n_55), .B1(n_85), .B2(n_102), .Y(n_84) );
AOI22xp33_ASAP7_75t_L g168 ( .A1(n_35), .A2(n_70), .B1(n_169), .B2(n_172), .Y(n_168) );
CKINVDCx20_ASAP7_75t_R g217 ( .A(n_36), .Y(n_217) );
CKINVDCx20_ASAP7_75t_R g233 ( .A(n_37), .Y(n_233) );
AOI22xp5_ASAP7_75t_L g511 ( .A1(n_38), .A2(n_73), .B1(n_512), .B2(n_513), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_38), .Y(n_512) );
OAI22xp5_ASAP7_75t_SL g516 ( .A1(n_39), .A2(n_72), .B1(n_517), .B2(n_518), .Y(n_516) );
INVx1_ASAP7_75t_L g518 ( .A(n_39), .Y(n_518) );
INVx1_ASAP7_75t_L g263 ( .A(n_40), .Y(n_263) );
CKINVDCx20_ASAP7_75t_R g135 ( .A(n_41), .Y(n_135) );
AO22x2_ASAP7_75t_L g90 ( .A1(n_43), .A2(n_65), .B1(n_91), .B2(n_92), .Y(n_90) );
INVxp67_ASAP7_75t_L g528 ( .A(n_43), .Y(n_528) );
CKINVDCx14_ASAP7_75t_R g250 ( .A(n_44), .Y(n_250) );
AOI22xp33_ASAP7_75t_SL g158 ( .A1(n_45), .A2(n_68), .B1(n_159), .B2(n_163), .Y(n_158) );
INVx1_ASAP7_75t_L g180 ( .A(n_46), .Y(n_180) );
INVx1_ASAP7_75t_L g214 ( .A(n_47), .Y(n_214) );
AOI22xp5_ASAP7_75t_L g79 ( .A1(n_48), .A2(n_80), .B1(n_81), .B2(n_174), .Y(n_79) );
CKINVDCx20_ASAP7_75t_R g174 ( .A(n_48), .Y(n_174) );
INVx1_ASAP7_75t_SL g325 ( .A(n_49), .Y(n_325) );
CKINVDCx20_ASAP7_75t_R g525 ( .A(n_50), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_51), .B(n_271), .Y(n_270) );
CKINVDCx20_ASAP7_75t_R g119 ( .A(n_52), .Y(n_119) );
INVx1_ASAP7_75t_L g314 ( .A(n_53), .Y(n_314) );
AO22x2_ASAP7_75t_L g95 ( .A1(n_54), .A2(n_71), .B1(n_91), .B2(n_96), .Y(n_95) );
AOI21xp5_ASAP7_75t_L g248 ( .A1(n_57), .A2(n_231), .B(n_249), .Y(n_248) );
AOI22xp5_ASAP7_75t_L g508 ( .A1(n_57), .A2(n_509), .B1(n_521), .B2(n_529), .Y(n_508) );
INVx1_ASAP7_75t_L g540 ( .A(n_57), .Y(n_540) );
CKINVDCx20_ASAP7_75t_R g318 ( .A(n_58), .Y(n_318) );
AOI21xp5_ASAP7_75t_L g275 ( .A1(n_59), .A2(n_231), .B(n_276), .Y(n_275) );
AOI21xp5_ASAP7_75t_L g229 ( .A1(n_60), .A2(n_230), .B(n_232), .Y(n_229) );
CKINVDCx16_ASAP7_75t_R g197 ( .A(n_61), .Y(n_197) );
INVx1_ASAP7_75t_L g277 ( .A(n_62), .Y(n_277) );
AOI21xp5_ASAP7_75t_L g261 ( .A1(n_63), .A2(n_231), .B(n_262), .Y(n_261) );
INVx1_ASAP7_75t_L g280 ( .A(n_64), .Y(n_280) );
INVx2_ASAP7_75t_L g212 ( .A(n_66), .Y(n_212) );
INVx1_ASAP7_75t_L g295 ( .A(n_67), .Y(n_295) );
A2O1A1Ixp33_ASAP7_75t_L g312 ( .A1(n_69), .A2(n_199), .B(n_313), .C(n_316), .Y(n_312) );
INVxp67_ASAP7_75t_L g517 ( .A(n_72), .Y(n_517) );
INVx1_ASAP7_75t_L g513 ( .A(n_73), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_74), .B(n_219), .Y(n_257) );
INVx1_ASAP7_75t_L g91 ( .A(n_75), .Y(n_91) );
INVx1_ASAP7_75t_L g93 ( .A(n_75), .Y(n_93) );
INVx2_ASAP7_75t_L g267 ( .A(n_76), .Y(n_267) );
AOI221xp5_ASAP7_75t_L g77 ( .A1(n_78), .A2(n_175), .B1(n_183), .B2(n_501), .C(n_505), .Y(n_77) );
CKINVDCx20_ASAP7_75t_R g78 ( .A(n_79), .Y(n_78) );
OAI322xp33_ASAP7_75t_L g505 ( .A1(n_80), .A2(n_506), .A3(n_507), .B1(n_508), .B2(n_535), .C1(n_538), .C2(n_539), .Y(n_505) );
INVx1_ASAP7_75t_L g80 ( .A(n_81), .Y(n_80) );
NAND2xp5_ASAP7_75t_SL g81 ( .A(n_82), .B(n_139), .Y(n_81) );
INVxp67_ASAP7_75t_L g506 ( .A(n_82), .Y(n_506) );
NOR3xp33_ASAP7_75t_L g82 ( .A(n_83), .B(n_118), .C(n_131), .Y(n_82) );
NAND2xp5_ASAP7_75t_L g83 ( .A(n_84), .B(n_106), .Y(n_83) );
BUFx6f_ASAP7_75t_L g85 ( .A(n_86), .Y(n_85) );
BUFx6f_ASAP7_75t_L g86 ( .A(n_87), .Y(n_86) );
AND2x2_ASAP7_75t_L g87 ( .A(n_88), .B(n_97), .Y(n_87) );
AND2x6_ASAP7_75t_L g123 ( .A(n_88), .B(n_124), .Y(n_123) );
AND2x4_ASAP7_75t_L g134 ( .A(n_88), .B(n_113), .Y(n_134) );
AND2x6_ASAP7_75t_L g142 ( .A(n_88), .B(n_143), .Y(n_142) );
AND2x2_ASAP7_75t_L g88 ( .A(n_89), .B(n_94), .Y(n_88) );
AND2x2_ASAP7_75t_L g130 ( .A(n_89), .B(n_95), .Y(n_130) );
INVx2_ASAP7_75t_L g89 ( .A(n_90), .Y(n_89) );
NAND2xp5_ASAP7_75t_L g105 ( .A(n_90), .B(n_95), .Y(n_105) );
AND2x2_ASAP7_75t_L g111 ( .A(n_90), .B(n_112), .Y(n_111) );
AND2x2_ASAP7_75t_L g152 ( .A(n_90), .B(n_99), .Y(n_152) );
INVx1_ASAP7_75t_L g92 ( .A(n_93), .Y(n_92) );
INVx1_ASAP7_75t_L g96 ( .A(n_93), .Y(n_96) );
INVx1_ASAP7_75t_L g94 ( .A(n_95), .Y(n_94) );
INVx1_ASAP7_75t_L g112 ( .A(n_95), .Y(n_112) );
INVx1_ASAP7_75t_L g151 ( .A(n_95), .Y(n_151) );
AND2x4_ASAP7_75t_L g103 ( .A(n_97), .B(n_104), .Y(n_103) );
AND2x4_ASAP7_75t_L g129 ( .A(n_97), .B(n_130), .Y(n_129) );
NAND2xp5_ASAP7_75t_L g138 ( .A(n_97), .B(n_111), .Y(n_138) );
AND2x2_ASAP7_75t_L g97 ( .A(n_98), .B(n_100), .Y(n_97) );
AND2x2_ASAP7_75t_L g113 ( .A(n_98), .B(n_101), .Y(n_113) );
OR2x2_ASAP7_75t_L g125 ( .A(n_98), .B(n_101), .Y(n_125) );
INVx2_ASAP7_75t_L g98 ( .A(n_99), .Y(n_98) );
AND2x2_ASAP7_75t_L g143 ( .A(n_99), .B(n_101), .Y(n_143) );
AND2x2_ASAP7_75t_L g150 ( .A(n_100), .B(n_151), .Y(n_150) );
INVx2_ASAP7_75t_L g100 ( .A(n_101), .Y(n_100) );
INVx1_ASAP7_75t_L g117 ( .A(n_101), .Y(n_117) );
BUFx2_ASAP7_75t_SL g102 ( .A(n_103), .Y(n_102) );
INVx1_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
OR2x6_ASAP7_75t_L g116 ( .A(n_105), .B(n_117), .Y(n_116) );
BUFx6f_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
INVx4_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
INVx8_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
AND2x2_ASAP7_75t_L g110 ( .A(n_111), .B(n_113), .Y(n_110) );
INVx1_ASAP7_75t_L g167 ( .A(n_112), .Y(n_167) );
AND2x6_ASAP7_75t_L g173 ( .A(n_113), .B(n_130), .Y(n_173) );
BUFx2_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
INVx6_ASAP7_75t_SL g115 ( .A(n_116), .Y(n_115) );
INVx1_ASAP7_75t_L g162 ( .A(n_117), .Y(n_162) );
OAI22xp5_ASAP7_75t_L g118 ( .A1(n_119), .A2(n_120), .B1(n_126), .B2(n_127), .Y(n_118) );
INVx1_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
INVx5_ASAP7_75t_SL g121 ( .A(n_122), .Y(n_121) );
INVx11_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
AND2x4_ASAP7_75t_L g171 ( .A(n_124), .B(n_130), .Y(n_171) );
INVx2_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
INVx4_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
BUFx6f_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
OAI22xp5_ASAP7_75t_L g131 ( .A1(n_132), .A2(n_133), .B1(n_135), .B2(n_136), .Y(n_131) );
INVx6_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
INVx1_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
INVxp67_ASAP7_75t_L g507 ( .A(n_139), .Y(n_507) );
NOR2xp33_ASAP7_75t_L g139 ( .A(n_140), .B(n_157), .Y(n_139) );
OAI21xp5_ASAP7_75t_SL g140 ( .A1(n_141), .A2(n_144), .B(n_145), .Y(n_140) );
INVx2_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
AND2x4_ASAP7_75t_L g166 ( .A(n_143), .B(n_167), .Y(n_166) );
INVx3_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx4_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
BUFx6f_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
AND2x4_ASAP7_75t_L g149 ( .A(n_150), .B(n_152), .Y(n_149) );
INVx1_ASAP7_75t_L g156 ( .A(n_151), .Y(n_156) );
AND2x4_ASAP7_75t_L g155 ( .A(n_152), .B(n_156), .Y(n_155) );
AND2x4_ASAP7_75t_L g161 ( .A(n_152), .B(n_162), .Y(n_161) );
BUFx4f_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_158), .B(n_168), .Y(n_157) );
INVx1_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx2_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVx1_ASAP7_75t_SL g164 ( .A(n_165), .Y(n_164) );
BUFx6f_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
INVx2_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
INVx4_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
BUFx2_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
CKINVDCx20_ASAP7_75t_R g175 ( .A(n_176), .Y(n_175) );
OR2x2_ASAP7_75t_SL g176 ( .A(n_177), .B(n_181), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
AND3x1_ASAP7_75t_SL g523 ( .A(n_178), .B(n_181), .C(n_524), .Y(n_523) );
AND2x2_ASAP7_75t_L g531 ( .A(n_178), .B(n_532), .Y(n_531) );
OAI21xp5_ASAP7_75t_L g536 ( .A1(n_178), .A2(n_503), .B(n_537), .Y(n_536) );
INVx1_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
NAND2xp5_ASAP7_75t_SL g537 ( .A(n_179), .B(n_182), .Y(n_537) );
HB1xp67_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
CKINVDCx20_ASAP7_75t_R g181 ( .A(n_182), .Y(n_181) );
HB1xp67_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
OR5x1_ASAP7_75t_L g184 ( .A(n_185), .B(n_395), .C(n_459), .D(n_475), .E(n_490), .Y(n_184) );
NAND4xp25_ASAP7_75t_L g185 ( .A(n_186), .B(n_329), .C(n_356), .D(n_379), .Y(n_185) );
AOI21xp5_ASAP7_75t_L g186 ( .A1(n_187), .A2(n_272), .B(n_283), .Y(n_186) );
NOR2xp33_ASAP7_75t_L g187 ( .A(n_188), .B(n_221), .Y(n_187) );
HB1xp67_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
INVx3_ASAP7_75t_SL g306 ( .A(n_189), .Y(n_306) );
AND2x4_ASAP7_75t_L g342 ( .A(n_189), .B(n_331), .Y(n_342) );
OR2x2_ASAP7_75t_L g352 ( .A(n_189), .B(n_308), .Y(n_352) );
OR2x2_ASAP7_75t_L g398 ( .A(n_189), .B(n_224), .Y(n_398) );
AND2x2_ASAP7_75t_L g412 ( .A(n_189), .B(n_307), .Y(n_412) );
AND2x2_ASAP7_75t_L g455 ( .A(n_189), .B(n_345), .Y(n_455) );
AND2x2_ASAP7_75t_L g462 ( .A(n_189), .B(n_319), .Y(n_462) );
AND2x2_ASAP7_75t_L g481 ( .A(n_189), .B(n_371), .Y(n_481) );
AND2x2_ASAP7_75t_L g499 ( .A(n_189), .B(n_341), .Y(n_499) );
OR2x6_ASAP7_75t_L g189 ( .A(n_190), .B(n_216), .Y(n_189) );
O2A1O1Ixp33_ASAP7_75t_L g190 ( .A1(n_191), .A2(n_197), .B(n_198), .C(n_211), .Y(n_190) );
OAI21xp5_ASAP7_75t_L g291 ( .A1(n_191), .A2(n_292), .B(n_293), .Y(n_291) );
OAI21xp5_ASAP7_75t_L g310 ( .A1(n_191), .A2(n_311), .B(n_312), .Y(n_310) );
NAND2x1p5_ASAP7_75t_L g191 ( .A(n_192), .B(n_196), .Y(n_191) );
AND2x4_ASAP7_75t_L g231 ( .A(n_192), .B(n_196), .Y(n_231) );
AND2x2_ASAP7_75t_L g192 ( .A(n_193), .B(n_195), .Y(n_192) );
INVx1_ASAP7_75t_L g209 ( .A(n_193), .Y(n_209) );
INVx1_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
INVx2_ASAP7_75t_L g200 ( .A(n_194), .Y(n_200) );
INVx1_ASAP7_75t_L g269 ( .A(n_194), .Y(n_269) );
INVx1_ASAP7_75t_L g201 ( .A(n_195), .Y(n_201) );
INVx3_ASAP7_75t_L g205 ( .A(n_195), .Y(n_205) );
BUFx6f_ASAP7_75t_L g207 ( .A(n_195), .Y(n_207) );
BUFx6f_ASAP7_75t_L g240 ( .A(n_195), .Y(n_240) );
BUFx3_ASAP7_75t_L g210 ( .A(n_196), .Y(n_210) );
INVx4_ASAP7_75t_SL g241 ( .A(n_196), .Y(n_241) );
INVx5_ASAP7_75t_L g234 ( .A(n_199), .Y(n_234) );
AND2x6_ASAP7_75t_L g199 ( .A(n_200), .B(n_201), .Y(n_199) );
BUFx3_ASAP7_75t_L g256 ( .A(n_200), .Y(n_256) );
BUFx6f_ASAP7_75t_L g327 ( .A(n_200), .Y(n_327) );
O2A1O1Ixp33_ASAP7_75t_L g202 ( .A1(n_203), .A2(n_204), .B(n_206), .C(n_208), .Y(n_202) );
OAI22xp33_ASAP7_75t_L g236 ( .A1(n_204), .A2(n_237), .B1(n_238), .B2(n_239), .Y(n_236) );
INVx5_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
NOR2xp33_ASAP7_75t_L g253 ( .A(n_205), .B(n_254), .Y(n_253) );
INVx2_ASAP7_75t_L g252 ( .A(n_207), .Y(n_252) );
INVx4_ASAP7_75t_L g265 ( .A(n_207), .Y(n_265) );
NOR2xp33_ASAP7_75t_L g503 ( .A(n_208), .B(n_504), .Y(n_503) );
INVx2_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
NAND2xp5_ASAP7_75t_SL g235 ( .A(n_209), .B(n_236), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_210), .B(n_503), .Y(n_502) );
INVx2_ASAP7_75t_L g245 ( .A(n_211), .Y(n_245) );
OA21x2_ASAP7_75t_L g247 ( .A1(n_211), .A2(n_248), .B(n_257), .Y(n_247) );
INVx1_ASAP7_75t_L g290 ( .A(n_211), .Y(n_290) );
AND2x2_ASAP7_75t_SL g211 ( .A(n_212), .B(n_213), .Y(n_211) );
AND2x2_ASAP7_75t_L g220 ( .A(n_212), .B(n_213), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_214), .B(n_215), .Y(n_213) );
NOR2xp33_ASAP7_75t_L g216 ( .A(n_217), .B(n_218), .Y(n_216) );
INVx3_ASAP7_75t_L g271 ( .A(n_218), .Y(n_271) );
NOR2xp33_ASAP7_75t_L g300 ( .A(n_218), .B(n_301), .Y(n_300) );
AO21x2_ASAP7_75t_L g309 ( .A1(n_218), .A2(n_310), .B(n_317), .Y(n_309) );
INVx4_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
HB1xp67_ASAP7_75t_L g260 ( .A(n_219), .Y(n_260) );
BUFx6f_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
INVx1_ASAP7_75t_L g227 ( .A(n_220), .Y(n_227) );
INVx1_ASAP7_75t_L g464 ( .A(n_221), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_222), .B(n_246), .Y(n_221) );
AND2x2_ASAP7_75t_L g374 ( .A(n_222), .B(n_307), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_222), .B(n_394), .Y(n_393) );
AOI32xp33_ASAP7_75t_L g407 ( .A1(n_222), .A2(n_408), .A3(n_411), .B1(n_413), .B2(n_417), .Y(n_407) );
AND2x2_ASAP7_75t_L g477 ( .A(n_222), .B(n_371), .Y(n_477) );
INVx2_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
INVx1_ASAP7_75t_SL g223 ( .A(n_224), .Y(n_223) );
AND2x2_ASAP7_75t_L g341 ( .A(n_224), .B(n_308), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_224), .B(n_351), .Y(n_350) );
AND2x2_ASAP7_75t_L g383 ( .A(n_224), .B(n_330), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_224), .B(n_462), .Y(n_461) );
AO21x2_ASAP7_75t_L g224 ( .A1(n_225), .A2(n_228), .B(n_242), .Y(n_224) );
INVx1_ASAP7_75t_L g346 ( .A(n_225), .Y(n_346) );
INVx1_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
INVx2_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
INVx1_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
OA21x2_ASAP7_75t_L g345 ( .A1(n_229), .A2(n_243), .B(n_346), .Y(n_345) );
BUFx2_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
O2A1O1Ixp33_ASAP7_75t_SL g232 ( .A1(n_233), .A2(n_234), .B(n_235), .C(n_241), .Y(n_232) );
O2A1O1Ixp33_ASAP7_75t_SL g249 ( .A1(n_234), .A2(n_241), .B(n_250), .C(n_251), .Y(n_249) );
O2A1O1Ixp33_ASAP7_75t_SL g262 ( .A1(n_234), .A2(n_241), .B(n_263), .C(n_264), .Y(n_262) );
O2A1O1Ixp33_ASAP7_75t_SL g276 ( .A1(n_234), .A2(n_241), .B(n_277), .C(n_278), .Y(n_276) );
O2A1O1Ixp33_ASAP7_75t_L g321 ( .A1(n_234), .A2(n_241), .B(n_322), .C(n_323), .Y(n_321) );
NOR2xp33_ASAP7_75t_L g266 ( .A(n_239), .B(n_267), .Y(n_266) );
NOR2xp33_ASAP7_75t_L g279 ( .A(n_239), .B(n_280), .Y(n_279) );
INVx4_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
INVx2_ASAP7_75t_L g297 ( .A(n_240), .Y(n_297) );
INVx1_ASAP7_75t_L g316 ( .A(n_241), .Y(n_316) );
INVx1_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
INVx1_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
NOR2xp33_ASAP7_75t_L g317 ( .A(n_245), .B(n_318), .Y(n_317) );
AND2x2_ASAP7_75t_L g348 ( .A(n_246), .B(n_287), .Y(n_348) );
AND2x2_ASAP7_75t_L g424 ( .A(n_246), .B(n_425), .Y(n_424) );
INVx1_ASAP7_75t_SL g496 ( .A(n_246), .Y(n_496) );
AND2x2_ASAP7_75t_L g246 ( .A(n_247), .B(n_258), .Y(n_246) );
OR2x2_ASAP7_75t_L g286 ( .A(n_247), .B(n_259), .Y(n_286) );
AND2x2_ASAP7_75t_L g303 ( .A(n_247), .B(n_304), .Y(n_303) );
NOR2xp33_ASAP7_75t_L g333 ( .A(n_247), .B(n_334), .Y(n_333) );
INVx2_ASAP7_75t_L g355 ( .A(n_247), .Y(n_355) );
AND2x2_ASAP7_75t_L g382 ( .A(n_247), .B(n_259), .Y(n_382) );
BUFx3_ASAP7_75t_L g385 ( .A(n_247), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_247), .B(n_360), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_247), .B(n_479), .Y(n_478) );
INVx2_ASAP7_75t_L g299 ( .A(n_255), .Y(n_299) );
INVx2_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
INVx1_ASAP7_75t_L g281 ( .A(n_256), .Y(n_281) );
INVx2_ASAP7_75t_L g336 ( .A(n_258), .Y(n_336) );
AND2x2_ASAP7_75t_L g354 ( .A(n_258), .B(n_334), .Y(n_354) );
INVx2_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
AND2x2_ASAP7_75t_L g365 ( .A(n_259), .B(n_274), .Y(n_365) );
HB1xp67_ASAP7_75t_L g378 ( .A(n_259), .Y(n_378) );
OA21x2_ASAP7_75t_L g259 ( .A1(n_260), .A2(n_261), .B(n_270), .Y(n_259) );
OA21x2_ASAP7_75t_L g274 ( .A1(n_260), .A2(n_275), .B(n_282), .Y(n_274) );
OA21x2_ASAP7_75t_L g319 ( .A1(n_260), .A2(n_320), .B(n_328), .Y(n_319) );
NOR2xp33_ASAP7_75t_L g324 ( .A(n_265), .B(n_325), .Y(n_324) );
INVx3_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
INVx1_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_273), .B(n_385), .Y(n_435) );
HB1xp67_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
INVx1_ASAP7_75t_SL g304 ( .A(n_274), .Y(n_304) );
NAND3xp33_ASAP7_75t_L g353 ( .A(n_274), .B(n_354), .C(n_355), .Y(n_353) );
OR2x2_ASAP7_75t_L g361 ( .A(n_274), .B(n_334), .Y(n_361) );
AND2x2_ASAP7_75t_L g381 ( .A(n_274), .B(n_334), .Y(n_381) );
AND2x2_ASAP7_75t_L g425 ( .A(n_274), .B(n_289), .Y(n_425) );
AOI21xp5_ASAP7_75t_L g283 ( .A1(n_284), .A2(n_302), .B(n_305), .Y(n_283) );
NAND2xp5_ASAP7_75t_SL g284 ( .A(n_285), .B(n_287), .Y(n_284) );
AND2x2_ASAP7_75t_L g500 ( .A(n_285), .B(n_425), .Y(n_500) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
OAI22xp5_ASAP7_75t_L g439 ( .A1(n_286), .A2(n_398), .B1(n_440), .B2(n_442), .Y(n_439) );
OR2x2_ASAP7_75t_L g446 ( .A(n_286), .B(n_361), .Y(n_446) );
OR2x2_ASAP7_75t_L g470 ( .A(n_286), .B(n_471), .Y(n_470) );
NOR2xp33_ASAP7_75t_L g483 ( .A(n_286), .B(n_390), .Y(n_483) );
AND2x2_ASAP7_75t_L g376 ( .A(n_287), .B(n_377), .Y(n_376) );
AOI21xp5_ASAP7_75t_L g463 ( .A1(n_287), .A2(n_449), .B(n_464), .Y(n_463) );
AOI32xp33_ASAP7_75t_L g484 ( .A1(n_287), .A2(n_374), .A3(n_485), .B1(n_487), .B2(n_488), .Y(n_484) );
OR2x2_ASAP7_75t_L g495 ( .A(n_287), .B(n_496), .Y(n_495) );
CKINVDCx16_ASAP7_75t_R g287 ( .A(n_288), .Y(n_287) );
OR2x2_ASAP7_75t_L g363 ( .A(n_288), .B(n_364), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_288), .B(n_377), .Y(n_442) );
BUFx3_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
INVx4_ASAP7_75t_L g334 ( .A(n_289), .Y(n_334) );
AND2x2_ASAP7_75t_L g400 ( .A(n_289), .B(n_365), .Y(n_400) );
AND3x2_ASAP7_75t_L g409 ( .A(n_289), .B(n_303), .C(n_410), .Y(n_409) );
AO21x2_ASAP7_75t_L g289 ( .A1(n_290), .A2(n_291), .B(n_300), .Y(n_289) );
O2A1O1Ixp5_ASAP7_75t_L g294 ( .A1(n_295), .A2(n_296), .B(n_298), .C(n_299), .Y(n_294) );
O2A1O1Ixp33_ASAP7_75t_L g313 ( .A1(n_296), .A2(n_299), .B(n_314), .C(n_315), .Y(n_313) );
HB1xp67_ASAP7_75t_L g504 ( .A(n_296), .Y(n_504) );
INVx2_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
AND2x2_ASAP7_75t_L g335 ( .A(n_304), .B(n_336), .Y(n_335) );
HB1xp67_ASAP7_75t_L g390 ( .A(n_304), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_304), .B(n_334), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_306), .B(n_307), .Y(n_305) );
AND2x2_ASAP7_75t_L g330 ( .A(n_306), .B(n_331), .Y(n_330) );
AND2x2_ASAP7_75t_L g370 ( .A(n_306), .B(n_371), .Y(n_370) );
AND2x2_ASAP7_75t_L g388 ( .A(n_306), .B(n_319), .Y(n_388) );
AND2x2_ASAP7_75t_L g406 ( .A(n_306), .B(n_308), .Y(n_406) );
OR2x2_ASAP7_75t_L g420 ( .A(n_306), .B(n_421), .Y(n_420) );
AND2x2_ASAP7_75t_L g466 ( .A(n_306), .B(n_394), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_307), .B(n_345), .Y(n_344) );
AND2x2_ASAP7_75t_L g307 ( .A(n_308), .B(n_319), .Y(n_307) );
AND2x2_ASAP7_75t_L g367 ( .A(n_308), .B(n_345), .Y(n_367) );
OR2x2_ASAP7_75t_L g421 ( .A(n_308), .B(n_345), .Y(n_421) );
AND2x2_ASAP7_75t_L g474 ( .A(n_308), .B(n_331), .Y(n_474) );
INVx2_ASAP7_75t_SL g308 ( .A(n_309), .Y(n_308) );
BUFx2_ASAP7_75t_L g372 ( .A(n_309), .Y(n_372) );
AND2x2_ASAP7_75t_L g394 ( .A(n_309), .B(n_319), .Y(n_394) );
INVx2_ASAP7_75t_L g331 ( .A(n_319), .Y(n_331) );
INVx1_ASAP7_75t_L g351 ( .A(n_319), .Y(n_351) );
INVx3_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
AOI211xp5_ASAP7_75t_L g329 ( .A1(n_330), .A2(n_332), .B(n_337), .C(n_349), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_330), .B(n_441), .Y(n_440) );
INVx1_ASAP7_75t_L g493 ( .A(n_330), .Y(n_493) );
AND2x2_ASAP7_75t_L g371 ( .A(n_331), .B(n_372), .Y(n_371) );
AND2x2_ASAP7_75t_L g332 ( .A(n_333), .B(n_335), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_334), .B(n_335), .Y(n_343) );
INVx1_ASAP7_75t_L g428 ( .A(n_334), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_334), .B(n_355), .Y(n_452) );
AND2x2_ASAP7_75t_L g468 ( .A(n_334), .B(n_382), .Y(n_468) );
NAND2xp5_ASAP7_75t_SL g450 ( .A(n_335), .B(n_451), .Y(n_450) );
INVx2_ASAP7_75t_L g359 ( .A(n_336), .Y(n_359) );
OAI22xp5_ASAP7_75t_L g337 ( .A1(n_338), .A2(n_343), .B1(n_344), .B2(n_347), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
NOR2xp33_ASAP7_75t_L g339 ( .A(n_340), .B(n_342), .Y(n_339) );
NOR2xp33_ASAP7_75t_L g492 ( .A(n_340), .B(n_493), .Y(n_492) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_341), .B(n_388), .Y(n_387) );
AND2x2_ASAP7_75t_L g366 ( .A(n_342), .B(n_367), .Y(n_366) );
AOI221xp5_ASAP7_75t_SL g431 ( .A1(n_342), .A2(n_384), .B1(n_432), .B2(n_437), .C(n_439), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_342), .B(n_405), .Y(n_438) );
INVx1_ASAP7_75t_L g498 ( .A(n_344), .Y(n_498) );
BUFx3_ASAP7_75t_L g405 ( .A(n_345), .Y(n_405) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
AOI21xp33_ASAP7_75t_SL g349 ( .A1(n_350), .A2(n_352), .B(n_353), .Y(n_349) );
INVx1_ASAP7_75t_L g414 ( .A(n_351), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_351), .B(n_405), .Y(n_458) );
INVx1_ASAP7_75t_L g415 ( .A(n_352), .Y(n_415) );
NAND2xp5_ASAP7_75t_SL g416 ( .A(n_352), .B(n_405), .Y(n_416) );
INVxp67_ASAP7_75t_L g436 ( .A(n_354), .Y(n_436) );
AND2x2_ASAP7_75t_L g377 ( .A(n_355), .B(n_378), .Y(n_377) );
O2A1O1Ixp33_ASAP7_75t_L g356 ( .A1(n_357), .A2(n_362), .B(n_366), .C(n_368), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_359), .B(n_360), .Y(n_358) );
INVx1_ASAP7_75t_SL g391 ( .A(n_359), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_360), .B(n_391), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_360), .B(n_382), .Y(n_433) );
INVx2_ASAP7_75t_SL g360 ( .A(n_361), .Y(n_360) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
OAI22xp5_ASAP7_75t_L g368 ( .A1(n_363), .A2(n_369), .B1(n_373), .B2(n_375), .Y(n_368) );
INVx1_ASAP7_75t_SL g364 ( .A(n_365), .Y(n_364) );
AND2x2_ASAP7_75t_L g384 ( .A(n_365), .B(n_385), .Y(n_384) );
AND2x2_ASAP7_75t_L g429 ( .A(n_365), .B(n_430), .Y(n_429) );
OAI21xp33_ASAP7_75t_L g432 ( .A1(n_367), .A2(n_433), .B(n_434), .Y(n_432) );
INVx1_ASAP7_75t_SL g369 ( .A(n_370), .Y(n_369) );
AOI221xp5_ASAP7_75t_L g379 ( .A1(n_371), .A2(n_380), .B1(n_383), .B2(n_384), .C(n_386), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_371), .B(n_405), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_371), .B(n_455), .Y(n_454) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g487 ( .A(n_377), .Y(n_487) );
INVxp67_ASAP7_75t_L g410 ( .A(n_378), .Y(n_410) );
INVx1_ASAP7_75t_L g417 ( .A(n_380), .Y(n_417) );
AND2x2_ASAP7_75t_L g380 ( .A(n_381), .B(n_382), .Y(n_380) );
AND2x2_ASAP7_75t_L g456 ( .A(n_381), .B(n_385), .Y(n_456) );
INVx1_ASAP7_75t_L g430 ( .A(n_385), .Y(n_430) );
NAND2xp5_ASAP7_75t_SL g460 ( .A(n_385), .B(n_400), .Y(n_460) );
OAI32xp33_ASAP7_75t_L g386 ( .A1(n_387), .A2(n_389), .A3(n_391), .B1(n_392), .B2(n_393), .Y(n_386) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVx2_ASAP7_75t_SL g399 ( .A(n_394), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_394), .B(n_426), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_394), .B(n_455), .Y(n_486) );
NAND2x1p5_ASAP7_75t_L g494 ( .A(n_394), .B(n_405), .Y(n_494) );
NAND5xp2_ASAP7_75t_L g395 ( .A(n_396), .B(n_418), .C(n_431), .D(n_443), .E(n_444), .Y(n_395) );
AOI221xp5_ASAP7_75t_L g396 ( .A1(n_397), .A2(n_400), .B1(n_401), .B2(n_403), .C(n_407), .Y(n_396) );
NOR2xp33_ASAP7_75t_L g397 ( .A(n_398), .B(n_399), .Y(n_397) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
NAND2xp33_ASAP7_75t_SL g422 ( .A(n_402), .B(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_405), .B(n_406), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_405), .B(n_474), .Y(n_473) );
AOI22xp33_ASAP7_75t_L g418 ( .A1(n_406), .A2(n_419), .B1(n_422), .B2(n_426), .Y(n_418) );
INVx2_ASAP7_75t_SL g408 ( .A(n_409), .Y(n_408) );
OAI211xp5_ASAP7_75t_SL g413 ( .A1(n_409), .A2(n_414), .B(n_415), .C(n_416), .Y(n_413) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx1_ASAP7_75t_SL g441 ( .A(n_421), .Y(n_441) );
INVx1_ASAP7_75t_SL g423 ( .A(n_424), .Y(n_423) );
INVx1_ASAP7_75t_SL g426 ( .A(n_427), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_428), .B(n_429), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_430), .B(n_479), .Y(n_489) );
OR2x2_ASAP7_75t_L g434 ( .A(n_435), .B(n_436), .Y(n_434) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
AOI222xp33_ASAP7_75t_L g444 ( .A1(n_445), .A2(n_447), .B1(n_449), .B2(n_453), .C1(n_456), .C2(n_457), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
OAI221xp5_ASAP7_75t_L g459 ( .A1(n_460), .A2(n_461), .B1(n_463), .B2(n_465), .C(n_467), .Y(n_459) );
INVx1_ASAP7_75t_SL g465 ( .A(n_466), .Y(n_465) );
OAI21xp33_ASAP7_75t_L g467 ( .A1(n_468), .A2(n_469), .B(n_472), .Y(n_467) );
INVx2_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
INVx1_ASAP7_75t_L g479 ( .A(n_471), .Y(n_479) );
INVx1_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
OAI221xp5_ASAP7_75t_L g475 ( .A1(n_476), .A2(n_478), .B1(n_480), .B2(n_482), .C(n_484), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
INVx1_ASAP7_75t_SL g480 ( .A(n_481), .Y(n_480) );
INVxp67_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
INVx1_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
INVx1_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
A2O1A1Ixp33_ASAP7_75t_L g490 ( .A1(n_491), .A2(n_494), .B(n_495), .C(n_497), .Y(n_490) );
INVxp67_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
OAI21xp33_ASAP7_75t_L g497 ( .A1(n_498), .A2(n_499), .B(n_500), .Y(n_497) );
CKINVDCx20_ASAP7_75t_R g501 ( .A(n_502), .Y(n_501) );
CKINVDCx20_ASAP7_75t_R g509 ( .A(n_510), .Y(n_509) );
AOI22xp5_ASAP7_75t_L g539 ( .A1(n_510), .A2(n_521), .B1(n_531), .B2(n_540), .Y(n_539) );
AOI22xp5_ASAP7_75t_L g510 ( .A1(n_511), .A2(n_514), .B1(n_519), .B2(n_520), .Y(n_510) );
CKINVDCx20_ASAP7_75t_R g519 ( .A(n_511), .Y(n_519) );
CKINVDCx20_ASAP7_75t_R g520 ( .A(n_514), .Y(n_520) );
INVx1_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
CKINVDCx20_ASAP7_75t_R g521 ( .A(n_522), .Y(n_521) );
CKINVDCx20_ASAP7_75t_R g522 ( .A(n_523), .Y(n_522) );
INVxp67_ASAP7_75t_L g534 ( .A(n_524), .Y(n_534) );
NOR2xp33_ASAP7_75t_L g526 ( .A(n_527), .B(n_528), .Y(n_526) );
CKINVDCx16_ASAP7_75t_R g529 ( .A(n_530), .Y(n_529) );
CKINVDCx20_ASAP7_75t_R g530 ( .A(n_531), .Y(n_530) );
CKINVDCx20_ASAP7_75t_R g532 ( .A(n_533), .Y(n_532) );
CKINVDCx16_ASAP7_75t_R g535 ( .A(n_536), .Y(n_535) );
endmodule