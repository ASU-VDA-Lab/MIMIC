module real_aes_7617_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_357;
wire n_287;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_725;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_527;
wire n_505;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_552;
wire n_602;
wire n_617;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_101;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_741;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g183 ( .A1(n_0), .A2(n_184), .B(n_185), .C(n_189), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_1), .B(n_179), .Y(n_190) );
NAND3xp33_ASAP7_75t_SL g104 ( .A(n_2), .B(n_105), .C(n_106), .Y(n_104) );
INVx1_ASAP7_75t_L g440 ( .A(n_2), .Y(n_440) );
NAND2xp5_ASAP7_75t_SL g261 ( .A(n_3), .B(n_144), .Y(n_261) );
AOI21xp5_ASAP7_75t_L g472 ( .A1(n_4), .A2(n_125), .B(n_473), .Y(n_472) );
A2O1A1Ixp33_ASAP7_75t_L g508 ( .A1(n_5), .A2(n_130), .B(n_135), .C(n_509), .Y(n_508) );
AOI21xp5_ASAP7_75t_L g229 ( .A1(n_6), .A2(n_125), .B(n_230), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_7), .B(n_179), .Y(n_479) );
AO21x2_ASAP7_75t_L g207 ( .A1(n_8), .A2(n_158), .B(n_208), .Y(n_207) );
AND2x6_ASAP7_75t_L g130 ( .A(n_9), .B(n_131), .Y(n_130) );
A2O1A1Ixp33_ASAP7_75t_L g197 ( .A1(n_10), .A2(n_130), .B(n_135), .C(n_198), .Y(n_197) );
INVx1_ASAP7_75t_L g534 ( .A(n_11), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g103 ( .A(n_12), .B(n_40), .Y(n_103) );
NOR2xp33_ASAP7_75t_L g441 ( .A(n_12), .B(n_40), .Y(n_441) );
NAND2xp5_ASAP7_75t_SL g511 ( .A(n_13), .B(n_188), .Y(n_511) );
INVx1_ASAP7_75t_L g154 ( .A(n_14), .Y(n_154) );
NAND2xp5_ASAP7_75t_SL g214 ( .A(n_15), .B(n_144), .Y(n_214) );
A2O1A1Ixp33_ASAP7_75t_L g518 ( .A1(n_16), .A2(n_145), .B(n_519), .C(n_521), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_17), .B(n_179), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_18), .B(n_172), .Y(n_563) );
A2O1A1Ixp33_ASAP7_75t_L g165 ( .A1(n_19), .A2(n_135), .B(n_166), .C(n_171), .Y(n_165) );
A2O1A1Ixp33_ASAP7_75t_L g498 ( .A1(n_20), .A2(n_187), .B(n_202), .C(n_499), .Y(n_498) );
NAND2xp5_ASAP7_75t_SL g464 ( .A(n_21), .B(n_188), .Y(n_464) );
OAI222xp33_ASAP7_75t_L g445 ( .A1(n_22), .A2(n_446), .B1(n_727), .B2(n_728), .C1(n_734), .C2(n_738), .Y(n_445) );
CKINVDCx20_ASAP7_75t_R g727 ( .A(n_22), .Y(n_727) );
NAND2xp5_ASAP7_75t_SL g486 ( .A(n_23), .B(n_188), .Y(n_486) );
CKINVDCx16_ASAP7_75t_R g460 ( .A(n_24), .Y(n_460) );
INVx1_ASAP7_75t_L g485 ( .A(n_25), .Y(n_485) );
A2O1A1Ixp33_ASAP7_75t_L g210 ( .A1(n_26), .A2(n_135), .B(n_171), .C(n_211), .Y(n_210) );
BUFx6f_ASAP7_75t_L g129 ( .A(n_27), .Y(n_129) );
CKINVDCx20_ASAP7_75t_R g507 ( .A(n_28), .Y(n_507) );
CKINVDCx20_ASAP7_75t_R g738 ( .A(n_29), .Y(n_738) );
INVx1_ASAP7_75t_L g561 ( .A(n_30), .Y(n_561) );
AOI21xp5_ASAP7_75t_L g180 ( .A1(n_31), .A2(n_125), .B(n_181), .Y(n_180) );
INVx2_ASAP7_75t_L g128 ( .A(n_32), .Y(n_128) );
A2O1A1Ixp33_ASAP7_75t_L g132 ( .A1(n_33), .A2(n_133), .B(n_138), .C(n_148), .Y(n_132) );
CKINVDCx20_ASAP7_75t_R g513 ( .A(n_34), .Y(n_513) );
A2O1A1Ixp33_ASAP7_75t_L g475 ( .A1(n_35), .A2(n_187), .B(n_476), .C(n_478), .Y(n_475) );
INVxp67_ASAP7_75t_L g562 ( .A(n_36), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_37), .B(n_213), .Y(n_212) );
CKINVDCx14_ASAP7_75t_R g474 ( .A(n_38), .Y(n_474) );
A2O1A1Ixp33_ASAP7_75t_L g483 ( .A1(n_39), .A2(n_135), .B(n_171), .C(n_484), .Y(n_483) );
A2O1A1Ixp33_ASAP7_75t_L g531 ( .A1(n_41), .A2(n_189), .B(n_532), .C(n_533), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_42), .B(n_164), .Y(n_163) );
CKINVDCx20_ASAP7_75t_R g205 ( .A(n_43), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_44), .B(n_144), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_45), .B(n_125), .Y(n_209) );
CKINVDCx20_ASAP7_75t_R g488 ( .A(n_46), .Y(n_488) );
CKINVDCx20_ASAP7_75t_R g443 ( .A(n_47), .Y(n_443) );
CKINVDCx20_ASAP7_75t_R g558 ( .A(n_48), .Y(n_558) );
A2O1A1Ixp33_ASAP7_75t_L g221 ( .A1(n_49), .A2(n_133), .B(n_148), .C(n_222), .Y(n_221) );
OAI22xp5_ASAP7_75t_L g115 ( .A1(n_50), .A2(n_116), .B1(n_117), .B2(n_435), .Y(n_115) );
CKINVDCx20_ASAP7_75t_R g116 ( .A(n_50), .Y(n_116) );
INVx1_ASAP7_75t_L g186 ( .A(n_51), .Y(n_186) );
INVx1_ASAP7_75t_L g223 ( .A(n_52), .Y(n_223) );
INVx1_ASAP7_75t_L g497 ( .A(n_53), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_54), .B(n_125), .Y(n_220) );
CKINVDCx20_ASAP7_75t_R g175 ( .A(n_55), .Y(n_175) );
CKINVDCx14_ASAP7_75t_R g530 ( .A(n_56), .Y(n_530) );
INVx1_ASAP7_75t_L g131 ( .A(n_57), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_58), .B(n_125), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_59), .B(n_179), .Y(n_237) );
A2O1A1Ixp33_ASAP7_75t_L g232 ( .A1(n_60), .A2(n_170), .B(n_233), .C(n_235), .Y(n_232) );
INVx1_ASAP7_75t_L g153 ( .A(n_61), .Y(n_153) );
INVx1_ASAP7_75t_SL g477 ( .A(n_62), .Y(n_477) );
CKINVDCx20_ASAP7_75t_R g113 ( .A(n_63), .Y(n_113) );
NAND2xp5_ASAP7_75t_SL g143 ( .A(n_64), .B(n_144), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_65), .B(n_179), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_66), .B(n_145), .Y(n_199) );
INVx1_ASAP7_75t_L g463 ( .A(n_67), .Y(n_463) );
CKINVDCx16_ASAP7_75t_R g182 ( .A(n_68), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_69), .B(n_141), .Y(n_167) );
A2O1A1Ixp33_ASAP7_75t_L g258 ( .A1(n_70), .A2(n_135), .B(n_148), .C(n_259), .Y(n_258) );
CKINVDCx16_ASAP7_75t_R g231 ( .A(n_71), .Y(n_231) );
INVx1_ASAP7_75t_L g108 ( .A(n_72), .Y(n_108) );
AOI21xp5_ASAP7_75t_L g528 ( .A1(n_73), .A2(n_125), .B(n_529), .Y(n_528) );
AOI22xp33_ASAP7_75t_L g99 ( .A1(n_74), .A2(n_100), .B1(n_109), .B2(n_741), .Y(n_99) );
CKINVDCx20_ASAP7_75t_R g467 ( .A(n_75), .Y(n_467) );
AOI21xp5_ASAP7_75t_L g515 ( .A1(n_76), .A2(n_125), .B(n_516), .Y(n_515) );
AOI21xp5_ASAP7_75t_L g556 ( .A1(n_77), .A2(n_164), .B(n_557), .Y(n_556) );
CKINVDCx16_ASAP7_75t_R g482 ( .A(n_78), .Y(n_482) );
INVx1_ASAP7_75t_L g517 ( .A(n_79), .Y(n_517) );
NAND2xp5_ASAP7_75t_SL g168 ( .A(n_80), .B(n_140), .Y(n_168) );
CKINVDCx20_ASAP7_75t_R g156 ( .A(n_81), .Y(n_156) );
AOI21xp5_ASAP7_75t_L g495 ( .A1(n_82), .A2(n_125), .B(n_496), .Y(n_495) );
INVx1_ASAP7_75t_L g520 ( .A(n_83), .Y(n_520) );
INVx2_ASAP7_75t_L g151 ( .A(n_84), .Y(n_151) );
INVx1_ASAP7_75t_L g510 ( .A(n_85), .Y(n_510) );
CKINVDCx20_ASAP7_75t_R g266 ( .A(n_86), .Y(n_266) );
NAND2xp5_ASAP7_75t_SL g200 ( .A(n_87), .B(n_188), .Y(n_200) );
INVx2_ASAP7_75t_L g105 ( .A(n_88), .Y(n_105) );
OR2x2_ASAP7_75t_L g437 ( .A(n_88), .B(n_438), .Y(n_437) );
OR2x2_ASAP7_75t_L g448 ( .A(n_88), .B(n_439), .Y(n_448) );
A2O1A1Ixp33_ASAP7_75t_L g461 ( .A1(n_89), .A2(n_135), .B(n_148), .C(n_462), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g124 ( .A(n_90), .B(n_125), .Y(n_124) );
INVx1_ASAP7_75t_L g139 ( .A(n_91), .Y(n_139) );
INVxp67_ASAP7_75t_L g236 ( .A(n_92), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_93), .B(n_158), .Y(n_535) );
INVx2_ASAP7_75t_L g500 ( .A(n_94), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g107 ( .A(n_95), .B(n_108), .Y(n_107) );
INVx1_ASAP7_75t_L g195 ( .A(n_96), .Y(n_195) );
INVx1_ASAP7_75t_L g260 ( .A(n_97), .Y(n_260) );
AND2x2_ASAP7_75t_L g225 ( .A(n_98), .B(n_150), .Y(n_225) );
INVx1_ASAP7_75t_SL g100 ( .A(n_101), .Y(n_100) );
INVx1_ASAP7_75t_L g742 ( .A(n_101), .Y(n_742) );
INVx1_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
NOR2xp33_ASAP7_75t_L g102 ( .A(n_103), .B(n_104), .Y(n_102) );
OR2x2_ASAP7_75t_L g450 ( .A(n_105), .B(n_439), .Y(n_450) );
NOR2x2_ASAP7_75t_L g737 ( .A(n_105), .B(n_438), .Y(n_737) );
INVx1_ASAP7_75t_SL g106 ( .A(n_107), .Y(n_106) );
OAI21x1_ASAP7_75t_SL g109 ( .A1(n_110), .A2(n_114), .B(n_444), .Y(n_109) );
BUFx2_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
BUFx2_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
INVx2_ASAP7_75t_SL g740 ( .A(n_112), .Y(n_740) );
INVx2_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
AOI21xp5_ASAP7_75t_L g114 ( .A1(n_115), .A2(n_436), .B(n_442), .Y(n_114) );
INVx2_ASAP7_75t_L g435 ( .A(n_117), .Y(n_435) );
AOI22xp5_ASAP7_75t_L g728 ( .A1(n_117), .A2(n_729), .B1(n_732), .B2(n_733), .Y(n_728) );
OR3x2_ASAP7_75t_L g117 ( .A(n_118), .B(n_349), .C(n_392), .Y(n_117) );
NAND5xp2_ASAP7_75t_L g118 ( .A(n_119), .B(n_276), .C(n_306), .D(n_323), .E(n_338), .Y(n_118) );
AOI221xp5_ASAP7_75t_SL g119 ( .A1(n_120), .A2(n_191), .B1(n_238), .B2(n_244), .C(n_248), .Y(n_119) );
AND2x2_ASAP7_75t_L g120 ( .A(n_121), .B(n_160), .Y(n_120) );
OR2x2_ASAP7_75t_L g253 ( .A(n_121), .B(n_254), .Y(n_253) );
AND2x2_ASAP7_75t_L g293 ( .A(n_121), .B(n_294), .Y(n_293) );
AND2x2_ASAP7_75t_L g311 ( .A(n_121), .B(n_312), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_121), .B(n_246), .Y(n_328) );
OR2x2_ASAP7_75t_L g340 ( .A(n_121), .B(n_341), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_121), .B(n_299), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_121), .B(n_373), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_121), .B(n_277), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_121), .B(n_285), .Y(n_391) );
AND2x2_ASAP7_75t_L g423 ( .A(n_121), .B(n_177), .Y(n_423) );
HB1xp67_ASAP7_75t_L g431 ( .A(n_121), .Y(n_431) );
INVx5_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_122), .B(n_246), .Y(n_245) );
AND2x2_ASAP7_75t_L g250 ( .A(n_122), .B(n_226), .Y(n_250) );
BUFx2_ASAP7_75t_L g273 ( .A(n_122), .Y(n_273) );
AND2x2_ASAP7_75t_L g302 ( .A(n_122), .B(n_161), .Y(n_302) );
AND2x2_ASAP7_75t_L g357 ( .A(n_122), .B(n_254), .Y(n_357) );
OR2x6_ASAP7_75t_L g122 ( .A(n_123), .B(n_155), .Y(n_122) );
AOI21xp5_ASAP7_75t_L g123 ( .A1(n_124), .A2(n_132), .B(n_150), .Y(n_123) );
BUFx2_ASAP7_75t_L g164 ( .A(n_125), .Y(n_164) );
AND2x4_ASAP7_75t_L g125 ( .A(n_126), .B(n_130), .Y(n_125) );
NAND2x1p5_ASAP7_75t_L g196 ( .A(n_126), .B(n_130), .Y(n_196) );
AND2x2_ASAP7_75t_L g126 ( .A(n_127), .B(n_129), .Y(n_126) );
INVx1_ASAP7_75t_L g170 ( .A(n_127), .Y(n_170) );
INVx1_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
INVx2_ASAP7_75t_L g136 ( .A(n_128), .Y(n_136) );
INVx1_ASAP7_75t_L g203 ( .A(n_128), .Y(n_203) );
INVx1_ASAP7_75t_L g137 ( .A(n_129), .Y(n_137) );
BUFx6f_ASAP7_75t_L g142 ( .A(n_129), .Y(n_142) );
INVx3_ASAP7_75t_L g145 ( .A(n_129), .Y(n_145) );
BUFx6f_ASAP7_75t_L g188 ( .A(n_129), .Y(n_188) );
INVx1_ASAP7_75t_L g213 ( .A(n_129), .Y(n_213) );
INVx4_ASAP7_75t_SL g149 ( .A(n_130), .Y(n_149) );
BUFx3_ASAP7_75t_L g171 ( .A(n_130), .Y(n_171) );
INVx2_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
O2A1O1Ixp33_ASAP7_75t_SL g181 ( .A1(n_134), .A2(n_149), .B(n_182), .C(n_183), .Y(n_181) );
O2A1O1Ixp33_ASAP7_75t_L g230 ( .A1(n_134), .A2(n_149), .B(n_231), .C(n_232), .Y(n_230) );
O2A1O1Ixp33_ASAP7_75t_L g473 ( .A1(n_134), .A2(n_149), .B(n_474), .C(n_475), .Y(n_473) );
O2A1O1Ixp33_ASAP7_75t_SL g496 ( .A1(n_134), .A2(n_149), .B(n_497), .C(n_498), .Y(n_496) );
O2A1O1Ixp33_ASAP7_75t_SL g516 ( .A1(n_134), .A2(n_149), .B(n_517), .C(n_518), .Y(n_516) );
O2A1O1Ixp33_ASAP7_75t_SL g529 ( .A1(n_134), .A2(n_149), .B(n_530), .C(n_531), .Y(n_529) );
O2A1O1Ixp33_ASAP7_75t_SL g557 ( .A1(n_134), .A2(n_149), .B(n_558), .C(n_559), .Y(n_557) );
INVx5_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
AND2x6_ASAP7_75t_L g135 ( .A(n_136), .B(n_137), .Y(n_135) );
BUFx3_ASAP7_75t_L g147 ( .A(n_136), .Y(n_147) );
BUFx6f_ASAP7_75t_L g263 ( .A(n_136), .Y(n_263) );
O2A1O1Ixp33_ASAP7_75t_L g138 ( .A1(n_139), .A2(n_140), .B(n_143), .C(n_146), .Y(n_138) );
O2A1O1Ixp33_ASAP7_75t_L g222 ( .A1(n_140), .A2(n_146), .B(n_223), .C(n_224), .Y(n_222) );
O2A1O1Ixp33_ASAP7_75t_L g462 ( .A1(n_140), .A2(n_463), .B(n_464), .C(n_465), .Y(n_462) );
O2A1O1Ixp5_ASAP7_75t_L g509 ( .A1(n_140), .A2(n_465), .B(n_510), .C(n_511), .Y(n_509) );
INVx2_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx2_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
INVx4_ASAP7_75t_L g234 ( .A(n_142), .Y(n_234) );
INVx2_ASAP7_75t_L g184 ( .A(n_144), .Y(n_184) );
NOR2xp33_ASAP7_75t_L g235 ( .A(n_144), .B(n_236), .Y(n_235) );
O2A1O1Ixp33_ASAP7_75t_L g484 ( .A1(n_144), .A2(n_169), .B(n_485), .C(n_486), .Y(n_484) );
OAI22xp33_ASAP7_75t_L g560 ( .A1(n_144), .A2(n_234), .B1(n_561), .B2(n_562), .Y(n_560) );
INVx5_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
NOR2xp33_ASAP7_75t_L g533 ( .A(n_145), .B(n_534), .Y(n_533) );
HB1xp67_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx2_ASAP7_75t_L g189 ( .A(n_147), .Y(n_189) );
INVx1_ASAP7_75t_L g521 ( .A(n_147), .Y(n_521) );
INVx1_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx2_ASAP7_75t_L g173 ( .A(n_150), .Y(n_173) );
INVx1_ASAP7_75t_L g176 ( .A(n_150), .Y(n_176) );
AOI21xp5_ASAP7_75t_L g219 ( .A1(n_150), .A2(n_220), .B(n_221), .Y(n_219) );
O2A1O1Ixp33_ASAP7_75t_L g481 ( .A1(n_150), .A2(n_196), .B(n_482), .C(n_483), .Y(n_481) );
OA21x2_ASAP7_75t_L g527 ( .A1(n_150), .A2(n_528), .B(n_535), .Y(n_527) );
AND2x2_ASAP7_75t_SL g150 ( .A(n_151), .B(n_152), .Y(n_150) );
AND2x2_ASAP7_75t_L g159 ( .A(n_151), .B(n_152), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_153), .B(n_154), .Y(n_152) );
NOR2xp33_ASAP7_75t_L g155 ( .A(n_156), .B(n_157), .Y(n_155) );
INVx3_ASAP7_75t_L g179 ( .A(n_157), .Y(n_179) );
AO21x2_ASAP7_75t_L g193 ( .A1(n_157), .A2(n_194), .B(n_204), .Y(n_193) );
AO21x2_ASAP7_75t_L g256 ( .A1(n_157), .A2(n_257), .B(n_265), .Y(n_256) );
NOR2xp33_ASAP7_75t_L g265 ( .A(n_157), .B(n_266), .Y(n_265) );
AO21x2_ASAP7_75t_L g458 ( .A1(n_157), .A2(n_459), .B(n_466), .Y(n_458) );
NOR2xp33_ASAP7_75t_L g487 ( .A(n_157), .B(n_488), .Y(n_487) );
NOR2xp33_ASAP7_75t_L g512 ( .A(n_157), .B(n_513), .Y(n_512) );
INVx4_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
AOI21xp5_ASAP7_75t_L g208 ( .A1(n_158), .A2(n_209), .B(n_210), .Y(n_208) );
HB1xp67_ASAP7_75t_L g228 ( .A(n_158), .Y(n_228) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
INVx1_ASAP7_75t_L g206 ( .A(n_159), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_160), .B(n_311), .Y(n_320) );
OAI32xp33_ASAP7_75t_L g334 ( .A1(n_160), .A2(n_270), .A3(n_335), .B1(n_336), .B2(n_337), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_160), .B(n_336), .Y(n_366) );
NOR2xp33_ASAP7_75t_L g377 ( .A(n_160), .B(n_253), .Y(n_377) );
INVx1_ASAP7_75t_SL g406 ( .A(n_160), .Y(n_406) );
NAND4xp25_ASAP7_75t_L g415 ( .A(n_160), .B(n_193), .C(n_357), .D(n_416), .Y(n_415) );
AND2x4_ASAP7_75t_L g160 ( .A(n_161), .B(n_177), .Y(n_160) );
INVx5_ASAP7_75t_L g247 ( .A(n_161), .Y(n_247) );
AND2x2_ASAP7_75t_L g277 ( .A(n_161), .B(n_178), .Y(n_277) );
HB1xp67_ASAP7_75t_L g356 ( .A(n_161), .Y(n_356) );
AND2x2_ASAP7_75t_L g426 ( .A(n_161), .B(n_373), .Y(n_426) );
OR2x6_ASAP7_75t_L g161 ( .A(n_162), .B(n_174), .Y(n_161) );
AOI21xp5_ASAP7_75t_SL g162 ( .A1(n_163), .A2(n_165), .B(n_172), .Y(n_162) );
AOI21xp5_ASAP7_75t_L g166 ( .A1(n_167), .A2(n_168), .B(n_169), .Y(n_166) );
INVx2_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
NAND2xp5_ASAP7_75t_SL g559 ( .A(n_170), .B(n_560), .Y(n_559) );
INVx1_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
NOR2xp33_ASAP7_75t_L g466 ( .A(n_173), .B(n_467), .Y(n_466) );
NOR2xp33_ASAP7_75t_L g174 ( .A(n_175), .B(n_176), .Y(n_174) );
AO21x2_ASAP7_75t_L g505 ( .A1(n_176), .A2(n_506), .B(n_512), .Y(n_505) );
AND2x4_ASAP7_75t_L g299 ( .A(n_177), .B(n_247), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_177), .B(n_309), .Y(n_308) );
AND2x2_ASAP7_75t_L g333 ( .A(n_177), .B(n_254), .Y(n_333) );
INVx2_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
AND2x2_ASAP7_75t_L g246 ( .A(n_178), .B(n_247), .Y(n_246) );
AND2x2_ASAP7_75t_L g285 ( .A(n_178), .B(n_256), .Y(n_285) );
AND2x2_ASAP7_75t_L g294 ( .A(n_178), .B(n_255), .Y(n_294) );
OA21x2_ASAP7_75t_L g178 ( .A1(n_179), .A2(n_180), .B(n_190), .Y(n_178) );
NOR2xp33_ASAP7_75t_L g185 ( .A(n_186), .B(n_187), .Y(n_185) );
NOR2xp33_ASAP7_75t_L g476 ( .A(n_187), .B(n_477), .Y(n_476) );
INVx4_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
INVx2_ASAP7_75t_L g532 ( .A(n_188), .Y(n_532) );
INVx2_ASAP7_75t_L g465 ( .A(n_189), .Y(n_465) );
AOI222xp33_ASAP7_75t_L g362 ( .A1(n_191), .A2(n_363), .B1(n_365), .B2(n_367), .C1(n_370), .C2(n_371), .Y(n_362) );
AND2x4_ASAP7_75t_L g191 ( .A(n_192), .B(n_215), .Y(n_191) );
AND2x2_ASAP7_75t_L g295 ( .A(n_192), .B(n_296), .Y(n_295) );
NAND3xp33_ASAP7_75t_L g412 ( .A(n_192), .B(n_273), .C(n_413), .Y(n_412) );
AND2x2_ASAP7_75t_L g192 ( .A(n_193), .B(n_207), .Y(n_192) );
INVx5_ASAP7_75t_SL g243 ( .A(n_193), .Y(n_243) );
OAI322xp33_ASAP7_75t_L g248 ( .A1(n_193), .A2(n_249), .A3(n_251), .B1(n_252), .B2(n_267), .C1(n_270), .C2(n_272), .Y(n_248) );
NAND2xp5_ASAP7_75t_SL g315 ( .A(n_193), .B(n_241), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_193), .B(n_227), .Y(n_421) );
OAI21xp5_ASAP7_75t_L g194 ( .A1(n_195), .A2(n_196), .B(n_197), .Y(n_194) );
OAI21xp5_ASAP7_75t_L g459 ( .A1(n_196), .A2(n_460), .B(n_461), .Y(n_459) );
OAI21xp5_ASAP7_75t_L g506 ( .A1(n_196), .A2(n_507), .B(n_508), .Y(n_506) );
AOI21xp5_ASAP7_75t_L g198 ( .A1(n_199), .A2(n_200), .B(n_201), .Y(n_198) );
AOI21xp5_ASAP7_75t_L g211 ( .A1(n_201), .A2(n_212), .B(n_214), .Y(n_211) );
INVx2_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
INVx3_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
NOR2xp33_ASAP7_75t_L g204 ( .A(n_205), .B(n_206), .Y(n_204) );
INVx2_ASAP7_75t_L g555 ( .A(n_206), .Y(n_555) );
INVx2_ASAP7_75t_L g241 ( .A(n_207), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_207), .B(n_217), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_215), .B(n_280), .Y(n_335) );
INVx2_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
OR2x2_ASAP7_75t_L g314 ( .A(n_216), .B(n_315), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_217), .B(n_226), .Y(n_216) );
OR2x2_ASAP7_75t_L g242 ( .A(n_217), .B(n_243), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_217), .B(n_250), .Y(n_249) );
OR2x2_ASAP7_75t_L g282 ( .A(n_217), .B(n_227), .Y(n_282) );
AND2x2_ASAP7_75t_L g305 ( .A(n_217), .B(n_241), .Y(n_305) );
NOR2xp33_ASAP7_75t_L g316 ( .A(n_217), .B(n_317), .Y(n_316) );
AND2x2_ASAP7_75t_L g321 ( .A(n_217), .B(n_280), .Y(n_321) );
AND2x2_ASAP7_75t_L g329 ( .A(n_217), .B(n_330), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_217), .B(n_289), .Y(n_379) );
INVx5_ASAP7_75t_SL g217 ( .A(n_218), .Y(n_217) );
AND2x2_ASAP7_75t_L g269 ( .A(n_218), .B(n_243), .Y(n_269) );
OR2x2_ASAP7_75t_L g270 ( .A(n_218), .B(n_271), .Y(n_270) );
AND2x2_ASAP7_75t_L g296 ( .A(n_218), .B(n_227), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_218), .B(n_343), .Y(n_384) );
OR2x2_ASAP7_75t_L g400 ( .A(n_218), .B(n_344), .Y(n_400) );
AND2x2_ASAP7_75t_SL g407 ( .A(n_218), .B(n_361), .Y(n_407) );
HB1xp67_ASAP7_75t_L g414 ( .A(n_218), .Y(n_414) );
OR2x6_ASAP7_75t_L g218 ( .A(n_219), .B(n_225), .Y(n_218) );
AND2x2_ASAP7_75t_L g268 ( .A(n_226), .B(n_269), .Y(n_268) );
AND2x2_ASAP7_75t_L g318 ( .A(n_226), .B(n_241), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_226), .B(n_243), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_226), .B(n_280), .Y(n_402) );
INVx3_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_227), .B(n_243), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_227), .B(n_241), .Y(n_290) );
OR2x2_ASAP7_75t_L g344 ( .A(n_227), .B(n_241), .Y(n_344) );
AND2x2_ASAP7_75t_L g361 ( .A(n_227), .B(n_240), .Y(n_361) );
INVxp67_ASAP7_75t_L g383 ( .A(n_227), .Y(n_383) );
AND2x2_ASAP7_75t_L g410 ( .A(n_227), .B(n_280), .Y(n_410) );
HB1xp67_ASAP7_75t_L g417 ( .A(n_227), .Y(n_417) );
OA21x2_ASAP7_75t_L g227 ( .A1(n_228), .A2(n_229), .B(n_237), .Y(n_227) );
OA21x2_ASAP7_75t_L g471 ( .A1(n_228), .A2(n_472), .B(n_479), .Y(n_471) );
OA21x2_ASAP7_75t_L g494 ( .A1(n_228), .A2(n_495), .B(n_501), .Y(n_494) );
OA21x2_ASAP7_75t_L g514 ( .A1(n_228), .A2(n_515), .B(n_522), .Y(n_514) );
O2A1O1Ixp33_ASAP7_75t_L g259 ( .A1(n_233), .A2(n_260), .B(n_261), .C(n_262), .Y(n_259) );
INVx1_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
NOR2xp33_ASAP7_75t_L g499 ( .A(n_234), .B(n_500), .Y(n_499) );
NOR2xp33_ASAP7_75t_L g519 ( .A(n_234), .B(n_520), .Y(n_519) );
INVx1_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
OR2x2_ASAP7_75t_L g239 ( .A(n_240), .B(n_242), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_240), .B(n_291), .Y(n_364) );
INVx1_ASAP7_75t_SL g240 ( .A(n_241), .Y(n_240) );
AND2x2_ASAP7_75t_L g280 ( .A(n_241), .B(n_243), .Y(n_280) );
OR2x2_ASAP7_75t_L g347 ( .A(n_241), .B(n_348), .Y(n_347) );
INVx2_ASAP7_75t_L g291 ( .A(n_242), .Y(n_291) );
OR2x2_ASAP7_75t_L g352 ( .A(n_242), .B(n_344), .Y(n_352) );
INVx1_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
INVx1_ASAP7_75t_L g251 ( .A(n_246), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_246), .B(n_311), .Y(n_310) );
OR2x2_ASAP7_75t_L g252 ( .A(n_247), .B(n_253), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_247), .B(n_275), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_247), .B(n_254), .Y(n_287) );
INVx2_ASAP7_75t_L g332 ( .A(n_247), .Y(n_332) );
AND2x2_ASAP7_75t_L g345 ( .A(n_247), .B(n_285), .Y(n_345) );
AND2x2_ASAP7_75t_L g370 ( .A(n_247), .B(n_294), .Y(n_370) );
INVx1_ASAP7_75t_L g322 ( .A(n_252), .Y(n_322) );
INVx2_ASAP7_75t_SL g309 ( .A(n_253), .Y(n_309) );
INVx1_ASAP7_75t_L g312 ( .A(n_254), .Y(n_312) );
INVx2_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
HB1xp67_ASAP7_75t_L g275 ( .A(n_255), .Y(n_275) );
INVx2_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
BUFx2_ASAP7_75t_L g373 ( .A(n_256), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_258), .B(n_264), .Y(n_257) );
HB1xp67_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
INVx3_ASAP7_75t_L g478 ( .A(n_263), .Y(n_478) );
INVx1_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
AND2x2_ASAP7_75t_L g342 ( .A(n_269), .B(n_343), .Y(n_342) );
INVx1_ASAP7_75t_L g348 ( .A(n_269), .Y(n_348) );
AOI22xp5_ASAP7_75t_L g350 ( .A1(n_269), .A2(n_351), .B1(n_353), .B2(n_358), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_269), .B(n_361), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_270), .B(n_364), .Y(n_363) );
INVx1_ASAP7_75t_SL g304 ( .A(n_271), .Y(n_304) );
OR2x2_ASAP7_75t_L g272 ( .A(n_273), .B(n_274), .Y(n_272) );
OR2x2_ASAP7_75t_L g286 ( .A(n_273), .B(n_287), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_273), .B(n_277), .Y(n_337) );
AND2x2_ASAP7_75t_L g360 ( .A(n_273), .B(n_361), .Y(n_360) );
BUFx2_ASAP7_75t_L g336 ( .A(n_275), .Y(n_336) );
AOI211xp5_ASAP7_75t_L g276 ( .A1(n_277), .A2(n_278), .B(n_283), .C(n_297), .Y(n_276) );
INVx1_ASAP7_75t_L g300 ( .A(n_277), .Y(n_300) );
OAI221xp5_ASAP7_75t_SL g408 ( .A1(n_277), .A2(n_409), .B1(n_411), .B2(n_412), .C(n_415), .Y(n_408) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_280), .B(n_281), .Y(n_279) );
INVx1_ASAP7_75t_L g427 ( .A(n_280), .Y(n_427) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
OR2x2_ASAP7_75t_L g376 ( .A(n_282), .B(n_315), .Y(n_376) );
A2O1A1Ixp33_ASAP7_75t_L g283 ( .A1(n_284), .A2(n_286), .B(n_288), .C(n_292), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_289), .B(n_291), .Y(n_288) );
INVx1_ASAP7_75t_SL g289 ( .A(n_290), .Y(n_289) );
OAI32xp33_ASAP7_75t_L g401 ( .A1(n_290), .A2(n_291), .A3(n_354), .B1(n_391), .B2(n_402), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_293), .B(n_295), .Y(n_292) );
AND2x2_ASAP7_75t_L g433 ( .A(n_293), .B(n_332), .Y(n_433) );
AND2x2_ASAP7_75t_L g380 ( .A(n_294), .B(n_332), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_294), .B(n_302), .Y(n_398) );
AOI31xp33_ASAP7_75t_SL g297 ( .A1(n_298), .A2(n_300), .A3(n_301), .B(n_303), .Y(n_297) );
INVxp67_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_299), .B(n_311), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_299), .B(n_309), .Y(n_396) );
AOI221xp5_ASAP7_75t_L g418 ( .A1(n_299), .A2(n_329), .B1(n_419), .B2(n_422), .C(n_424), .Y(n_418) );
CKINVDCx16_ASAP7_75t_R g301 ( .A(n_302), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_304), .B(n_305), .Y(n_303) );
AND2x2_ASAP7_75t_L g324 ( .A(n_304), .B(n_325), .Y(n_324) );
AOI222xp33_ASAP7_75t_L g306 ( .A1(n_307), .A2(n_313), .B1(n_316), .B2(n_319), .C1(n_321), .C2(n_322), .Y(n_306) );
NAND2xp5_ASAP7_75t_SL g307 ( .A(n_308), .B(n_310), .Y(n_307) );
INVx1_ASAP7_75t_L g389 ( .A(n_308), .Y(n_389) );
INVx1_ASAP7_75t_L g411 ( .A(n_311), .Y(n_411) );
INVx2_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
OAI22xp5_ASAP7_75t_L g424 ( .A1(n_314), .A2(n_425), .B1(n_427), .B2(n_428), .Y(n_424) );
INVx1_ASAP7_75t_L g330 ( .A(n_315), .Y(n_330) );
INVx1_ASAP7_75t_SL g317 ( .A(n_318), .Y(n_317) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
AOI221xp5_ASAP7_75t_L g323 ( .A1(n_324), .A2(n_327), .B1(n_329), .B2(n_331), .C(n_334), .Y(n_323) );
INVx1_ASAP7_75t_SL g325 ( .A(n_326), .Y(n_325) );
OR2x2_ASAP7_75t_L g368 ( .A(n_326), .B(n_369), .Y(n_368) );
OR2x2_ASAP7_75t_L g420 ( .A(n_326), .B(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
INVx1_ASAP7_75t_L g395 ( .A(n_331), .Y(n_395) );
AND2x2_ASAP7_75t_L g331 ( .A(n_332), .B(n_333), .Y(n_331) );
INVx1_ASAP7_75t_L g359 ( .A(n_332), .Y(n_359) );
INVx1_ASAP7_75t_L g341 ( .A(n_333), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_336), .B(n_423), .Y(n_428) );
AOI22xp33_ASAP7_75t_L g338 ( .A1(n_339), .A2(n_342), .B1(n_345), .B2(n_346), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
INVx1_ASAP7_75t_SL g343 ( .A(n_344), .Y(n_343) );
INVx1_ASAP7_75t_SL g432 ( .A(n_345), .Y(n_432) );
INVxp33_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
NOR2xp33_ASAP7_75t_L g390 ( .A(n_347), .B(n_391), .Y(n_390) );
OAI32xp33_ASAP7_75t_L g381 ( .A1(n_348), .A2(n_382), .A3(n_383), .B1(n_384), .B2(n_385), .Y(n_381) );
NAND4xp25_ASAP7_75t_L g349 ( .A(n_350), .B(n_362), .C(n_374), .D(n_386), .Y(n_349) );
INVx1_ASAP7_75t_SL g351 ( .A(n_352), .Y(n_351) );
NAND2xp33_ASAP7_75t_SL g353 ( .A(n_354), .B(n_355), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_356), .B(n_357), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_357), .B(n_406), .Y(n_405) );
AND2x2_ASAP7_75t_L g358 ( .A(n_359), .B(n_360), .Y(n_358) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
CKINVDCx16_ASAP7_75t_R g367 ( .A(n_368), .Y(n_367) );
AOI221xp5_ASAP7_75t_L g403 ( .A1(n_371), .A2(n_387), .B1(n_404), .B2(n_407), .C(n_408), .Y(n_403) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
AND2x2_ASAP7_75t_L g422 ( .A(n_373), .B(n_423), .Y(n_422) );
AOI221xp5_ASAP7_75t_L g374 ( .A1(n_375), .A2(n_377), .B1(n_378), .B2(n_380), .C(n_381), .Y(n_374) );
INVx1_ASAP7_75t_SL g375 ( .A(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
NOR2xp33_ASAP7_75t_L g413 ( .A(n_383), .B(n_414), .Y(n_413) );
AOI21xp5_ASAP7_75t_L g386 ( .A1(n_387), .A2(n_389), .B(n_390), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
NAND4xp25_ASAP7_75t_L g392 ( .A(n_393), .B(n_403), .C(n_418), .D(n_429), .Y(n_392) );
O2A1O1Ixp33_ASAP7_75t_L g393 ( .A1(n_394), .A2(n_397), .B(n_399), .C(n_401), .Y(n_393) );
NAND2xp5_ASAP7_75t_SL g394 ( .A(n_395), .B(n_396), .Y(n_394) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVxp67_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx1_ASAP7_75t_SL g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g434 ( .A(n_421), .Y(n_434) );
INVx2_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
OAI21xp5_ASAP7_75t_L g429 ( .A1(n_430), .A2(n_433), .B(n_434), .Y(n_429) );
NOR2xp33_ASAP7_75t_L g430 ( .A(n_431), .B(n_432), .Y(n_430) );
AOI22xp5_ASAP7_75t_L g446 ( .A1(n_435), .A2(n_447), .B1(n_449), .B2(n_451), .Y(n_446) );
NOR2xp33_ASAP7_75t_SL g442 ( .A(n_436), .B(n_443), .Y(n_442) );
HB1xp67_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx2_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
AND2x2_ASAP7_75t_L g439 ( .A(n_440), .B(n_441), .Y(n_439) );
OAI21xp5_ASAP7_75t_SL g444 ( .A1(n_442), .A2(n_445), .B(n_739), .Y(n_444) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx1_ASAP7_75t_L g731 ( .A(n_448), .Y(n_731) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx6_ASAP7_75t_L g732 ( .A(n_450), .Y(n_732) );
INVx3_ASAP7_75t_L g733 ( .A(n_451), .Y(n_733) );
AND2x2_ASAP7_75t_SL g451 ( .A(n_452), .B(n_682), .Y(n_451) );
NOR4xp25_ASAP7_75t_L g452 ( .A(n_453), .B(n_619), .C(n_653), .D(n_669), .Y(n_452) );
NAND4xp25_ASAP7_75t_SL g453 ( .A(n_454), .B(n_548), .C(n_583), .D(n_599), .Y(n_453) );
AOI222xp33_ASAP7_75t_L g454 ( .A1(n_455), .A2(n_489), .B1(n_523), .B2(n_536), .C1(n_541), .C2(n_547), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
AOI31xp33_ASAP7_75t_L g715 ( .A1(n_456), .A2(n_716), .A3(n_717), .B(n_719), .Y(n_715) );
OR2x2_ASAP7_75t_L g456 ( .A(n_457), .B(n_468), .Y(n_456) );
AND2x2_ASAP7_75t_L g690 ( .A(n_457), .B(n_470), .Y(n_690) );
BUFx2_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx2_ASAP7_75t_SL g540 ( .A(n_458), .Y(n_540) );
AND2x2_ASAP7_75t_L g547 ( .A(n_458), .B(n_480), .Y(n_547) );
AND2x2_ASAP7_75t_L g604 ( .A(n_458), .B(n_471), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_468), .B(n_634), .Y(n_633) );
INVx3_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
NOR2xp33_ASAP7_75t_L g567 ( .A(n_469), .B(n_568), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_469), .B(n_551), .Y(n_594) );
AND2x2_ASAP7_75t_L g687 ( .A(n_469), .B(n_627), .Y(n_687) );
OAI321xp33_ASAP7_75t_L g721 ( .A1(n_469), .A2(n_540), .A3(n_694), .B1(n_722), .B2(n_724), .C(n_725), .Y(n_721) );
NAND4xp25_ASAP7_75t_L g725 ( .A(n_469), .B(n_526), .C(n_634), .D(n_726), .Y(n_725) );
AND2x4_ASAP7_75t_L g469 ( .A(n_470), .B(n_480), .Y(n_469) );
AND2x2_ASAP7_75t_L g589 ( .A(n_470), .B(n_538), .Y(n_589) );
AND2x2_ASAP7_75t_L g608 ( .A(n_470), .B(n_540), .Y(n_608) );
INVx2_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
AND2x2_ASAP7_75t_L g539 ( .A(n_471), .B(n_540), .Y(n_539) );
AND2x2_ASAP7_75t_L g564 ( .A(n_471), .B(n_480), .Y(n_564) );
AND2x2_ASAP7_75t_L g650 ( .A(n_471), .B(n_538), .Y(n_650) );
INVx3_ASAP7_75t_SL g538 ( .A(n_480), .Y(n_538) );
AND2x2_ASAP7_75t_L g582 ( .A(n_480), .B(n_569), .Y(n_582) );
OR2x2_ASAP7_75t_L g615 ( .A(n_480), .B(n_540), .Y(n_615) );
HB1xp67_ASAP7_75t_L g622 ( .A(n_480), .Y(n_622) );
AND2x2_ASAP7_75t_L g651 ( .A(n_480), .B(n_539), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_480), .B(n_624), .Y(n_666) );
AND2x2_ASAP7_75t_L g698 ( .A(n_480), .B(n_690), .Y(n_698) );
AND2x2_ASAP7_75t_L g707 ( .A(n_480), .B(n_552), .Y(n_707) );
OR2x6_ASAP7_75t_L g480 ( .A(n_481), .B(n_487), .Y(n_480) );
INVx1_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_491), .B(n_502), .Y(n_490) );
INVx1_ASAP7_75t_SL g675 ( .A(n_491), .Y(n_675) );
INVx2_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
AND2x2_ASAP7_75t_L g543 ( .A(n_492), .B(n_544), .Y(n_543) );
INVx2_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
AND2x2_ASAP7_75t_L g525 ( .A(n_493), .B(n_504), .Y(n_525) );
AND2x2_ASAP7_75t_L g611 ( .A(n_493), .B(n_527), .Y(n_611) );
INVx2_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
AND2x2_ASAP7_75t_L g581 ( .A(n_494), .B(n_514), .Y(n_581) );
OR2x2_ASAP7_75t_L g592 ( .A(n_494), .B(n_527), .Y(n_592) );
AND2x2_ASAP7_75t_L g618 ( .A(n_494), .B(n_527), .Y(n_618) );
HB1xp67_ASAP7_75t_L g663 ( .A(n_494), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_502), .B(n_618), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_502), .B(n_675), .Y(n_674) );
INVx2_ASAP7_75t_SL g502 ( .A(n_503), .Y(n_502) );
OR2x2_ASAP7_75t_L g591 ( .A(n_503), .B(n_592), .Y(n_591) );
AOI322xp5_ASAP7_75t_L g677 ( .A1(n_503), .A2(n_581), .A3(n_587), .B1(n_618), .B2(n_668), .C1(n_678), .C2(n_680), .Y(n_677) );
OR2x2_ASAP7_75t_L g503 ( .A(n_504), .B(n_514), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_504), .B(n_526), .Y(n_546) );
NOR2xp33_ASAP7_75t_L g574 ( .A(n_504), .B(n_527), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_504), .B(n_544), .Y(n_598) );
AND2x2_ASAP7_75t_L g652 ( .A(n_504), .B(n_618), .Y(n_652) );
INVx1_ASAP7_75t_L g656 ( .A(n_504), .Y(n_656) );
AND2x2_ASAP7_75t_L g668 ( .A(n_504), .B(n_514), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_504), .B(n_543), .Y(n_700) );
INVx4_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
AND2x2_ASAP7_75t_L g565 ( .A(n_505), .B(n_514), .Y(n_565) );
BUFx3_ASAP7_75t_L g579 ( .A(n_505), .Y(n_579) );
AND3x2_ASAP7_75t_L g661 ( .A(n_505), .B(n_641), .C(n_662), .Y(n_661) );
NAND3xp33_ASAP7_75t_L g524 ( .A(n_514), .B(n_525), .C(n_526), .Y(n_524) );
INVx1_ASAP7_75t_SL g544 ( .A(n_514), .Y(n_544) );
HB1xp67_ASAP7_75t_L g646 ( .A(n_514), .Y(n_646) );
INVx1_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
AND2x2_ASAP7_75t_L g640 ( .A(n_525), .B(n_641), .Y(n_640) );
INVxp67_ASAP7_75t_L g647 ( .A(n_525), .Y(n_647) );
AND2x2_ASAP7_75t_L g685 ( .A(n_526), .B(n_663), .Y(n_685) );
INVx2_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
BUFx3_ASAP7_75t_L g566 ( .A(n_527), .Y(n_566) );
AND2x2_ASAP7_75t_L g641 ( .A(n_527), .B(n_544), .Y(n_641) );
INVx1_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_538), .B(n_539), .Y(n_537) );
OR2x2_ASAP7_75t_L g585 ( .A(n_538), .B(n_586), .Y(n_585) );
AND2x2_ASAP7_75t_L g704 ( .A(n_538), .B(n_604), .Y(n_704) );
AND2x2_ASAP7_75t_L g718 ( .A(n_538), .B(n_540), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_539), .B(n_552), .Y(n_659) );
AND2x2_ASAP7_75t_L g706 ( .A(n_539), .B(n_707), .Y(n_706) );
AND2x2_ASAP7_75t_L g569 ( .A(n_540), .B(n_570), .Y(n_569) );
OR2x2_ASAP7_75t_L g586 ( .A(n_540), .B(n_552), .Y(n_586) );
INVx1_ASAP7_75t_L g596 ( .A(n_540), .Y(n_596) );
AND2x2_ASAP7_75t_L g627 ( .A(n_540), .B(n_552), .Y(n_627) );
INVx1_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
OAI221xp5_ASAP7_75t_L g669 ( .A1(n_542), .A2(n_670), .B1(n_674), .B2(n_676), .C(n_677), .Y(n_669) );
NAND2xp5_ASAP7_75t_SL g542 ( .A(n_543), .B(n_545), .Y(n_542) );
AND2x2_ASAP7_75t_L g573 ( .A(n_543), .B(n_574), .Y(n_573) );
INVx1_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
NOR2xp33_ASAP7_75t_L g723 ( .A(n_546), .B(n_580), .Y(n_723) );
AOI322xp5_ASAP7_75t_L g548 ( .A1(n_549), .A2(n_565), .A3(n_566), .B1(n_567), .B2(n_573), .C1(n_575), .C2(n_582), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_551), .B(n_564), .Y(n_550) );
NAND2x1p5_ASAP7_75t_L g603 ( .A(n_551), .B(n_604), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_551), .B(n_614), .Y(n_613) );
O2A1O1Ixp33_ASAP7_75t_L g637 ( .A1(n_551), .A2(n_564), .B(n_638), .C(n_639), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_551), .B(n_650), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_551), .B(n_608), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_551), .B(n_690), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_551), .B(n_718), .Y(n_717) );
BUFx3_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_552), .B(n_589), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_552), .B(n_596), .Y(n_595) );
OR2x2_ASAP7_75t_L g679 ( .A(n_552), .B(n_566), .Y(n_679) );
OA21x2_ASAP7_75t_L g552 ( .A1(n_553), .A2(n_556), .B(n_563), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
AO21x2_ASAP7_75t_L g570 ( .A1(n_554), .A2(n_571), .B(n_572), .Y(n_570) );
INVx1_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
INVx1_ASAP7_75t_L g571 ( .A(n_556), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_563), .Y(n_572) );
INVx1_ASAP7_75t_L g654 ( .A(n_564), .Y(n_654) );
OAI31xp33_ASAP7_75t_L g664 ( .A1(n_564), .A2(n_589), .A3(n_665), .B(n_667), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_564), .B(n_570), .Y(n_716) );
INVx1_ASAP7_75t_SL g577 ( .A(n_565), .Y(n_577) );
AND2x2_ASAP7_75t_L g610 ( .A(n_565), .B(n_611), .Y(n_610) );
AND2x2_ASAP7_75t_L g691 ( .A(n_565), .B(n_692), .Y(n_691) );
OR2x2_ASAP7_75t_L g576 ( .A(n_566), .B(n_577), .Y(n_576) );
INVx1_ASAP7_75t_L g601 ( .A(n_566), .Y(n_601) );
AND2x2_ASAP7_75t_L g628 ( .A(n_566), .B(n_581), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_566), .B(n_646), .Y(n_645) );
AND2x2_ASAP7_75t_L g720 ( .A(n_566), .B(n_668), .Y(n_720) );
NOR2xp33_ASAP7_75t_L g711 ( .A(n_568), .B(n_638), .Y(n_711) );
INVx1_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
AND2x2_ASAP7_75t_L g607 ( .A(n_570), .B(n_608), .Y(n_607) );
INVx1_ASAP7_75t_SL g625 ( .A(n_570), .Y(n_625) );
NAND2xp33_ASAP7_75t_SL g575 ( .A(n_576), .B(n_578), .Y(n_575) );
OAI211xp5_ASAP7_75t_SL g619 ( .A1(n_577), .A2(n_620), .B(n_626), .C(n_642), .Y(n_619) );
OR2x2_ASAP7_75t_L g694 ( .A(n_577), .B(n_675), .Y(n_694) );
OR2x2_ASAP7_75t_L g578 ( .A(n_579), .B(n_580), .Y(n_578) );
CKINVDCx16_ASAP7_75t_R g631 ( .A(n_579), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_579), .B(n_685), .Y(n_684) );
INVx1_ASAP7_75t_SL g580 ( .A(n_581), .Y(n_580) );
AND2x2_ASAP7_75t_L g600 ( .A(n_581), .B(n_601), .Y(n_600) );
O2A1O1Ixp33_ASAP7_75t_L g583 ( .A1(n_584), .A2(n_587), .B(n_590), .C(n_593), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
INVx1_ASAP7_75t_SL g634 ( .A(n_586), .Y(n_634) );
INVx1_ASAP7_75t_SL g587 ( .A(n_588), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_589), .B(n_627), .Y(n_632) );
INVx1_ASAP7_75t_L g638 ( .A(n_589), .Y(n_638) );
INVx1_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
OR2x2_ASAP7_75t_L g597 ( .A(n_592), .B(n_598), .Y(n_597) );
OR2x2_ASAP7_75t_L g630 ( .A(n_592), .B(n_631), .Y(n_630) );
INVx1_ASAP7_75t_L g692 ( .A(n_592), .Y(n_692) );
AOI21xp33_ASAP7_75t_SL g593 ( .A1(n_594), .A2(n_595), .B(n_597), .Y(n_593) );
AOI21xp5_ASAP7_75t_L g605 ( .A1(n_595), .A2(n_606), .B(n_609), .Y(n_605) );
AOI211xp5_ASAP7_75t_L g599 ( .A1(n_600), .A2(n_602), .B(n_605), .C(n_612), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_600), .B(n_656), .Y(n_655) );
INVx1_ASAP7_75t_SL g602 ( .A(n_603), .Y(n_602) );
NOR2xp33_ASAP7_75t_L g693 ( .A(n_603), .B(n_694), .Y(n_693) );
INVx2_ASAP7_75t_SL g616 ( .A(n_604), .Y(n_616) );
OAI21xp5_ASAP7_75t_L g671 ( .A1(n_606), .A2(n_672), .B(n_673), .Y(n_671) );
INVx1_ASAP7_75t_SL g606 ( .A(n_607), .Y(n_606) );
INVx1_ASAP7_75t_SL g609 ( .A(n_610), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_611), .B(n_624), .Y(n_623) );
INVx1_ASAP7_75t_SL g636 ( .A(n_611), .Y(n_636) );
AOI21xp33_ASAP7_75t_SL g612 ( .A1(n_613), .A2(n_616), .B(n_617), .Y(n_612) );
INVx1_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
AND2x2_ASAP7_75t_L g667 ( .A(n_618), .B(n_668), .Y(n_667) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
NOR2xp33_ASAP7_75t_L g621 ( .A(n_622), .B(n_623), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_624), .B(n_650), .Y(n_676) );
AND2x2_ASAP7_75t_L g689 ( .A(n_624), .B(n_690), .Y(n_689) );
AND2x2_ASAP7_75t_L g703 ( .A(n_624), .B(n_704), .Y(n_703) );
AND2x2_ASAP7_75t_L g713 ( .A(n_624), .B(n_651), .Y(n_713) );
INVx2_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
AOI211xp5_ASAP7_75t_L g626 ( .A1(n_627), .A2(n_628), .B(n_629), .C(n_637), .Y(n_626) );
INVx1_ASAP7_75t_L g673 ( .A(n_627), .Y(n_673) );
OAI22xp33_ASAP7_75t_L g629 ( .A1(n_630), .A2(n_632), .B1(n_633), .B2(n_635), .Y(n_629) );
OR2x2_ASAP7_75t_L g635 ( .A(n_631), .B(n_636), .Y(n_635) );
NAND2xp5_ASAP7_75t_SL g714 ( .A(n_631), .B(n_692), .Y(n_714) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
INVx1_ASAP7_75t_L g708 ( .A(n_641), .Y(n_708) );
AOI22xp33_ASAP7_75t_L g642 ( .A1(n_643), .A2(n_648), .B1(n_651), .B2(n_652), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
OR2x2_ASAP7_75t_L g644 ( .A(n_645), .B(n_647), .Y(n_644) );
INVx1_ASAP7_75t_L g726 ( .A(n_646), .Y(n_726) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
INVx1_ASAP7_75t_L g672 ( .A(n_650), .Y(n_672) );
OAI211xp5_ASAP7_75t_SL g653 ( .A1(n_654), .A2(n_655), .B(n_657), .C(n_664), .Y(n_653) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
NOR2xp33_ASAP7_75t_L g658 ( .A(n_659), .B(n_660), .Y(n_658) );
INVx2_ASAP7_75t_SL g660 ( .A(n_661), .Y(n_660) );
INVxp67_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
INVxp67_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
NOR2xp33_ASAP7_75t_L g678 ( .A(n_672), .B(n_679), .Y(n_678) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
NOR5xp2_ASAP7_75t_L g682 ( .A(n_683), .B(n_701), .C(n_709), .D(n_715), .E(n_721), .Y(n_682) );
OAI211xp5_ASAP7_75t_SL g683 ( .A1(n_684), .A2(n_686), .B(n_688), .C(n_695), .Y(n_683) );
INVxp67_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
AOI21xp5_ASAP7_75t_L g688 ( .A1(n_689), .A2(n_691), .B(n_693), .Y(n_688) );
OAI21xp33_ASAP7_75t_L g695 ( .A1(n_696), .A2(n_698), .B(n_699), .Y(n_695) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
NOR2xp33_ASAP7_75t_L g710 ( .A(n_698), .B(n_711), .Y(n_710) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
AOI21xp33_ASAP7_75t_L g701 ( .A1(n_702), .A2(n_705), .B(n_708), .Y(n_701) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
INVx1_ASAP7_75t_SL g724 ( .A(n_704), .Y(n_724) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
AOI21xp5_ASAP7_75t_L g709 ( .A1(n_710), .A2(n_712), .B(n_714), .Y(n_709) );
INVx1_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
INVx1_ASAP7_75t_SL g729 ( .A(n_730), .Y(n_729) );
INVx2_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
INVx1_ASAP7_75t_SL g734 ( .A(n_735), .Y(n_734) );
INVx1_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
INVx2_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
INVx2_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
INVx1_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
endmodule