module fake_jpeg_21106_n_173 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_173);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_173;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx14_ASAP7_75t_R g15 ( 
.A(n_0),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx1_ASAP7_75t_SL g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_22),
.B(n_5),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_32),
.B(n_39),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

AND2x2_ASAP7_75t_SL g34 ( 
.A(n_22),
.B(n_0),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_34),
.B(n_27),
.Y(n_47)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

BUFx4f_ASAP7_75t_SL g37 ( 
.A(n_27),
.Y(n_37)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_19),
.B(n_4),
.Y(n_39)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_47),
.B(n_33),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g48 ( 
.A(n_37),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_48),
.B(n_49),
.Y(n_65)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

INVx4_ASAP7_75t_SL g60 ( 
.A(n_50),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_31),
.A2(n_24),
.B1(n_26),
.B2(n_15),
.Y(n_51)
);

AO22x1_ASAP7_75t_SL g57 ( 
.A1(n_51),
.A2(n_53),
.B1(n_49),
.B2(n_35),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_32),
.B(n_19),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_54),
.B(n_29),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_55),
.B(n_27),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_29),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_56),
.B(n_25),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_57),
.A2(n_40),
.B1(n_43),
.B2(n_44),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_L g58 ( 
.A1(n_47),
.A2(n_34),
.B(n_38),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_58),
.B(n_61),
.Y(n_87)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_59),
.Y(n_83)
);

AO22x1_ASAP7_75t_SL g61 ( 
.A1(n_53),
.A2(n_34),
.B1(n_37),
.B2(n_40),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_62),
.B(n_64),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_46),
.B(n_34),
.C(n_36),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_63),
.B(n_67),
.Y(n_95)
);

FAx1_ASAP7_75t_SL g64 ( 
.A(n_45),
.B(n_34),
.CI(n_37),
.CON(n_64),
.SN(n_64)
);

INVxp33_ASAP7_75t_L g84 ( 
.A(n_66),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_50),
.B(n_25),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_68),
.B(n_70),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_69),
.B(n_72),
.Y(n_78)
);

AOI21xp33_ASAP7_75t_L g70 ( 
.A1(n_55),
.A2(n_18),
.B(n_21),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_52),
.Y(n_71)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_71),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_52),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_42),
.B(n_36),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_73),
.B(n_74),
.Y(n_89)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_52),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_41),
.B(n_36),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_75),
.B(n_76),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_43),
.B(n_18),
.Y(n_76)
);

AND2x4_ASAP7_75t_SL g79 ( 
.A(n_61),
.B(n_41),
.Y(n_79)
);

AO22x1_ASAP7_75t_L g98 ( 
.A1(n_79),
.A2(n_82),
.B1(n_73),
.B2(n_61),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_62),
.B(n_21),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_80),
.B(n_90),
.Y(n_99)
);

INVxp33_ASAP7_75t_L g88 ( 
.A(n_65),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_88),
.B(n_93),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_60),
.B(n_24),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_75),
.Y(n_91)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_91),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_59),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_92),
.B(n_94),
.Y(n_101)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_71),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_60),
.B(n_17),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_58),
.A2(n_33),
.B1(n_26),
.B2(n_44),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_96),
.B(n_57),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_98),
.A2(n_103),
.B1(n_82),
.B2(n_97),
.Y(n_114)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_83),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_100),
.B(n_109),
.Y(n_127)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_83),
.Y(n_102)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_102),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_95),
.B(n_67),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_105),
.B(n_106),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_95),
.B(n_63),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_87),
.B(n_91),
.C(n_96),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_107),
.B(n_111),
.C(n_112),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_87),
.B(n_64),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_108),
.B(n_85),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_78),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_79),
.A2(n_81),
.B1(n_74),
.B2(n_93),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_110),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_79),
.B(n_64),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_79),
.B(n_72),
.C(n_57),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_89),
.A2(n_0),
.B(n_1),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_113),
.A2(n_86),
.B(n_15),
.Y(n_122)
);

NAND3xp33_ASAP7_75t_SL g139 ( 
.A(n_114),
.B(n_126),
.C(n_98),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_104),
.B(n_78),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_115),
.B(n_117),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_101),
.B(n_85),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_103),
.A2(n_89),
.B1(n_77),
.B2(n_92),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_119),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_121),
.B(n_124),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_122),
.A2(n_28),
.B(n_20),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_102),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_107),
.A2(n_86),
.B1(n_84),
.B2(n_81),
.Y(n_125)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_125),
.Y(n_130)
);

NOR2x1_ASAP7_75t_L g126 ( 
.A(n_113),
.B(n_28),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_99),
.B(n_27),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_128),
.B(n_112),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_123),
.B(n_106),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_129),
.B(n_132),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_123),
.B(n_105),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_133),
.B(n_138),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_120),
.B(n_111),
.C(n_108),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_134),
.B(n_135),
.C(n_119),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_125),
.B(n_120),
.Y(n_135)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_139),
.Y(n_148)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_118),
.Y(n_140)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_140),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_141),
.B(n_132),
.C(n_30),
.Y(n_151)
);

AOI322xp5_ASAP7_75t_L g143 ( 
.A1(n_130),
.A2(n_117),
.A3(n_121),
.B1(n_127),
.B2(n_114),
.C1(n_116),
.C2(n_122),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_143),
.A2(n_144),
.B(n_6),
.Y(n_152)
);

AOI322xp5_ASAP7_75t_L g144 ( 
.A1(n_136),
.A2(n_98),
.A3(n_126),
.B1(n_118),
.B2(n_124),
.C1(n_30),
.C2(n_23),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_136),
.A2(n_131),
.B1(n_129),
.B2(n_135),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_146),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_134),
.A2(n_17),
.B1(n_30),
.B2(n_23),
.Y(n_149)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_149),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_146),
.B(n_137),
.Y(n_150)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_150),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_151),
.B(n_154),
.C(n_149),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_152),
.B(n_153),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_145),
.B(n_141),
.C(n_147),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_148),
.A2(n_4),
.B(n_9),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_156),
.A2(n_9),
.B(n_10),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_154),
.B(n_145),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_157),
.B(n_158),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_151),
.B(n_142),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_159),
.B(n_155),
.Y(n_165)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_160),
.Y(n_164)
);

OR2x2_ASAP7_75t_L g163 ( 
.A(n_161),
.B(n_142),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_163),
.A2(n_2),
.B1(n_3),
.B2(n_14),
.Y(n_168)
);

OAI21xp33_ASAP7_75t_L g167 ( 
.A1(n_165),
.A2(n_162),
.B(n_157),
.Y(n_167)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_167),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_168),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_166),
.B(n_2),
.C(n_3),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_171),
.A2(n_164),
.B(n_169),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_172),
.B(n_170),
.Y(n_173)
);


endmodule