module fake_jpeg_26205_n_271 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_271);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_271;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_127;
wire n_154;
wire n_76;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_155;
wire n_118;
wire n_258;
wire n_96;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx16f_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

CKINVDCx16_ASAP7_75t_R g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_7),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_10),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_0),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_18),
.B(n_8),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_38),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_18),
.B(n_0),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_36),
.B(n_41),
.Y(n_48)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_18),
.B(n_0),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_26),
.B(n_34),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_39),
.B(n_40),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_26),
.B(n_1),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_26),
.B(n_34),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_43),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_36),
.A2(n_30),
.B1(n_31),
.B2(n_32),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_46),
.A2(n_63),
.B1(n_40),
.B2(n_24),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_36),
.A2(n_30),
.B1(n_31),
.B2(n_32),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_47),
.A2(n_33),
.B1(n_28),
.B2(n_27),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

INVx13_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_51),
.B(n_54),
.Y(n_81)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx2_ASAP7_75t_SL g76 ( 
.A(n_52),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_37),
.A2(n_31),
.B1(n_30),
.B2(n_29),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_53),
.Y(n_84)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_38),
.B(n_35),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_55),
.B(n_24),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_56),
.Y(n_69)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_58),
.Y(n_68)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_59),
.Y(n_80)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_60),
.Y(n_64)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

AO22x1_ASAP7_75t_L g83 ( 
.A1(n_61),
.A2(n_22),
.B1(n_28),
.B2(n_27),
.Y(n_83)
);

OAI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_41),
.A2(n_29),
.B1(n_24),
.B2(n_34),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_55),
.B(n_17),
.Y(n_65)
);

A2O1A1Ixp33_ASAP7_75t_L g120 ( 
.A1(n_65),
.A2(n_57),
.B(n_22),
.C(n_4),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_46),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_67),
.B(n_70),
.Y(n_101)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_60),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_56),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_71),
.B(n_74),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_72),
.B(n_83),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_73),
.B(n_89),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_54),
.B(n_25),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_62),
.B(n_25),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_75),
.B(n_91),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_56),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_77),
.Y(n_118)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_60),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_78),
.B(n_79),
.Y(n_116)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_45),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_48),
.B(n_33),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_82),
.B(n_87),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_61),
.A2(n_33),
.B1(n_28),
.B2(n_27),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_85),
.A2(n_86),
.B1(n_20),
.B2(n_19),
.Y(n_111)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_45),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_48),
.B(n_23),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_88),
.B(n_94),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_56),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_49),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_90),
.B(n_92),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_50),
.B(n_23),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_50),
.B(n_23),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_61),
.A2(n_22),
.B(n_2),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_93),
.A2(n_84),
.B(n_65),
.Y(n_103)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_49),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_51),
.B(n_21),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_95),
.B(n_1),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_51),
.Y(n_96)
);

HB1xp67_ASAP7_75t_L g102 ( 
.A(n_96),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_44),
.A2(n_21),
.B1(n_20),
.B2(n_19),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_97),
.A2(n_73),
.B1(n_92),
.B2(n_72),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_58),
.Y(n_98)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_98),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_59),
.B(n_21),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_99),
.B(n_16),
.Y(n_126)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_52),
.Y(n_100)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_100),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_103),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_67),
.A2(n_57),
.B1(n_44),
.B2(n_20),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_106),
.A2(n_113),
.B1(n_114),
.B2(n_123),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_66),
.Y(n_110)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_110),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_111),
.A2(n_121),
.B1(n_109),
.B2(n_97),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_65),
.A2(n_19),
.B(n_2),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_112),
.A2(n_120),
.B(n_5),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_93),
.A2(n_57),
.B1(n_44),
.B2(n_22),
.Y(n_114)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_68),
.Y(n_117)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_117),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_86),
.A2(n_22),
.B1(n_3),
.B2(n_4),
.Y(n_121)
);

CKINVDCx14_ASAP7_75t_R g149 ( 
.A(n_122),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_82),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_88),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_124),
.A2(n_123),
.B1(n_113),
.B2(n_126),
.Y(n_148)
);

CKINVDCx14_ASAP7_75t_R g150 ( 
.A(n_126),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_115),
.A2(n_85),
.B1(n_83),
.B2(n_64),
.Y(n_129)
);

CKINVDCx14_ASAP7_75t_R g159 ( 
.A(n_129),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_119),
.B(n_83),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_130),
.B(n_131),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_119),
.B(n_81),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_133),
.A2(n_136),
.B1(n_147),
.B2(n_107),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_115),
.A2(n_70),
.B1(n_78),
.B2(n_64),
.Y(n_135)
);

HAxp5_ASAP7_75t_SL g172 ( 
.A(n_135),
.B(n_146),
.CON(n_172),
.SN(n_172)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_101),
.A2(n_94),
.B1(n_79),
.B2(n_87),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_116),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_137),
.B(n_139),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_109),
.B(n_81),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_138),
.B(n_151),
.Y(n_179)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_116),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_103),
.B(n_96),
.C(n_90),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_140),
.B(n_155),
.C(n_108),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_105),
.B(n_99),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_141),
.B(n_127),
.Y(n_158)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_101),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_142),
.B(n_144),
.Y(n_170)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_106),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_104),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_145),
.B(n_148),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_115),
.A2(n_66),
.B1(n_68),
.B2(n_80),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_105),
.B(n_80),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_102),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_152),
.B(n_154),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_107),
.B(n_89),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_153),
.B(n_156),
.Y(n_182)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_118),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_104),
.B(n_100),
.C(n_77),
.Y(n_155)
);

AO22x1_ASAP7_75t_SL g156 ( 
.A1(n_114),
.A2(n_76),
.B1(n_71),
.B2(n_69),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_157),
.B(n_173),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_158),
.B(n_163),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_152),
.B(n_118),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_143),
.A2(n_112),
.B(n_120),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_SL g203 ( 
.A(n_164),
.B(n_168),
.Y(n_203)
);

AO22x2_ASAP7_75t_SL g165 ( 
.A1(n_129),
.A2(n_111),
.B1(n_121),
.B2(n_110),
.Y(n_165)
);

OA21x2_ASAP7_75t_L g196 ( 
.A1(n_165),
.A2(n_146),
.B(n_132),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_151),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_166),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_141),
.B(n_124),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_167),
.B(n_171),
.Y(n_202)
);

A2O1A1O1Ixp25_ASAP7_75t_L g168 ( 
.A1(n_135),
.A2(n_126),
.B(n_122),
.C(n_76),
.D(n_125),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_133),
.A2(n_122),
.B1(n_108),
.B2(n_76),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_169),
.A2(n_178),
.B1(n_139),
.B2(n_137),
.Y(n_192)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_136),
.Y(n_171)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_147),
.Y(n_173)
);

AOI322xp5_ASAP7_75t_SL g174 ( 
.A1(n_149),
.A2(n_5),
.A3(n_6),
.B1(n_7),
.B2(n_8),
.C1(n_9),
.C2(n_11),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_174),
.B(n_175),
.Y(n_193)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_153),
.Y(n_175)
);

HB1xp67_ASAP7_75t_L g176 ( 
.A(n_155),
.Y(n_176)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_176),
.Y(n_184)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_156),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_177),
.B(n_110),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_144),
.A2(n_142),
.B1(n_128),
.B2(n_156),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_180),
.B(n_128),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_180),
.B(n_140),
.C(n_138),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_183),
.B(n_188),
.C(n_191),
.Y(n_211)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_181),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_187),
.B(n_198),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_160),
.B(n_131),
.C(n_130),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_172),
.Y(n_189)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_189),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_181),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_190),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_192),
.A2(n_165),
.B1(n_194),
.B2(n_169),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_165),
.A2(n_154),
.B1(n_156),
.B2(n_150),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_194),
.A2(n_196),
.B1(n_182),
.B2(n_171),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_160),
.B(n_179),
.C(n_159),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_197),
.B(n_164),
.C(n_175),
.Y(n_217)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_170),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_166),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_199),
.B(n_201),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_161),
.B(n_148),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_200),
.B(n_204),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_179),
.B(n_178),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_185),
.A2(n_177),
.B1(n_165),
.B2(n_173),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_205),
.A2(n_214),
.B1(n_220),
.B2(n_219),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_191),
.B(n_157),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_207),
.B(n_215),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_195),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_208),
.A2(n_202),
.B(n_192),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_210),
.A2(n_216),
.B1(n_132),
.B2(n_134),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_196),
.A2(n_182),
.B(n_170),
.Y(n_214)
);

A2O1A1Ixp33_ASAP7_75t_SL g234 ( 
.A1(n_214),
.A2(n_9),
.B(n_12),
.C(n_13),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_183),
.B(n_203),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_217),
.B(n_189),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_203),
.B(n_162),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_218),
.B(n_200),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_184),
.B(n_162),
.C(n_167),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_220),
.B(n_187),
.C(n_197),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_184),
.A2(n_158),
.B(n_168),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_221),
.B(n_196),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_223),
.B(n_229),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_224),
.B(n_225),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_211),
.B(n_204),
.C(n_188),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_226),
.B(n_227),
.Y(n_236)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_212),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_228),
.B(n_230),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_206),
.A2(n_186),
.B(n_193),
.Y(n_230)
);

NOR3xp33_ASAP7_75t_SL g231 ( 
.A(n_208),
.B(n_125),
.C(n_12),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_231),
.B(n_12),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_232),
.A2(n_233),
.B1(n_205),
.B2(n_213),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_216),
.A2(n_134),
.B1(n_117),
.B2(n_69),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_234),
.B(n_218),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_235),
.A2(n_209),
.B1(n_207),
.B2(n_217),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_237),
.B(n_240),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_239),
.B(n_245),
.Y(n_247)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_231),
.Y(n_240)
);

INVx6_ASAP7_75t_L g242 ( 
.A(n_224),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_242),
.A2(n_223),
.B1(n_215),
.B2(n_234),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_226),
.A2(n_234),
.B1(n_211),
.B2(n_229),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_243),
.B(n_244),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_239),
.B(n_222),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_248),
.B(n_254),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_L g249 ( 
.A1(n_236),
.A2(n_238),
.B(n_242),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_249),
.B(n_250),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_246),
.B(n_222),
.C(n_209),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_251),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_241),
.B(n_234),
.Y(n_254)
);

OR2x2_ASAP7_75t_L g255 ( 
.A(n_252),
.B(n_245),
.Y(n_255)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_255),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_253),
.A2(n_246),
.B1(n_241),
.B2(n_16),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_258),
.A2(n_260),
.B1(n_14),
.B2(n_250),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_254),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_259),
.B(n_247),
.Y(n_262)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_262),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_257),
.B(n_247),
.C(n_248),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_263),
.B(n_264),
.Y(n_265)
);

NAND2xp33_ASAP7_75t_SL g266 ( 
.A(n_261),
.B(n_255),
.Y(n_266)
);

NAND3xp33_ASAP7_75t_SL g269 ( 
.A(n_266),
.B(n_256),
.C(n_263),
.Y(n_269)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_265),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_268),
.B(n_269),
.C(n_267),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_270),
.B(n_256),
.Y(n_271)
);


endmodule