module fake_jpeg_2871_n_132 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_132);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_132;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_5),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_6),
.Y(n_14)
);

INVx3_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_4),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_12),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_24),
.Y(n_28)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_24),
.Y(n_29)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_25),
.Y(n_30)
);

INVx3_ASAP7_75t_SL g49 ( 
.A(n_30),
.Y(n_49)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_25),
.Y(n_31)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_31),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_22),
.B(n_0),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_32),
.B(n_27),
.Y(n_52)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_34),
.B(n_35),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_16),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_26),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_37),
.A2(n_15),
.B1(n_17),
.B2(n_16),
.Y(n_45)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_40),
.B(n_36),
.Y(n_58)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

BUFx2_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_45),
.A2(n_21),
.B1(n_20),
.B2(n_19),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_32),
.B(n_23),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_46),
.B(n_53),
.Y(n_72)
);

AO21x1_ASAP7_75t_L g48 ( 
.A1(n_30),
.A2(n_23),
.B(n_18),
.Y(n_48)
);

OR2x2_ASAP7_75t_L g71 ( 
.A(n_48),
.B(n_1),
.Y(n_71)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_51),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_52),
.B(n_13),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_40),
.B(n_21),
.Y(n_53)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

CKINVDCx14_ASAP7_75t_R g60 ( 
.A(n_58),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_59),
.B(n_61),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_41),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_55),
.A2(n_37),
.B1(n_17),
.B2(n_13),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_62),
.A2(n_64),
.B1(n_68),
.B2(n_71),
.Y(n_82)
);

AND2x6_ASAP7_75t_L g65 ( 
.A(n_52),
.B(n_9),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_65),
.B(n_66),
.Y(n_77)
);

NOR2x1_ASAP7_75t_L g66 ( 
.A(n_48),
.B(n_20),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_55),
.A2(n_19),
.B1(n_14),
.B2(n_3),
.Y(n_67)
);

INVx1_ASAP7_75t_SL g85 ( 
.A(n_67),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_42),
.A2(n_14),
.B1(n_2),
.B2(n_1),
.Y(n_68)
);

INVx13_ASAP7_75t_L g73 ( 
.A(n_54),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_73),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g74 ( 
.A1(n_47),
.A2(n_43),
.B(n_42),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_74),
.B(n_49),
.Y(n_80)
);

CKINVDCx5p33_ASAP7_75t_R g75 ( 
.A(n_51),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_75),
.B(n_47),
.Y(n_83)
);

XOR2xp5_ASAP7_75t_L g78 ( 
.A(n_72),
.B(n_43),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_78),
.B(n_69),
.C(n_71),
.Y(n_90)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_63),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_79),
.B(n_83),
.Y(n_92)
);

AOI21xp33_ASAP7_75t_SL g100 ( 
.A1(n_80),
.A2(n_88),
.B(n_75),
.Y(n_100)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_74),
.Y(n_81)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_81),
.Y(n_93)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_63),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_84),
.B(n_89),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_60),
.B(n_49),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g91 ( 
.A(n_87),
.B(n_70),
.Y(n_91)
);

OAI32xp33_ASAP7_75t_L g88 ( 
.A1(n_62),
.A2(n_49),
.A3(n_44),
.B1(n_57),
.B2(n_56),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_69),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_90),
.B(n_96),
.C(n_64),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_91),
.B(n_70),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_76),
.B(n_61),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_95),
.B(n_97),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_78),
.B(n_87),
.C(n_81),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_86),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_77),
.B(n_66),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_98),
.B(n_99),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_89),
.B(n_65),
.Y(n_99)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_100),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_93),
.A2(n_80),
.B1(n_82),
.B2(n_88),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_102),
.B(n_104),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_94),
.Y(n_105)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_105),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_92),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_106),
.B(n_90),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_91),
.B(n_79),
.Y(n_108)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_108),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_109),
.B(n_96),
.Y(n_112)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_111),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_112),
.B(n_114),
.C(n_104),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_109),
.B(n_100),
.C(n_70),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_115),
.B(n_105),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_116),
.B(n_119),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_113),
.A2(n_106),
.B1(n_102),
.B2(n_107),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_118),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_110),
.A2(n_107),
.B1(n_101),
.B2(n_85),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_120),
.A2(n_117),
.B(n_112),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_123),
.A2(n_124),
.B(n_85),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_120),
.A2(n_103),
.B(n_114),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_121),
.B(n_108),
.Y(n_125)
);

NOR3xp33_ASAP7_75t_L g128 ( 
.A(n_125),
.B(n_126),
.C(n_127),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_122),
.B(n_68),
.Y(n_127)
);

AOI322xp5_ASAP7_75t_L g129 ( 
.A1(n_125),
.A2(n_73),
.A3(n_50),
.B1(n_9),
.B2(n_11),
.C1(n_8),
.C2(n_7),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_129),
.B(n_7),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_130),
.A2(n_128),
.B1(n_50),
.B2(n_56),
.Y(n_131)
);

OR2x2_ASAP7_75t_L g132 ( 
.A(n_131),
.B(n_57),
.Y(n_132)
);


endmodule