module real_aes_7911_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_766;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_754;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_769;
wire n_434;
wire n_502;
wire n_505;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_756;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_735;
wire n_728;
wire n_713;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_481;
wire n_148;
wire n_498;
wire n_765;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g512 ( .A1(n_0), .A2(n_176), .B(n_513), .C(n_516), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_1), .B(n_508), .Y(n_517) );
INVx1_ASAP7_75t_L g111 ( .A(n_2), .Y(n_111) );
INVx1_ASAP7_75t_L g174 ( .A(n_3), .Y(n_174) );
NAND2xp5_ASAP7_75t_SL g581 ( .A(n_4), .B(n_177), .Y(n_581) );
OAI22xp5_ASAP7_75t_SL g129 ( .A1(n_5), .A2(n_130), .B1(n_133), .B2(n_134), .Y(n_129) );
CKINVDCx20_ASAP7_75t_R g134 ( .A(n_5), .Y(n_134) );
AOI21xp5_ASAP7_75t_L g551 ( .A1(n_6), .A2(n_476), .B(n_552), .Y(n_551) );
AO21x2_ASAP7_75t_L g530 ( .A1(n_7), .A2(n_184), .B(n_531), .Y(n_530) );
AOI22xp33_ASAP7_75t_L g230 ( .A1(n_8), .A2(n_38), .B1(n_164), .B2(n_212), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_9), .B(n_184), .Y(n_192) );
AND2x6_ASAP7_75t_L g179 ( .A(n_10), .B(n_180), .Y(n_179) );
A2O1A1Ixp33_ASAP7_75t_L g524 ( .A1(n_11), .A2(n_179), .B(n_481), .C(n_525), .Y(n_524) );
OAI22xp5_ASAP7_75t_L g130 ( .A1(n_12), .A2(n_42), .B1(n_131), .B2(n_132), .Y(n_130) );
CKINVDCx20_ASAP7_75t_R g131 ( .A(n_12), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_13), .B(n_39), .Y(n_109) );
NOR2xp33_ASAP7_75t_L g126 ( .A(n_13), .B(n_39), .Y(n_126) );
INVx1_ASAP7_75t_L g158 ( .A(n_14), .Y(n_158) );
INVx1_ASAP7_75t_L g155 ( .A(n_15), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_16), .B(n_160), .Y(n_221) );
NAND2xp5_ASAP7_75t_SL g536 ( .A(n_17), .B(n_177), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_18), .B(n_151), .Y(n_258) );
AO32x2_ASAP7_75t_L g228 ( .A1(n_19), .A2(n_150), .A3(n_184), .B1(n_203), .B2(n_229), .Y(n_228) );
AOI222xp33_ASAP7_75t_SL g128 ( .A1(n_20), .A2(n_129), .B1(n_135), .B2(n_754), .C1(n_755), .C2(n_757), .Y(n_128) );
NAND2xp5_ASAP7_75t_SL g225 ( .A(n_21), .B(n_164), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_22), .B(n_151), .Y(n_181) );
AOI22xp33_ASAP7_75t_L g231 ( .A1(n_23), .A2(n_57), .B1(n_164), .B2(n_212), .Y(n_231) );
CKINVDCx20_ASAP7_75t_R g127 ( .A(n_24), .Y(n_127) );
AOI22xp33_ASAP7_75t_SL g214 ( .A1(n_25), .A2(n_84), .B1(n_160), .B2(n_164), .Y(n_214) );
NAND2xp5_ASAP7_75t_SL g244 ( .A(n_26), .B(n_164), .Y(n_244) );
A2O1A1Ixp33_ASAP7_75t_L g498 ( .A1(n_27), .A2(n_203), .B(n_481), .C(n_499), .Y(n_498) );
A2O1A1Ixp33_ASAP7_75t_L g533 ( .A1(n_28), .A2(n_203), .B(n_481), .C(n_534), .Y(n_533) );
BUFx6f_ASAP7_75t_L g169 ( .A(n_29), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_30), .B(n_205), .Y(n_204) );
AOI21xp5_ASAP7_75t_L g509 ( .A1(n_31), .A2(n_476), .B(n_510), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_32), .B(n_205), .Y(n_246) );
INVx2_ASAP7_75t_L g162 ( .A(n_33), .Y(n_162) );
A2O1A1Ixp33_ASAP7_75t_L g478 ( .A1(n_34), .A2(n_479), .B(n_483), .C(n_489), .Y(n_478) );
NAND2xp5_ASAP7_75t_SL g196 ( .A(n_35), .B(n_164), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_36), .B(n_205), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_37), .B(n_223), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_40), .B(n_497), .Y(n_496) );
CKINVDCx20_ASAP7_75t_R g529 ( .A(n_41), .Y(n_529) );
INVx1_ASAP7_75t_L g132 ( .A(n_42), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_43), .B(n_177), .Y(n_546) );
OAI22xp5_ASAP7_75t_SL g767 ( .A1(n_44), .A2(n_768), .B1(n_770), .B2(n_771), .Y(n_767) );
CKINVDCx20_ASAP7_75t_R g770 ( .A(n_44), .Y(n_770) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_45), .B(n_476), .Y(n_532) );
OAI22xp5_ASAP7_75t_SL g137 ( .A1(n_46), .A2(n_138), .B1(n_139), .B2(n_460), .Y(n_137) );
INVx1_ASAP7_75t_L g460 ( .A(n_46), .Y(n_460) );
OAI22xp5_ASAP7_75t_SL g768 ( .A1(n_46), .A2(n_48), .B1(n_460), .B2(n_769), .Y(n_768) );
A2O1A1Ixp33_ASAP7_75t_L g543 ( .A1(n_47), .A2(n_479), .B(n_489), .C(n_544), .Y(n_543) );
CKINVDCx20_ASAP7_75t_R g769 ( .A(n_48), .Y(n_769) );
NAND2xp5_ASAP7_75t_SL g187 ( .A(n_49), .B(n_164), .Y(n_187) );
INVx1_ASAP7_75t_L g514 ( .A(n_50), .Y(n_514) );
AOI22xp33_ASAP7_75t_L g211 ( .A1(n_51), .A2(n_93), .B1(n_212), .B2(n_213), .Y(n_211) );
INVx1_ASAP7_75t_L g545 ( .A(n_52), .Y(n_545) );
NAND2xp5_ASAP7_75t_SL g190 ( .A(n_53), .B(n_164), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_54), .B(n_164), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_55), .B(n_476), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_56), .B(n_172), .Y(n_191) );
AOI22xp33_ASAP7_75t_SL g256 ( .A1(n_58), .A2(n_62), .B1(n_160), .B2(n_164), .Y(n_256) );
CKINVDCx20_ASAP7_75t_R g504 ( .A(n_59), .Y(n_504) );
NAND2xp5_ASAP7_75t_SL g200 ( .A(n_60), .B(n_164), .Y(n_200) );
NAND2xp5_ASAP7_75t_SL g220 ( .A(n_61), .B(n_164), .Y(n_220) );
INVx1_ASAP7_75t_L g180 ( .A(n_63), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_64), .B(n_476), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_65), .B(n_508), .Y(n_557) );
A2O1A1Ixp33_ASAP7_75t_L g554 ( .A1(n_66), .A2(n_166), .B(n_172), .C(n_555), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_67), .B(n_164), .Y(n_175) );
INVx1_ASAP7_75t_L g154 ( .A(n_68), .Y(n_154) );
AOI22xp33_ASAP7_75t_L g104 ( .A1(n_69), .A2(n_105), .B1(n_115), .B2(n_775), .Y(n_104) );
OAI22xp33_ASAP7_75t_SL g764 ( .A1(n_70), .A2(n_765), .B1(n_772), .B2(n_773), .Y(n_764) );
CKINVDCx20_ASAP7_75t_R g772 ( .A(n_70), .Y(n_772) );
CKINVDCx20_ASAP7_75t_R g120 ( .A(n_71), .Y(n_120) );
NAND2xp5_ASAP7_75t_SL g487 ( .A(n_72), .B(n_177), .Y(n_487) );
AO32x2_ASAP7_75t_L g209 ( .A1(n_73), .A2(n_184), .A3(n_203), .B1(n_210), .B2(n_215), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_74), .B(n_178), .Y(n_526) );
INVx1_ASAP7_75t_L g199 ( .A(n_75), .Y(n_199) );
INVx1_ASAP7_75t_L g241 ( .A(n_76), .Y(n_241) );
CKINVDCx16_ASAP7_75t_R g511 ( .A(n_77), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_78), .B(n_486), .Y(n_500) );
A2O1A1Ixp33_ASAP7_75t_L g578 ( .A1(n_79), .A2(n_481), .B(n_489), .C(n_579), .Y(n_578) );
NAND2xp5_ASAP7_75t_SL g242 ( .A(n_80), .B(n_160), .Y(n_242) );
CKINVDCx16_ASAP7_75t_R g553 ( .A(n_81), .Y(n_553) );
INVx1_ASAP7_75t_L g114 ( .A(n_82), .Y(n_114) );
NAND2xp5_ASAP7_75t_SL g501 ( .A(n_83), .B(n_485), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_85), .B(n_212), .Y(n_226) );
CKINVDCx20_ASAP7_75t_R g492 ( .A(n_86), .Y(n_492) );
NAND2xp5_ASAP7_75t_SL g245 ( .A(n_87), .B(n_160), .Y(n_245) );
INVx2_ASAP7_75t_L g152 ( .A(n_88), .Y(n_152) );
CKINVDCx20_ASAP7_75t_R g585 ( .A(n_89), .Y(n_585) );
NAND2xp5_ASAP7_75t_SL g527 ( .A(n_90), .B(n_202), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_91), .B(n_160), .Y(n_188) );
NAND3xp33_ASAP7_75t_SL g110 ( .A(n_92), .B(n_111), .C(n_112), .Y(n_110) );
OR2x2_ASAP7_75t_L g123 ( .A(n_92), .B(n_124), .Y(n_123) );
OR2x2_ASAP7_75t_L g463 ( .A(n_92), .B(n_125), .Y(n_463) );
INVx2_ASAP7_75t_L g467 ( .A(n_92), .Y(n_467) );
AOI22xp33_ASAP7_75t_L g255 ( .A1(n_94), .A2(n_103), .B1(n_160), .B2(n_161), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_95), .B(n_476), .Y(n_475) );
INVx1_ASAP7_75t_L g484 ( .A(n_96), .Y(n_484) );
INVxp67_ASAP7_75t_L g556 ( .A(n_97), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_98), .B(n_160), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g113 ( .A(n_99), .B(n_114), .Y(n_113) );
INVx1_ASAP7_75t_L g522 ( .A(n_100), .Y(n_522) );
INVx1_ASAP7_75t_L g580 ( .A(n_101), .Y(n_580) );
AND2x2_ASAP7_75t_L g547 ( .A(n_102), .B(n_205), .Y(n_547) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
CKINVDCx20_ASAP7_75t_R g775 ( .A(n_107), .Y(n_775) );
CKINVDCx12_ASAP7_75t_R g107 ( .A(n_108), .Y(n_107) );
OR2x2_ASAP7_75t_L g108 ( .A(n_109), .B(n_110), .Y(n_108) );
AND2x2_ASAP7_75t_L g125 ( .A(n_111), .B(n_126), .Y(n_125) );
INVx1_ASAP7_75t_SL g112 ( .A(n_113), .Y(n_112) );
BUFx3_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
AOI22xp5_ASAP7_75t_L g116 ( .A1(n_117), .A2(n_128), .B1(n_760), .B2(n_763), .Y(n_116) );
NOR2xp33_ASAP7_75t_L g117 ( .A(n_118), .B(n_121), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx2_ASAP7_75t_L g762 ( .A(n_120), .Y(n_762) );
AOI21xp5_ASAP7_75t_L g763 ( .A1(n_121), .A2(n_764), .B(n_774), .Y(n_763) );
NOR2xp33_ASAP7_75t_SL g121 ( .A(n_122), .B(n_127), .Y(n_121) );
HB1xp67_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
HB1xp67_ASAP7_75t_L g774 ( .A(n_123), .Y(n_774) );
NOR2x2_ASAP7_75t_L g759 ( .A(n_124), .B(n_467), .Y(n_759) );
INVx2_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
OR2x2_ASAP7_75t_L g466 ( .A(n_125), .B(n_467), .Y(n_466) );
INVx1_ASAP7_75t_L g754 ( .A(n_129), .Y(n_754) );
CKINVDCx14_ASAP7_75t_R g133 ( .A(n_130), .Y(n_133) );
OAI22x1_ASAP7_75t_SL g135 ( .A1(n_136), .A2(n_461), .B1(n_464), .B2(n_468), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
OAI22xp5_ASAP7_75t_SL g755 ( .A1(n_137), .A2(n_461), .B1(n_466), .B2(n_756), .Y(n_755) );
OAI22xp5_ASAP7_75t_SL g765 ( .A1(n_138), .A2(n_139), .B1(n_766), .B2(n_767), .Y(n_765) );
INVx1_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
AND2x2_ASAP7_75t_SL g139 ( .A(n_140), .B(n_426), .Y(n_139) );
NOR3xp33_ASAP7_75t_L g140 ( .A(n_141), .B(n_330), .C(n_414), .Y(n_140) );
NAND4xp25_ASAP7_75t_L g141 ( .A(n_142), .B(n_273), .C(n_295), .D(n_311), .Y(n_141) );
AOI221xp5_ASAP7_75t_L g142 ( .A1(n_143), .A2(n_206), .B1(n_232), .B2(n_251), .C(n_259), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g144 ( .A(n_145), .B(n_182), .Y(n_144) );
NAND2xp5_ASAP7_75t_SL g285 ( .A(n_145), .B(n_251), .Y(n_285) );
NAND4xp25_ASAP7_75t_L g325 ( .A(n_145), .B(n_313), .C(n_326), .D(n_328), .Y(n_325) );
INVxp67_ASAP7_75t_L g442 ( .A(n_145), .Y(n_442) );
INVx3_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
OR2x2_ASAP7_75t_L g324 ( .A(n_146), .B(n_262), .Y(n_324) );
AND2x2_ASAP7_75t_L g348 ( .A(n_146), .B(n_182), .Y(n_348) );
INVx2_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
AND2x2_ASAP7_75t_L g315 ( .A(n_147), .B(n_250), .Y(n_315) );
AND2x2_ASAP7_75t_L g355 ( .A(n_147), .B(n_336), .Y(n_355) );
AND2x2_ASAP7_75t_L g372 ( .A(n_147), .B(n_373), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_147), .B(n_183), .Y(n_396) );
INVx2_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
AND2x2_ASAP7_75t_L g249 ( .A(n_148), .B(n_250), .Y(n_249) );
AND2x2_ASAP7_75t_L g267 ( .A(n_148), .B(n_268), .Y(n_267) );
AND2x2_ASAP7_75t_L g279 ( .A(n_148), .B(n_183), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_148), .B(n_193), .Y(n_301) );
OA21x2_ASAP7_75t_L g148 ( .A1(n_149), .A2(n_156), .B(n_181), .Y(n_148) );
OA21x2_ASAP7_75t_L g193 ( .A1(n_149), .A2(n_194), .B(n_204), .Y(n_193) );
INVx2_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
NOR2xp33_ASAP7_75t_L g528 ( .A(n_150), .B(n_529), .Y(n_528) );
INVx1_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
BUFx6f_ASAP7_75t_L g184 ( .A(n_151), .Y(n_184) );
AND2x2_ASAP7_75t_L g151 ( .A(n_152), .B(n_153), .Y(n_151) );
AND2x2_ASAP7_75t_SL g205 ( .A(n_152), .B(n_153), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g153 ( .A(n_154), .B(n_155), .Y(n_153) );
OAI21xp5_ASAP7_75t_L g156 ( .A1(n_157), .A2(n_170), .B(n_179), .Y(n_156) );
O2A1O1Ixp33_ASAP7_75t_L g157 ( .A1(n_158), .A2(n_159), .B(n_163), .C(n_166), .Y(n_157) );
AOI21xp5_ASAP7_75t_L g525 ( .A1(n_159), .A2(n_526), .B(n_527), .Y(n_525) );
AOI21xp5_ASAP7_75t_L g534 ( .A1(n_159), .A2(n_535), .B(n_536), .Y(n_534) );
INVx2_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
INVx3_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
INVx2_ASAP7_75t_L g165 ( .A(n_162), .Y(n_165) );
INVx1_ASAP7_75t_L g173 ( .A(n_162), .Y(n_173) );
INVx3_ASAP7_75t_L g240 ( .A(n_164), .Y(n_240) );
HB1xp67_ASAP7_75t_L g582 ( .A(n_164), .Y(n_582) );
BUFx6f_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
INVx1_ASAP7_75t_L g212 ( .A(n_165), .Y(n_212) );
BUFx3_ASAP7_75t_L g213 ( .A(n_165), .Y(n_213) );
AND2x6_ASAP7_75t_L g481 ( .A(n_165), .B(n_482), .Y(n_481) );
O2A1O1Ixp33_ASAP7_75t_L g579 ( .A1(n_166), .A2(n_580), .B(n_581), .C(n_582), .Y(n_579) );
INVx1_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
AOI21xp5_ASAP7_75t_L g243 ( .A1(n_167), .A2(n_244), .B(n_245), .Y(n_243) );
INVx4_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
INVx2_ASAP7_75t_L g486 ( .A(n_168), .Y(n_486) );
BUFx6f_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
INVx3_ASAP7_75t_L g178 ( .A(n_169), .Y(n_178) );
BUFx6f_ASAP7_75t_L g202 ( .A(n_169), .Y(n_202) );
INVx1_ASAP7_75t_L g223 ( .A(n_169), .Y(n_223) );
AND2x2_ASAP7_75t_L g477 ( .A(n_169), .B(n_173), .Y(n_477) );
INVx1_ASAP7_75t_L g482 ( .A(n_169), .Y(n_482) );
O2A1O1Ixp33_ASAP7_75t_L g170 ( .A1(n_171), .A2(n_174), .B(n_175), .C(n_176), .Y(n_170) );
O2A1O1Ixp5_ASAP7_75t_L g198 ( .A1(n_171), .A2(n_199), .B(n_200), .C(n_201), .Y(n_198) );
AOI21xp5_ASAP7_75t_L g499 ( .A1(n_171), .A2(n_500), .B(n_501), .Y(n_499) );
INVx2_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
AOI21xp5_ASAP7_75t_L g189 ( .A1(n_176), .A2(n_190), .B(n_191), .Y(n_189) );
OAI22xp5_ASAP7_75t_L g229 ( .A1(n_176), .A2(n_202), .B1(n_230), .B2(n_231), .Y(n_229) );
OAI22xp5_ASAP7_75t_L g254 ( .A1(n_176), .A2(n_202), .B1(n_255), .B2(n_256), .Y(n_254) );
INVx2_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
AOI21xp5_ASAP7_75t_L g186 ( .A1(n_177), .A2(n_187), .B(n_188), .Y(n_186) );
AOI21xp5_ASAP7_75t_L g195 ( .A1(n_177), .A2(n_196), .B(n_197), .Y(n_195) );
O2A1O1Ixp5_ASAP7_75t_SL g239 ( .A1(n_177), .A2(n_240), .B(n_241), .C(n_242), .Y(n_239) );
NOR2xp33_ASAP7_75t_L g555 ( .A(n_177), .B(n_556), .Y(n_555) );
INVx5_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
OAI22xp5_ASAP7_75t_SL g210 ( .A1(n_178), .A2(n_202), .B1(n_211), .B2(n_214), .Y(n_210) );
OAI21xp5_ASAP7_75t_L g185 ( .A1(n_179), .A2(n_186), .B(n_189), .Y(n_185) );
BUFx3_ASAP7_75t_L g203 ( .A(n_179), .Y(n_203) );
OAI21xp5_ASAP7_75t_L g218 ( .A1(n_179), .A2(n_219), .B(n_224), .Y(n_218) );
OAI21xp5_ASAP7_75t_L g238 ( .A1(n_179), .A2(n_239), .B(n_243), .Y(n_238) );
AND2x4_ASAP7_75t_L g476 ( .A(n_179), .B(n_477), .Y(n_476) );
INVx4_ASAP7_75t_SL g490 ( .A(n_179), .Y(n_490) );
NAND2x1p5_ASAP7_75t_L g523 ( .A(n_179), .B(n_477), .Y(n_523) );
AND2x2_ASAP7_75t_L g282 ( .A(n_182), .B(n_283), .Y(n_282) );
AOI221xp5_ASAP7_75t_L g331 ( .A1(n_182), .A2(n_332), .B1(n_335), .B2(n_337), .C(n_341), .Y(n_331) );
AND2x2_ASAP7_75t_L g390 ( .A(n_182), .B(n_355), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_182), .B(n_372), .Y(n_424) );
AND2x2_ASAP7_75t_L g182 ( .A(n_183), .B(n_193), .Y(n_182) );
INVx3_ASAP7_75t_L g250 ( .A(n_183), .Y(n_250) );
AND2x2_ASAP7_75t_L g299 ( .A(n_183), .B(n_300), .Y(n_299) );
AND2x2_ASAP7_75t_L g353 ( .A(n_183), .B(n_268), .Y(n_353) );
AND2x2_ASAP7_75t_L g411 ( .A(n_183), .B(n_412), .Y(n_411) );
OA21x2_ASAP7_75t_L g183 ( .A1(n_184), .A2(n_185), .B(n_192), .Y(n_183) );
INVx4_ASAP7_75t_L g253 ( .A(n_184), .Y(n_253) );
AOI21xp5_ASAP7_75t_L g531 ( .A1(n_184), .A2(n_532), .B(n_533), .Y(n_531) );
HB1xp67_ASAP7_75t_L g550 ( .A(n_184), .Y(n_550) );
AND2x2_ASAP7_75t_L g251 ( .A(n_193), .B(n_252), .Y(n_251) );
INVx2_ASAP7_75t_L g268 ( .A(n_193), .Y(n_268) );
INVx1_ASAP7_75t_L g323 ( .A(n_193), .Y(n_323) );
HB1xp67_ASAP7_75t_L g329 ( .A(n_193), .Y(n_329) );
AND2x2_ASAP7_75t_L g374 ( .A(n_193), .B(n_250), .Y(n_374) );
OR2x2_ASAP7_75t_L g413 ( .A(n_193), .B(n_252), .Y(n_413) );
OAI21xp5_ASAP7_75t_L g194 ( .A1(n_195), .A2(n_198), .B(n_203), .Y(n_194) );
AOI21xp5_ASAP7_75t_L g224 ( .A1(n_201), .A2(n_225), .B(n_226), .Y(n_224) );
INVx2_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
INVx4_ASAP7_75t_L g515 ( .A(n_202), .Y(n_515) );
NAND3xp33_ASAP7_75t_L g272 ( .A(n_203), .B(n_253), .C(n_254), .Y(n_272) );
INVx2_ASAP7_75t_L g215 ( .A(n_205), .Y(n_215) );
OA21x2_ASAP7_75t_L g217 ( .A1(n_205), .A2(n_218), .B(n_227), .Y(n_217) );
OA21x2_ASAP7_75t_L g237 ( .A1(n_205), .A2(n_238), .B(n_246), .Y(n_237) );
AOI21xp5_ASAP7_75t_L g474 ( .A1(n_205), .A2(n_475), .B(n_478), .Y(n_474) );
INVx1_ASAP7_75t_L g505 ( .A(n_205), .Y(n_505) );
AOI21xp5_ASAP7_75t_L g541 ( .A1(n_205), .A2(n_542), .B(n_543), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_206), .B(n_293), .Y(n_292) );
AND2x2_ASAP7_75t_L g206 ( .A(n_207), .B(n_216), .Y(n_206) );
AND2x2_ASAP7_75t_L g409 ( .A(n_207), .B(n_406), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_207), .B(n_391), .Y(n_441) );
BUFx2_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
AND2x2_ASAP7_75t_L g340 ( .A(n_208), .B(n_264), .Y(n_340) );
AND2x2_ASAP7_75t_L g389 ( .A(n_208), .B(n_235), .Y(n_389) );
INVx1_ASAP7_75t_L g435 ( .A(n_208), .Y(n_435) );
INVx1_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
BUFx6f_ASAP7_75t_L g248 ( .A(n_209), .Y(n_248) );
AND2x2_ASAP7_75t_L g290 ( .A(n_209), .B(n_264), .Y(n_290) );
INVx1_ASAP7_75t_L g307 ( .A(n_209), .Y(n_307) );
AND2x2_ASAP7_75t_L g313 ( .A(n_209), .B(n_228), .Y(n_313) );
HB1xp67_ASAP7_75t_L g488 ( .A(n_213), .Y(n_488) );
INVx2_ASAP7_75t_L g516 ( .A(n_213), .Y(n_516) );
INVx1_ASAP7_75t_L g502 ( .A(n_215), .Y(n_502) );
AND2x2_ASAP7_75t_L g381 ( .A(n_216), .B(n_289), .Y(n_381) );
INVx2_ASAP7_75t_L g446 ( .A(n_216), .Y(n_446) );
AND2x2_ASAP7_75t_L g216 ( .A(n_217), .B(n_228), .Y(n_216) );
AND2x2_ASAP7_75t_L g263 ( .A(n_217), .B(n_264), .Y(n_263) );
OR2x2_ASAP7_75t_L g276 ( .A(n_217), .B(n_236), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_217), .B(n_235), .Y(n_304) );
INVx1_ASAP7_75t_L g310 ( .A(n_217), .Y(n_310) );
INVx1_ASAP7_75t_L g327 ( .A(n_217), .Y(n_327) );
HB1xp67_ASAP7_75t_L g339 ( .A(n_217), .Y(n_339) );
INVx2_ASAP7_75t_L g407 ( .A(n_217), .Y(n_407) );
AOI21xp5_ASAP7_75t_L g219 ( .A1(n_220), .A2(n_221), .B(n_222), .Y(n_219) );
INVx1_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
INVx2_ASAP7_75t_L g264 ( .A(n_228), .Y(n_264) );
BUFx2_ASAP7_75t_L g361 ( .A(n_228), .Y(n_361) );
AND2x2_ASAP7_75t_L g406 ( .A(n_228), .B(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_234), .B(n_247), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_234), .B(n_343), .Y(n_342) );
AOI21xp5_ASAP7_75t_L g429 ( .A1(n_234), .A2(n_405), .B(n_419), .Y(n_429) );
AND2x2_ASAP7_75t_L g454 ( .A(n_234), .B(n_340), .Y(n_454) );
BUFx2_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
INVx2_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
INVx1_ASAP7_75t_L g376 ( .A(n_236), .Y(n_376) );
AND2x2_ASAP7_75t_L g405 ( .A(n_236), .B(n_406), .Y(n_405) );
INVx2_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
HB1xp67_ASAP7_75t_L g289 ( .A(n_237), .Y(n_289) );
INVx2_ASAP7_75t_L g308 ( .A(n_237), .Y(n_308) );
OR2x2_ASAP7_75t_L g309 ( .A(n_237), .B(n_310), .Y(n_309) );
AND2x2_ASAP7_75t_L g247 ( .A(n_248), .B(n_249), .Y(n_247) );
INVx2_ASAP7_75t_L g262 ( .A(n_248), .Y(n_262) );
OR2x2_ASAP7_75t_L g275 ( .A(n_248), .B(n_276), .Y(n_275) );
AND2x2_ASAP7_75t_L g343 ( .A(n_248), .B(n_339), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_248), .B(n_439), .Y(n_438) );
OR2x2_ASAP7_75t_L g444 ( .A(n_248), .B(n_445), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_248), .B(n_381), .Y(n_456) );
AND2x2_ASAP7_75t_L g335 ( .A(n_249), .B(n_336), .Y(n_335) );
AND2x2_ASAP7_75t_L g358 ( .A(n_249), .B(n_251), .Y(n_358) );
INVx2_ASAP7_75t_L g270 ( .A(n_250), .Y(n_270) );
AND2x2_ASAP7_75t_L g298 ( .A(n_250), .B(n_271), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_250), .B(n_323), .Y(n_379) );
AND2x2_ASAP7_75t_L g293 ( .A(n_251), .B(n_294), .Y(n_293) );
INVx1_ASAP7_75t_L g440 ( .A(n_251), .Y(n_440) );
AND2x2_ASAP7_75t_L g452 ( .A(n_251), .B(n_315), .Y(n_452) );
AND2x2_ASAP7_75t_L g278 ( .A(n_252), .B(n_268), .Y(n_278) );
INVx1_ASAP7_75t_L g373 ( .A(n_252), .Y(n_373) );
AO21x1_ASAP7_75t_L g252 ( .A1(n_253), .A2(n_254), .B(n_257), .Y(n_252) );
NOR2xp33_ASAP7_75t_L g491 ( .A(n_253), .B(n_492), .Y(n_491) );
INVx3_ASAP7_75t_L g508 ( .A(n_253), .Y(n_508) );
AO21x2_ASAP7_75t_L g520 ( .A1(n_253), .A2(n_521), .B(n_528), .Y(n_520) );
AO21x2_ASAP7_75t_L g576 ( .A1(n_253), .A2(n_577), .B(n_584), .Y(n_576) );
NOR2xp33_ASAP7_75t_L g584 ( .A(n_253), .B(n_585), .Y(n_584) );
INVx1_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
AND2x4_ASAP7_75t_L g271 ( .A(n_258), .B(n_272), .Y(n_271) );
INVxp67_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_261), .B(n_265), .Y(n_260) );
AND2x2_ASAP7_75t_L g261 ( .A(n_262), .B(n_263), .Y(n_261) );
NOR2xp33_ASAP7_75t_L g318 ( .A(n_262), .B(n_309), .Y(n_318) );
OR2x2_ASAP7_75t_L g450 ( .A(n_262), .B(n_451), .Y(n_450) );
AND2x2_ASAP7_75t_L g367 ( .A(n_263), .B(n_308), .Y(n_367) );
AND2x2_ASAP7_75t_L g375 ( .A(n_263), .B(n_376), .Y(n_375) );
AND2x2_ASAP7_75t_L g434 ( .A(n_263), .B(n_435), .Y(n_434) );
AND2x2_ASAP7_75t_L g458 ( .A(n_263), .B(n_305), .Y(n_458) );
NOR2xp67_ASAP7_75t_L g416 ( .A(n_264), .B(n_417), .Y(n_416) );
OR2x2_ASAP7_75t_L g445 ( .A(n_264), .B(n_308), .Y(n_445) );
INVx1_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
NAND2x1p5_ASAP7_75t_L g266 ( .A(n_267), .B(n_269), .Y(n_266) );
AND2x2_ASAP7_75t_L g297 ( .A(n_267), .B(n_298), .Y(n_297) );
INVxp67_ASAP7_75t_L g459 ( .A(n_267), .Y(n_459) );
NOR2x1_ASAP7_75t_L g269 ( .A(n_270), .B(n_271), .Y(n_269) );
INVx1_ASAP7_75t_L g294 ( .A(n_270), .Y(n_294) );
AND2x2_ASAP7_75t_L g345 ( .A(n_270), .B(n_278), .Y(n_345) );
NOR2xp33_ASAP7_75t_L g439 ( .A(n_270), .B(n_413), .Y(n_439) );
INVx2_ASAP7_75t_L g284 ( .A(n_271), .Y(n_284) );
INVx3_ASAP7_75t_L g336 ( .A(n_271), .Y(n_336) );
OR2x2_ASAP7_75t_L g364 ( .A(n_271), .B(n_365), .Y(n_364) );
AOI311xp33_ASAP7_75t_L g273 ( .A1(n_274), .A2(n_277), .A3(n_279), .B(n_280), .C(n_291), .Y(n_273) );
O2A1O1Ixp33_ASAP7_75t_L g311 ( .A1(n_274), .A2(n_312), .B(n_314), .C(n_316), .Y(n_311) );
INVx2_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
INVx2_ASAP7_75t_SL g296 ( .A(n_276), .Y(n_296) );
INVx2_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
AND2x2_ASAP7_75t_L g314 ( .A(n_278), .B(n_315), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_278), .B(n_294), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_278), .B(n_279), .Y(n_447) );
AND2x2_ASAP7_75t_L g369 ( .A(n_279), .B(n_283), .Y(n_369) );
AOI21xp33_ASAP7_75t_L g280 ( .A1(n_281), .A2(n_285), .B(n_286), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
AND2x2_ASAP7_75t_L g427 ( .A(n_283), .B(n_315), .Y(n_427) );
INVx2_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
NOR2xp33_ASAP7_75t_L g300 ( .A(n_284), .B(n_301), .Y(n_300) );
INVx1_ASAP7_75t_L g321 ( .A(n_284), .Y(n_321) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
AND2x2_ASAP7_75t_L g287 ( .A(n_288), .B(n_290), .Y(n_287) );
AND2x2_ASAP7_75t_L g312 ( .A(n_288), .B(n_313), .Y(n_312) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
INVx1_ASAP7_75t_L g357 ( .A(n_290), .Y(n_357) );
AND2x4_ASAP7_75t_L g419 ( .A(n_290), .B(n_388), .Y(n_419) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
AOI222xp33_ASAP7_75t_L g370 ( .A1(n_293), .A2(n_359), .B1(n_371), .B2(n_375), .C1(n_377), .C2(n_381), .Y(n_370) );
A2O1A1Ixp33_ASAP7_75t_L g295 ( .A1(n_296), .A2(n_297), .B(n_299), .C(n_302), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_296), .B(n_340), .Y(n_363) );
INVx1_ASAP7_75t_L g385 ( .A(n_298), .Y(n_385) );
INVx1_ASAP7_75t_L g319 ( .A(n_300), .Y(n_319) );
OR2x2_ASAP7_75t_L g384 ( .A(n_301), .B(n_385), .Y(n_384) );
OAI21xp33_ASAP7_75t_SL g302 ( .A1(n_303), .A2(n_305), .B(n_309), .Y(n_302) );
NAND3xp33_ASAP7_75t_L g320 ( .A(n_303), .B(n_321), .C(n_322), .Y(n_320) );
AOI21xp5_ASAP7_75t_L g418 ( .A1(n_303), .A2(n_340), .B(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
INVx1_ASAP7_75t_SL g305 ( .A(n_306), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_307), .B(n_308), .Y(n_306) );
HB1xp67_ASAP7_75t_L g360 ( .A(n_307), .Y(n_360) );
AND2x2_ASAP7_75t_SL g326 ( .A(n_308), .B(n_327), .Y(n_326) );
INVx1_ASAP7_75t_L g417 ( .A(n_308), .Y(n_417) );
HB1xp67_ASAP7_75t_L g433 ( .A(n_308), .Y(n_433) );
INVx2_ASAP7_75t_L g391 ( .A(n_309), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_313), .B(n_334), .Y(n_333) );
INVx2_ASAP7_75t_L g365 ( .A(n_315), .Y(n_365) );
OAI221xp5_ASAP7_75t_L g316 ( .A1(n_317), .A2(n_319), .B1(n_320), .B2(n_324), .C(n_325), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
NAND2xp5_ASAP7_75t_SL g398 ( .A(n_319), .B(n_399), .Y(n_398) );
INVx1_ASAP7_75t_SL g453 ( .A(n_319), .Y(n_453) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
INVx2_ASAP7_75t_L g334 ( .A(n_326), .Y(n_334) );
NOR2xp33_ASAP7_75t_L g356 ( .A(n_326), .B(n_357), .Y(n_356) );
AND2x2_ASAP7_75t_L g392 ( .A(n_326), .B(n_340), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_326), .B(n_402), .Y(n_401) );
AND2x2_ASAP7_75t_L g425 ( .A(n_326), .B(n_360), .Y(n_425) );
BUFx3_ASAP7_75t_L g388 ( .A(n_327), .Y(n_388) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
NAND5xp2_ASAP7_75t_L g330 ( .A(n_331), .B(n_349), .C(n_370), .D(n_382), .E(n_397), .Y(n_330) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
AOI32xp33_ASAP7_75t_L g422 ( .A1(n_334), .A2(n_361), .A3(n_377), .B1(n_423), .B2(n_425), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_336), .B(n_395), .Y(n_394) );
AND2x2_ASAP7_75t_L g337 ( .A(n_338), .B(n_340), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
INVx1_ASAP7_75t_SL g346 ( .A(n_340), .Y(n_346) );
OAI22xp5_ASAP7_75t_L g341 ( .A1(n_342), .A2(n_344), .B1(n_346), .B2(n_347), .Y(n_341) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
INVx1_ASAP7_75t_SL g347 ( .A(n_348), .Y(n_347) );
AOI221xp5_ASAP7_75t_L g349 ( .A1(n_350), .A2(n_356), .B1(n_358), .B2(n_359), .C(n_362), .Y(n_349) );
INVx2_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
OR2x2_ASAP7_75t_L g351 ( .A(n_352), .B(n_354), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
AND2x2_ASAP7_75t_L g421 ( .A(n_353), .B(n_372), .Y(n_421) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
AOI221xp5_ASAP7_75t_L g436 ( .A1(n_358), .A2(n_419), .B1(n_437), .B2(n_442), .C(n_443), .Y(n_436) );
AND2x2_ASAP7_75t_L g359 ( .A(n_360), .B(n_361), .Y(n_359) );
INVx2_ASAP7_75t_L g402 ( .A(n_361), .Y(n_402) );
OAI22xp5_ASAP7_75t_L g362 ( .A1(n_363), .A2(n_364), .B1(n_366), .B2(n_368), .Y(n_362) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
INVx1_ASAP7_75t_SL g368 ( .A(n_369), .Y(n_368) );
AND2x2_ASAP7_75t_L g371 ( .A(n_372), .B(n_374), .Y(n_371) );
INVx1_ASAP7_75t_L g380 ( .A(n_372), .Y(n_380) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
OR2x2_ASAP7_75t_L g378 ( .A(n_379), .B(n_380), .Y(n_378) );
AOI222xp33_ASAP7_75t_L g382 ( .A1(n_383), .A2(n_386), .B1(n_390), .B2(n_391), .C1(n_392), .C2(n_393), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
AND2x2_ASAP7_75t_L g386 ( .A(n_387), .B(n_389), .Y(n_386) );
INVxp67_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
OAI22xp33_ASAP7_75t_L g437 ( .A1(n_391), .A2(n_438), .B1(n_440), .B2(n_441), .Y(n_437) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx1_ASAP7_75t_SL g395 ( .A(n_396), .Y(n_395) );
AOI21xp5_ASAP7_75t_L g397 ( .A1(n_398), .A2(n_400), .B(n_403), .Y(n_397) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
AOI21xp33_ASAP7_75t_L g403 ( .A1(n_404), .A2(n_408), .B(n_410), .Y(n_403) );
INVx2_ASAP7_75t_SL g404 ( .A(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g451 ( .A(n_406), .Y(n_451) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_SL g412 ( .A(n_413), .Y(n_412) );
A2O1A1Ixp33_ASAP7_75t_L g414 ( .A1(n_415), .A2(n_418), .B(n_420), .C(n_422), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
AOI211xp5_ASAP7_75t_L g426 ( .A1(n_427), .A2(n_428), .B(n_430), .C(n_455), .Y(n_426) );
CKINVDCx16_ASAP7_75t_R g431 ( .A(n_427), .Y(n_431) );
INVxp67_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
OAI211xp5_ASAP7_75t_L g430 ( .A1(n_431), .A2(n_432), .B(n_436), .C(n_448), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_433), .B(n_434), .Y(n_432) );
AOI21xp33_ASAP7_75t_L g443 ( .A1(n_444), .A2(n_446), .B(n_447), .Y(n_443) );
AOI22xp5_ASAP7_75t_L g448 ( .A1(n_449), .A2(n_452), .B1(n_453), .B2(n_454), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
AOI21xp33_ASAP7_75t_L g455 ( .A1(n_456), .A2(n_457), .B(n_459), .Y(n_455) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx2_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx2_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx2_ASAP7_75t_L g756 ( .A(n_468), .Y(n_756) );
OR3x2_ASAP7_75t_L g468 ( .A(n_469), .B(n_668), .C(n_711), .Y(n_468) );
NAND5xp2_ASAP7_75t_L g469 ( .A(n_470), .B(n_595), .C(n_625), .D(n_642), .E(n_657), .Y(n_469) );
AOI221xp5_ASAP7_75t_SL g470 ( .A1(n_471), .A2(n_518), .B1(n_558), .B2(n_564), .C(n_568), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_472), .B(n_493), .Y(n_471) );
OR2x2_ASAP7_75t_L g573 ( .A(n_472), .B(n_574), .Y(n_573) );
AND2x2_ASAP7_75t_L g612 ( .A(n_472), .B(n_613), .Y(n_612) );
AND2x2_ASAP7_75t_L g630 ( .A(n_472), .B(n_631), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_472), .B(n_566), .Y(n_647) );
OR2x2_ASAP7_75t_L g659 ( .A(n_472), .B(n_660), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_472), .B(n_618), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_472), .B(n_692), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_472), .B(n_596), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_472), .B(n_604), .Y(n_710) );
AND2x2_ASAP7_75t_L g742 ( .A(n_472), .B(n_506), .Y(n_742) );
HB1xp67_ASAP7_75t_L g750 ( .A(n_472), .Y(n_750) );
INVx5_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_473), .B(n_566), .Y(n_565) );
AND2x2_ASAP7_75t_L g570 ( .A(n_473), .B(n_548), .Y(n_570) );
BUFx2_ASAP7_75t_L g592 ( .A(n_473), .Y(n_592) );
AND2x2_ASAP7_75t_L g621 ( .A(n_473), .B(n_494), .Y(n_621) );
AND2x2_ASAP7_75t_L g676 ( .A(n_473), .B(n_574), .Y(n_676) );
OR2x6_ASAP7_75t_L g473 ( .A(n_474), .B(n_491), .Y(n_473) );
BUFx2_ASAP7_75t_L g497 ( .A(n_476), .Y(n_497) );
INVx2_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
O2A1O1Ixp33_ASAP7_75t_SL g510 ( .A1(n_480), .A2(n_490), .B(n_511), .C(n_512), .Y(n_510) );
O2A1O1Ixp33_ASAP7_75t_L g552 ( .A1(n_480), .A2(n_490), .B(n_553), .C(n_554), .Y(n_552) );
INVx5_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
O2A1O1Ixp33_ASAP7_75t_L g483 ( .A1(n_484), .A2(n_485), .B(n_487), .C(n_488), .Y(n_483) );
O2A1O1Ixp33_ASAP7_75t_L g544 ( .A1(n_485), .A2(n_488), .B(n_545), .C(n_546), .Y(n_544) );
INVx2_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
INVx1_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_493), .B(n_630), .Y(n_639) );
OAI32xp33_ASAP7_75t_L g653 ( .A1(n_493), .A2(n_589), .A3(n_654), .B1(n_655), .B2(n_656), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_493), .B(n_655), .Y(n_685) );
NOR2xp33_ASAP7_75t_L g696 ( .A(n_493), .B(n_573), .Y(n_696) );
INVx1_ASAP7_75t_SL g725 ( .A(n_493), .Y(n_725) );
NAND4xp25_ASAP7_75t_L g734 ( .A(n_493), .B(n_520), .C(n_676), .D(n_735), .Y(n_734) );
AND2x4_ASAP7_75t_L g493 ( .A(n_494), .B(n_506), .Y(n_493) );
INVx5_ASAP7_75t_L g567 ( .A(n_494), .Y(n_567) );
AND2x2_ASAP7_75t_L g596 ( .A(n_494), .B(n_507), .Y(n_596) );
HB1xp67_ASAP7_75t_L g675 ( .A(n_494), .Y(n_675) );
AND2x2_ASAP7_75t_L g745 ( .A(n_494), .B(n_692), .Y(n_745) );
OR2x6_ASAP7_75t_L g494 ( .A(n_495), .B(n_503), .Y(n_494) );
AOI21xp5_ASAP7_75t_SL g495 ( .A1(n_496), .A2(n_498), .B(n_502), .Y(n_495) );
NOR2xp33_ASAP7_75t_L g503 ( .A(n_504), .B(n_505), .Y(n_503) );
AND2x4_ASAP7_75t_L g618 ( .A(n_506), .B(n_567), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_506), .B(n_628), .Y(n_627) );
AND2x2_ASAP7_75t_L g652 ( .A(n_506), .B(n_574), .Y(n_652) );
INVx2_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
AND2x2_ASAP7_75t_L g566 ( .A(n_507), .B(n_567), .Y(n_566) );
AND2x2_ASAP7_75t_L g604 ( .A(n_507), .B(n_576), .Y(n_604) );
AND2x2_ASAP7_75t_L g613 ( .A(n_507), .B(n_575), .Y(n_613) );
OA21x2_ASAP7_75t_L g507 ( .A1(n_508), .A2(n_509), .B(n_517), .Y(n_507) );
NOR2xp33_ASAP7_75t_L g513 ( .A(n_514), .B(n_515), .Y(n_513) );
AOI222xp33_ASAP7_75t_L g681 ( .A1(n_518), .A2(n_682), .B1(n_684), .B2(n_686), .C1(n_689), .C2(n_690), .Y(n_681) );
AND2x4_ASAP7_75t_L g518 ( .A(n_519), .B(n_537), .Y(n_518) );
AND2x2_ASAP7_75t_L g614 ( .A(n_519), .B(n_615), .Y(n_614) );
NAND3xp33_ASAP7_75t_L g731 ( .A(n_519), .B(n_592), .C(n_732), .Y(n_731) );
AND2x2_ASAP7_75t_L g519 ( .A(n_520), .B(n_530), .Y(n_519) );
INVx5_ASAP7_75t_SL g563 ( .A(n_520), .Y(n_563) );
OAI322xp33_ASAP7_75t_L g568 ( .A1(n_520), .A2(n_569), .A3(n_571), .B1(n_572), .B2(n_586), .C1(n_589), .C2(n_591), .Y(n_568) );
NAND2xp5_ASAP7_75t_SL g634 ( .A(n_520), .B(n_561), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g740 ( .A(n_520), .B(n_549), .Y(n_740) );
OAI21xp5_ASAP7_75t_L g521 ( .A1(n_522), .A2(n_523), .B(n_524), .Y(n_521) );
INVx2_ASAP7_75t_L g561 ( .A(n_530), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_530), .B(n_539), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_537), .B(n_599), .Y(n_654) );
INVx2_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
OR2x2_ASAP7_75t_L g633 ( .A(n_538), .B(n_634), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_539), .B(n_548), .Y(n_538) );
OR2x2_ASAP7_75t_L g562 ( .A(n_539), .B(n_563), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_539), .B(n_570), .Y(n_569) );
OR2x2_ASAP7_75t_L g601 ( .A(n_539), .B(n_549), .Y(n_601) );
AND2x2_ASAP7_75t_L g624 ( .A(n_539), .B(n_561), .Y(n_624) );
NOR2xp33_ASAP7_75t_L g635 ( .A(n_539), .B(n_636), .Y(n_635) );
AND2x2_ASAP7_75t_L g640 ( .A(n_539), .B(n_599), .Y(n_640) );
AND2x2_ASAP7_75t_L g648 ( .A(n_539), .B(n_649), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_539), .B(n_608), .Y(n_698) );
INVx5_ASAP7_75t_SL g539 ( .A(n_540), .Y(n_539) );
AND2x2_ASAP7_75t_L g588 ( .A(n_540), .B(n_563), .Y(n_588) );
OR2x2_ASAP7_75t_L g589 ( .A(n_540), .B(n_590), .Y(n_589) );
AND2x2_ASAP7_75t_L g615 ( .A(n_540), .B(n_549), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_540), .B(n_662), .Y(n_703) );
OR2x2_ASAP7_75t_L g719 ( .A(n_540), .B(n_663), .Y(n_719) );
AND2x2_ASAP7_75t_SL g726 ( .A(n_540), .B(n_680), .Y(n_726) );
HB1xp67_ASAP7_75t_L g733 ( .A(n_540), .Y(n_733) );
OR2x6_ASAP7_75t_L g540 ( .A(n_541), .B(n_547), .Y(n_540) );
AND2x2_ASAP7_75t_L g587 ( .A(n_548), .B(n_588), .Y(n_587) );
AND2x2_ASAP7_75t_L g637 ( .A(n_548), .B(n_561), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_548), .B(n_563), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_548), .B(n_599), .Y(n_721) );
INVx3_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_549), .B(n_563), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_549), .B(n_561), .Y(n_609) );
OR2x2_ASAP7_75t_L g663 ( .A(n_549), .B(n_561), .Y(n_663) );
AND2x2_ASAP7_75t_L g680 ( .A(n_549), .B(n_560), .Y(n_680) );
INVxp67_ASAP7_75t_L g702 ( .A(n_549), .Y(n_702) );
AND2x2_ASAP7_75t_L g729 ( .A(n_549), .B(n_599), .Y(n_729) );
HB1xp67_ASAP7_75t_L g736 ( .A(n_549), .Y(n_736) );
OA21x2_ASAP7_75t_L g549 ( .A1(n_550), .A2(n_551), .B(n_557), .Y(n_549) );
INVx1_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
OR2x2_ASAP7_75t_L g559 ( .A(n_560), .B(n_562), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_560), .B(n_610), .Y(n_683) );
INVx1_ASAP7_75t_SL g560 ( .A(n_561), .Y(n_560) );
AND2x2_ASAP7_75t_L g599 ( .A(n_561), .B(n_563), .Y(n_599) );
OR2x2_ASAP7_75t_L g666 ( .A(n_561), .B(n_667), .Y(n_666) );
INVx2_ASAP7_75t_L g610 ( .A(n_562), .Y(n_610) );
OR2x2_ASAP7_75t_L g671 ( .A(n_562), .B(n_663), .Y(n_671) );
INVx1_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
INVx1_ASAP7_75t_L g571 ( .A(n_566), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_566), .B(n_630), .Y(n_629) );
OR2x2_ASAP7_75t_L g572 ( .A(n_567), .B(n_573), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_567), .B(n_594), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_567), .B(n_574), .Y(n_606) );
INVx2_ASAP7_75t_L g651 ( .A(n_567), .Y(n_651) );
AND2x2_ASAP7_75t_L g664 ( .A(n_567), .B(n_604), .Y(n_664) );
AND2x2_ASAP7_75t_L g689 ( .A(n_567), .B(n_613), .Y(n_689) );
INVx1_ASAP7_75t_L g641 ( .A(n_572), .Y(n_641) );
INVx2_ASAP7_75t_SL g628 ( .A(n_573), .Y(n_628) );
INVx1_ASAP7_75t_L g631 ( .A(n_574), .Y(n_631) );
INVx2_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
HB1xp67_ASAP7_75t_L g594 ( .A(n_575), .Y(n_594) );
INVx2_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
BUFx2_ASAP7_75t_L g692 ( .A(n_576), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_578), .B(n_583), .Y(n_577) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
AND2x2_ASAP7_75t_L g661 ( .A(n_588), .B(n_662), .Y(n_661) );
INVx1_ASAP7_75t_L g667 ( .A(n_588), .Y(n_667) );
AOI22xp5_ASAP7_75t_L g669 ( .A1(n_588), .A2(n_670), .B1(n_672), .B2(n_677), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_588), .B(n_680), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_589), .B(n_683), .Y(n_682) );
INVx1_ASAP7_75t_SL g623 ( .A(n_590), .Y(n_623) );
OR2x2_ASAP7_75t_L g591 ( .A(n_592), .B(n_593), .Y(n_591) );
OR2x2_ASAP7_75t_L g605 ( .A(n_592), .B(n_606), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_592), .B(n_596), .Y(n_656) );
AND2x2_ASAP7_75t_L g679 ( .A(n_592), .B(n_680), .Y(n_679) );
BUFx2_ASAP7_75t_L g655 ( .A(n_594), .Y(n_655) );
AOI211xp5_ASAP7_75t_L g595 ( .A1(n_596), .A2(n_597), .B(n_602), .C(n_616), .Y(n_595) );
INVx1_ASAP7_75t_L g619 ( .A(n_596), .Y(n_619) );
OAI221xp5_ASAP7_75t_SL g727 ( .A1(n_596), .A2(n_728), .B1(n_730), .B2(n_731), .C(n_734), .Y(n_727) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_599), .B(n_600), .Y(n_598) );
INVx1_ASAP7_75t_L g746 ( .A(n_599), .Y(n_746) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
OR2x2_ASAP7_75t_L g695 ( .A(n_601), .B(n_634), .Y(n_695) );
A2O1A1Ixp33_ASAP7_75t_L g602 ( .A1(n_603), .A2(n_605), .B(n_607), .C(n_611), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_608), .B(n_610), .Y(n_607) );
INVx1_ASAP7_75t_SL g608 ( .A(n_609), .Y(n_608) );
OAI32xp33_ASAP7_75t_L g720 ( .A1(n_609), .A2(n_610), .A3(n_673), .B1(n_710), .B2(n_721), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_612), .B(n_614), .Y(n_611) );
AND2x2_ASAP7_75t_L g752 ( .A(n_612), .B(n_651), .Y(n_752) );
AND2x2_ASAP7_75t_L g699 ( .A(n_613), .B(n_651), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_613), .B(n_621), .Y(n_717) );
AOI31xp33_ASAP7_75t_SL g616 ( .A1(n_617), .A2(n_619), .A3(n_620), .B(n_622), .Y(n_616) );
INVxp67_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_618), .B(n_630), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_618), .B(n_628), .Y(n_715) );
AOI221xp5_ASAP7_75t_L g737 ( .A1(n_618), .A2(n_648), .B1(n_738), .B2(n_741), .C(n_743), .Y(n_737) );
CKINVDCx16_ASAP7_75t_R g620 ( .A(n_621), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_623), .B(n_624), .Y(n_622) );
AND2x2_ASAP7_75t_L g643 ( .A(n_623), .B(n_644), .Y(n_643) );
AOI222xp33_ASAP7_75t_L g625 ( .A1(n_626), .A2(n_632), .B1(n_635), .B2(n_638), .C1(n_640), .C2(n_641), .Y(n_625) );
NAND2xp5_ASAP7_75t_SL g626 ( .A(n_627), .B(n_629), .Y(n_626) );
INVx1_ASAP7_75t_L g708 ( .A(n_627), .Y(n_708) );
INVx1_ASAP7_75t_L g730 ( .A(n_630), .Y(n_730) );
INVx2_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
OAI22xp5_ASAP7_75t_L g743 ( .A1(n_633), .A2(n_744), .B1(n_746), .B2(n_747), .Y(n_743) );
INVx1_ASAP7_75t_L g649 ( .A(n_634), .Y(n_649) );
INVx1_ASAP7_75t_SL g636 ( .A(n_637), .Y(n_636) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
AOI221xp5_ASAP7_75t_L g642 ( .A1(n_643), .A2(n_646), .B1(n_648), .B2(n_650), .C(n_653), .Y(n_642) );
INVx1_ASAP7_75t_SL g644 ( .A(n_645), .Y(n_644) );
OR2x2_ASAP7_75t_L g687 ( .A(n_645), .B(n_688), .Y(n_687) );
OR2x2_ASAP7_75t_L g739 ( .A(n_645), .B(n_740), .Y(n_739) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
INVx1_ASAP7_75t_L g714 ( .A(n_650), .Y(n_714) );
AND2x2_ASAP7_75t_L g650 ( .A(n_651), .B(n_652), .Y(n_650) );
INVx1_ASAP7_75t_L g678 ( .A(n_651), .Y(n_678) );
INVx1_ASAP7_75t_L g660 ( .A(n_652), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g747 ( .A(n_655), .B(n_742), .Y(n_747) );
AOI22xp33_ASAP7_75t_L g657 ( .A1(n_658), .A2(n_661), .B1(n_664), .B2(n_665), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
INVx1_ASAP7_75t_SL g662 ( .A(n_663), .Y(n_662) );
INVx1_ASAP7_75t_SL g751 ( .A(n_664), .Y(n_751) );
INVxp33_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
NOR2xp33_ASAP7_75t_L g709 ( .A(n_666), .B(n_710), .Y(n_709) );
OAI32xp33_ASAP7_75t_L g700 ( .A1(n_667), .A2(n_701), .A3(n_702), .B1(n_703), .B2(n_704), .Y(n_700) );
NAND4xp25_ASAP7_75t_L g668 ( .A(n_669), .B(n_681), .C(n_693), .D(n_705), .Y(n_668) );
INVx1_ASAP7_75t_SL g670 ( .A(n_671), .Y(n_670) );
NAND2xp33_ASAP7_75t_SL g672 ( .A(n_673), .B(n_674), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_675), .B(n_676), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_676), .B(n_725), .Y(n_724) );
AND2x2_ASAP7_75t_L g677 ( .A(n_678), .B(n_679), .Y(n_677) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
CKINVDCx16_ASAP7_75t_R g686 ( .A(n_687), .Y(n_686) );
AOI221xp5_ASAP7_75t_L g722 ( .A1(n_690), .A2(n_706), .B1(n_723), .B2(n_726), .C(n_727), .Y(n_722) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
AND2x2_ASAP7_75t_L g741 ( .A(n_692), .B(n_742), .Y(n_741) );
AOI221xp5_ASAP7_75t_L g693 ( .A1(n_694), .A2(n_696), .B1(n_697), .B2(n_699), .C(n_700), .Y(n_693) );
INVx1_ASAP7_75t_SL g694 ( .A(n_695), .Y(n_694) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
NOR2xp33_ASAP7_75t_L g732 ( .A(n_702), .B(n_733), .Y(n_732) );
AOI21xp5_ASAP7_75t_L g705 ( .A1(n_706), .A2(n_708), .B(n_709), .Y(n_705) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
NAND4xp25_ASAP7_75t_L g711 ( .A(n_712), .B(n_722), .C(n_737), .D(n_748), .Y(n_711) );
O2A1O1Ixp33_ASAP7_75t_L g712 ( .A1(n_713), .A2(n_716), .B(n_718), .C(n_720), .Y(n_712) );
NAND2xp5_ASAP7_75t_SL g713 ( .A(n_714), .B(n_715), .Y(n_713) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVxp67_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx1_ASAP7_75t_SL g728 ( .A(n_729), .Y(n_728) );
INVx1_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
INVx1_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
INVx1_ASAP7_75t_L g753 ( .A(n_740), .Y(n_753) );
INVx2_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
OAI21xp5_ASAP7_75t_L g748 ( .A1(n_749), .A2(n_752), .B(n_753), .Y(n_748) );
NOR2xp33_ASAP7_75t_L g749 ( .A(n_750), .B(n_751), .Y(n_749) );
INVx2_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
INVx2_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
INVx1_ASAP7_75t_SL g760 ( .A(n_761), .Y(n_760) );
BUFx2_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
INVx1_ASAP7_75t_L g773 ( .A(n_765), .Y(n_773) );
INVx1_ASAP7_75t_L g766 ( .A(n_767), .Y(n_766) );
CKINVDCx20_ASAP7_75t_R g771 ( .A(n_768), .Y(n_771) );
endmodule