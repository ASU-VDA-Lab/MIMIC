module fake_jpeg_19372_n_181 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_181);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_181;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_93;
wire n_91;
wire n_54;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx13_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_10),
.B(n_14),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_13),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx16f_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

INVxp33_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_7),
.Y(n_34)
);

BUFx12_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

OAI22xp33_ASAP7_75t_L g36 ( 
.A1(n_26),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_36),
.A2(n_30),
.B1(n_28),
.B2(n_23),
.Y(n_70)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_38),
.B(n_39),
.Y(n_54)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_19),
.B(n_0),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_41),
.B(n_46),
.Y(n_61)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

INVx2_ASAP7_75t_SL g43 ( 
.A(n_17),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_43),
.B(n_44),
.Y(n_55)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_21),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_45),
.B(n_48),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_19),
.B(n_22),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_47),
.Y(n_52)
);

INVx13_ASAP7_75t_L g48 ( 
.A(n_17),
.Y(n_48)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_18),
.Y(n_49)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_45),
.A2(n_33),
.B1(n_23),
.B2(n_28),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_50),
.A2(n_62),
.B1(n_70),
.B2(n_43),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_46),
.B(n_19),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_53),
.B(n_66),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_41),
.B(n_20),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_57),
.B(n_59),
.Y(n_82)
);

BUFx8_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_58),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_41),
.B(n_20),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_37),
.A2(n_34),
.B1(n_24),
.B2(n_21),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_38),
.B(n_31),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_44),
.B(n_31),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_42),
.A2(n_30),
.B1(n_28),
.B2(n_23),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_67),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_39),
.B(n_34),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_68),
.B(n_27),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_48),
.B(n_24),
.Y(n_69)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_37),
.Y(n_71)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_71),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_43),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_72),
.B(n_55),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_L g73 ( 
.A1(n_61),
.A2(n_30),
.B(n_21),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_73),
.A2(n_93),
.B(n_55),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_51),
.Y(n_74)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_74),
.Y(n_107)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_75),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_76),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_77),
.B(n_91),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_61),
.B(n_22),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_79),
.B(n_88),
.Y(n_102)
);

AND2x6_ASAP7_75t_L g81 ( 
.A(n_56),
.B(n_48),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_81),
.B(n_95),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_64),
.B(n_25),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_83),
.B(n_32),
.Y(n_105)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_63),
.Y(n_84)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_84),
.Y(n_104)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_52),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_86),
.Y(n_98)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_63),
.Y(n_87)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_87),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_57),
.B(n_59),
.Y(n_88)
);

CKINVDCx14_ASAP7_75t_R g114 ( 
.A(n_89),
.Y(n_114)
);

OR2x2_ASAP7_75t_L g91 ( 
.A(n_69),
.B(n_49),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_62),
.Y(n_92)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_92),
.Y(n_109)
);

A2O1A1Ixp33_ASAP7_75t_L g93 ( 
.A1(n_56),
.A2(n_25),
.B(n_35),
.C(n_32),
.Y(n_93)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_51),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_70),
.A2(n_54),
.B1(n_68),
.B2(n_39),
.Y(n_95)
);

AO22x1_ASAP7_75t_L g99 ( 
.A1(n_81),
.A2(n_72),
.B1(n_58),
.B2(n_54),
.Y(n_99)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_99),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_91),
.B(n_49),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_100),
.A2(n_80),
.B(n_87),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_86),
.Y(n_103)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_103),
.Y(n_126)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_74),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_111),
.B(n_90),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_78),
.B(n_32),
.Y(n_112)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_112),
.Y(n_130)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_75),
.Y(n_113)
);

INVx1_ASAP7_75t_SL g133 ( 
.A(n_113),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_114),
.A2(n_95),
.B1(n_89),
.B2(n_92),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_115),
.A2(n_117),
.B1(n_132),
.B2(n_108),
.Y(n_142)
);

NOR2x1_ASAP7_75t_L g116 ( 
.A(n_96),
.B(n_93),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_116),
.B(n_118),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_110),
.A2(n_85),
.B1(n_79),
.B2(n_73),
.Y(n_117)
);

OR2x2_ASAP7_75t_L g118 ( 
.A(n_101),
.B(n_77),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_102),
.B(n_110),
.C(n_99),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_119),
.B(n_121),
.C(n_125),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_102),
.B(n_88),
.Y(n_121)
);

NOR4xp25_ASAP7_75t_L g122 ( 
.A(n_105),
.B(n_85),
.C(n_82),
.D(n_80),
.Y(n_122)
);

MAJx2_ASAP7_75t_L g149 ( 
.A(n_122),
.B(n_123),
.C(n_124),
.Y(n_149)
);

XOR2x2_ASAP7_75t_L g123 ( 
.A(n_99),
.B(n_82),
.Y(n_123)
);

XNOR2x1_ASAP7_75t_L g124 ( 
.A(n_100),
.B(n_101),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_106),
.B(n_71),
.C(n_84),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_127),
.A2(n_109),
.B(n_104),
.Y(n_136)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_128),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_106),
.B(n_60),
.C(n_65),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_129),
.B(n_131),
.C(n_107),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_100),
.B(n_60),
.C(n_65),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_109),
.A2(n_90),
.B1(n_94),
.B2(n_52),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_130),
.B(n_103),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_135),
.B(n_138),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_136),
.A2(n_137),
.B(n_141),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_120),
.A2(n_113),
.B(n_97),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_126),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_117),
.A2(n_108),
.B(n_97),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_142),
.A2(n_116),
.B1(n_115),
.B2(n_124),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_123),
.A2(n_104),
.B(n_111),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_143),
.A2(n_58),
.B(n_17),
.Y(n_154)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_132),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_144),
.B(n_146),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_118),
.B(n_98),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_145),
.B(n_147),
.Y(n_158)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_125),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_129),
.B(n_98),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_133),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_151),
.B(n_152),
.Y(n_161)
);

OAI321xp33_ASAP7_75t_L g152 ( 
.A1(n_141),
.A2(n_131),
.A3(n_133),
.B1(n_40),
.B2(n_35),
.C(n_32),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_140),
.B(n_40),
.C(n_58),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_149),
.A2(n_16),
.B(n_15),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_159),
.B(n_139),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_155),
.A2(n_142),
.B1(n_144),
.B2(n_134),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_160),
.B(n_162),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_153),
.A2(n_134),
.B1(n_148),
.B2(n_137),
.Y(n_162)
);

A2O1A1Ixp33_ASAP7_75t_SL g163 ( 
.A1(n_154),
.A2(n_143),
.B(n_136),
.C(n_149),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_163),
.B(n_2),
.Y(n_169)
);

NAND3xp33_ASAP7_75t_L g164 ( 
.A(n_157),
.B(n_139),
.C(n_150),
.Y(n_164)
);

AOI31xp67_ASAP7_75t_L g172 ( 
.A1(n_164),
.A2(n_166),
.A3(n_167),
.B(n_5),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_165),
.B(n_5),
.Y(n_171)
);

XOR2x2_ASAP7_75t_L g166 ( 
.A(n_156),
.B(n_1),
.Y(n_166)
);

OAI21x1_ASAP7_75t_L g167 ( 
.A1(n_158),
.A2(n_16),
.B(n_15),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_169),
.A2(n_163),
.B(n_8),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_161),
.B(n_2),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_170),
.B(n_171),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_172),
.A2(n_166),
.B(n_163),
.Y(n_173)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_173),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_168),
.A2(n_163),
.B1(n_7),
.B2(n_8),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_174),
.B(n_175),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_178),
.B(n_176),
.C(n_9),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_179),
.B(n_177),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_180),
.B(n_179),
.Y(n_181)
);


endmodule