module fake_jpeg_4506_n_345 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_345);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_345;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx16_ASAP7_75t_R g17 ( 
.A(n_12),
.Y(n_17)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx8_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_16),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx12_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_35),
.B(n_36),
.Y(n_49)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_37),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_39),
.B(n_43),
.Y(n_54)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

BUFx2_ASAP7_75t_SL g58 ( 
.A(n_40),
.Y(n_58)
);

INVx6_ASAP7_75t_SL g41 ( 
.A(n_24),
.Y(n_41)
);

CKINVDCx14_ASAP7_75t_R g53 ( 
.A(n_41),
.Y(n_53)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_44),
.B(n_45),
.Y(n_70)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_22),
.Y(n_45)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_46),
.A2(n_18),
.B1(n_28),
.B2(n_31),
.Y(n_56)
);

BUFx24_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

INVx1_ASAP7_75t_SL g69 ( 
.A(n_47),
.Y(n_69)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_50),
.Y(n_99)
);

INVx6_ASAP7_75t_SL g51 ( 
.A(n_41),
.Y(n_51)
);

CKINVDCx14_ASAP7_75t_R g79 ( 
.A(n_51),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_47),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_52),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_46),
.A2(n_18),
.B1(n_31),
.B2(n_28),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_55),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_56),
.A2(n_59),
.B1(n_61),
.B2(n_44),
.Y(n_78)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

HB1xp67_ASAP7_75t_L g87 ( 
.A(n_57),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_39),
.A2(n_18),
.B1(n_17),
.B2(n_20),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_42),
.A2(n_20),
.B1(n_29),
.B2(n_25),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_60),
.A2(n_21),
.B1(n_27),
.B2(n_19),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_39),
.A2(n_17),
.B1(n_29),
.B2(n_27),
.Y(n_61)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_62),
.Y(n_85)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_63),
.Y(n_93)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_64),
.B(n_67),
.Y(n_90)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_66),
.Y(n_89)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_68),
.Y(n_86)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_72),
.Y(n_98)
);

INVx1_ASAP7_75t_SL g73 ( 
.A(n_38),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_73),
.B(n_24),
.Y(n_77)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_38),
.Y(n_74)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_74),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_77),
.B(n_69),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_78),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_60),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_80),
.Y(n_102)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_48),
.Y(n_81)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_81),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_82),
.A2(n_44),
.B1(n_74),
.B2(n_71),
.Y(n_105)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_48),
.Y(n_83)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_83),
.Y(n_106)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_58),
.Y(n_84)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_84),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_58),
.Y(n_88)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_88),
.Y(n_101)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_51),
.Y(n_91)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_91),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_49),
.B(n_25),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_92),
.B(n_70),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_50),
.A2(n_46),
.B1(n_35),
.B2(n_40),
.Y(n_94)
);

INVx1_ASAP7_75t_SL g116 ( 
.A(n_94),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_70),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_95),
.B(n_54),
.Y(n_109)
);

OAI32xp33_ASAP7_75t_L g97 ( 
.A1(n_55),
.A2(n_36),
.A3(n_19),
.B1(n_21),
.B2(n_46),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_97),
.B(n_54),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_100),
.B(n_109),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_105),
.A2(n_122),
.B1(n_83),
.B2(n_76),
.Y(n_132)
);

NOR2x1_ASAP7_75t_R g107 ( 
.A(n_97),
.B(n_46),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_107),
.A2(n_118),
.B(n_24),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_90),
.B(n_49),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_108),
.B(n_127),
.Y(n_136)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_87),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_110),
.Y(n_154)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_82),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_111),
.B(n_114),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_112),
.B(n_113),
.Y(n_130)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_88),
.Y(n_114)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_87),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_115),
.B(n_120),
.Y(n_148)
);

AND2x4_ASAP7_75t_SL g118 ( 
.A(n_80),
.B(n_52),
.Y(n_118)
);

OAI22xp33_ASAP7_75t_L g119 ( 
.A1(n_96),
.A2(n_71),
.B1(n_72),
.B2(n_68),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_119),
.A2(n_126),
.B1(n_65),
.B2(n_73),
.Y(n_150)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_90),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_92),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_121),
.B(n_123),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_95),
.A2(n_44),
.B1(n_37),
.B2(n_43),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_77),
.Y(n_123)
);

INVxp33_ASAP7_75t_L g124 ( 
.A(n_81),
.Y(n_124)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_124),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_75),
.B(n_67),
.C(n_64),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_125),
.B(n_53),
.C(n_79),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_75),
.A2(n_43),
.B1(n_37),
.B2(n_66),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_77),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_110),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_129),
.Y(n_159)
);

O2A1O1Ixp33_ASAP7_75t_L g131 ( 
.A1(n_118),
.A2(n_84),
.B(n_71),
.C(n_43),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_131),
.A2(n_122),
.B(n_117),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_132),
.A2(n_135),
.B1(n_155),
.B2(n_151),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_107),
.A2(n_37),
.B1(n_62),
.B2(n_57),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_133),
.A2(n_138),
.B1(n_142),
.B2(n_146),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_111),
.A2(n_63),
.B1(n_98),
.B2(n_86),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_137),
.B(n_151),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_118),
.A2(n_86),
.B1(n_98),
.B2(n_35),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_120),
.B(n_93),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_139),
.B(n_141),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_108),
.B(n_93),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_102),
.A2(n_35),
.B1(n_85),
.B2(n_79),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_127),
.B(n_36),
.C(n_85),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_143),
.B(n_121),
.C(n_104),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_128),
.A2(n_91),
.B1(n_40),
.B2(n_99),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_145),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_113),
.A2(n_40),
.B1(n_76),
.B2(n_99),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_147),
.A2(n_101),
.B(n_106),
.Y(n_178)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_103),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_149),
.B(n_155),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_150),
.A2(n_65),
.B1(n_89),
.B2(n_30),
.Y(n_183)
);

OR2x2_ASAP7_75t_L g151 ( 
.A(n_119),
.B(n_38),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_103),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_153),
.Y(n_167)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_126),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_100),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_156),
.B(n_157),
.Y(n_187)
);

BUFx8_ASAP7_75t_L g157 ( 
.A(n_124),
.Y(n_157)
);

OR2x2_ASAP7_75t_L g158 ( 
.A(n_134),
.B(n_105),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_158),
.B(n_176),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_160),
.A2(n_164),
.B1(n_166),
.B2(n_131),
.Y(n_188)
);

AND2x2_ASAP7_75t_SL g162 ( 
.A(n_130),
.B(n_125),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_162),
.A2(n_171),
.B(n_172),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_165),
.B(n_169),
.C(n_175),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_151),
.A2(n_116),
.B1(n_112),
.B2(n_115),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_146),
.B(n_112),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_139),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_170),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_147),
.A2(n_116),
.B(n_114),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_144),
.A2(n_136),
.B(n_141),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_136),
.B(n_47),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_173),
.B(n_174),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_SL g174 ( 
.A(n_130),
.B(n_47),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_130),
.B(n_47),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_148),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_130),
.B(n_69),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_177),
.B(n_138),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_178),
.A2(n_184),
.B(n_157),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_137),
.B(n_101),
.C(n_38),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_179),
.B(n_129),
.C(n_140),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_142),
.B(n_13),
.Y(n_180)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_180),
.Y(n_210)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_148),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_181),
.B(n_182),
.Y(n_193)
);

CKINVDCx14_ASAP7_75t_R g182 ( 
.A(n_135),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_183),
.A2(n_167),
.B1(n_159),
.B2(n_158),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_144),
.A2(n_33),
.B(n_89),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_188),
.A2(n_199),
.B(n_208),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_160),
.A2(n_133),
.B1(n_131),
.B2(n_156),
.Y(n_189)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_189),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_190),
.B(n_198),
.C(n_213),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_163),
.B(n_143),
.Y(n_194)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_194),
.Y(n_234)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_163),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_195),
.B(n_205),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_168),
.A2(n_132),
.B1(n_134),
.B2(n_145),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_197),
.A2(n_203),
.B1(n_161),
.B2(n_166),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_185),
.A2(n_152),
.B1(n_140),
.B2(n_150),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_186),
.A2(n_152),
.B1(n_153),
.B2(n_154),
.Y(n_200)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_200),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_201),
.A2(n_204),
.B1(n_176),
.B2(n_183),
.Y(n_225)
);

XOR2x2_ASAP7_75t_L g202 ( 
.A(n_162),
.B(n_174),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_202),
.B(n_30),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_168),
.A2(n_157),
.B1(n_149),
.B2(n_65),
.Y(n_203)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_187),
.Y(n_205)
);

NAND3xp33_ASAP7_75t_L g207 ( 
.A(n_162),
.B(n_157),
.C(n_24),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_207),
.B(n_32),
.Y(n_239)
);

XNOR2x2_ASAP7_75t_L g208 ( 
.A(n_177),
.B(n_24),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_186),
.A2(n_89),
.B1(n_34),
.B2(n_26),
.Y(n_209)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_209),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_167),
.B(n_34),
.Y(n_212)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_212),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_169),
.B(n_33),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_175),
.B(n_33),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_214),
.B(n_165),
.C(n_179),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_159),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_215),
.B(n_0),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_217),
.B(n_221),
.C(n_222),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_218),
.A2(n_225),
.B1(n_188),
.B2(n_200),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_197),
.A2(n_186),
.B1(n_172),
.B2(n_164),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_220),
.A2(n_224),
.B1(n_199),
.B2(n_201),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_196),
.B(n_171),
.C(n_170),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_196),
.B(n_178),
.C(n_184),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_213),
.B(n_173),
.C(n_181),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_223),
.B(n_241),
.C(n_242),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_208),
.A2(n_185),
.B1(n_211),
.B2(n_202),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_206),
.B(n_32),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_226),
.B(n_230),
.Y(n_249)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_229),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_206),
.B(n_32),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_193),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_231),
.B(n_240),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_192),
.B(n_32),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_232),
.B(n_226),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_205),
.B(n_34),
.Y(n_233)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_233),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_195),
.B(n_0),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_237),
.B(n_1),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_191),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_238),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_239),
.B(n_210),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_192),
.B(n_34),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_243),
.A2(n_252),
.B1(n_217),
.B2(n_230),
.Y(n_269)
);

INVxp67_ASAP7_75t_SL g244 ( 
.A(n_218),
.Y(n_244)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_244),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_246),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_247),
.B(n_248),
.Y(n_274)
);

CKINVDCx16_ASAP7_75t_R g248 ( 
.A(n_228),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_251),
.B(n_254),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_227),
.A2(n_189),
.B1(n_203),
.B2(n_209),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_236),
.B(n_194),
.Y(n_253)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_253),
.Y(n_272)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_255),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_SL g256 ( 
.A(n_220),
.B(n_190),
.Y(n_256)
);

MAJx2_ASAP7_75t_L g284 ( 
.A(n_256),
.B(n_262),
.C(n_4),
.Y(n_284)
);

XOR2x2_ASAP7_75t_L g257 ( 
.A(n_219),
.B(n_198),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_257),
.A2(n_263),
.B(n_265),
.Y(n_282)
);

CKINVDCx16_ASAP7_75t_R g258 ( 
.A(n_242),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_258),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_234),
.B(n_235),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_259),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_SL g262 ( 
.A(n_241),
.B(n_214),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_219),
.B(n_26),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_222),
.A2(n_221),
.B1(n_224),
.B2(n_232),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_264),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_277)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_223),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_256),
.B(n_216),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_267),
.B(n_268),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_257),
.B(n_216),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_269),
.A2(n_281),
.B1(n_268),
.B2(n_267),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_250),
.B(n_1),
.C(n_2),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_276),
.B(n_277),
.C(n_278),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_250),
.B(n_1),
.C(n_2),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_254),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_279),
.A2(n_11),
.B1(n_15),
.B2(n_14),
.Y(n_296)
);

AND2x2_ASAP7_75t_L g280 ( 
.A(n_259),
.B(n_3),
.Y(n_280)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_280),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_284),
.B(n_262),
.C(n_255),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_264),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_285),
.A2(n_11),
.B1(n_15),
.B2(n_14),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g313 ( 
.A1(n_288),
.A2(n_292),
.B(n_299),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_273),
.B(n_265),
.C(n_261),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_290),
.B(n_291),
.C(n_294),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_273),
.B(n_261),
.C(n_266),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_271),
.B(n_245),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_272),
.B(n_245),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_293),
.B(n_301),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_282),
.B(n_251),
.C(n_249),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_270),
.A2(n_260),
.B1(n_249),
.B2(n_6),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_295),
.A2(n_296),
.B1(n_285),
.B2(n_277),
.Y(n_302)
);

HB1xp67_ASAP7_75t_L g297 ( 
.A(n_280),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_297),
.B(n_300),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_298),
.B(n_284),
.Y(n_307)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_280),
.Y(n_299)
);

OR2x2_ASAP7_75t_L g300 ( 
.A(n_283),
.B(n_4),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_302),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_287),
.B(n_269),
.C(n_278),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_305),
.B(n_294),
.C(n_288),
.Y(n_317)
);

HB1xp67_ASAP7_75t_L g306 ( 
.A(n_300),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_306),
.B(n_312),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_307),
.B(n_308),
.Y(n_318)
);

XNOR2x1_ASAP7_75t_L g308 ( 
.A(n_287),
.B(n_279),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_289),
.B(n_275),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_309),
.B(n_5),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_290),
.B(n_276),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_310),
.B(n_5),
.C(n_8),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_295),
.A2(n_274),
.B1(n_6),
.B2(n_7),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_286),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_314),
.B(n_301),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_291),
.B(n_9),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_315),
.B(n_286),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_316),
.B(n_321),
.Y(n_331)
);

AND2x2_ASAP7_75t_L g326 ( 
.A(n_317),
.B(n_323),
.Y(n_326)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_308),
.Y(n_319)
);

AOI22xp33_ASAP7_75t_SL g327 ( 
.A1(n_319),
.A2(n_322),
.B1(n_9),
.B2(n_13),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_SL g322 ( 
.A1(n_311),
.A2(n_9),
.B(n_12),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_324),
.B(n_303),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_L g337 ( 
.A1(n_327),
.A2(n_329),
.B(n_330),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_328),
.B(n_332),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_322),
.B(n_313),
.Y(n_329)
);

OR2x2_ASAP7_75t_L g330 ( 
.A(n_325),
.B(n_307),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_SL g332 ( 
.A(n_320),
.B(n_318),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_SL g333 ( 
.A(n_318),
.B(n_310),
.Y(n_333)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_333),
.Y(n_336)
);

NOR2xp67_ASAP7_75t_SL g335 ( 
.A(n_326),
.B(n_317),
.Y(n_335)
);

MAJx2_ASAP7_75t_L g339 ( 
.A(n_335),
.B(n_333),
.C(n_304),
.Y(n_339)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_331),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_338),
.B(n_304),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_339),
.B(n_340),
.C(n_305),
.Y(n_341)
);

NOR3xp33_ASAP7_75t_L g342 ( 
.A(n_341),
.B(n_336),
.C(n_337),
.Y(n_342)
);

BUFx24_ASAP7_75t_SL g343 ( 
.A(n_342),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_SL g344 ( 
.A1(n_343),
.A2(n_334),
.B(n_16),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g345 ( 
.A(n_344),
.B(n_8),
.Y(n_345)
);


endmodule