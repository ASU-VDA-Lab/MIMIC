module fake_jpeg_13259_n_526 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_526);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_526;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx12_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx2_ASAP7_75t_R g32 ( 
.A(n_11),
.Y(n_32)
);

BUFx12_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

BUFx12_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_4),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

INVx13_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_9),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g46 ( 
.A(n_9),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_8),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_13),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_32),
.B(n_15),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_50),
.B(n_54),
.Y(n_109)
);

INVx4_ASAP7_75t_SL g51 ( 
.A(n_44),
.Y(n_51)
);

INVx13_ASAP7_75t_L g159 ( 
.A(n_51),
.Y(n_159)
);

INVx2_ASAP7_75t_SL g52 ( 
.A(n_41),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_52),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_19),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_53),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_32),
.B(n_15),
.Y(n_54)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g118 ( 
.A(n_55),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_32),
.B(n_15),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_56),
.B(n_82),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_32),
.B(n_14),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_57),
.B(n_62),
.Y(n_152)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_29),
.Y(n_58)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_58),
.Y(n_102)
);

INVx13_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

INVx6_ASAP7_75t_SL g131 ( 
.A(n_59),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_19),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_60),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_19),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_61),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_17),
.B(n_13),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_25),
.Y(n_63)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_63),
.Y(n_105)
);

OR2x2_ASAP7_75t_L g64 ( 
.A(n_47),
.B(n_13),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_64),
.B(n_76),
.Y(n_123)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_65),
.Y(n_140)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_23),
.Y(n_66)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_66),
.Y(n_100)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_67),
.Y(n_112)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

HB1xp67_ASAP7_75t_L g153 ( 
.A(n_68),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_19),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_69),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_70),
.Y(n_128)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_49),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_71),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_72),
.Y(n_137)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_25),
.Y(n_73)
);

INVx5_ASAP7_75t_L g158 ( 
.A(n_73),
.Y(n_158)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_43),
.Y(n_74)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_74),
.Y(n_134)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_25),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_75),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_30),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_17),
.B(n_12),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_77),
.B(n_78),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_46),
.B(n_12),
.Y(n_78)
);

INVx11_ASAP7_75t_L g79 ( 
.A(n_42),
.Y(n_79)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_79),
.Y(n_107)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_29),
.Y(n_80)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_80),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_47),
.B(n_12),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_81),
.B(n_8),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_18),
.B(n_10),
.Y(n_82)
);

BUFx5_ASAP7_75t_L g83 ( 
.A(n_28),
.Y(n_83)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_83),
.Y(n_117)
);

INVx4_ASAP7_75t_SL g84 ( 
.A(n_42),
.Y(n_84)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_84),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_45),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_85),
.Y(n_149)
);

INVx11_ASAP7_75t_L g86 ( 
.A(n_28),
.Y(n_86)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_86),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_45),
.Y(n_87)
);

INVx6_ASAP7_75t_L g127 ( 
.A(n_87),
.Y(n_127)
);

BUFx4f_ASAP7_75t_L g88 ( 
.A(n_41),
.Y(n_88)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_88),
.Y(n_111)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_18),
.Y(n_89)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_89),
.Y(n_113)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_48),
.Y(n_90)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_90),
.Y(n_114)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_23),
.Y(n_91)
);

HB1xp67_ASAP7_75t_L g157 ( 
.A(n_91),
.Y(n_157)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_49),
.Y(n_92)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_92),
.Y(n_120)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_43),
.Y(n_93)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_93),
.Y(n_124)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_23),
.Y(n_94)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_94),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_49),
.Y(n_95)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_95),
.Y(n_129)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_18),
.Y(n_96)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_96),
.Y(n_135)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_41),
.Y(n_97)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_97),
.Y(n_139)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_41),
.Y(n_98)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_98),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_48),
.B(n_24),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_99),
.B(n_24),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_104),
.B(n_136),
.Y(n_185)
);

AND2x2_ASAP7_75t_SL g115 ( 
.A(n_82),
.B(n_38),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_115),
.B(n_123),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_52),
.A2(n_22),
.B1(n_36),
.B2(n_35),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_116),
.A2(n_132),
.B(n_148),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_58),
.B(n_31),
.C(n_27),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_121),
.B(n_150),
.Y(n_174)
);

AOI21xp33_ASAP7_75t_L g130 ( 
.A1(n_62),
.A2(n_37),
.B(n_26),
.Y(n_130)
);

AOI21xp33_ASAP7_75t_L g191 ( 
.A1(n_130),
.A2(n_147),
.B(n_84),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_52),
.A2(n_22),
.B1(n_36),
.B2(n_35),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_64),
.B(n_26),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_77),
.A2(n_40),
.B1(n_21),
.B2(n_49),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_138),
.A2(n_40),
.B1(n_21),
.B2(n_72),
.Y(n_196)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_90),
.Y(n_141)
);

INVx1_ASAP7_75t_SL g201 ( 
.A(n_141),
.Y(n_201)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_80),
.Y(n_144)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_144),
.Y(n_161)
);

AOI21xp33_ASAP7_75t_L g147 ( 
.A1(n_65),
.A2(n_37),
.B(n_16),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_73),
.A2(n_36),
.B1(n_35),
.B2(n_22),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_97),
.B(n_16),
.C(n_20),
.Y(n_150)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_89),
.Y(n_151)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_151),
.Y(n_177)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_96),
.Y(n_154)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_154),
.Y(n_186)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_88),
.Y(n_155)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_155),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_156),
.B(n_145),
.Y(n_180)
);

INVx3_ASAP7_75t_SL g160 ( 
.A(n_131),
.Y(n_160)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_160),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_153),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_162),
.B(n_176),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_L g163 ( 
.A1(n_114),
.A2(n_92),
.B1(n_71),
.B2(n_70),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_163),
.A2(n_179),
.B1(n_182),
.B2(n_203),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_109),
.A2(n_63),
.B1(n_66),
.B2(n_94),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g211 ( 
.A(n_164),
.Y(n_211)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_103),
.Y(n_165)
);

INVx4_ASAP7_75t_L g234 ( 
.A(n_165),
.Y(n_234)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_103),
.Y(n_166)
);

INVx1_ASAP7_75t_SL g235 ( 
.A(n_166),
.Y(n_235)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_107),
.Y(n_168)
);

INVx5_ASAP7_75t_L g222 ( 
.A(n_168),
.Y(n_222)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_119),
.Y(n_169)
);

BUFx3_ASAP7_75t_L g233 ( 
.A(n_169),
.Y(n_233)
);

AOI32xp33_ASAP7_75t_L g170 ( 
.A1(n_101),
.A2(n_86),
.A3(n_76),
.B1(n_55),
.B2(n_79),
.Y(n_170)
);

AOI21xp33_ASAP7_75t_L g217 ( 
.A1(n_170),
.A2(n_83),
.B(n_88),
.Y(n_217)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_107),
.Y(n_171)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_171),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_115),
.A2(n_152),
.B1(n_91),
.B2(n_117),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_172),
.Y(n_220)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_119),
.Y(n_173)
);

BUFx3_ASAP7_75t_L g238 ( 
.A(n_173),
.Y(n_238)
);

BUFx2_ASAP7_75t_L g175 ( 
.A(n_105),
.Y(n_175)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_175),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_157),
.Y(n_176)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_113),
.Y(n_178)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_178),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_148),
.A2(n_53),
.B1(n_60),
.B2(n_61),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_180),
.B(n_192),
.Y(n_224)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_112),
.Y(n_181)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_181),
.Y(n_245)
);

OAI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_116),
.A2(n_69),
.B1(n_95),
.B2(n_87),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_183),
.B(n_38),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_117),
.A2(n_93),
.B1(n_67),
.B2(n_74),
.Y(n_184)
);

OAI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_184),
.A2(n_196),
.B1(n_140),
.B2(n_142),
.Y(n_214)
);

HB1xp67_ASAP7_75t_L g187 ( 
.A(n_125),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_187),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_102),
.B(n_31),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_188),
.B(n_198),
.Y(n_227)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_146),
.Y(n_189)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_189),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_105),
.A2(n_75),
.B1(n_27),
.B2(n_20),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_190),
.A2(n_207),
.B1(n_140),
.B2(n_142),
.Y(n_213)
);

NOR2x1_ASAP7_75t_R g210 ( 
.A(n_191),
.B(n_200),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_106),
.B(n_98),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_135),
.Y(n_193)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_193),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_128),
.Y(n_194)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_194),
.Y(n_228)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_111),
.Y(n_195)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_195),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_139),
.B(n_68),
.Y(n_198)
);

INVx3_ASAP7_75t_SL g199 ( 
.A(n_146),
.Y(n_199)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_199),
.Y(n_240)
);

AND2x4_ASAP7_75t_L g200 ( 
.A(n_143),
.B(n_28),
.Y(n_200)
);

CKINVDCx14_ASAP7_75t_R g202 ( 
.A(n_159),
.Y(n_202)
);

CKINVDCx14_ASAP7_75t_R g225 ( 
.A(n_202),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_132),
.A2(n_85),
.B1(n_21),
.B2(n_40),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_128),
.Y(n_204)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_204),
.Y(n_244)
);

BUFx2_ASAP7_75t_L g205 ( 
.A(n_158),
.Y(n_205)
);

BUFx24_ASAP7_75t_L g239 ( 
.A(n_205),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_100),
.B(n_38),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_206),
.B(n_38),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_158),
.A2(n_38),
.B1(n_51),
.B2(n_59),
.Y(n_207)
);

BUFx12_ASAP7_75t_L g208 ( 
.A(n_159),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_208),
.Y(n_232)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_120),
.Y(n_209)
);

OR2x2_ASAP7_75t_L g215 ( 
.A(n_209),
.B(n_112),
.Y(n_215)
);

OAI21xp33_ASAP7_75t_SL g252 ( 
.A1(n_213),
.A2(n_236),
.B(n_247),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_214),
.A2(n_200),
.B1(n_201),
.B2(n_160),
.Y(n_253)
);

INVx1_ASAP7_75t_SL g251 ( 
.A(n_215),
.Y(n_251)
);

AND2x2_ASAP7_75t_L g256 ( 
.A(n_217),
.B(n_200),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_183),
.B(n_124),
.C(n_129),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_226),
.B(n_167),
.C(n_161),
.Y(n_284)
);

OR2x2_ASAP7_75t_L g230 ( 
.A(n_188),
.B(n_134),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_230),
.A2(n_208),
.B(n_195),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_179),
.A2(n_134),
.B1(n_127),
.B2(n_118),
.Y(n_236)
);

XNOR2x1_ASAP7_75t_L g275 ( 
.A(n_237),
.B(n_39),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_241),
.B(n_173),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_203),
.A2(n_127),
.B1(n_133),
.B2(n_108),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_243),
.A2(n_197),
.B1(n_184),
.B2(n_196),
.Y(n_249)
);

AOI32xp33_ASAP7_75t_L g246 ( 
.A1(n_172),
.A2(n_118),
.A3(n_133),
.B1(n_126),
.B2(n_122),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_SL g264 ( 
.A1(n_246),
.A2(n_164),
.B(n_199),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_SL g247 ( 
.A1(n_197),
.A2(n_118),
.B1(n_108),
.B2(n_126),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_249),
.A2(n_241),
.B1(n_210),
.B2(n_243),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_227),
.B(n_174),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_250),
.B(n_279),
.Y(n_292)
);

OA21x2_ASAP7_75t_L g309 ( 
.A1(n_253),
.A2(n_166),
.B(n_239),
.Y(n_309)
);

AOI22xp33_ASAP7_75t_L g254 ( 
.A1(n_211),
.A2(n_201),
.B1(n_189),
.B2(n_205),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g295 ( 
.A(n_254),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_220),
.A2(n_211),
.B1(n_227),
.B2(n_221),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_255),
.A2(n_257),
.B1(n_258),
.B2(n_186),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_256),
.A2(n_264),
.B(n_274),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_220),
.A2(n_183),
.B1(n_200),
.B2(n_198),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_221),
.A2(n_209),
.B1(n_193),
.B2(n_178),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_224),
.B(n_185),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_259),
.B(n_260),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_230),
.B(n_162),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_212),
.Y(n_261)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_261),
.Y(n_285)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_212),
.Y(n_262)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_262),
.Y(n_287)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_248),
.Y(n_263)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_263),
.Y(n_289)
);

AOI22xp33_ASAP7_75t_L g265 ( 
.A1(n_246),
.A2(n_149),
.B1(n_137),
.B2(n_122),
.Y(n_265)
);

CKINVDCx16_ASAP7_75t_R g315 ( 
.A(n_265),
.Y(n_315)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_248),
.Y(n_266)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_266),
.Y(n_300)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_231),
.Y(n_267)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_267),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_216),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_268),
.B(n_276),
.Y(n_286)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_231),
.Y(n_269)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_269),
.Y(n_307)
);

INVx3_ASAP7_75t_L g270 ( 
.A(n_218),
.Y(n_270)
);

INVx4_ASAP7_75t_L g313 ( 
.A(n_270),
.Y(n_313)
);

AOI22xp33_ASAP7_75t_L g271 ( 
.A1(n_240),
.A2(n_149),
.B1(n_137),
.B2(n_110),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_271),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_237),
.B(n_226),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_272),
.B(n_284),
.C(n_275),
.Y(n_293)
);

AND2x2_ASAP7_75t_L g273 ( 
.A(n_230),
.B(n_216),
.Y(n_273)
);

INVx1_ASAP7_75t_SL g306 ( 
.A(n_273),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_275),
.B(n_235),
.Y(n_294)
);

CKINVDCx14_ASAP7_75t_R g276 ( 
.A(n_225),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_240),
.Y(n_277)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_277),
.Y(n_308)
);

INVx3_ASAP7_75t_L g278 ( 
.A(n_218),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_278),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_210),
.B(n_161),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_219),
.Y(n_280)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_280),
.Y(n_310)
);

BUFx3_ASAP7_75t_L g281 ( 
.A(n_242),
.Y(n_281)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_281),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_224),
.B(n_169),
.Y(n_282)
);

CKINVDCx14_ASAP7_75t_R g314 ( 
.A(n_282),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_283),
.B(n_232),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_288),
.A2(n_299),
.B1(n_316),
.B2(n_277),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_293),
.B(n_312),
.C(n_283),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_294),
.B(n_312),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_SL g322 ( 
.A(n_296),
.B(n_303),
.Y(n_322)
);

OAI22x1_ASAP7_75t_SL g297 ( 
.A1(n_255),
.A2(n_215),
.B1(n_219),
.B2(n_245),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_297),
.A2(n_311),
.B1(n_251),
.B2(n_279),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_L g298 ( 
.A1(n_274),
.A2(n_215),
.B(n_223),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_L g336 ( 
.A1(n_298),
.A2(n_301),
.B(n_269),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_249),
.A2(n_244),
.B1(n_228),
.B2(n_223),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_L g301 ( 
.A1(n_273),
.A2(n_232),
.B(n_235),
.Y(n_301)
);

AOI322xp5_ASAP7_75t_L g303 ( 
.A1(n_268),
.A2(n_245),
.A3(n_222),
.B1(n_242),
.B2(n_229),
.C1(n_238),
.C2(n_233),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_250),
.B(n_244),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_305),
.B(n_267),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_SL g354 ( 
.A1(n_309),
.A2(n_239),
.B(n_208),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_272),
.B(n_167),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_256),
.A2(n_228),
.B1(n_110),
.B2(n_204),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_273),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_317),
.B(n_251),
.Y(n_320)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_320),
.Y(n_358)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_285),
.Y(n_321)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_321),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_286),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_323),
.B(n_326),
.Y(n_360)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_285),
.Y(n_324)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_324),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_L g355 ( 
.A1(n_325),
.A2(n_329),
.B1(n_345),
.B2(n_346),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_304),
.B(n_260),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_L g327 ( 
.A1(n_315),
.A2(n_258),
.B1(n_253),
.B2(n_257),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_327),
.A2(n_328),
.B1(n_334),
.B2(n_339),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_L g328 ( 
.A1(n_288),
.A2(n_264),
.B1(n_252),
.B2(n_282),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_311),
.A2(n_256),
.B1(n_284),
.B2(n_261),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_SL g359 ( 
.A(n_330),
.B(n_294),
.Y(n_359)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_289),
.Y(n_331)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_331),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_332),
.B(n_308),
.C(n_316),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_314),
.B(n_259),
.Y(n_333)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_333),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_305),
.B(n_280),
.Y(n_335)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_335),
.Y(n_383)
);

INVxp67_ASAP7_75t_L g380 ( 
.A(n_336),
.Y(n_380)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_337),
.Y(n_386)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_289),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_338),
.B(n_341),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_L g339 ( 
.A1(n_299),
.A2(n_263),
.B1(n_266),
.B2(n_262),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_292),
.A2(n_278),
.B1(n_270),
.B2(n_194),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_340),
.A2(n_343),
.B1(n_347),
.B2(n_348),
.Y(n_385)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_300),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_317),
.B(n_281),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g363 ( 
.A(n_342),
.B(n_344),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_292),
.A2(n_238),
.B1(n_233),
.B2(n_234),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_290),
.Y(n_344)
);

INVx1_ASAP7_75t_SL g345 ( 
.A(n_309),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_306),
.A2(n_175),
.B1(n_234),
.B2(n_181),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_306),
.A2(n_229),
.B1(n_222),
.B2(n_186),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_293),
.A2(n_177),
.B1(n_239),
.B2(n_165),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_297),
.A2(n_239),
.B1(n_177),
.B2(n_168),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_L g367 ( 
.A1(n_349),
.A2(n_350),
.B1(n_351),
.B2(n_353),
.Y(n_367)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_300),
.Y(n_350)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_290),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_308),
.B(n_0),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_352),
.Y(n_357)
);

INVxp67_ASAP7_75t_L g353 ( 
.A(n_301),
.Y(n_353)
);

AOI21xp5_ASAP7_75t_L g376 ( 
.A1(n_354),
.A2(n_313),
.B(n_318),
.Y(n_376)
);

XOR2xp5_ASAP7_75t_L g356 ( 
.A(n_330),
.B(n_319),
.Y(n_356)
);

XOR2xp5_ASAP7_75t_L g399 ( 
.A(n_356),
.B(n_372),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_SL g418 ( 
.A(n_359),
.B(n_368),
.Y(n_418)
);

A2O1A1O1Ixp25_ASAP7_75t_L g361 ( 
.A1(n_336),
.A2(n_319),
.B(n_298),
.C(n_307),
.D(n_302),
.Y(n_361)
);

OAI21xp5_ASAP7_75t_SL g410 ( 
.A1(n_361),
.A2(n_376),
.B(n_33),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_365),
.B(n_371),
.C(n_375),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_SL g368 ( 
.A(n_332),
.B(n_309),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_325),
.A2(n_295),
.B1(n_291),
.B2(n_302),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_L g389 ( 
.A1(n_369),
.A2(n_381),
.B1(n_387),
.B2(n_324),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_L g370 ( 
.A1(n_333),
.A2(n_291),
.B1(n_295),
.B2(n_307),
.Y(n_370)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_370),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_329),
.B(n_310),
.C(n_287),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_326),
.B(n_310),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_320),
.B(n_287),
.Y(n_373)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_373),
.B(n_374),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_328),
.B(n_337),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_348),
.B(n_318),
.C(n_290),
.Y(n_375)
);

XOR2xp5_ASAP7_75t_L g377 ( 
.A(n_335),
.B(n_313),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_377),
.B(n_384),
.C(n_39),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_345),
.A2(n_171),
.B1(n_1),
.B2(n_2),
.Y(n_381)
);

OA22x2_ASAP7_75t_L g382 ( 
.A1(n_349),
.A2(n_11),
.B1(n_10),
.B2(n_2),
.Y(n_382)
);

INVxp67_ASAP7_75t_L g391 ( 
.A(n_382),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_342),
.B(n_34),
.C(n_30),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_322),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_387)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_389),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_L g390 ( 
.A(n_368),
.B(n_334),
.Y(n_390)
);

XOR2xp5_ASAP7_75t_L g434 ( 
.A(n_390),
.B(n_397),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_360),
.B(n_323),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_SL g441 ( 
.A(n_392),
.B(n_407),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_379),
.A2(n_322),
.B1(n_346),
.B2(n_350),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_L g433 ( 
.A1(n_394),
.A2(n_404),
.B1(n_381),
.B2(n_387),
.Y(n_433)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_378),
.Y(n_395)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_395),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_356),
.B(n_327),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_366),
.B(n_343),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_398),
.Y(n_427)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_383),
.Y(n_400)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_400),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_365),
.B(n_339),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_401),
.B(n_402),
.C(n_403),
.Y(n_429)
);

XNOR2x1_ASAP7_75t_L g402 ( 
.A(n_374),
.B(n_340),
.Y(n_402)
);

XNOR2xp5_ASAP7_75t_L g403 ( 
.A(n_359),
.B(n_347),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_SL g404 ( 
.A1(n_379),
.A2(n_338),
.B1(n_331),
.B2(n_321),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_L g405 ( 
.A1(n_385),
.A2(n_341),
.B1(n_352),
.B2(n_354),
.Y(n_405)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_405),
.Y(n_442)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_358),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_406),
.B(n_411),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_363),
.Y(n_407)
);

AOI21x1_ASAP7_75t_SL g408 ( 
.A1(n_376),
.A2(n_351),
.B(n_344),
.Y(n_408)
);

OAI21xp5_ASAP7_75t_SL g438 ( 
.A1(n_408),
.A2(n_382),
.B(n_3),
.Y(n_438)
);

INVxp67_ASAP7_75t_L g409 ( 
.A(n_375),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_409),
.B(n_413),
.Y(n_419)
);

AOI21xp5_ASAP7_75t_L g443 ( 
.A1(n_410),
.A2(n_39),
.B(n_33),
.Y(n_443)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_362),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_SL g412 ( 
.A(n_372),
.B(n_10),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_412),
.B(n_384),
.Y(n_435)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_364),
.Y(n_413)
);

HB1xp67_ASAP7_75t_L g414 ( 
.A(n_367),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_414),
.B(n_355),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_L g416 ( 
.A(n_371),
.B(n_34),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_416),
.B(n_417),
.C(n_380),
.Y(n_430)
);

AND2x2_ASAP7_75t_L g420 ( 
.A(n_404),
.B(n_377),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_420),
.B(n_435),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_SL g422 ( 
.A1(n_393),
.A2(n_386),
.B1(n_380),
.B2(n_385),
.Y(n_422)
);

AOI22xp5_ASAP7_75t_SL g462 ( 
.A1(n_422),
.A2(n_431),
.B1(n_439),
.B2(n_4),
.Y(n_462)
);

BUFx4f_ASAP7_75t_SL g425 ( 
.A(n_408),
.Y(n_425)
);

HB1xp67_ASAP7_75t_L g445 ( 
.A(n_425),
.Y(n_445)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_426),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_L g451 ( 
.A(n_430),
.B(n_403),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_SL g431 ( 
.A1(n_391),
.A2(n_357),
.B1(n_361),
.B2(n_369),
.Y(n_431)
);

AOI21xp5_ASAP7_75t_L g432 ( 
.A1(n_410),
.A2(n_373),
.B(n_388),
.Y(n_432)
);

AOI21xp5_ASAP7_75t_L g455 ( 
.A1(n_432),
.A2(n_436),
.B(n_11),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_L g448 ( 
.A1(n_433),
.A2(n_440),
.B1(n_417),
.B2(n_416),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_SL g436 ( 
.A(n_409),
.B(n_382),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_391),
.B(n_382),
.Y(n_437)
);

AND2x2_ASAP7_75t_L g460 ( 
.A(n_437),
.B(n_438),
.Y(n_460)
);

OAI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_402),
.A2(n_394),
.B1(n_396),
.B2(n_390),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_415),
.A2(n_11),
.B1(n_3),
.B2(n_4),
.Y(n_440)
);

XOR2xp5_ASAP7_75t_L g452 ( 
.A(n_443),
.B(n_33),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_429),
.B(n_396),
.C(n_401),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_446),
.B(n_448),
.Y(n_465)
);

MAJx2_ASAP7_75t_L g447 ( 
.A(n_429),
.B(n_397),
.C(n_418),
.Y(n_447)
);

AOI21xp5_ASAP7_75t_SL g477 ( 
.A1(n_447),
.A2(n_446),
.B(n_461),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_SL g449 ( 
.A(n_419),
.B(n_418),
.C(n_399),
.Y(n_449)
);

BUFx24_ASAP7_75t_SL g467 ( 
.A(n_449),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_434),
.B(n_415),
.C(n_399),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_450),
.B(n_451),
.Y(n_481)
);

XOR2xp5_ASAP7_75t_L g472 ( 
.A(n_452),
.B(n_461),
.Y(n_472)
);

BUFx24_ASAP7_75t_SL g453 ( 
.A(n_441),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_453),
.B(n_456),
.Y(n_468)
);

AOI21xp5_ASAP7_75t_L g466 ( 
.A1(n_455),
.A2(n_459),
.B(n_443),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_SL g456 ( 
.A(n_423),
.B(n_0),
.Y(n_456)
);

BUFx24_ASAP7_75t_SL g457 ( 
.A(n_423),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_457),
.B(n_458),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_434),
.B(n_34),
.C(n_30),
.Y(n_458)
);

AOI21xp5_ASAP7_75t_L g459 ( 
.A1(n_419),
.A2(n_33),
.B(n_30),
.Y(n_459)
);

XOR2xp5_ASAP7_75t_L g461 ( 
.A(n_439),
.B(n_33),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_SL g470 ( 
.A1(n_462),
.A2(n_433),
.B1(n_440),
.B2(n_424),
.Y(n_470)
);

OAI22xp5_ASAP7_75t_L g463 ( 
.A1(n_442),
.A2(n_30),
.B1(n_34),
.B2(n_6),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_463),
.Y(n_464)
);

HB1xp67_ASAP7_75t_L g495 ( 
.A(n_466),
.Y(n_495)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_445),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_469),
.B(n_471),
.Y(n_483)
);

AOI22xp5_ASAP7_75t_L g482 ( 
.A1(n_470),
.A2(n_431),
.B1(n_427),
.B2(n_420),
.Y(n_482)
);

OAI321xp33_ASAP7_75t_L g471 ( 
.A1(n_444),
.A2(n_437),
.A3(n_426),
.B1(n_421),
.B2(n_436),
.C(n_442),
.Y(n_471)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_454),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_473),
.B(n_475),
.Y(n_487)
);

XOR2xp5_ASAP7_75t_L g474 ( 
.A(n_450),
.B(n_422),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_L g496 ( 
.A(n_474),
.B(n_472),
.Y(n_496)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_460),
.Y(n_475)
);

BUFx2_ASAP7_75t_L g476 ( 
.A(n_460),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_476),
.B(n_478),
.Y(n_491)
);

XNOR2xp5_ASAP7_75t_L g493 ( 
.A(n_477),
.B(n_447),
.Y(n_493)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_458),
.Y(n_478)
);

AND2x2_ASAP7_75t_L g480 ( 
.A(n_452),
.B(n_421),
.Y(n_480)
);

INVxp67_ASAP7_75t_L g488 ( 
.A(n_480),
.Y(n_488)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_482),
.Y(n_502)
);

AOI22xp5_ASAP7_75t_L g484 ( 
.A1(n_476),
.A2(n_427),
.B1(n_424),
.B2(n_420),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_484),
.B(n_485),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_465),
.B(n_428),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_468),
.B(n_425),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_SL g506 ( 
.A(n_486),
.B(n_489),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_481),
.B(n_425),
.Y(n_489)
);

AOI22xp5_ASAP7_75t_L g490 ( 
.A1(n_470),
.A2(n_430),
.B1(n_425),
.B2(n_432),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_SL g500 ( 
.A(n_490),
.B(n_496),
.Y(n_500)
);

XOR2xp5_ASAP7_75t_L g492 ( 
.A(n_474),
.B(n_477),
.Y(n_492)
);

AND2x2_ASAP7_75t_L g503 ( 
.A(n_492),
.B(n_493),
.Y(n_503)
);

XOR2xp5_ASAP7_75t_L g494 ( 
.A(n_480),
.B(n_438),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_494),
.B(n_472),
.Y(n_497)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_497),
.Y(n_512)
);

NAND2xp33_ASAP7_75t_SL g499 ( 
.A(n_483),
.B(n_464),
.Y(n_499)
);

OAI21xp5_ASAP7_75t_L g513 ( 
.A1(n_499),
.A2(n_501),
.B(n_504),
.Y(n_513)
);

OAI21xp5_ASAP7_75t_L g501 ( 
.A1(n_487),
.A2(n_491),
.B(n_467),
.Y(n_501)
);

OAI21xp5_ASAP7_75t_SL g504 ( 
.A1(n_488),
.A2(n_479),
.B(n_466),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_492),
.B(n_435),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_505),
.B(n_507),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_496),
.B(n_4),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_SL g508 ( 
.A(n_488),
.B(n_5),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_508),
.B(n_6),
.Y(n_515)
);

OAI22xp5_ASAP7_75t_L g509 ( 
.A1(n_498),
.A2(n_495),
.B1(n_494),
.B2(n_34),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_509),
.B(n_511),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_SL g510 ( 
.A(n_506),
.B(n_5),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_510),
.B(n_515),
.Y(n_517)
);

FAx1_ASAP7_75t_SL g511 ( 
.A(n_499),
.B(n_6),
.CI(n_7),
.CON(n_511),
.SN(n_511)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_500),
.B(n_6),
.Y(n_516)
);

OAI21x1_ASAP7_75t_SL g520 ( 
.A1(n_516),
.A2(n_503),
.B(n_7),
.Y(n_520)
);

MAJx2_ASAP7_75t_L g518 ( 
.A(n_512),
.B(n_503),
.C(n_502),
.Y(n_518)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_518),
.Y(n_521)
);

CKINVDCx20_ASAP7_75t_R g522 ( 
.A(n_520),
.Y(n_522)
);

AOI21x1_ASAP7_75t_L g523 ( 
.A1(n_521),
.A2(n_513),
.B(n_519),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_523),
.B(n_522),
.C(n_516),
.Y(n_524)
);

OAI21xp5_ASAP7_75t_L g525 ( 
.A1(n_524),
.A2(n_514),
.B(n_517),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_525),
.B(n_511),
.C(n_7),
.Y(n_526)
);


endmodule