module fake_jpeg_23149_n_88 (n_13, n_21, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_88);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_88;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_24;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_17),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_7),
.B(n_10),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_21),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_12),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_11),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_6),
.B(n_1),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_15),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_3),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_6),
.B(n_5),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_14),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_35),
.A2(n_5),
.B1(n_1),
.B2(n_2),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_44),
.B(n_49),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_47),
.B(n_53),
.Y(n_64)
);

AOI21xp5_ASAP7_75t_L g48 ( 
.A1(n_29),
.A2(n_2),
.B(n_26),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_42),
.B(n_41),
.Y(n_49)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_26),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_51),
.B(n_52),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_27),
.B(n_36),
.Y(n_52)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_28),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_22),
.B(n_33),
.Y(n_54)
);

AOI21xp33_ASAP7_75t_L g62 ( 
.A1(n_54),
.A2(n_55),
.B(n_56),
.Y(n_62)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_24),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_31),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_28),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_25),
.A2(n_32),
.B1(n_37),
.B2(n_43),
.Y(n_59)
);

HAxp5_ASAP7_75t_SL g60 ( 
.A(n_23),
.B(n_39),
.CON(n_60),
.SN(n_60)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_34),
.B(n_38),
.Y(n_61)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_64),
.Y(n_70)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_70),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_68),
.B(n_59),
.C(n_58),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_L g78 ( 
.A1(n_71),
.A2(n_74),
.B(n_60),
.Y(n_78)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_63),
.Y(n_72)
);

AO21x2_ASAP7_75t_L g76 ( 
.A1(n_72),
.A2(n_73),
.B(n_51),
.Y(n_76)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_63),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_62),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_76),
.B(n_77),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_72),
.A2(n_67),
.B1(n_66),
.B2(n_60),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_L g79 ( 
.A(n_78),
.B(n_58),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_79),
.A2(n_57),
.B(n_58),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_80),
.A2(n_76),
.B1(n_75),
.B2(n_50),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_SL g83 ( 
.A1(n_81),
.A2(n_82),
.B(n_65),
.Y(n_83)
);

XOR2xp5_ASAP7_75t_L g85 ( 
.A(n_83),
.B(n_84),
.Y(n_85)
);

XNOR2x1_ASAP7_75t_L g84 ( 
.A(n_82),
.B(n_23),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_85),
.A2(n_65),
.B1(n_39),
.B2(n_69),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g87 ( 
.A1(n_86),
.A2(n_69),
.B(n_23),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_87),
.B(n_61),
.Y(n_88)
);


endmodule