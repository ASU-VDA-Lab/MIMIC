module real_aes_8501_n_77 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_77);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_77;
wire n_480;
wire n_113;
wire n_476;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_522;
wire n_485;
wire n_222;
wire n_287;
wire n_503;
wire n_357;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_341;
wire n_232;
wire n_460;
wire n_401;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_320;
wire n_260;
wire n_97;
wire n_186;
wire n_138;
wire n_379;
wire n_374;
wire n_453;
wire n_235;
wire n_399;
wire n_378;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_145;
wire n_415;
wire n_227;
wire n_519;
wire n_92;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_292;
wire n_400;
wire n_116;
wire n_94;
wire n_289;
wire n_462;
wire n_280;
wire n_333;
wire n_213;
wire n_478;
wire n_356;
wire n_408;
wire n_184;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_530;
wire n_104;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_506;
wire n_513;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_164;
wire n_231;
wire n_102;
wire n_454;
wire n_122;
wire n_443;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_204;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_331;
wire n_93;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_323;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_368;
wire n_502;
wire n_527;
wire n_505;
wire n_434;
wire n_250;
wire n_85;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_402;
wire n_87;
wire n_171;
wire n_78;
wire n_531;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_501;
wire n_488;
wire n_251;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_95;
wire n_188;
wire n_430;
wire n_269;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_158;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_109;
wire n_203;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_526;
wire n_155;
wire n_243;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_446;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_524;
wire n_219;
wire n_180;
wire n_212;
wire n_210;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_103;
wire n_166;
wire n_224;
wire n_151;
wire n_130;
wire n_253;
wire n_459;
wire n_99;
wire n_440;
wire n_525;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_305;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_465;
wire n_473;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_340;
wire n_483;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_206;
wire n_307;
wire n_500;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_264;
wire n_237;
wire n_91;
AOI22xp5_ASAP7_75t_SL g160 ( .A1(n_0), .A2(n_21), .B1(n_161), .B2(n_164), .Y(n_160) );
A2O1A1Ixp33_ASAP7_75t_L g272 ( .A1(n_1), .A2(n_189), .B(n_192), .C(n_273), .Y(n_272) );
INVx1_ASAP7_75t_L g532 ( .A(n_1), .Y(n_532) );
AOI21xp5_ASAP7_75t_L g299 ( .A1(n_2), .A2(n_222), .B(n_300), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_3), .B(n_289), .Y(n_308) );
INVx1_ASAP7_75t_L g175 ( .A(n_4), .Y(n_175) );
AND2x6_ASAP7_75t_L g189 ( .A(n_4), .B(n_173), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_4), .B(n_526), .Y(n_525) );
INVx1_ASAP7_75t_L g263 ( .A(n_5), .Y(n_263) );
NAND2xp5_ASAP7_75t_SL g275 ( .A(n_6), .B(n_200), .Y(n_275) );
AOI22xp5_ASAP7_75t_SL g154 ( .A1(n_7), .A2(n_76), .B1(n_155), .B2(n_157), .Y(n_154) );
AO22x2_ASAP7_75t_L g88 ( .A1(n_8), .A2(n_28), .B1(n_89), .B2(n_90), .Y(n_88) );
INVx1_ASAP7_75t_L g208 ( .A(n_9), .Y(n_208) );
A2O1A1Ixp33_ASAP7_75t_L g284 ( .A1(n_10), .A2(n_198), .B(n_285), .C(n_287), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_11), .B(n_289), .Y(n_288) );
AOI22xp5_ASAP7_75t_SL g137 ( .A1(n_12), .A2(n_43), .B1(n_138), .B2(n_141), .Y(n_137) );
AO22x2_ASAP7_75t_L g92 ( .A1(n_13), .A2(n_30), .B1(n_89), .B2(n_93), .Y(n_92) );
AOI22xp5_ASAP7_75t_L g506 ( .A1(n_14), .A2(n_23), .B1(n_507), .B2(n_508), .Y(n_506) );
INVx1_ASAP7_75t_L g508 ( .A(n_14), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_15), .B(n_234), .Y(n_233) );
A2O1A1Ixp33_ASAP7_75t_L g317 ( .A1(n_16), .A2(n_303), .B(n_318), .C(n_320), .Y(n_317) );
AOI22xp5_ASAP7_75t_L g509 ( .A1(n_16), .A2(n_510), .B1(n_511), .B2(n_512), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_16), .Y(n_510) );
NAND2xp5_ASAP7_75t_SL g245 ( .A(n_17), .B(n_200), .Y(n_245) );
NAND2xp5_ASAP7_75t_SL g199 ( .A(n_18), .B(n_200), .Y(n_199) );
CKINVDCx16_ASAP7_75t_R g239 ( .A(n_19), .Y(n_239) );
INVx1_ASAP7_75t_L g196 ( .A(n_20), .Y(n_196) );
BUFx6f_ASAP7_75t_L g188 ( .A(n_22), .Y(n_188) );
INVxp67_ASAP7_75t_L g507 ( .A(n_23), .Y(n_507) );
CKINVDCx20_ASAP7_75t_R g271 ( .A(n_24), .Y(n_271) );
AOI22xp33_ASAP7_75t_SL g127 ( .A1(n_25), .A2(n_71), .B1(n_128), .B2(n_132), .Y(n_127) );
INVx1_ASAP7_75t_L g228 ( .A(n_26), .Y(n_228) );
INVx2_ASAP7_75t_L g187 ( .A(n_27), .Y(n_187) );
CKINVDCx20_ASAP7_75t_R g277 ( .A(n_29), .Y(n_277) );
OAI221xp5_ASAP7_75t_L g518 ( .A1(n_30), .A2(n_45), .B1(n_55), .B2(n_519), .C(n_520), .Y(n_518) );
INVxp67_ASAP7_75t_L g521 ( .A(n_30), .Y(n_521) );
NAND2xp5_ASAP7_75t_SL g120 ( .A(n_31), .B(n_121), .Y(n_120) );
A2O1A1Ixp33_ASAP7_75t_L g302 ( .A1(n_32), .A2(n_303), .B(n_304), .C(n_306), .Y(n_302) );
INVxp67_ASAP7_75t_L g229 ( .A(n_33), .Y(n_229) );
A2O1A1Ixp33_ASAP7_75t_L g191 ( .A1(n_34), .A2(n_192), .B(n_195), .C(n_203), .Y(n_191) );
CKINVDCx14_ASAP7_75t_R g301 ( .A(n_35), .Y(n_301) );
A2O1A1Ixp33_ASAP7_75t_L g260 ( .A1(n_36), .A2(n_247), .B(n_261), .C(n_262), .Y(n_260) );
AOI22xp33_ASAP7_75t_SL g100 ( .A1(n_37), .A2(n_52), .B1(n_101), .B2(n_109), .Y(n_100) );
CKINVDCx20_ASAP7_75t_R g210 ( .A(n_38), .Y(n_210) );
CKINVDCx20_ASAP7_75t_R g224 ( .A(n_39), .Y(n_224) );
OAI22xp5_ASAP7_75t_SL g512 ( .A1(n_40), .A2(n_44), .B1(n_513), .B2(n_514), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_40), .Y(n_513) );
INVx1_ASAP7_75t_L g316 ( .A(n_41), .Y(n_316) );
CKINVDCx20_ASAP7_75t_R g99 ( .A(n_42), .Y(n_99) );
INVx1_ASAP7_75t_L g514 ( .A(n_44), .Y(n_514) );
AO22x2_ASAP7_75t_L g96 ( .A1(n_45), .A2(n_66), .B1(n_89), .B2(n_93), .Y(n_96) );
INVxp67_ASAP7_75t_L g522 ( .A(n_45), .Y(n_522) );
CKINVDCx14_ASAP7_75t_R g259 ( .A(n_46), .Y(n_259) );
AOI22xp5_ASAP7_75t_SL g143 ( .A1(n_47), .A2(n_64), .B1(n_144), .B2(n_149), .Y(n_143) );
INVx1_ASAP7_75t_L g173 ( .A(n_48), .Y(n_173) );
INVx1_ASAP7_75t_L g207 ( .A(n_49), .Y(n_207) );
INVx1_ASAP7_75t_SL g305 ( .A(n_50), .Y(n_305) );
CKINVDCx20_ASAP7_75t_R g519 ( .A(n_51), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_53), .B(n_289), .Y(n_322) );
INVx1_ASAP7_75t_L g242 ( .A(n_54), .Y(n_242) );
AO22x2_ASAP7_75t_L g98 ( .A1(n_55), .A2(n_70), .B1(n_89), .B2(n_90), .Y(n_98) );
AOI22xp5_ASAP7_75t_SL g79 ( .A1(n_56), .A2(n_80), .B1(n_81), .B2(n_167), .Y(n_79) );
CKINVDCx20_ASAP7_75t_R g167 ( .A(n_56), .Y(n_167) );
AOI21xp5_ASAP7_75t_L g257 ( .A1(n_57), .A2(n_222), .B(n_258), .Y(n_257) );
CKINVDCx20_ASAP7_75t_R g251 ( .A(n_58), .Y(n_251) );
AOI21xp5_ASAP7_75t_L g281 ( .A1(n_59), .A2(n_222), .B(n_282), .Y(n_281) );
AOI21xp5_ASAP7_75t_L g220 ( .A1(n_60), .A2(n_221), .B(n_223), .Y(n_220) );
CKINVDCx16_ASAP7_75t_R g190 ( .A(n_61), .Y(n_190) );
INVx1_ASAP7_75t_L g283 ( .A(n_62), .Y(n_283) );
AOI21xp5_ASAP7_75t_L g314 ( .A1(n_63), .A2(n_222), .B(n_315), .Y(n_314) );
INVx1_ASAP7_75t_L g286 ( .A(n_65), .Y(n_286) );
INVx2_ASAP7_75t_L g205 ( .A(n_67), .Y(n_205) );
INVx1_ASAP7_75t_L g274 ( .A(n_68), .Y(n_274) );
AOI22xp5_ASAP7_75t_L g503 ( .A1(n_68), .A2(n_504), .B1(n_517), .B2(n_523), .Y(n_503) );
A2O1A1Ixp33_ASAP7_75t_L g240 ( .A1(n_69), .A2(n_192), .B(n_241), .C(n_249), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_72), .B(n_212), .Y(n_264) );
INVx1_ASAP7_75t_L g89 ( .A(n_73), .Y(n_89) );
INVx1_ASAP7_75t_L g91 ( .A(n_73), .Y(n_91) );
INVx2_ASAP7_75t_L g319 ( .A(n_74), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g113 ( .A(n_75), .B(n_114), .Y(n_113) );
AOI221xp5_ASAP7_75t_L g77 ( .A1(n_78), .A2(n_168), .B1(n_176), .B2(n_501), .C(n_502), .Y(n_77) );
CKINVDCx20_ASAP7_75t_R g78 ( .A(n_79), .Y(n_78) );
OAI322xp33_ASAP7_75t_L g502 ( .A1(n_80), .A2(n_503), .A3(n_527), .B1(n_528), .B2(n_529), .C1(n_532), .C2(n_533), .Y(n_502) );
CKINVDCx14_ASAP7_75t_R g80 ( .A(n_81), .Y(n_80) );
HB1xp67_ASAP7_75t_L g81 ( .A(n_82), .Y(n_81) );
NAND3x1_ASAP7_75t_L g82 ( .A(n_83), .B(n_136), .C(n_153), .Y(n_82) );
INVxp67_ASAP7_75t_L g528 ( .A(n_83), .Y(n_528) );
NOR2x1_ASAP7_75t_L g83 ( .A(n_84), .B(n_112), .Y(n_83) );
OAI21xp5_ASAP7_75t_SL g84 ( .A1(n_85), .A2(n_99), .B(n_100), .Y(n_84) );
INVx4_ASAP7_75t_L g85 ( .A(n_86), .Y(n_85) );
AND2x6_ASAP7_75t_L g86 ( .A(n_87), .B(n_94), .Y(n_86) );
AND2x4_ASAP7_75t_L g133 ( .A(n_87), .B(n_134), .Y(n_133) );
AND2x2_ASAP7_75t_L g87 ( .A(n_88), .B(n_92), .Y(n_87) );
AND2x2_ASAP7_75t_L g108 ( .A(n_88), .B(n_96), .Y(n_108) );
INVx2_ASAP7_75t_L g118 ( .A(n_88), .Y(n_118) );
INVx1_ASAP7_75t_L g90 ( .A(n_91), .Y(n_90) );
INVx1_ASAP7_75t_L g93 ( .A(n_91), .Y(n_93) );
INVx2_ASAP7_75t_L g107 ( .A(n_92), .Y(n_107) );
AND2x2_ASAP7_75t_L g117 ( .A(n_92), .B(n_118), .Y(n_117) );
OR2x2_ASAP7_75t_L g126 ( .A(n_92), .B(n_118), .Y(n_126) );
INVx1_ASAP7_75t_L g131 ( .A(n_92), .Y(n_131) );
AND2x2_ASAP7_75t_L g139 ( .A(n_94), .B(n_140), .Y(n_139) );
AND2x6_ASAP7_75t_L g163 ( .A(n_94), .B(n_125), .Y(n_163) );
AND2x4_ASAP7_75t_L g166 ( .A(n_94), .B(n_117), .Y(n_166) );
AND2x2_ASAP7_75t_L g94 ( .A(n_95), .B(n_97), .Y(n_94) );
AND2x2_ASAP7_75t_L g119 ( .A(n_95), .B(n_98), .Y(n_119) );
INVx2_ASAP7_75t_L g95 ( .A(n_96), .Y(n_95) );
AND2x2_ASAP7_75t_L g148 ( .A(n_96), .B(n_135), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_96), .B(n_98), .Y(n_152) );
INVx1_ASAP7_75t_L g97 ( .A(n_98), .Y(n_97) );
INVx1_ASAP7_75t_L g106 ( .A(n_98), .Y(n_106) );
INVx1_ASAP7_75t_L g135 ( .A(n_98), .Y(n_135) );
INVx3_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
INVx4_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
BUFx6f_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
AND2x4_ASAP7_75t_L g104 ( .A(n_105), .B(n_108), .Y(n_104) );
AND2x2_ASAP7_75t_L g105 ( .A(n_106), .B(n_107), .Y(n_105) );
INVx1_ASAP7_75t_L g111 ( .A(n_106), .Y(n_111) );
AND2x2_ASAP7_75t_L g140 ( .A(n_107), .B(n_118), .Y(n_140) );
AND2x4_ASAP7_75t_L g110 ( .A(n_108), .B(n_111), .Y(n_110) );
AND2x4_ASAP7_75t_L g129 ( .A(n_108), .B(n_130), .Y(n_129) );
BUFx12f_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
NAND3xp33_ASAP7_75t_L g112 ( .A(n_113), .B(n_120), .C(n_127), .Y(n_112) );
INVx1_ASAP7_75t_SL g114 ( .A(n_115), .Y(n_114) );
INVx1_ASAP7_75t_SL g115 ( .A(n_116), .Y(n_115) );
AND2x6_ASAP7_75t_L g116 ( .A(n_117), .B(n_119), .Y(n_116) );
AND2x2_ASAP7_75t_L g147 ( .A(n_117), .B(n_148), .Y(n_147) );
AND2x4_ASAP7_75t_L g124 ( .A(n_119), .B(n_125), .Y(n_124) );
AND2x4_ASAP7_75t_L g142 ( .A(n_119), .B(n_140), .Y(n_142) );
BUFx6f_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
INVx5_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
INVx4_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
INVx2_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
BUFx3_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
INVx1_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
OR2x6_ASAP7_75t_L g151 ( .A(n_131), .B(n_152), .Y(n_151) );
BUFx2_ASAP7_75t_SL g132 ( .A(n_133), .Y(n_132) );
INVx1_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
AND2x2_ASAP7_75t_L g136 ( .A(n_137), .B(n_143), .Y(n_136) );
NAND4xp25_ASAP7_75t_L g527 ( .A(n_137), .B(n_143), .C(n_154), .D(n_160), .Y(n_527) );
BUFx2_ASAP7_75t_SL g138 ( .A(n_139), .Y(n_138) );
AND2x2_ASAP7_75t_L g156 ( .A(n_140), .B(n_148), .Y(n_156) );
AND2x4_ASAP7_75t_L g158 ( .A(n_140), .B(n_159), .Y(n_158) );
BUFx3_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
BUFx2_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx4_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx8_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
BUFx2_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx6_ASAP7_75t_SL g150 ( .A(n_151), .Y(n_150) );
INVx1_ASAP7_75t_L g159 ( .A(n_152), .Y(n_159) );
AND2x2_ASAP7_75t_L g153 ( .A(n_154), .B(n_160), .Y(n_153) );
BUFx3_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
BUFx2_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx2_ASAP7_75t_SL g161 ( .A(n_162), .Y(n_161) );
INVx11_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
INVx2_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
INVx6_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
CKINVDCx20_ASAP7_75t_R g168 ( .A(n_169), .Y(n_168) );
OR2x2_ASAP7_75t_SL g169 ( .A(n_170), .B(n_174), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
AND3x1_ASAP7_75t_SL g517 ( .A(n_171), .B(n_174), .C(n_518), .Y(n_517) );
AND2x2_ASAP7_75t_L g523 ( .A(n_171), .B(n_524), .Y(n_523) );
OAI21xp5_ASAP7_75t_L g530 ( .A1(n_171), .A2(n_192), .B(n_531), .Y(n_530) );
INVx1_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
NAND2xp5_ASAP7_75t_SL g531 ( .A(n_172), .B(n_175), .Y(n_531) );
HB1xp67_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
CKINVDCx20_ASAP7_75t_R g174 ( .A(n_175), .Y(n_174) );
HB1xp67_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
OR4x2_ASAP7_75t_L g177 ( .A(n_178), .B(n_391), .C(n_438), .D(n_478), .Y(n_177) );
NAND3xp33_ASAP7_75t_SL g178 ( .A(n_179), .B(n_337), .C(n_366), .Y(n_178) );
AOI211xp5_ASAP7_75t_L g179 ( .A1(n_180), .A2(n_252), .B(n_290), .C(n_330), .Y(n_179) );
O2A1O1Ixp33_ASAP7_75t_L g366 ( .A1(n_180), .A2(n_350), .B(n_367), .C(n_371), .Y(n_366) );
INVx1_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_182), .B(n_214), .Y(n_181) );
NAND2xp5_ASAP7_75t_SL g328 ( .A(n_182), .B(n_329), .Y(n_328) );
INVx3_ASAP7_75t_SL g333 ( .A(n_182), .Y(n_333) );
HB1xp67_ASAP7_75t_L g345 ( .A(n_182), .Y(n_345) );
AND2x4_ASAP7_75t_L g349 ( .A(n_182), .B(n_297), .Y(n_349) );
AND2x2_ASAP7_75t_L g360 ( .A(n_182), .B(n_237), .Y(n_360) );
OR2x2_ASAP7_75t_L g384 ( .A(n_182), .B(n_293), .Y(n_384) );
AND2x2_ASAP7_75t_L g397 ( .A(n_182), .B(n_298), .Y(n_397) );
AND2x2_ASAP7_75t_L g437 ( .A(n_182), .B(n_423), .Y(n_437) );
AND2x2_ASAP7_75t_L g444 ( .A(n_182), .B(n_407), .Y(n_444) );
AND2x2_ASAP7_75t_L g474 ( .A(n_182), .B(n_215), .Y(n_474) );
OR2x6_ASAP7_75t_L g182 ( .A(n_183), .B(n_209), .Y(n_182) );
O2A1O1Ixp33_ASAP7_75t_L g183 ( .A1(n_184), .A2(n_190), .B(n_191), .C(n_204), .Y(n_183) );
OAI21xp5_ASAP7_75t_L g238 ( .A1(n_184), .A2(n_239), .B(n_240), .Y(n_238) );
OAI21xp5_ASAP7_75t_L g270 ( .A1(n_184), .A2(n_271), .B(n_272), .Y(n_270) );
NAND2x1p5_ASAP7_75t_L g184 ( .A(n_185), .B(n_189), .Y(n_184) );
AND2x4_ASAP7_75t_L g222 ( .A(n_185), .B(n_189), .Y(n_222) );
AND2x2_ASAP7_75t_L g185 ( .A(n_186), .B(n_188), .Y(n_185) );
INVx1_ASAP7_75t_L g202 ( .A(n_186), .Y(n_202) );
INVx1_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
INVx2_ASAP7_75t_L g193 ( .A(n_187), .Y(n_193) );
INVx1_ASAP7_75t_L g321 ( .A(n_187), .Y(n_321) );
INVx1_ASAP7_75t_L g194 ( .A(n_188), .Y(n_194) );
INVx3_ASAP7_75t_L g198 ( .A(n_188), .Y(n_198) );
BUFx6f_ASAP7_75t_L g200 ( .A(n_188), .Y(n_200) );
BUFx6f_ASAP7_75t_L g231 ( .A(n_188), .Y(n_231) );
BUFx3_ASAP7_75t_L g203 ( .A(n_189), .Y(n_203) );
INVx4_ASAP7_75t_SL g232 ( .A(n_189), .Y(n_232) );
INVx5_ASAP7_75t_L g225 ( .A(n_192), .Y(n_225) );
AND2x2_ASAP7_75t_L g501 ( .A(n_192), .B(n_203), .Y(n_501) );
AND2x6_ASAP7_75t_L g192 ( .A(n_193), .B(n_194), .Y(n_192) );
BUFx3_ASAP7_75t_L g248 ( .A(n_193), .Y(n_248) );
BUFx6f_ASAP7_75t_L g307 ( .A(n_193), .Y(n_307) );
O2A1O1Ixp33_ASAP7_75t_L g195 ( .A1(n_196), .A2(n_197), .B(n_199), .C(n_201), .Y(n_195) );
OAI22xp33_ASAP7_75t_L g227 ( .A1(n_197), .A2(n_228), .B1(n_229), .B2(n_230), .Y(n_227) );
INVx5_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
NOR2xp33_ASAP7_75t_L g262 ( .A(n_198), .B(n_263), .Y(n_262) );
INVx2_ASAP7_75t_L g261 ( .A(n_200), .Y(n_261) );
INVx4_ASAP7_75t_L g303 ( .A(n_200), .Y(n_303) );
INVx2_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
NAND2xp5_ASAP7_75t_SL g226 ( .A(n_202), .B(n_227), .Y(n_226) );
INVx2_ASAP7_75t_L g235 ( .A(n_204), .Y(n_235) );
OA21x2_ASAP7_75t_L g256 ( .A1(n_204), .A2(n_257), .B(n_264), .Y(n_256) );
INVx1_ASAP7_75t_L g269 ( .A(n_204), .Y(n_269) );
AND2x2_ASAP7_75t_SL g204 ( .A(n_205), .B(n_206), .Y(n_204) );
AND2x2_ASAP7_75t_L g213 ( .A(n_205), .B(n_206), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_207), .B(n_208), .Y(n_206) );
NOR2xp33_ASAP7_75t_L g209 ( .A(n_210), .B(n_211), .Y(n_209) );
AO21x2_ASAP7_75t_L g237 ( .A1(n_211), .A2(n_238), .B(n_250), .Y(n_237) );
NOR2xp33_ASAP7_75t_L g276 ( .A(n_211), .B(n_277), .Y(n_276) );
INVx3_ASAP7_75t_L g289 ( .A(n_211), .Y(n_289) );
INVx4_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
HB1xp67_ASAP7_75t_L g280 ( .A(n_212), .Y(n_280) );
BUFx6f_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
INVx1_ASAP7_75t_L g219 ( .A(n_213), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_214), .B(n_401), .Y(n_413) );
AND2x2_ASAP7_75t_L g214 ( .A(n_215), .B(n_236), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_215), .B(n_344), .Y(n_343) );
OR2x2_ASAP7_75t_L g351 ( .A(n_215), .B(n_236), .Y(n_351) );
BUFx3_ASAP7_75t_L g359 ( .A(n_215), .Y(n_359) );
OR2x2_ASAP7_75t_L g380 ( .A(n_215), .B(n_255), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_215), .B(n_401), .Y(n_491) );
OA21x2_ASAP7_75t_L g215 ( .A1(n_216), .A2(n_220), .B(n_233), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
AO21x2_ASAP7_75t_L g293 ( .A1(n_217), .A2(n_294), .B(n_295), .Y(n_293) );
INVx1_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
INVx2_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
INVx1_ASAP7_75t_L g294 ( .A(n_220), .Y(n_294) );
BUFx2_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
O2A1O1Ixp33_ASAP7_75t_SL g223 ( .A1(n_224), .A2(n_225), .B(n_226), .C(n_232), .Y(n_223) );
O2A1O1Ixp33_ASAP7_75t_SL g258 ( .A1(n_225), .A2(n_232), .B(n_259), .C(n_260), .Y(n_258) );
O2A1O1Ixp33_ASAP7_75t_SL g282 ( .A1(n_225), .A2(n_232), .B(n_283), .C(n_284), .Y(n_282) );
O2A1O1Ixp33_ASAP7_75t_L g300 ( .A1(n_225), .A2(n_232), .B(n_301), .C(n_302), .Y(n_300) );
O2A1O1Ixp33_ASAP7_75t_SL g315 ( .A1(n_225), .A2(n_232), .B(n_316), .C(n_317), .Y(n_315) );
NOR2xp33_ASAP7_75t_L g285 ( .A(n_230), .B(n_286), .Y(n_285) );
NOR2xp33_ASAP7_75t_L g318 ( .A(n_230), .B(n_319), .Y(n_318) );
INVx4_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
INVx2_ASAP7_75t_L g244 ( .A(n_231), .Y(n_244) );
INVx1_ASAP7_75t_L g249 ( .A(n_232), .Y(n_249) );
INVx1_ASAP7_75t_L g295 ( .A(n_233), .Y(n_295) );
INVx1_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
NOR2xp33_ASAP7_75t_L g250 ( .A(n_235), .B(n_251), .Y(n_250) );
AND2x2_ASAP7_75t_L g296 ( .A(n_236), .B(n_297), .Y(n_296) );
INVx1_ASAP7_75t_L g344 ( .A(n_236), .Y(n_344) );
AND2x2_ASAP7_75t_L g407 ( .A(n_236), .B(n_298), .Y(n_407) );
AOI221xp5_ASAP7_75t_L g409 ( .A1(n_236), .A2(n_410), .B1(n_412), .B2(n_414), .C(n_415), .Y(n_409) );
AND2x2_ASAP7_75t_L g423 ( .A(n_236), .B(n_293), .Y(n_423) );
AND2x2_ASAP7_75t_L g449 ( .A(n_236), .B(n_333), .Y(n_449) );
INVx2_ASAP7_75t_SL g236 ( .A(n_237), .Y(n_236) );
AND2x2_ASAP7_75t_L g329 ( .A(n_237), .B(n_298), .Y(n_329) );
BUFx2_ASAP7_75t_L g463 ( .A(n_237), .Y(n_463) );
O2A1O1Ixp33_ASAP7_75t_L g241 ( .A1(n_242), .A2(n_243), .B(n_245), .C(n_246), .Y(n_241) );
O2A1O1Ixp5_ASAP7_75t_L g273 ( .A1(n_243), .A2(n_246), .B(n_274), .C(n_275), .Y(n_273) );
INVx2_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
INVx2_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
INVx2_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
INVx1_ASAP7_75t_L g287 ( .A(n_248), .Y(n_287) );
INVx1_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
OAI32xp33_ASAP7_75t_L g429 ( .A1(n_253), .A2(n_390), .A3(n_404), .B1(n_430), .B2(n_431), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_254), .B(n_265), .Y(n_253) );
AND2x2_ASAP7_75t_L g370 ( .A(n_254), .B(n_312), .Y(n_370) );
INVx1_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
OR2x2_ASAP7_75t_L g352 ( .A(n_255), .B(n_353), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_255), .B(n_363), .Y(n_362) );
AND2x2_ASAP7_75t_L g424 ( .A(n_255), .B(n_312), .Y(n_424) );
AND2x2_ASAP7_75t_L g435 ( .A(n_255), .B(n_327), .Y(n_435) );
BUFx3_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
OR2x2_ASAP7_75t_L g336 ( .A(n_256), .B(n_313), .Y(n_336) );
AND2x2_ASAP7_75t_L g340 ( .A(n_256), .B(n_313), .Y(n_340) );
AND2x2_ASAP7_75t_L g375 ( .A(n_256), .B(n_326), .Y(n_375) );
AND2x2_ASAP7_75t_L g382 ( .A(n_256), .B(n_278), .Y(n_382) );
OAI211xp5_ASAP7_75t_L g387 ( .A1(n_256), .A2(n_333), .B(n_344), .C(n_388), .Y(n_387) );
INVx2_ASAP7_75t_L g441 ( .A(n_256), .Y(n_441) );
NOR2xp33_ASAP7_75t_L g452 ( .A(n_256), .B(n_267), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_265), .B(n_324), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_265), .B(n_340), .Y(n_430) );
INVx1_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
OR2x2_ASAP7_75t_L g335 ( .A(n_266), .B(n_336), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_267), .B(n_278), .Y(n_266) );
AND2x2_ASAP7_75t_L g327 ( .A(n_267), .B(n_279), .Y(n_327) );
OR2x2_ASAP7_75t_L g342 ( .A(n_267), .B(n_279), .Y(n_342) );
AND2x2_ASAP7_75t_L g365 ( .A(n_267), .B(n_326), .Y(n_365) );
INVx1_ASAP7_75t_L g369 ( .A(n_267), .Y(n_369) );
AND2x2_ASAP7_75t_L g388 ( .A(n_267), .B(n_325), .Y(n_388) );
OAI22xp33_ASAP7_75t_L g398 ( .A1(n_267), .A2(n_353), .B1(n_399), .B2(n_400), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_267), .B(n_441), .Y(n_465) );
AND2x2_ASAP7_75t_L g480 ( .A(n_267), .B(n_340), .Y(n_480) );
INVx4_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
BUFx3_ASAP7_75t_L g310 ( .A(n_268), .Y(n_310) );
AND2x2_ASAP7_75t_L g354 ( .A(n_268), .B(n_279), .Y(n_354) );
AND2x2_ASAP7_75t_L g356 ( .A(n_268), .B(n_312), .Y(n_356) );
AND3x2_ASAP7_75t_L g418 ( .A(n_268), .B(n_382), .C(n_419), .Y(n_418) );
AO21x2_ASAP7_75t_L g268 ( .A1(n_269), .A2(n_270), .B(n_276), .Y(n_268) );
AOI22xp5_ASAP7_75t_L g533 ( .A1(n_274), .A2(n_505), .B1(n_517), .B2(n_523), .Y(n_533) );
AND2x2_ASAP7_75t_L g453 ( .A(n_278), .B(n_325), .Y(n_453) );
INVx1_ASAP7_75t_SL g278 ( .A(n_279), .Y(n_278) );
AND2x2_ASAP7_75t_L g312 ( .A(n_279), .B(n_313), .Y(n_312) );
HB1xp67_ASAP7_75t_L g363 ( .A(n_279), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_279), .B(n_324), .Y(n_386) );
NAND3xp33_ASAP7_75t_L g493 ( .A(n_279), .B(n_365), .C(n_441), .Y(n_493) );
OA21x2_ASAP7_75t_L g279 ( .A1(n_280), .A2(n_281), .B(n_288), .Y(n_279) );
OA21x2_ASAP7_75t_L g298 ( .A1(n_280), .A2(n_299), .B(n_308), .Y(n_298) );
OA21x2_ASAP7_75t_L g313 ( .A1(n_280), .A2(n_314), .B(n_322), .Y(n_313) );
OAI22xp5_ASAP7_75t_L g290 ( .A1(n_291), .A2(n_309), .B1(n_323), .B2(n_328), .Y(n_290) );
INVx1_ASAP7_75t_SL g291 ( .A(n_292), .Y(n_291) );
AND2x2_ASAP7_75t_L g292 ( .A(n_293), .B(n_296), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_293), .B(n_390), .Y(n_389) );
INVx1_ASAP7_75t_SL g405 ( .A(n_293), .Y(n_405) );
OAI31xp33_ASAP7_75t_L g421 ( .A1(n_296), .A2(n_422), .A3(n_423), .B(n_424), .Y(n_421) );
AND2x2_ASAP7_75t_L g446 ( .A(n_296), .B(n_333), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_296), .B(n_359), .Y(n_492) );
AND2x2_ASAP7_75t_L g401 ( .A(n_297), .B(n_333), .Y(n_401) );
AND2x2_ASAP7_75t_L g462 ( .A(n_297), .B(n_463), .Y(n_462) );
INVx2_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
AND2x2_ASAP7_75t_L g332 ( .A(n_298), .B(n_333), .Y(n_332) );
INVx1_ASAP7_75t_L g390 ( .A(n_298), .Y(n_390) );
NOR2xp33_ASAP7_75t_L g304 ( .A(n_303), .B(n_305), .Y(n_304) );
INVx3_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
OR2x2_ASAP7_75t_L g309 ( .A(n_310), .B(n_311), .Y(n_309) );
CKINVDCx16_ASAP7_75t_R g411 ( .A(n_310), .Y(n_411) );
NOR2xp33_ASAP7_75t_L g464 ( .A(n_311), .B(n_465), .Y(n_464) );
INVx1_ASAP7_75t_SL g311 ( .A(n_312), .Y(n_311) );
AOI221x1_ASAP7_75t_SL g378 ( .A1(n_312), .A2(n_379), .B1(n_381), .B2(n_383), .C(n_385), .Y(n_378) );
INVx2_ASAP7_75t_L g326 ( .A(n_313), .Y(n_326) );
HB1xp67_ASAP7_75t_L g420 ( .A(n_313), .Y(n_420) );
INVx3_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
INVx1_ASAP7_75t_L g408 ( .A(n_323), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_324), .B(n_327), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_324), .B(n_341), .Y(n_433) );
INVx1_ASAP7_75t_SL g496 ( .A(n_324), .Y(n_496) );
INVx2_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
INVx2_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
AND2x2_ASAP7_75t_L g414 ( .A(n_327), .B(n_340), .Y(n_414) );
INVx1_ASAP7_75t_L g482 ( .A(n_328), .Y(n_482) );
NOR2xp33_ASAP7_75t_L g495 ( .A(n_328), .B(n_411), .Y(n_495) );
INVx2_ASAP7_75t_SL g334 ( .A(n_329), .Y(n_334) );
AND2x2_ASAP7_75t_L g377 ( .A(n_329), .B(n_333), .Y(n_377) );
NOR2xp33_ASAP7_75t_L g383 ( .A(n_329), .B(n_384), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_329), .B(n_404), .Y(n_431) );
AOI21xp33_ASAP7_75t_SL g330 ( .A1(n_331), .A2(n_334), .B(n_335), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_332), .B(n_404), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_332), .B(n_359), .Y(n_500) );
OR2x2_ASAP7_75t_L g372 ( .A(n_333), .B(n_351), .Y(n_372) );
AND2x2_ASAP7_75t_L g471 ( .A(n_333), .B(n_462), .Y(n_471) );
OAI22xp5_ASAP7_75t_SL g346 ( .A1(n_334), .A2(n_347), .B1(n_352), .B2(n_355), .Y(n_346) );
NOR2xp33_ASAP7_75t_L g379 ( .A(n_334), .B(n_380), .Y(n_379) );
OR2x2_ASAP7_75t_L g394 ( .A(n_336), .B(n_342), .Y(n_394) );
INVx1_ASAP7_75t_L g458 ( .A(n_336), .Y(n_458) );
AOI311xp33_ASAP7_75t_L g337 ( .A1(n_338), .A2(n_343), .A3(n_345), .B(n_346), .C(n_357), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_340), .B(n_341), .Y(n_339) );
AOI221xp5_ASAP7_75t_L g484 ( .A1(n_341), .A2(n_473), .B1(n_485), .B2(n_488), .C(n_490), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_341), .B(n_496), .Y(n_498) );
INVx2_ASAP7_75t_SL g341 ( .A(n_342), .Y(n_341) );
INVx1_ASAP7_75t_L g395 ( .A(n_343), .Y(n_395) );
AOI211xp5_ASAP7_75t_L g385 ( .A1(n_344), .A2(n_386), .B(n_387), .C(n_389), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_348), .B(n_350), .Y(n_347) );
O2A1O1Ixp33_ASAP7_75t_SL g454 ( .A1(n_348), .A2(n_350), .B(n_455), .C(n_456), .Y(n_454) );
INVx3_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_349), .B(n_423), .Y(n_489) );
INVx1_ASAP7_75t_SL g350 ( .A(n_351), .Y(n_350) );
OAI221xp5_ASAP7_75t_L g371 ( .A1(n_352), .A2(n_372), .B1(n_373), .B2(n_376), .C(n_378), .Y(n_371) );
INVx1_ASAP7_75t_SL g353 ( .A(n_354), .Y(n_353) );
AND2x2_ASAP7_75t_L g374 ( .A(n_354), .B(n_375), .Y(n_374) );
AND2x2_ASAP7_75t_L g457 ( .A(n_354), .B(n_458), .Y(n_457) );
INVx1_ASAP7_75t_SL g355 ( .A(n_356), .Y(n_355) );
NOR2xp33_ASAP7_75t_L g357 ( .A(n_358), .B(n_361), .Y(n_357) );
A2O1A1Ixp33_ASAP7_75t_L g415 ( .A1(n_358), .A2(n_416), .B(n_417), .C(n_421), .Y(n_415) );
NAND2xp5_ASAP7_75t_SL g358 ( .A(n_359), .B(n_360), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_359), .B(n_449), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_359), .B(n_462), .Y(n_461) );
OR2x2_ASAP7_75t_L g361 ( .A(n_362), .B(n_364), .Y(n_361) );
INVxp67_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
AND2x2_ASAP7_75t_L g381 ( .A(n_365), .B(n_382), .Y(n_381) );
INVx1_ASAP7_75t_SL g367 ( .A(n_368), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_369), .B(n_370), .Y(n_368) );
NOR2xp33_ASAP7_75t_L g440 ( .A(n_369), .B(n_441), .Y(n_440) );
INVx1_ASAP7_75t_L g483 ( .A(n_372), .Y(n_483) );
INVx1_ASAP7_75t_SL g373 ( .A(n_374), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_375), .B(n_404), .Y(n_403) );
AND2x2_ASAP7_75t_L g410 ( .A(n_375), .B(n_411), .Y(n_410) );
INVx1_ASAP7_75t_SL g487 ( .A(n_375), .Y(n_487) );
INVx1_ASAP7_75t_SL g376 ( .A(n_377), .Y(n_376) );
AND2x2_ASAP7_75t_L g428 ( .A(n_377), .B(n_404), .Y(n_428) );
INVx1_ASAP7_75t_SL g422 ( .A(n_384), .Y(n_422) );
INVx1_ASAP7_75t_L g399 ( .A(n_390), .Y(n_399) );
NAND3xp33_ASAP7_75t_SL g391 ( .A(n_392), .B(n_409), .C(n_425), .Y(n_391) );
AOI322xp5_ASAP7_75t_L g392 ( .A1(n_393), .A2(n_395), .A3(n_396), .B1(n_398), .B2(n_402), .C1(n_406), .C2(n_408), .Y(n_392) );
AOI211xp5_ASAP7_75t_L g445 ( .A1(n_393), .A2(n_446), .B(n_447), .C(n_454), .Y(n_445) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
OAI22xp5_ASAP7_75t_L g447 ( .A1(n_396), .A2(n_417), .B1(n_448), .B2(n_450), .Y(n_447) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
AND2x2_ASAP7_75t_L g406 ( .A(n_404), .B(n_407), .Y(n_406) );
AND2x2_ASAP7_75t_L g443 ( .A(n_404), .B(n_444), .Y(n_443) );
AOI32xp33_ASAP7_75t_L g494 ( .A1(n_404), .A2(n_495), .A3(n_496), .B1(n_497), .B2(n_499), .Y(n_494) );
INVx2_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g416 ( .A(n_407), .Y(n_416) );
AOI221xp5_ASAP7_75t_L g459 ( .A1(n_407), .A2(n_460), .B1(n_464), .B2(n_466), .C(n_469), .Y(n_459) );
AND2x2_ASAP7_75t_L g473 ( .A(n_407), .B(n_474), .Y(n_473) );
AND2x2_ASAP7_75t_L g476 ( .A(n_411), .B(n_477), .Y(n_476) );
OR2x2_ASAP7_75t_L g486 ( .A(n_411), .B(n_487), .Y(n_486) );
INVxp67_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx2_ASAP7_75t_SL g417 ( .A(n_418), .Y(n_417) );
INVxp67_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
AND2x2_ASAP7_75t_L g477 ( .A(n_420), .B(n_441), .Y(n_477) );
AOI211xp5_ASAP7_75t_L g425 ( .A1(n_426), .A2(n_428), .B(n_429), .C(n_432), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
AOI21xp33_ASAP7_75t_L g432 ( .A1(n_433), .A2(n_434), .B(n_436), .Y(n_432) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
OAI211xp5_ASAP7_75t_SL g438 ( .A1(n_439), .A2(n_442), .B(n_445), .C(n_459), .Y(n_438) );
INVxp67_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
AND2x2_ASAP7_75t_L g451 ( .A(n_452), .B(n_453), .Y(n_451) );
NAND2xp5_ASAP7_75t_SL g467 ( .A(n_453), .B(n_468), .Y(n_467) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVx1_ASAP7_75t_L g468 ( .A(n_465), .Y(n_468) );
INVx1_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
AOI21xp33_ASAP7_75t_L g469 ( .A1(n_470), .A2(n_472), .B(n_475), .Y(n_469) );
INVx1_ASAP7_75t_SL g470 ( .A(n_471), .Y(n_470) );
INVx1_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
INVx1_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
OAI211xp5_ASAP7_75t_SL g478 ( .A1(n_479), .A2(n_481), .B(n_484), .C(n_494), .Y(n_478) );
CKINVDCx20_ASAP7_75t_R g479 ( .A(n_480), .Y(n_479) );
NOR2xp33_ASAP7_75t_L g481 ( .A(n_482), .B(n_483), .Y(n_481) );
INVx1_ASAP7_75t_SL g485 ( .A(n_486), .Y(n_485) );
INVx1_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
AOI21xp33_ASAP7_75t_L g490 ( .A1(n_491), .A2(n_492), .B(n_493), .Y(n_490) );
INVx1_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
INVx1_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
CKINVDCx20_ASAP7_75t_R g504 ( .A(n_505), .Y(n_504) );
AOI22xp5_ASAP7_75t_L g505 ( .A1(n_506), .A2(n_509), .B1(n_515), .B2(n_516), .Y(n_505) );
CKINVDCx20_ASAP7_75t_R g515 ( .A(n_506), .Y(n_515) );
CKINVDCx20_ASAP7_75t_R g516 ( .A(n_509), .Y(n_516) );
INVx1_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
INVxp67_ASAP7_75t_L g526 ( .A(n_518), .Y(n_526) );
NOR2xp33_ASAP7_75t_L g520 ( .A(n_521), .B(n_522), .Y(n_520) );
CKINVDCx20_ASAP7_75t_R g524 ( .A(n_525), .Y(n_524) );
CKINVDCx20_ASAP7_75t_R g529 ( .A(n_530), .Y(n_529) );
endmodule