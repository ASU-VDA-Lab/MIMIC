module fake_netlist_6_77_n_370 (n_52, n_16, n_1, n_91, n_46, n_18, n_21, n_88, n_3, n_98, n_39, n_63, n_73, n_4, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_77, n_106, n_92, n_42, n_96, n_8, n_90, n_24, n_105, n_54, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_100, n_13, n_11, n_17, n_23, n_20, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_45, n_34, n_70, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_55, n_94, n_97, n_108, n_58, n_64, n_48, n_65, n_25, n_40, n_93, n_80, n_41, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_72, n_89, n_103, n_111, n_60, n_35, n_12, n_69, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_370);

input n_52;
input n_16;
input n_1;
input n_91;
input n_46;
input n_18;
input n_21;
input n_88;
input n_3;
input n_98;
input n_39;
input n_63;
input n_73;
input n_4;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_77;
input n_106;
input n_92;
input n_42;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_54;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_100;
input n_13;
input n_11;
input n_17;
input n_23;
input n_20;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_45;
input n_34;
input n_70;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_55;
input n_94;
input n_97;
input n_108;
input n_58;
input n_64;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_41;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_12;
input n_69;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_370;

wire n_326;
wire n_256;
wire n_209;
wire n_367;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_148;
wire n_226;
wire n_208;
wire n_161;
wire n_316;
wire n_304;
wire n_212;
wire n_144;
wire n_365;
wire n_125;
wire n_168;
wire n_297;
wire n_342;
wire n_358;
wire n_160;
wire n_131;
wire n_188;
wire n_310;
wire n_186;
wire n_245;
wire n_368;
wire n_350;
wire n_142;
wire n_143;
wire n_180;
wire n_349;
wire n_233;
wire n_255;
wire n_284;
wire n_140;
wire n_337;
wire n_214;
wire n_246;
wire n_289;
wire n_181;
wire n_182;
wire n_238;
wire n_202;
wire n_320;
wire n_327;
wire n_369;
wire n_280;
wire n_287;
wire n_353;
wire n_230;
wire n_141;
wire n_200;
wire n_176;
wire n_114;
wire n_198;
wire n_222;
wire n_179;
wire n_248;
wire n_300;
wire n_229;
wire n_305;
wire n_173;
wire n_250;
wire n_314;
wire n_183;
wire n_338;
wire n_360;
wire n_119;
wire n_235;
wire n_147;
wire n_191;
wire n_340;
wire n_344;
wire n_167;
wire n_174;
wire n_127;
wire n_153;
wire n_156;
wire n_145;
wire n_133;
wire n_189;
wire n_213;
wire n_294;
wire n_302;
wire n_129;
wire n_197;
wire n_137;
wire n_343;
wire n_155;
wire n_122;
wire n_218;
wire n_234;
wire n_236;
wire n_172;
wire n_270;
wire n_239;
wire n_126;
wire n_290;
wire n_220;
wire n_118;
wire n_224;
wire n_196;
wire n_352;
wire n_366;
wire n_272;
wire n_185;
wire n_348;
wire n_293;
wire n_334;
wire n_232;
wire n_163;
wire n_330;
wire n_298;
wire n_281;
wire n_258;
wire n_154;
wire n_260;
wire n_265;
wire n_313;
wire n_279;
wire n_252;
wire n_228;
wire n_356;
wire n_166;
wire n_184;
wire n_216;
wire n_363;
wire n_323;
wire n_152;
wire n_321;
wire n_331;
wire n_227;
wire n_132;
wire n_204;
wire n_261;
wire n_312;
wire n_130;
wire n_164;
wire n_292;
wire n_121;
wire n_307;
wire n_291;
wire n_219;
wire n_357;
wire n_150;
wire n_264;
wire n_263;
wire n_325;
wire n_329;
wire n_237;
wire n_244;
wire n_243;
wire n_124;
wire n_282;
wire n_116;
wire n_211;
wire n_175;
wire n_117;
wire n_322;
wire n_345;
wire n_231;
wire n_354;
wire n_240;
wire n_139;
wire n_319;
wire n_134;
wire n_273;
wire n_311;
wire n_253;
wire n_123;
wire n_136;
wire n_249;
wire n_201;
wire n_159;
wire n_157;
wire n_162;
wire n_115;
wire n_128;
wire n_241;
wire n_275;
wire n_276;
wire n_221;
wire n_146;
wire n_318;
wire n_303;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_346;
wire n_277;
wire n_113;
wire n_199;
wire n_138;
wire n_266;
wire n_296;
wire n_268;
wire n_271;
wire n_158;
wire n_217;
wire n_210;
wire n_299;
wire n_206;
wire n_333;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_355;
wire n_317;
wire n_149;
wire n_347;
wire n_328;
wire n_195;
wire n_285;
wire n_257;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_242;
wire n_324;
wire n_335;
wire n_205;
wire n_120;
wire n_251;
wire n_301;
wire n_274;
wire n_151;
wire n_267;
wire n_339;
wire n_315;
wire n_288;
wire n_135;
wire n_165;
wire n_351;
wire n_259;
wire n_177;
wire n_364;
wire n_295;
wire n_190;
wire n_262;
wire n_187;
wire n_361;
wire n_170;
wire n_332;
wire n_336;
wire n_194;
wire n_171;
wire n_192;
wire n_169;
wire n_283;

CKINVDCx5p33_ASAP7_75t_R g113 ( 
.A(n_61),
.Y(n_113)
);

CKINVDCx5p33_ASAP7_75t_R g114 ( 
.A(n_28),
.Y(n_114)
);

HB1xp67_ASAP7_75t_L g115 ( 
.A(n_90),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_103),
.Y(n_116)
);

INVxp67_ASAP7_75t_SL g117 ( 
.A(n_68),
.Y(n_117)
);

BUFx2_ASAP7_75t_L g118 ( 
.A(n_31),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_59),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_79),
.Y(n_120)
);

CKINVDCx5p33_ASAP7_75t_R g121 ( 
.A(n_94),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_29),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_84),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_107),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g125 ( 
.A(n_100),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_39),
.Y(n_126)
);

CKINVDCx5p33_ASAP7_75t_R g127 ( 
.A(n_15),
.Y(n_127)
);

CKINVDCx5p33_ASAP7_75t_R g128 ( 
.A(n_10),
.Y(n_128)
);

CKINVDCx5p33_ASAP7_75t_R g129 ( 
.A(n_41),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_74),
.Y(n_130)
);

CKINVDCx5p33_ASAP7_75t_R g131 ( 
.A(n_16),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_32),
.Y(n_132)
);

INVx1_ASAP7_75t_SL g133 ( 
.A(n_1),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g134 ( 
.A(n_92),
.Y(n_134)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_7),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_104),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_56),
.B(n_48),
.Y(n_137)
);

INVxp33_ASAP7_75t_L g138 ( 
.A(n_40),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_44),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_34),
.Y(n_140)
);

CKINVDCx5p33_ASAP7_75t_R g141 ( 
.A(n_54),
.Y(n_141)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_112),
.Y(n_142)
);

BUFx2_ASAP7_75t_L g143 ( 
.A(n_111),
.Y(n_143)
);

CKINVDCx5p33_ASAP7_75t_R g144 ( 
.A(n_77),
.Y(n_144)
);

CKINVDCx5p33_ASAP7_75t_R g145 ( 
.A(n_93),
.Y(n_145)
);

CKINVDCx5p33_ASAP7_75t_R g146 ( 
.A(n_55),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_14),
.Y(n_147)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_105),
.Y(n_148)
);

CKINVDCx5p33_ASAP7_75t_R g149 ( 
.A(n_70),
.Y(n_149)
);

INVx1_ASAP7_75t_SL g150 ( 
.A(n_51),
.Y(n_150)
);

INVxp67_ASAP7_75t_SL g151 ( 
.A(n_85),
.Y(n_151)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_58),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_80),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_72),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_45),
.Y(n_155)
);

INVx1_ASAP7_75t_SL g156 ( 
.A(n_43),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_11),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_2),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_75),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_1),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_23),
.Y(n_161)
);

BUFx10_ASAP7_75t_L g162 ( 
.A(n_5),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_47),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_50),
.Y(n_164)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_35),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_110),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_33),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_18),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_98),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_63),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_116),
.Y(n_171)
);

AND2x4_ASAP7_75t_L g172 ( 
.A(n_125),
.B(n_0),
.Y(n_172)
);

OAI21x1_ASAP7_75t_L g173 ( 
.A1(n_148),
.A2(n_57),
.B(n_108),
.Y(n_173)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_134),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_119),
.Y(n_175)
);

INVx5_ASAP7_75t_L g176 ( 
.A(n_122),
.Y(n_176)
);

CKINVDCx6p67_ASAP7_75t_R g177 ( 
.A(n_162),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_113),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_122),
.Y(n_179)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_162),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_122),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_148),
.B(n_0),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_120),
.Y(n_183)
);

HB1xp67_ASAP7_75t_L g184 ( 
.A(n_133),
.Y(n_184)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_158),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_123),
.Y(n_186)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_124),
.Y(n_187)
);

HB1xp67_ASAP7_75t_L g188 ( 
.A(n_133),
.Y(n_188)
);

OAI21x1_ASAP7_75t_L g189 ( 
.A1(n_135),
.A2(n_60),
.B(n_106),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_126),
.Y(n_190)
);

HB1xp67_ASAP7_75t_L g191 ( 
.A(n_160),
.Y(n_191)
);

OAI21xp33_ASAP7_75t_L g192 ( 
.A1(n_182),
.A2(n_138),
.B(n_115),
.Y(n_192)
);

OR2x2_ASAP7_75t_L g193 ( 
.A(n_184),
.B(n_118),
.Y(n_193)
);

OR2x2_ASAP7_75t_L g194 ( 
.A(n_184),
.B(n_143),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_171),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_179),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_175),
.Y(n_197)
);

NAND3xp33_ASAP7_75t_L g198 ( 
.A(n_182),
.B(n_188),
.C(n_190),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_179),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_179),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_183),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_178),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_185),
.B(n_150),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_186),
.Y(n_204)
);

BUFx4f_ASAP7_75t_L g205 ( 
.A(n_179),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_187),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_180),
.B(n_150),
.Y(n_207)
);

OR2x2_ASAP7_75t_L g208 ( 
.A(n_188),
.B(n_2),
.Y(n_208)
);

INVx5_ASAP7_75t_L g209 ( 
.A(n_181),
.Y(n_209)
);

INVx2_ASAP7_75t_SL g210 ( 
.A(n_180),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_181),
.Y(n_211)
);

NAND3xp33_ASAP7_75t_L g212 ( 
.A(n_172),
.B(n_137),
.C(n_124),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_181),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_174),
.B(n_114),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_177),
.Y(n_215)
);

BUFx3_ASAP7_75t_L g216 ( 
.A(n_185),
.Y(n_216)
);

BUFx2_ASAP7_75t_L g217 ( 
.A(n_191),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_195),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_203),
.B(n_191),
.Y(n_219)
);

AND2x6_ASAP7_75t_SL g220 ( 
.A(n_214),
.B(n_172),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_192),
.B(n_156),
.Y(n_221)
);

AND3x1_ASAP7_75t_L g222 ( 
.A(n_192),
.B(n_136),
.C(n_154),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_214),
.B(n_176),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_210),
.B(n_147),
.Y(n_224)
);

OR2x6_ASAP7_75t_L g225 ( 
.A(n_217),
.B(n_130),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_193),
.Y(n_226)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_196),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_212),
.B(n_176),
.Y(n_228)
);

BUFx12f_ASAP7_75t_L g229 ( 
.A(n_215),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_198),
.B(n_207),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_198),
.B(n_163),
.Y(n_231)
);

AOI221xp5_ASAP7_75t_L g232 ( 
.A1(n_208),
.A2(n_140),
.B1(n_170),
.B2(n_155),
.C(n_161),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_205),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_212),
.B(n_176),
.Y(n_234)
);

AND2x6_ASAP7_75t_L g235 ( 
.A(n_216),
.B(n_139),
.Y(n_235)
);

AND2x2_ASAP7_75t_L g236 ( 
.A(n_194),
.B(n_176),
.Y(n_236)
);

OAI22xp33_ASAP7_75t_L g237 ( 
.A1(n_197),
.A2(n_167),
.B1(n_168),
.B2(n_132),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_211),
.B(n_181),
.Y(n_238)
);

O2A1O1Ixp5_ASAP7_75t_L g239 ( 
.A1(n_201),
.A2(n_142),
.B(n_165),
.C(n_152),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_213),
.B(n_121),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_202),
.A2(n_145),
.B1(n_127),
.B2(n_169),
.Y(n_241)
);

OAI22xp33_ASAP7_75t_L g242 ( 
.A1(n_204),
.A2(n_149),
.B1(n_128),
.B2(n_129),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_205),
.B(n_131),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_199),
.Y(n_244)
);

BUFx5_ASAP7_75t_L g245 ( 
.A(n_206),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_200),
.B(n_141),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_209),
.B(n_144),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_219),
.B(n_146),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_228),
.A2(n_173),
.B(n_209),
.Y(n_249)
);

AND2x2_ASAP7_75t_L g250 ( 
.A(n_226),
.B(n_153),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_221),
.A2(n_164),
.B1(n_157),
.B2(n_159),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_230),
.A2(n_151),
.B1(n_117),
.B2(n_166),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_233),
.B(n_222),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_231),
.A2(n_218),
.B1(n_236),
.B2(n_234),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_223),
.B(n_139),
.Y(n_255)
);

O2A1O1Ixp33_ASAP7_75t_L g256 ( 
.A1(n_237),
.A2(n_232),
.B(n_239),
.C(n_242),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_245),
.B(n_139),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_224),
.B(n_3),
.Y(n_258)
);

INVx3_ASAP7_75t_L g259 ( 
.A(n_227),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_241),
.A2(n_189),
.B1(n_62),
.B2(n_64),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_233),
.B(n_3),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_240),
.A2(n_53),
.B(n_102),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_245),
.B(n_52),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_L g264 ( 
.A1(n_245),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_220),
.B(n_8),
.Y(n_265)
);

AND2x4_ASAP7_75t_L g266 ( 
.A(n_225),
.B(n_9),
.Y(n_266)
);

OAI21xp33_ASAP7_75t_L g267 ( 
.A1(n_246),
.A2(n_12),
.B(n_13),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_238),
.A2(n_17),
.B(n_19),
.Y(n_268)
);

OR2x6_ASAP7_75t_L g269 ( 
.A(n_229),
.B(n_20),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_245),
.B(n_21),
.Y(n_270)
);

NAND3xp33_ASAP7_75t_SL g271 ( 
.A(n_243),
.B(n_22),
.C(n_24),
.Y(n_271)
);

O2A1O1Ixp33_ASAP7_75t_L g272 ( 
.A1(n_247),
.A2(n_25),
.B(n_26),
.C(n_27),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_244),
.A2(n_30),
.B(n_36),
.Y(n_273)
);

INVx6_ASAP7_75t_L g274 ( 
.A(n_235),
.Y(n_274)
);

INVx3_ASAP7_75t_L g275 ( 
.A(n_259),
.Y(n_275)
);

INVx2_ASAP7_75t_SL g276 ( 
.A(n_250),
.Y(n_276)
);

INVxp67_ASAP7_75t_SL g277 ( 
.A(n_254),
.Y(n_277)
);

INVx5_ASAP7_75t_L g278 ( 
.A(n_274),
.Y(n_278)
);

OAI21x1_ASAP7_75t_L g279 ( 
.A1(n_249),
.A2(n_270),
.B(n_263),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_261),
.Y(n_280)
);

AOI21x1_ASAP7_75t_L g281 ( 
.A1(n_257),
.A2(n_235),
.B(n_38),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_248),
.B(n_37),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_253),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_255),
.A2(n_42),
.B(n_46),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_251),
.Y(n_285)
);

INVx3_ASAP7_75t_L g286 ( 
.A(n_274),
.Y(n_286)
);

OAI21x1_ASAP7_75t_L g287 ( 
.A1(n_260),
.A2(n_109),
.B(n_65),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_L g288 ( 
.A1(n_256),
.A2(n_49),
.B(n_66),
.Y(n_288)
);

AND2x4_ASAP7_75t_L g289 ( 
.A(n_266),
.B(n_67),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_252),
.Y(n_290)
);

A2O1A1Ixp33_ASAP7_75t_L g291 ( 
.A1(n_258),
.A2(n_69),
.B(n_71),
.C(n_73),
.Y(n_291)
);

NAND3xp33_ASAP7_75t_SL g292 ( 
.A(n_265),
.B(n_76),
.C(n_78),
.Y(n_292)
);

AND2x6_ASAP7_75t_L g293 ( 
.A(n_271),
.B(n_81),
.Y(n_293)
);

BUFx2_ASAP7_75t_L g294 ( 
.A(n_277),
.Y(n_294)
);

INVx3_ASAP7_75t_L g295 ( 
.A(n_281),
.Y(n_295)
);

OA21x2_ASAP7_75t_L g296 ( 
.A1(n_288),
.A2(n_267),
.B(n_262),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_283),
.A2(n_264),
.B1(n_269),
.B2(n_272),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_276),
.Y(n_298)
);

OAI21x1_ASAP7_75t_L g299 ( 
.A1(n_279),
.A2(n_273),
.B(n_268),
.Y(n_299)
);

INVx1_ASAP7_75t_SL g300 ( 
.A(n_275),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_282),
.A2(n_269),
.B(n_83),
.Y(n_301)
);

AOI21xp33_ASAP7_75t_L g302 ( 
.A1(n_290),
.A2(n_82),
.B(n_86),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_280),
.B(n_87),
.Y(n_303)
);

NOR2x1_ASAP7_75t_SL g304 ( 
.A(n_292),
.B(n_101),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_275),
.Y(n_305)
);

AO21x2_ASAP7_75t_L g306 ( 
.A1(n_287),
.A2(n_88),
.B(n_89),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_294),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_294),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_295),
.Y(n_309)
);

BUFx3_ASAP7_75t_L g310 ( 
.A(n_300),
.Y(n_310)
);

AND2x2_ASAP7_75t_L g311 ( 
.A(n_298),
.B(n_289),
.Y(n_311)
);

BUFx6f_ASAP7_75t_L g312 ( 
.A(n_305),
.Y(n_312)
);

OR2x2_ASAP7_75t_L g313 ( 
.A(n_303),
.B(n_285),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_295),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_297),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_309),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_309),
.Y(n_317)
);

INVx8_ASAP7_75t_L g318 ( 
.A(n_311),
.Y(n_318)
);

AND2x2_ASAP7_75t_L g319 ( 
.A(n_307),
.B(n_289),
.Y(n_319)
);

AND2x2_ASAP7_75t_L g320 ( 
.A(n_308),
.B(n_313),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_314),
.Y(n_321)
);

OR2x2_ASAP7_75t_L g322 ( 
.A(n_310),
.B(n_301),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_312),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_312),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_314),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_315),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_312),
.Y(n_327)
);

INVx2_ASAP7_75t_SL g328 ( 
.A(n_327),
.Y(n_328)
);

HB1xp67_ASAP7_75t_L g329 ( 
.A(n_326),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_326),
.Y(n_330)
);

AND2x2_ASAP7_75t_L g331 ( 
.A(n_320),
.B(n_310),
.Y(n_331)
);

AND2x4_ASAP7_75t_L g332 ( 
.A(n_327),
.B(n_312),
.Y(n_332)
);

INVx3_ASAP7_75t_L g333 ( 
.A(n_316),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_L g334 ( 
.A1(n_322),
.A2(n_296),
.B(n_302),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_317),
.Y(n_335)
);

BUFx2_ASAP7_75t_L g336 ( 
.A(n_318),
.Y(n_336)
);

OR2x2_ASAP7_75t_SL g337 ( 
.A(n_323),
.B(n_296),
.Y(n_337)
);

AND2x2_ASAP7_75t_L g338 ( 
.A(n_319),
.B(n_304),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_318),
.B(n_293),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_335),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_333),
.Y(n_341)
);

INVx3_ASAP7_75t_L g342 ( 
.A(n_331),
.Y(n_342)
);

OR2x2_ASAP7_75t_L g343 ( 
.A(n_337),
.B(n_324),
.Y(n_343)
);

AND2x2_ASAP7_75t_L g344 ( 
.A(n_328),
.B(n_325),
.Y(n_344)
);

OR2x2_ASAP7_75t_L g345 ( 
.A(n_329),
.B(n_321),
.Y(n_345)
);

NAND2x1_ASAP7_75t_L g346 ( 
.A(n_341),
.B(n_330),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_342),
.B(n_338),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_340),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_348),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_346),
.Y(n_350)
);

AOI221xp5_ASAP7_75t_L g351 ( 
.A1(n_349),
.A2(n_347),
.B1(n_343),
.B2(n_334),
.C(n_344),
.Y(n_351)
);

A2O1A1Ixp33_ASAP7_75t_L g352 ( 
.A1(n_350),
.A2(n_343),
.B(n_291),
.C(n_336),
.Y(n_352)
);

OAI22xp33_ASAP7_75t_L g353 ( 
.A1(n_351),
.A2(n_345),
.B1(n_339),
.B2(n_328),
.Y(n_353)
);

A2O1A1Ixp33_ASAP7_75t_L g354 ( 
.A1(n_352),
.A2(n_284),
.B(n_332),
.C(n_329),
.Y(n_354)
);

NOR3xp33_ASAP7_75t_L g355 ( 
.A(n_354),
.B(n_332),
.C(n_333),
.Y(n_355)
);

NOR2x1_ASAP7_75t_L g356 ( 
.A(n_353),
.B(n_332),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_356),
.B(n_333),
.Y(n_357)
);

NOR2xp67_ASAP7_75t_L g358 ( 
.A(n_357),
.B(n_355),
.Y(n_358)
);

AND2x2_ASAP7_75t_L g359 ( 
.A(n_358),
.B(n_278),
.Y(n_359)
);

XNOR2x1_ASAP7_75t_L g360 ( 
.A(n_359),
.B(n_286),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_359),
.Y(n_361)
);

OAI31xp33_ASAP7_75t_L g362 ( 
.A1(n_361),
.A2(n_293),
.A3(n_295),
.B(n_278),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_360),
.B(n_91),
.Y(n_363)
);

AOI22xp33_ASAP7_75t_L g364 ( 
.A1(n_363),
.A2(n_293),
.B1(n_306),
.B2(n_296),
.Y(n_364)
);

NAND3xp33_ASAP7_75t_L g365 ( 
.A(n_362),
.B(n_278),
.C(n_96),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_365),
.B(n_95),
.Y(n_366)
);

AND2x2_ASAP7_75t_L g367 ( 
.A(n_364),
.B(n_97),
.Y(n_367)
);

NAND2xp33_ASAP7_75t_L g368 ( 
.A(n_366),
.B(n_293),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_368),
.B(n_367),
.Y(n_369)
);

AOI22xp33_ASAP7_75t_L g370 ( 
.A1(n_369),
.A2(n_306),
.B1(n_299),
.B2(n_99),
.Y(n_370)
);


endmodule