module fake_jpeg_13650_n_68 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_68);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_68;

wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_51;
wire n_47;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_44;
wire n_26;
wire n_38;
wire n_36;
wire n_62;
wire n_25;
wire n_31;
wire n_56;
wire n_67;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;
wire n_66;

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_4),
.Y(n_23)
);

INVx11_ASAP7_75t_SL g24 ( 
.A(n_6),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_14),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_25),
.Y(n_28)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_21),
.B(n_26),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_30),
.B(n_31),
.Y(n_40)
);

INVx1_ASAP7_75t_SL g31 ( 
.A(n_22),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_27),
.B(n_0),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_32),
.B(n_35),
.Y(n_42)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_33),
.B(n_36),
.Y(n_38)
);

INVx6_ASAP7_75t_SL g34 ( 
.A(n_24),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_23),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

INVx1_ASAP7_75t_SL g50 ( 
.A(n_37),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_44),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_42),
.B(n_38),
.C(n_43),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_46),
.B(n_51),
.C(n_2),
.Y(n_56)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_48),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_40),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_49),
.B(n_52),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_11),
.C(n_17),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_42),
.B(n_1),
.Y(n_52)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_47),
.Y(n_55)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_55),
.Y(n_59)
);

XOR2xp5_ASAP7_75t_L g61 ( 
.A(n_56),
.B(n_58),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_50),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_57)
);

CKINVDCx14_ASAP7_75t_R g60 ( 
.A(n_57),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_45),
.B(n_10),
.Y(n_58)
);

OAI21xp5_ASAP7_75t_L g62 ( 
.A1(n_60),
.A2(n_53),
.B(n_54),
.Y(n_62)
);

BUFx24_ASAP7_75t_SL g63 ( 
.A(n_62),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_63),
.B(n_59),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_64),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_65),
.Y(n_66)
);

HB1xp67_ASAP7_75t_L g67 ( 
.A(n_66),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_67),
.B(n_61),
.Y(n_68)
);


endmodule