module real_jpeg_24848_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_312;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_0),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_2),
.A2(n_56),
.B1(n_71),
.B2(n_72),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_2),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_2),
.A2(n_40),
.B1(n_41),
.B2(n_71),
.Y(n_153)
);

OAI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_2),
.A2(n_63),
.B1(n_66),
.B2(n_71),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_2),
.A2(n_27),
.B1(n_28),
.B2(n_71),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_4),
.A2(n_27),
.B1(n_28),
.B2(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_4),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_4),
.A2(n_35),
.B1(n_40),
.B2(n_41),
.Y(n_89)
);

INVx8_ASAP7_75t_SL g65 ( 
.A(n_5),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_6),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_6),
.B(n_62),
.Y(n_176)
);

O2A1O1Ixp33_ASAP7_75t_L g218 ( 
.A1(n_6),
.A2(n_66),
.B(n_80),
.C(n_219),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_L g231 ( 
.A1(n_6),
.A2(n_63),
.B1(n_66),
.B2(n_157),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_6),
.B(n_28),
.C(n_44),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_L g242 ( 
.A1(n_6),
.A2(n_40),
.B1(n_41),
.B2(n_157),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_6),
.A2(n_25),
.B(n_253),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_6),
.B(n_123),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_7),
.A2(n_56),
.B1(n_59),
.B2(n_60),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_7),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_7),
.A2(n_60),
.B1(n_63),
.B2(n_66),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_7),
.A2(n_40),
.B1(n_41),
.B2(n_60),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_L g178 ( 
.A1(n_7),
.A2(n_27),
.B1(n_28),
.B2(n_60),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_8),
.A2(n_63),
.B1(n_66),
.B2(n_147),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_8),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_8),
.A2(n_58),
.B1(n_59),
.B2(n_147),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_L g228 ( 
.A1(n_8),
.A2(n_40),
.B1(n_41),
.B2(n_147),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_8),
.A2(n_27),
.B1(n_28),
.B2(n_147),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_9),
.A2(n_40),
.B1(n_41),
.B2(n_49),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_9),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_9),
.A2(n_27),
.B1(n_28),
.B2(n_49),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_9),
.A2(n_49),
.B1(n_63),
.B2(n_66),
.Y(n_125)
);

BUFx5_ASAP7_75t_L g80 ( 
.A(n_10),
.Y(n_80)
);

INVx13_ASAP7_75t_L g58 ( 
.A(n_11),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_12),
.A2(n_63),
.B1(n_66),
.B2(n_84),
.Y(n_83)
);

CKINVDCx14_ASAP7_75t_R g84 ( 
.A(n_12),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_12),
.A2(n_40),
.B1(n_41),
.B2(n_84),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_12),
.A2(n_59),
.B1(n_84),
.B2(n_132),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_12),
.A2(n_27),
.B1(n_28),
.B2(n_84),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_13),
.A2(n_59),
.B1(n_107),
.B2(n_108),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_13),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_13),
.A2(n_63),
.B1(n_66),
.B2(n_107),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_13),
.A2(n_40),
.B1(n_41),
.B2(n_107),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_L g247 ( 
.A1(n_13),
.A2(n_27),
.B1(n_28),
.B2(n_107),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_14),
.A2(n_39),
.B1(n_40),
.B2(n_41),
.Y(n_38)
);

CKINVDCx16_ASAP7_75t_R g39 ( 
.A(n_14),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_14),
.A2(n_39),
.B1(n_63),
.B2(n_66),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_14),
.A2(n_27),
.B1(n_28),
.B2(n_39),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_16),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_16),
.A2(n_26),
.B1(n_163),
.B2(n_165),
.Y(n_162)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_16),
.Y(n_179)
);

INVx6_ASAP7_75t_L g196 ( 
.A(n_16),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_16),
.A2(n_26),
.B1(n_244),
.B2(n_246),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_136),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_134),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_112),
.Y(n_20)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_21),
.B(n_112),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_75),
.C(n_91),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_22),
.A2(n_75),
.B1(n_76),
.B2(n_314),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_22),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_51),
.Y(n_22)
);

AOI21xp33_ASAP7_75t_L g113 ( 
.A1(n_23),
.A2(n_24),
.B(n_53),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_36),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_24),
.A2(n_52),
.B1(n_53),
.B2(n_54),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_24),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_24),
.A2(n_36),
.B1(n_37),
.B2(n_52),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_32),
.B(n_34),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_25),
.A2(n_34),
.B1(n_96),
.B2(n_97),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_25),
.A2(n_164),
.B1(n_178),
.B2(n_179),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_25),
.A2(n_96),
.B1(n_193),
.B2(n_194),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_25),
.A2(n_247),
.B(n_253),
.Y(n_267)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_26),
.B(n_222),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_30),
.Y(n_26)
);

OA22x2_ASAP7_75t_L g47 ( 
.A1(n_27),
.A2(n_28),
.B1(n_44),
.B2(n_46),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_27),
.B(n_251),
.Y(n_250)
);

INVx6_ASAP7_75t_SL g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_31),
.Y(n_33)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_37),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_42),
.B1(n_48),
.B2(n_50),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_38),
.A2(n_42),
.B1(n_50),
.B2(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_SL g41 ( 
.A(n_40),
.Y(n_41)
);

OAI22xp33_ASAP7_75t_L g43 ( 
.A1(n_40),
.A2(n_41),
.B1(n_44),
.B2(n_46),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_40),
.A2(n_41),
.B1(n_80),
.B2(n_81),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_40),
.B(n_239),
.Y(n_238)
);

OAI21xp33_ASAP7_75t_L g219 ( 
.A1(n_41),
.A2(n_81),
.B(n_157),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_42),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_42),
.A2(n_50),
.B(n_128),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_42),
.B(n_153),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_42),
.A2(n_50),
.B1(n_214),
.B2(n_227),
.Y(n_226)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_47),
.Y(n_42)
);

INVx13_ASAP7_75t_L g46 ( 
.A(n_44),
.Y(n_46)
);

BUFx24_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_47),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_47),
.A2(n_87),
.B1(n_88),
.B2(n_89),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_47),
.A2(n_151),
.B(n_152),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_47),
.A2(n_87),
.B1(n_101),
.B2(n_151),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_47),
.B(n_157),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_L g266 ( 
.A1(n_47),
.A2(n_152),
.B(n_228),
.Y(n_266)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_48),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_50),
.B(n_153),
.Y(n_215)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_61),
.B(n_68),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_55),
.A2(n_61),
.B1(n_109),
.B2(n_131),
.Y(n_130)
);

INVx8_ASAP7_75t_L g156 ( 
.A(n_56),
.Y(n_156)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

OAI22xp33_ASAP7_75t_L g74 ( 
.A1(n_57),
.A2(n_58),
.B1(n_65),
.B2(n_67),
.Y(n_74)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_58),
.Y(n_59)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_58),
.Y(n_72)
);

INVx8_ASAP7_75t_L g169 ( 
.A(n_58),
.Y(n_169)
);

INVx11_ASAP7_75t_L g132 ( 
.A(n_59),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_61),
.B(n_74),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_61),
.B(n_70),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_61),
.A2(n_68),
.B(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_62),
.A2(n_73),
.B1(n_106),
.B2(n_188),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_63),
.A2(n_65),
.B1(n_66),
.B2(n_67),
.Y(n_62)
);

INVx5_ASAP7_75t_SL g66 ( 
.A(n_63),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_63),
.A2(n_66),
.B1(n_80),
.B2(n_81),
.Y(n_82)
);

A2O1A1Ixp33_ASAP7_75t_L g167 ( 
.A1(n_63),
.A2(n_67),
.B(n_158),
.C(n_168),
.Y(n_167)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_65),
.Y(n_67)
);

NAND3xp33_ASAP7_75t_SL g168 ( 
.A(n_65),
.B(n_66),
.C(n_169),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_73),
.Y(n_68)
);

CKINVDCx14_ASAP7_75t_R g69 ( 
.A(n_70),
.Y(n_69)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_72),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_72),
.B(n_157),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_73),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_73),
.A2(n_111),
.B(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_86),
.B(n_90),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_77),
.B(n_86),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_78),
.A2(n_79),
.B1(n_83),
.B2(n_85),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_78),
.A2(n_79),
.B1(n_83),
.B2(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_78),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_78),
.A2(n_184),
.B(n_185),
.Y(n_183)
);

OAI21xp33_ASAP7_75t_L g230 ( 
.A1(n_78),
.A2(n_185),
.B(n_231),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_82),
.Y(n_78)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_79),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_79),
.A2(n_172),
.B(n_173),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g297 ( 
.A1(n_79),
.A2(n_103),
.B(n_173),
.Y(n_297)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_80),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_85),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_87),
.A2(n_213),
.B(n_215),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_87),
.A2(n_215),
.B(n_242),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_89),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_90),
.A2(n_115),
.B1(n_116),
.B2(n_117),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_90),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_91),
.A2(n_92),
.B1(n_313),
.B2(n_315),
.Y(n_312)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_102),
.C(n_104),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_93),
.A2(n_94),
.B1(n_307),
.B2(n_308),
.Y(n_306)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_98),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_95),
.A2(n_98),
.B1(n_99),
.B2(n_290),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_95),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_97),
.B(n_157),
.Y(n_251)
);

INVx3_ASAP7_75t_L g254 ( 
.A(n_97),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g256 ( 
.A1(n_97),
.A2(n_221),
.B(n_245),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_99),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_SL g308 ( 
.A(n_102),
.B(n_104),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_109),
.B(n_110),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_114),
.Y(n_112)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_118),
.A2(n_119),
.B1(n_130),
.B2(n_133),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_120),
.A2(n_126),
.B1(n_127),
.B2(n_129),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_120),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_122),
.B1(n_123),
.B2(n_124),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_122),
.A2(n_123),
.B1(n_146),
.B2(n_148),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_122),
.B(n_174),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_123),
.B(n_174),
.Y(n_185)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_130),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_135),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_137),
.A2(n_311),
.B(n_317),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_138),
.A2(n_301),
.B(n_310),
.Y(n_137)
);

O2A1O1Ixp33_ASAP7_75t_SL g138 ( 
.A1(n_139),
.A2(n_200),
.B(n_284),
.C(n_300),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_180),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_140),
.B(n_180),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_159),
.C(n_170),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_141),
.A2(n_142),
.B1(n_279),
.B2(n_280),
.Y(n_278)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_154),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_145),
.B1(n_149),
.B2(n_150),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_145),
.B(n_149),
.C(n_154),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_146),
.Y(n_172)
);

CKINVDCx14_ASAP7_75t_R g184 ( 
.A(n_148),
.Y(n_184)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

OAI21xp33_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_157),
.B(n_158),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_159),
.A2(n_160),
.B1(n_170),
.B2(n_281),
.Y(n_280)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_161),
.A2(n_162),
.B1(n_166),
.B2(n_167),
.Y(n_160)
);

CKINVDCx14_ASAP7_75t_R g161 ( 
.A(n_162),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_162),
.B(n_166),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_165),
.Y(n_193)
);

CKINVDCx14_ASAP7_75t_R g166 ( 
.A(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_170),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_175),
.C(n_177),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_171),
.B(n_208),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_175),
.A2(n_176),
.B1(n_177),
.B2(n_209),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_177),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_178),
.A2(n_179),
.B(n_221),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_181),
.A2(n_189),
.B1(n_190),
.B2(n_199),
.Y(n_180)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_181),
.Y(n_199)
);

BUFx24_ASAP7_75t_SL g319 ( 
.A(n_181),
.Y(n_319)
);

FAx1_ASAP7_75t_SL g181 ( 
.A(n_182),
.B(n_183),
.CI(n_186),
.CON(n_181),
.SN(n_181)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_182),
.B(n_183),
.C(n_186),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_SL g190 ( 
.A(n_191),
.B(n_198),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_191),
.B(n_198),
.C(n_199),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_197),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_192),
.B(n_197),
.Y(n_298)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_202),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_203),
.A2(n_277),
.B(n_283),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_204),
.A2(n_232),
.B(n_276),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_205),
.B(n_224),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_205),
.B(n_224),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_206),
.A2(n_207),
.B1(n_210),
.B2(n_223),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_206),
.B(n_212),
.C(n_216),
.Y(n_282)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_210),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_211),
.A2(n_212),
.B1(n_216),
.B2(n_217),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_214),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_217),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_220),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_SL g225 ( 
.A(n_218),
.B(n_220),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_222),
.B(n_254),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_226),
.C(n_229),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_225),
.B(n_272),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_226),
.A2(n_229),
.B1(n_230),
.B2(n_273),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_226),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_233),
.A2(n_270),
.B(n_275),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_234),
.A2(n_260),
.B(n_269),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_235),
.A2(n_248),
.B(n_259),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_236),
.B(n_243),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_236),
.B(n_243),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_237),
.A2(n_238),
.B1(n_240),
.B2(n_241),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_238),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_238),
.B(n_240),
.Y(n_268)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

CKINVDCx16_ASAP7_75t_R g244 ( 
.A(n_245),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_249),
.A2(n_255),
.B(n_258),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_252),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_256),
.B(n_257),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_256),
.B(n_257),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_261),
.B(n_268),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_261),
.B(n_268),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_267),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_263),
.A2(n_264),
.B1(n_265),
.B2(n_266),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_263),
.B(n_266),
.C(n_267),
.Y(n_274)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_271),
.B(n_274),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_271),
.B(n_274),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_278),
.B(n_282),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_278),
.B(n_282),
.Y(n_283)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_285),
.B(n_299),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_285),
.B(n_299),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_287),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_286),
.B(n_289),
.C(n_291),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_288),
.A2(n_289),
.B1(n_291),
.B2(n_292),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_298),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_294),
.A2(n_295),
.B1(n_296),
.B2(n_297),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_295),
.B(n_296),
.C(n_298),
.Y(n_309)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_303),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_302),
.B(n_303),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_309),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_306),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_305),
.B(n_306),
.C(n_309),
.Y(n_316)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_312),
.B(n_316),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_312),
.B(n_316),
.Y(n_317)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_313),
.Y(n_315)
);


endmodule