module fake_jpeg_9326_n_283 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_283);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_283;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_282;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_8),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_11),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_7),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_8),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_41),
.Y(n_44)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

BUFx24_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

CKINVDCx14_ASAP7_75t_R g53 ( 
.A(n_39),
.Y(n_53)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_40),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_26),
.B(n_15),
.Y(n_41)
);

AOI21xp33_ASAP7_75t_L g42 ( 
.A1(n_19),
.A2(n_1),
.B(n_2),
.Y(n_42)
);

A2O1A1Ixp33_ASAP7_75t_L g52 ( 
.A1(n_42),
.A2(n_19),
.B(n_25),
.C(n_31),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_L g43 ( 
.A1(n_40),
.A2(n_24),
.B1(n_30),
.B2(n_21),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_43),
.A2(n_16),
.B1(n_21),
.B2(n_30),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_41),
.B(n_24),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_45),
.B(n_58),
.Y(n_65)
);

INVx13_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_48),
.B(n_50),
.Y(n_68)
);

OAI21xp33_ASAP7_75t_L g49 ( 
.A1(n_42),
.A2(n_12),
.B(n_10),
.Y(n_49)
);

CKINVDCx14_ASAP7_75t_R g82 ( 
.A(n_49),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_33),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_52),
.B(n_54),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_36),
.B(n_33),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_35),
.B(n_22),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_55),
.B(n_56),
.Y(n_86)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_40),
.Y(n_58)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_60),
.Y(n_78)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_61),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_35),
.B(n_33),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_62),
.B(n_64),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_34),
.B(n_24),
.Y(n_64)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

BUFx2_ASAP7_75t_SL g115 ( 
.A(n_67),
.Y(n_115)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_69),
.B(n_71),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_48),
.A2(n_27),
.B1(n_22),
.B2(n_32),
.Y(n_70)
);

OAI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_70),
.A2(n_72),
.B1(n_77),
.B2(n_19),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_64),
.Y(n_71)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_74),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_52),
.B(n_22),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_76),
.A2(n_65),
.B(n_75),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_59),
.A2(n_27),
.B1(n_32),
.B2(n_31),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_50),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_80),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_54),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_81),
.Y(n_113)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_46),
.Y(n_83)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_83),
.Y(n_103)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_60),
.Y(n_84)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_84),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_52),
.A2(n_40),
.B1(n_35),
.B2(n_27),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_85),
.A2(n_88),
.B1(n_29),
.B2(n_25),
.Y(n_108)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_57),
.Y(n_87)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_87),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_43),
.A2(n_16),
.B1(n_21),
.B2(n_30),
.Y(n_88)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_57),
.Y(n_89)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_89),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g90 ( 
.A1(n_44),
.A2(n_16),
.B(n_39),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g99 ( 
.A(n_90),
.B(n_53),
.Y(n_99)
);

AOI32xp33_ASAP7_75t_L g91 ( 
.A1(n_73),
.A2(n_44),
.A3(n_62),
.B1(n_55),
.B2(n_63),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_91),
.A2(n_78),
.B(n_23),
.Y(n_129)
);

A2O1A1Ixp33_ASAP7_75t_L g92 ( 
.A1(n_73),
.A2(n_45),
.B(n_53),
.C(n_31),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_92),
.B(n_104),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_82),
.A2(n_51),
.B1(n_58),
.B2(n_61),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_93),
.A2(n_97),
.B1(n_100),
.B2(n_105),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_71),
.B(n_51),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_95),
.B(n_98),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_82),
.A2(n_61),
.B1(n_63),
.B2(n_59),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_75),
.B(n_37),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_99),
.B(n_106),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_85),
.A2(n_56),
.B1(n_59),
.B2(n_63),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_102),
.B(n_17),
.Y(n_133)
);

A2O1A1Ixp33_ASAP7_75t_L g104 ( 
.A1(n_76),
.A2(n_25),
.B(n_26),
.C(n_29),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_76),
.A2(n_34),
.B1(n_37),
.B2(n_28),
.Y(n_105)
);

A2O1A1Ixp33_ASAP7_75t_L g107 ( 
.A1(n_65),
.A2(n_32),
.B(n_29),
.C(n_26),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_107),
.B(n_114),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_108),
.A2(n_89),
.B1(n_87),
.B2(n_78),
.Y(n_132)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_86),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_112),
.B(n_116),
.Y(n_119)
);

A2O1A1Ixp33_ASAP7_75t_L g114 ( 
.A1(n_68),
.A2(n_90),
.B(n_86),
.C(n_88),
.Y(n_114)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_72),
.Y(n_116)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_94),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_121),
.B(n_125),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_99),
.B(n_68),
.C(n_79),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_122),
.B(n_123),
.C(n_109),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_106),
.B(n_37),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_115),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_116),
.A2(n_67),
.B1(n_69),
.B2(n_84),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_126),
.A2(n_133),
.B1(n_111),
.B2(n_66),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_98),
.B(n_79),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_127),
.B(n_135),
.Y(n_152)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_94),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_128),
.B(n_132),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_129),
.A2(n_137),
.B(n_139),
.Y(n_144)
);

INVx2_ASAP7_75t_SL g131 ( 
.A(n_115),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_131),
.B(n_141),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_108),
.A2(n_83),
.B1(n_74),
.B2(n_66),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_134),
.A2(n_113),
.B1(n_96),
.B2(n_111),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_95),
.B(n_112),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_114),
.B(n_57),
.Y(n_136)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_136),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_91),
.A2(n_20),
.B(n_23),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_103),
.B(n_66),
.Y(n_138)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_138),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_92),
.A2(n_20),
.B(n_23),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_105),
.B(n_39),
.Y(n_140)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_140),
.Y(n_149)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_93),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_100),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_142),
.B(n_143),
.Y(n_170)
);

INVx5_ASAP7_75t_L g143 ( 
.A(n_101),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_130),
.B(n_104),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_145),
.B(n_150),
.C(n_156),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_138),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_148),
.B(n_154),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_151),
.A2(n_158),
.B1(n_159),
.B2(n_160),
.Y(n_181)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_119),
.Y(n_154)
);

AO22x1_ASAP7_75t_L g155 ( 
.A1(n_141),
.A2(n_142),
.B1(n_136),
.B2(n_117),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_155),
.B(n_158),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_130),
.B(n_104),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_123),
.B(n_107),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_157),
.B(n_164),
.C(n_118),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_126),
.Y(n_158)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_119),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_161),
.B(n_162),
.Y(n_178)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_135),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_163),
.A2(n_166),
.B1(n_132),
.B2(n_149),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_122),
.B(n_39),
.Y(n_164)
);

OAI22xp33_ASAP7_75t_L g165 ( 
.A1(n_121),
.A2(n_110),
.B1(n_109),
.B2(n_103),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_165),
.A2(n_166),
.B1(n_171),
.B2(n_134),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_133),
.A2(n_110),
.B1(n_101),
.B2(n_28),
.Y(n_166)
);

INVx13_ASAP7_75t_L g167 ( 
.A(n_131),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_167),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_128),
.B(n_10),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_168),
.B(n_169),
.Y(n_188)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_127),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_140),
.A2(n_28),
.B1(n_17),
.B2(n_20),
.Y(n_171)
);

BUFx24_ASAP7_75t_SL g174 ( 
.A(n_145),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_174),
.B(n_175),
.Y(n_207)
);

HB1xp67_ASAP7_75t_L g175 ( 
.A(n_167),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g213 ( 
.A(n_177),
.Y(n_213)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_153),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_179),
.B(n_180),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_170),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_181),
.A2(n_189),
.B1(n_191),
.B2(n_196),
.Y(n_199)
);

A2O1A1O1Ixp25_ASAP7_75t_L g182 ( 
.A1(n_144),
.A2(n_137),
.B(n_129),
.C(n_139),
.D(n_120),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_182),
.B(n_144),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_148),
.Y(n_183)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_183),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_184),
.B(n_186),
.C(n_156),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_165),
.Y(n_185)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_185),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_150),
.B(n_164),
.Y(n_186)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_187),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_146),
.A2(n_120),
.B1(n_117),
.B2(n_125),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_152),
.B(n_118),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_190),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_155),
.A2(n_124),
.B1(n_131),
.B2(n_143),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_152),
.B(n_124),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_192),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_157),
.B(n_143),
.Y(n_193)
);

FAx1_ASAP7_75t_SL g202 ( 
.A(n_193),
.B(n_171),
.CI(n_23),
.CON(n_202),
.SN(n_202)
);

NOR2x1_ASAP7_75t_L g194 ( 
.A(n_151),
.B(n_20),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g215 ( 
.A(n_194),
.B(n_8),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_155),
.A2(n_17),
.B1(n_23),
.B2(n_39),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_SL g220 ( 
.A(n_197),
.B(n_202),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_200),
.B(n_209),
.C(n_210),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_172),
.A2(n_147),
.B(n_163),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_201),
.A2(n_199),
.B(n_208),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_186),
.B(n_39),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_203),
.B(n_206),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_176),
.B(n_23),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_172),
.A2(n_17),
.B1(n_2),
.B2(n_3),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_208),
.A2(n_218),
.B1(n_177),
.B2(n_188),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_176),
.B(n_1),
.C(n_2),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_193),
.B(n_7),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_184),
.B(n_1),
.C(n_3),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_214),
.B(n_217),
.Y(n_223)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_215),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_191),
.B(n_7),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_181),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_213),
.A2(n_189),
.B1(n_196),
.B2(n_194),
.Y(n_222)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_222),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_212),
.A2(n_190),
.B1(n_180),
.B2(n_195),
.Y(n_224)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_224),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_225),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_199),
.A2(n_182),
.B1(n_178),
.B2(n_173),
.Y(n_226)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_226),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_216),
.Y(n_227)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_227),
.Y(n_240)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_201),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_228),
.B(n_231),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g244 ( 
.A1(n_229),
.A2(n_215),
.B(n_214),
.Y(n_244)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_217),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_211),
.A2(n_173),
.B1(n_183),
.B2(n_11),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_232),
.A2(n_209),
.B1(n_11),
.B2(n_13),
.Y(n_246)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_218),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_233),
.B(n_234),
.Y(n_247)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_205),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_210),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_235),
.A2(n_204),
.B1(n_198),
.B2(n_202),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_237),
.A2(n_244),
.B1(n_248),
.B2(n_14),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_226),
.A2(n_197),
.B1(n_200),
.B2(n_202),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_243),
.A2(n_220),
.B1(n_227),
.B2(n_219),
.Y(n_251)
);

A2O1A1Ixp33_ASAP7_75t_SL g245 ( 
.A1(n_222),
.A2(n_215),
.B(n_203),
.C(n_206),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_SL g249 ( 
.A1(n_245),
.A2(n_220),
.B1(n_224),
.B2(n_225),
.Y(n_249)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_246),
.Y(n_256)
);

AOI21xp33_ASAP7_75t_L g248 ( 
.A1(n_221),
.A2(n_207),
.B(n_9),
.Y(n_248)
);

XNOR2x1_ASAP7_75t_L g266 ( 
.A(n_249),
.B(n_245),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_240),
.B(n_230),
.C(n_219),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_250),
.B(n_252),
.C(n_253),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_251),
.B(n_237),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_240),
.B(n_230),
.C(n_223),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_243),
.B(n_223),
.C(n_9),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_239),
.B(n_9),
.C(n_13),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_254),
.B(n_14),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_238),
.A2(n_14),
.B1(n_4),
.B2(n_5),
.Y(n_255)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_255),
.Y(n_262)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_257),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_247),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_L g260 ( 
.A1(n_258),
.A2(n_259),
.B(n_236),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_L g259 ( 
.A1(n_242),
.A2(n_241),
.B(n_244),
.Y(n_259)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_260),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_261),
.B(n_265),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_263),
.B(n_245),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_254),
.B(n_3),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_266),
.A2(n_258),
.B(n_253),
.Y(n_271)
);

BUFx2_ASAP7_75t_L g269 ( 
.A(n_266),
.Y(n_269)
);

OR2x2_ASAP7_75t_L g275 ( 
.A(n_269),
.B(n_273),
.Y(n_275)
);

AO21x1_ASAP7_75t_L g276 ( 
.A1(n_271),
.A2(n_272),
.B(n_267),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_L g272 ( 
.A1(n_267),
.A2(n_252),
.B(n_250),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_270),
.A2(n_269),
.B1(n_264),
.B2(n_256),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_274),
.A2(n_276),
.B(n_277),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_268),
.A2(n_262),
.B(n_245),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_275),
.A2(n_4),
.B(n_6),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_SL g280 ( 
.A1(n_279),
.A2(n_4),
.B(n_6),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_280),
.A2(n_278),
.B(n_6),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_281),
.B(n_6),
.Y(n_282)
);

HB1xp67_ASAP7_75t_L g283 ( 
.A(n_282),
.Y(n_283)
);


endmodule