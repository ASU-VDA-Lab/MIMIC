module fake_jpeg_194_n_714 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_714);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_714;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_696;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_686;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_678;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_699;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_713;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_701;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_672;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_688;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_689;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_704;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_698;
wire n_195;
wire n_450;
wire n_557;
wire n_681;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_694;
wire n_692;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_668;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_682;
wire n_305;
wire n_161;
wire n_441;
wire n_697;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_710;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_679;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_691;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_676;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_709;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_670;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_708;
wire n_467;
wire n_683;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_690;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_693;
wire n_674;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_703;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_684;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_680;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_695;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_702;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_687;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_707;
wire n_232;
wire n_527;
wire n_482;
wire n_673;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_705;
wire n_665;
wire n_706;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_677;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_700;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_671;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_669;
wire n_524;
wire n_402;
wire n_563;
wire n_685;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_712;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_711;
wire n_462;
wire n_167;
wire n_675;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_11),
.B(n_14),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_19),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx6_ASAP7_75t_SL g30 ( 
.A(n_15),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

BUFx8_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_12),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_11),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_13),
.Y(n_47)
);

BUFx10_ASAP7_75t_L g48 ( 
.A(n_6),
.Y(n_48)
);

BUFx12_ASAP7_75t_L g49 ( 
.A(n_10),
.Y(n_49)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_19),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_11),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_15),
.Y(n_52)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_19),
.Y(n_53)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_15),
.Y(n_54)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_6),
.Y(n_55)
);

BUFx16f_ASAP7_75t_L g56 ( 
.A(n_12),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_6),
.Y(n_57)
);

BUFx10_ASAP7_75t_L g58 ( 
.A(n_12),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_19),
.B(n_12),
.Y(n_59)
);

INVx13_ASAP7_75t_L g60 ( 
.A(n_9),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_22),
.B(n_7),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_61),
.B(n_79),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_21),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_62),
.Y(n_164)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_51),
.Y(n_63)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_63),
.Y(n_135)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_64),
.Y(n_146)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

INVx2_ASAP7_75t_SL g216 ( 
.A(n_65),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_21),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_66),
.Y(n_179)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_55),
.Y(n_67)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_67),
.Y(n_148)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

INVx1_ASAP7_75t_SL g226 ( 
.A(n_68),
.Y(n_226)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_51),
.Y(n_69)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_69),
.Y(n_156)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_21),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_70),
.Y(n_186)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_55),
.Y(n_71)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_71),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_30),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g172 ( 
.A(n_72),
.Y(n_172)
);

BUFx5_ASAP7_75t_L g73 ( 
.A(n_30),
.Y(n_73)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_73),
.Y(n_138)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_24),
.Y(n_74)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_74),
.Y(n_136)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_36),
.Y(n_75)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_75),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_21),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_76),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_28),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_77),
.Y(n_229)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_30),
.Y(n_78)
);

BUFx2_ASAP7_75t_L g224 ( 
.A(n_78),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_22),
.B(n_18),
.Y(n_79)
);

INVx11_ASAP7_75t_L g80 ( 
.A(n_38),
.Y(n_80)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_80),
.Y(n_162)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_34),
.Y(n_81)
);

INVx5_ASAP7_75t_L g141 ( 
.A(n_81),
.Y(n_141)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_24),
.Y(n_82)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_82),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_28),
.Y(n_83)
);

INVx6_ASAP7_75t_L g144 ( 
.A(n_83),
.Y(n_144)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_36),
.Y(n_84)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_84),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_28),
.Y(n_85)
);

INVx3_ASAP7_75t_SL g208 ( 
.A(n_85),
.Y(n_208)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_46),
.Y(n_86)
);

INVx5_ASAP7_75t_L g170 ( 
.A(n_86),
.Y(n_170)
);

BUFx12f_ASAP7_75t_L g87 ( 
.A(n_38),
.Y(n_87)
);

INVx8_ASAP7_75t_L g158 ( 
.A(n_87),
.Y(n_158)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_55),
.Y(n_88)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_88),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_59),
.B(n_18),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_89),
.B(n_102),
.Y(n_183)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_50),
.Y(n_90)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_90),
.Y(n_198)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_28),
.Y(n_91)
);

INVx5_ASAP7_75t_L g173 ( 
.A(n_91),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_39),
.Y(n_92)
);

INVx5_ASAP7_75t_L g184 ( 
.A(n_92),
.Y(n_184)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_50),
.Y(n_93)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_93),
.Y(n_199)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_50),
.Y(n_94)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_94),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_39),
.Y(n_95)
);

INVx5_ASAP7_75t_L g187 ( 
.A(n_95),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_56),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_96),
.B(n_134),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_39),
.Y(n_97)
);

INVx5_ASAP7_75t_L g204 ( 
.A(n_97),
.Y(n_204)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_25),
.Y(n_98)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_98),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_34),
.Y(n_99)
);

INVx5_ASAP7_75t_L g217 ( 
.A(n_99),
.Y(n_217)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_52),
.Y(n_100)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_100),
.Y(n_215)
);

BUFx12f_ASAP7_75t_L g101 ( 
.A(n_38),
.Y(n_101)
);

INVx5_ASAP7_75t_L g218 ( 
.A(n_101),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_59),
.B(n_7),
.Y(n_102)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_39),
.Y(n_103)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_103),
.Y(n_165)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_46),
.Y(n_104)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_104),
.Y(n_168)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_25),
.Y(n_105)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_105),
.Y(n_142)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_34),
.Y(n_106)
);

INVx4_ASAP7_75t_L g210 ( 
.A(n_106),
.Y(n_210)
);

INVx3_ASAP7_75t_SL g107 ( 
.A(n_38),
.Y(n_107)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_107),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_43),
.Y(n_108)
);

BUFx12f_ASAP7_75t_L g206 ( 
.A(n_108),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_43),
.Y(n_109)
);

BUFx12f_ASAP7_75t_L g211 ( 
.A(n_109),
.Y(n_211)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_29),
.Y(n_110)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_110),
.Y(n_185)
);

INVx11_ASAP7_75t_L g111 ( 
.A(n_38),
.Y(n_111)
);

INVx4_ASAP7_75t_L g219 ( 
.A(n_111),
.Y(n_219)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_52),
.Y(n_112)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_112),
.Y(n_150)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_52),
.Y(n_113)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_113),
.Y(n_152)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_53),
.Y(n_114)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_114),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_31),
.B(n_45),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_115),
.B(n_120),
.Y(n_188)
);

INVx8_ASAP7_75t_L g116 ( 
.A(n_46),
.Y(n_116)
);

INVx3_ASAP7_75t_L g220 ( 
.A(n_116),
.Y(n_220)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_56),
.Y(n_117)
);

INVx4_ASAP7_75t_L g222 ( 
.A(n_117),
.Y(n_222)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_53),
.Y(n_118)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_118),
.Y(n_180)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_53),
.Y(n_119)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_119),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_31),
.B(n_40),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_43),
.Y(n_121)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_121),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_33),
.B(n_8),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_122),
.B(n_10),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_43),
.Y(n_123)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_123),
.Y(n_228)
);

INVx8_ASAP7_75t_L g124 ( 
.A(n_46),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g190 ( 
.A(n_124),
.B(n_128),
.Y(n_190)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_44),
.Y(n_125)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_125),
.Y(n_193)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_47),
.Y(n_126)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_126),
.Y(n_203)
);

BUFx12_ASAP7_75t_L g127 ( 
.A(n_56),
.Y(n_127)
);

CKINVDCx14_ASAP7_75t_R g230 ( 
.A(n_127),
.Y(n_230)
);

INVx8_ASAP7_75t_L g128 ( 
.A(n_46),
.Y(n_128)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_56),
.Y(n_129)
);

NAND2xp33_ASAP7_75t_SL g157 ( 
.A(n_129),
.B(n_133),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_47),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_130),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_47),
.Y(n_131)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_131),
.Y(n_205)
);

BUFx5_ASAP7_75t_L g132 ( 
.A(n_56),
.Y(n_132)
);

INVx5_ASAP7_75t_SL g169 ( 
.A(n_132),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_47),
.Y(n_133)
);

INVx8_ASAP7_75t_L g134 ( 
.A(n_35),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_70),
.A2(n_35),
.B1(n_41),
.B2(n_20),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_145),
.A2(n_175),
.B1(n_221),
.B2(n_162),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_87),
.A2(n_54),
.B1(n_35),
.B2(n_57),
.Y(n_149)
);

OA22x2_ASAP7_75t_L g283 ( 
.A1(n_149),
.A2(n_154),
.B1(n_155),
.B2(n_174),
.Y(n_283)
);

AOI22xp33_ASAP7_75t_L g151 ( 
.A1(n_62),
.A2(n_35),
.B1(n_57),
.B2(n_26),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_151),
.A2(n_196),
.B1(n_202),
.B2(n_207),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_87),
.A2(n_54),
.B1(n_26),
.B2(n_40),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_101),
.A2(n_54),
.B1(n_33),
.B2(n_45),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_72),
.B(n_42),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_159),
.B(n_161),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_78),
.B(n_20),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_91),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_163),
.B(n_166),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_117),
.B(n_41),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_101),
.B(n_42),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g310 ( 
.A(n_167),
.B(n_171),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_81),
.B(n_37),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_110),
.A2(n_37),
.B1(n_23),
.B2(n_32),
.Y(n_174)
);

OAI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_66),
.A2(n_32),
.B1(n_23),
.B2(n_58),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_99),
.B(n_11),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_177),
.B(n_178),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_67),
.B(n_13),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_106),
.B(n_13),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_182),
.B(n_191),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_71),
.B(n_16),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_192),
.B(n_194),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_107),
.B(n_16),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_103),
.A2(n_58),
.B1(n_27),
.B2(n_48),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_76),
.B(n_58),
.C(n_27),
.Y(n_200)
);

AND2x2_ASAP7_75t_L g234 ( 
.A(n_200),
.B(n_133),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_86),
.B(n_16),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_201),
.B(n_225),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_77),
.A2(n_58),
.B1(n_27),
.B2(n_48),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_L g207 ( 
.A1(n_83),
.A2(n_48),
.B1(n_58),
.B2(n_27),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_85),
.A2(n_58),
.B1(n_27),
.B2(n_48),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_209),
.A2(n_131),
.B(n_130),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_126),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_213),
.B(n_134),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_L g214 ( 
.A1(n_92),
.A2(n_48),
.B1(n_27),
.B2(n_60),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_214),
.A2(n_231),
.B1(n_0),
.B2(n_1),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_95),
.A2(n_48),
.B1(n_29),
.B2(n_60),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_97),
.B(n_18),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_108),
.A2(n_60),
.B1(n_49),
.B2(n_29),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_109),
.B(n_18),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_232),
.B(n_0),
.Y(n_270)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_136),
.Y(n_233)
);

INVx1_ASAP7_75t_SL g327 ( 
.A(n_233),
.Y(n_327)
);

AND2x2_ASAP7_75t_L g332 ( 
.A(n_234),
.B(n_264),
.Y(n_332)
);

CKINVDCx16_ASAP7_75t_R g236 ( 
.A(n_224),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g348 ( 
.A(n_236),
.B(n_271),
.Y(n_348)
);

INVx6_ASAP7_75t_L g238 ( 
.A(n_164),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g338 ( 
.A(n_238),
.Y(n_338)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_239),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_230),
.Y(n_240)
);

NAND3xp33_ASAP7_75t_L g379 ( 
.A(n_240),
.B(n_259),
.C(n_270),
.Y(n_379)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_203),
.Y(n_241)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_241),
.Y(n_322)
);

INVx11_ASAP7_75t_L g242 ( 
.A(n_206),
.Y(n_242)
);

INVx4_ASAP7_75t_L g333 ( 
.A(n_242),
.Y(n_333)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_137),
.Y(n_244)
);

INVx1_ASAP7_75t_SL g368 ( 
.A(n_244),
.Y(n_368)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_205),
.Y(n_247)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_247),
.Y(n_325)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_140),
.Y(n_249)
);

INVx1_ASAP7_75t_SL g376 ( 
.A(n_249),
.Y(n_376)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_142),
.Y(n_250)
);

INVx1_ASAP7_75t_SL g378 ( 
.A(n_250),
.Y(n_378)
);

OAI21xp33_ASAP7_75t_L g335 ( 
.A1(n_251),
.A2(n_265),
.B(n_267),
.Y(n_335)
);

BUFx3_ASAP7_75t_L g252 ( 
.A(n_218),
.Y(n_252)
);

INVxp67_ASAP7_75t_SL g356 ( 
.A(n_252),
.Y(n_356)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_143),
.Y(n_253)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_253),
.Y(n_340)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_193),
.Y(n_254)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_254),
.Y(n_349)
);

INVx2_ASAP7_75t_SL g255 ( 
.A(n_147),
.Y(n_255)
);

INVx2_ASAP7_75t_SL g355 ( 
.A(n_255),
.Y(n_355)
);

INVx5_ASAP7_75t_L g256 ( 
.A(n_158),
.Y(n_256)
);

INVx4_ASAP7_75t_L g346 ( 
.A(n_256),
.Y(n_346)
);

OAI22xp33_ASAP7_75t_SL g257 ( 
.A1(n_151),
.A2(n_121),
.B1(n_123),
.B2(n_127),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_257),
.A2(n_207),
.B1(n_160),
.B2(n_214),
.Y(n_324)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_165),
.Y(n_258)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_258),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_224),
.Y(n_259)
);

INVx4_ASAP7_75t_L g260 ( 
.A(n_158),
.Y(n_260)
);

INVx4_ASAP7_75t_L g370 ( 
.A(n_260),
.Y(n_370)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_165),
.Y(n_261)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_261),
.Y(n_341)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_150),
.Y(n_262)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_262),
.Y(n_351)
);

INVx3_ASAP7_75t_SL g263 ( 
.A(n_190),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g366 ( 
.A(n_263),
.Y(n_366)
);

AND2x2_ASAP7_75t_L g265 ( 
.A(n_188),
.B(n_128),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_208),
.Y(n_266)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_266),
.Y(n_342)
);

OAI21xp33_ASAP7_75t_L g267 ( 
.A1(n_157),
.A2(n_16),
.B(n_9),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_139),
.B(n_124),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_268),
.B(n_285),
.Y(n_321)
);

AOI22xp33_ASAP7_75t_SL g269 ( 
.A1(n_138),
.A2(n_104),
.B1(n_116),
.B2(n_49),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_SL g326 ( 
.A1(n_269),
.A2(n_294),
.B1(n_305),
.B2(n_307),
.Y(n_326)
);

CKINVDCx14_ASAP7_75t_R g271 ( 
.A(n_190),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_183),
.B(n_189),
.Y(n_272)
);

NOR2xp67_ASAP7_75t_R g365 ( 
.A(n_272),
.B(n_282),
.Y(n_365)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_152),
.Y(n_273)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_273),
.Y(n_353)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_208),
.Y(n_274)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_274),
.Y(n_357)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_135),
.Y(n_275)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_275),
.Y(n_381)
);

INVx4_ASAP7_75t_SL g276 ( 
.A(n_185),
.Y(n_276)
);

INVx4_ASAP7_75t_SL g360 ( 
.A(n_276),
.Y(n_360)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_176),
.Y(n_277)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_277),
.Y(n_362)
);

HB1xp67_ASAP7_75t_L g278 ( 
.A(n_216),
.Y(n_278)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_278),
.Y(n_364)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_180),
.Y(n_279)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_279),
.Y(n_367)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_181),
.Y(n_280)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_280),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_195),
.B(n_9),
.Y(n_282)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_146),
.Y(n_284)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_284),
.Y(n_380)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_174),
.Y(n_285)
);

OA22x2_ASAP7_75t_L g286 ( 
.A1(n_209),
.A2(n_49),
.B1(n_1),
.B2(n_2),
.Y(n_286)
);

AO22x1_ASAP7_75t_L g374 ( 
.A1(n_286),
.A2(n_172),
.B1(n_204),
.B2(n_187),
.Y(n_374)
);

INVx4_ASAP7_75t_L g287 ( 
.A(n_218),
.Y(n_287)
);

INVx3_ASAP7_75t_L g369 ( 
.A(n_287),
.Y(n_369)
);

INVx3_ASAP7_75t_L g288 ( 
.A(n_170),
.Y(n_288)
);

INVx3_ASAP7_75t_L g375 ( 
.A(n_288),
.Y(n_375)
);

CKINVDCx14_ASAP7_75t_R g289 ( 
.A(n_169),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_289),
.B(n_293),
.Y(n_323)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_156),
.Y(n_290)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_290),
.Y(n_344)
);

INVx4_ASAP7_75t_L g291 ( 
.A(n_170),
.Y(n_291)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_291),
.Y(n_373)
);

INVx5_ASAP7_75t_L g292 ( 
.A(n_141),
.Y(n_292)
);

BUFx6f_ASAP7_75t_L g354 ( 
.A(n_292),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_198),
.B(n_9),
.Y(n_293)
);

AOI22xp33_ASAP7_75t_SL g294 ( 
.A1(n_138),
.A2(n_49),
.B1(n_1),
.B2(n_2),
.Y(n_294)
);

INVx5_ASAP7_75t_L g295 ( 
.A(n_141),
.Y(n_295)
);

AND2x2_ASAP7_75t_L g361 ( 
.A(n_295),
.B(n_297),
.Y(n_361)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_197),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_296),
.B(n_298),
.Y(n_328)
);

INVx3_ASAP7_75t_L g297 ( 
.A(n_222),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_199),
.Y(n_298)
);

INVx3_ASAP7_75t_L g299 ( 
.A(n_222),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_299),
.B(n_300),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_212),
.A2(n_49),
.B(n_1),
.Y(n_300)
);

CKINVDCx16_ASAP7_75t_R g301 ( 
.A(n_169),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_301),
.B(n_302),
.Y(n_358)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_210),
.Y(n_302)
);

INVx4_ASAP7_75t_L g303 ( 
.A(n_168),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_303),
.B(n_306),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_175),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g319 ( 
.A1(n_304),
.A2(n_311),
.B1(n_294),
.B2(n_149),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_172),
.B(n_0),
.Y(n_306)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_210),
.Y(n_307)
);

AND2x2_ASAP7_75t_L g308 ( 
.A(n_226),
.B(n_3),
.Y(n_308)
);

NAND2xp33_ASAP7_75t_SL g320 ( 
.A(n_308),
.B(n_313),
.Y(n_320)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_215),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_309),
.B(n_312),
.Y(n_337)
);

AOI22xp33_ASAP7_75t_SL g311 ( 
.A1(n_185),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_223),
.Y(n_312)
);

AND2x2_ASAP7_75t_L g313 ( 
.A(n_226),
.B(n_3),
.Y(n_313)
);

INVx4_ASAP7_75t_L g314 ( 
.A(n_168),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_314),
.B(n_315),
.Y(n_345)
);

INVx5_ASAP7_75t_L g315 ( 
.A(n_217),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g316 ( 
.A(n_216),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_316),
.B(n_317),
.Y(n_347)
);

HB1xp67_ASAP7_75t_L g317 ( 
.A(n_148),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_234),
.B(n_265),
.C(n_263),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_318),
.B(n_148),
.C(n_153),
.Y(n_423)
);

AOI22xp33_ASAP7_75t_SL g409 ( 
.A1(n_319),
.A2(n_302),
.B1(n_258),
.B2(n_295),
.Y(n_409)
);

AND2x2_ASAP7_75t_L g390 ( 
.A(n_324),
.B(n_374),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_L g329 ( 
.A1(n_237),
.A2(n_264),
.B1(n_245),
.B2(n_235),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g403 ( 
.A1(n_329),
.A2(n_352),
.B1(n_288),
.B2(n_312),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_285),
.A2(n_304),
.B1(n_267),
.B2(n_286),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_L g429 ( 
.A1(n_330),
.A2(n_339),
.B1(n_343),
.B2(n_377),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_286),
.A2(n_200),
.B1(n_228),
.B2(n_223),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_286),
.A2(n_228),
.B1(n_186),
.B2(n_173),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_246),
.B(n_173),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_350),
.B(n_372),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_L g352 ( 
.A1(n_243),
.A2(n_154),
.B1(n_155),
.B2(n_144),
.Y(n_352)
);

AOI32xp33_ASAP7_75t_L g363 ( 
.A1(n_310),
.A2(n_162),
.A3(n_219),
.B1(n_217),
.B2(n_153),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_363),
.B(n_283),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_281),
.B(n_313),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_283),
.A2(n_186),
.B1(n_229),
.B2(n_227),
.Y(n_377)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_337),
.Y(n_382)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_382),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_334),
.B(n_248),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_SL g462 ( 
.A(n_383),
.B(n_385),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_332),
.A2(n_283),
.B1(n_269),
.B2(n_144),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g435 ( 
.A1(n_384),
.A2(n_400),
.B1(n_403),
.B2(n_412),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_SL g385 ( 
.A(n_350),
.B(n_284),
.Y(n_385)
);

CKINVDCx16_ASAP7_75t_R g386 ( 
.A(n_361),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_386),
.B(n_387),
.Y(n_459)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_337),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_355),
.Y(n_388)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_388),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_L g391 ( 
.A(n_318),
.B(n_255),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_391),
.B(n_423),
.C(n_431),
.Y(n_456)
);

OR2x2_ASAP7_75t_L g450 ( 
.A(n_392),
.B(n_417),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_SL g393 ( 
.A(n_372),
.B(n_323),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_SL g465 ( 
.A(n_393),
.B(n_401),
.Y(n_465)
);

CKINVDCx16_ASAP7_75t_R g394 ( 
.A(n_361),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_394),
.B(n_407),
.Y(n_463)
);

INVx3_ASAP7_75t_L g395 ( 
.A(n_354),
.Y(n_395)
);

INVx4_ASAP7_75t_L g468 ( 
.A(n_395),
.Y(n_468)
);

XOR2x1_ASAP7_75t_SL g396 ( 
.A(n_332),
.B(n_335),
.Y(n_396)
);

OAI21xp5_ASAP7_75t_L g446 ( 
.A1(n_396),
.A2(n_398),
.B(n_410),
.Y(n_446)
);

AND2x2_ASAP7_75t_SL g397 ( 
.A(n_332),
.B(n_308),
.Y(n_397)
);

CKINVDCx16_ASAP7_75t_R g461 ( 
.A(n_397),
.Y(n_461)
);

OAI21xp5_ASAP7_75t_L g398 ( 
.A1(n_321),
.A2(n_283),
.B(n_311),
.Y(n_398)
);

AO21x2_ASAP7_75t_SL g399 ( 
.A1(n_374),
.A2(n_276),
.B(n_314),
.Y(n_399)
);

OA22x2_ASAP7_75t_L g469 ( 
.A1(n_399),
.A2(n_346),
.B1(n_333),
.B2(n_375),
.Y(n_469)
);

OAI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_339),
.A2(n_164),
.B1(n_179),
.B2(n_227),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_SL g401 ( 
.A(n_340),
.B(n_290),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_320),
.B(n_275),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_402),
.B(n_418),
.Y(n_434)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_355),
.Y(n_404)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_404),
.Y(n_442)
);

AOI22xp33_ASAP7_75t_L g405 ( 
.A1(n_331),
.A2(n_247),
.B1(n_241),
.B2(n_261),
.Y(n_405)
);

AOI22xp33_ASAP7_75t_SL g452 ( 
.A1(n_405),
.A2(n_360),
.B1(n_368),
.B2(n_378),
.Y(n_452)
);

AOI22x1_ASAP7_75t_SL g406 ( 
.A1(n_330),
.A2(n_291),
.B1(n_303),
.B2(n_307),
.Y(n_406)
);

CKINVDCx16_ASAP7_75t_R g467 ( 
.A(n_406),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_328),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_342),
.Y(n_408)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_408),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_L g444 ( 
.A1(n_409),
.A2(n_386),
.B1(n_394),
.B2(n_411),
.Y(n_444)
);

OAI21xp5_ASAP7_75t_L g410 ( 
.A1(n_379),
.A2(n_316),
.B(n_297),
.Y(n_410)
);

CKINVDCx16_ASAP7_75t_R g411 ( 
.A(n_361),
.Y(n_411)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_411),
.Y(n_454)
);

OAI22x1_ASAP7_75t_SL g412 ( 
.A1(n_377),
.A2(n_242),
.B1(n_260),
.B2(n_219),
.Y(n_412)
);

INVx1_ASAP7_75t_SL g413 ( 
.A(n_360),
.Y(n_413)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_413),
.Y(n_473)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_355),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_SL g466 ( 
.A(n_414),
.B(n_415),
.Y(n_466)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_347),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_345),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_416),
.B(n_325),
.Y(n_475)
);

AOI22xp5_ASAP7_75t_SL g417 ( 
.A1(n_374),
.A2(n_315),
.B1(n_292),
.B2(n_256),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_347),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_359),
.B(n_299),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_419),
.B(n_421),
.Y(n_439)
);

HB1xp67_ASAP7_75t_L g420 ( 
.A(n_364),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_420),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_320),
.B(n_345),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_325),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_422),
.B(n_424),
.Y(n_445)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_342),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_SL g425 ( 
.A1(n_343),
.A2(n_179),
.B1(n_229),
.B2(n_184),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_L g470 ( 
.A1(n_425),
.A2(n_427),
.B1(n_274),
.B2(n_266),
.Y(n_470)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_357),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_426),
.B(n_428),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_SL g427 ( 
.A1(n_326),
.A2(n_184),
.B1(n_204),
.B2(n_187),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_357),
.Y(n_428)
);

CKINVDCx16_ASAP7_75t_R g430 ( 
.A(n_358),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_430),
.B(n_432),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_366),
.B(n_348),
.C(n_351),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_365),
.B(n_238),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_SL g436 ( 
.A1(n_403),
.A2(n_324),
.B1(n_365),
.B2(n_366),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_436),
.B(n_437),
.Y(n_491)
);

A2O1A1Ixp33_ASAP7_75t_L g437 ( 
.A1(n_432),
.A2(n_373),
.B(n_344),
.C(n_362),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_SL g441 ( 
.A1(n_415),
.A2(n_368),
.B1(n_327),
.B2(n_378),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_441),
.B(n_449),
.Y(n_508)
);

AOI21xp5_ASAP7_75t_L g443 ( 
.A1(n_398),
.A2(n_333),
.B(n_356),
.Y(n_443)
);

AOI21xp5_ASAP7_75t_L g496 ( 
.A1(n_443),
.A2(n_402),
.B(n_390),
.Y(n_496)
);

AOI22xp5_ASAP7_75t_SL g476 ( 
.A1(n_444),
.A2(n_384),
.B1(n_429),
.B2(n_399),
.Y(n_476)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_419),
.Y(n_447)
);

CKINVDCx14_ASAP7_75t_R g487 ( 
.A(n_447),
.Y(n_487)
);

A2O1A1Ixp33_ASAP7_75t_L g449 ( 
.A1(n_399),
.A2(n_373),
.B(n_344),
.C(n_367),
.Y(n_449)
);

OAI22xp33_ASAP7_75t_SL g477 ( 
.A1(n_452),
.A2(n_470),
.B1(n_417),
.B2(n_399),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_385),
.Y(n_453)
);

AND2x2_ASAP7_75t_L g480 ( 
.A(n_453),
.B(n_469),
.Y(n_480)
);

OAI22xp5_ASAP7_75t_SL g455 ( 
.A1(n_418),
.A2(n_327),
.B1(n_376),
.B2(n_338),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_455),
.B(n_460),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_391),
.B(n_371),
.C(n_353),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_458),
.B(n_471),
.C(n_396),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_387),
.B(n_376),
.Y(n_460)
);

OAI22xp5_ASAP7_75t_SL g464 ( 
.A1(n_416),
.A2(n_338),
.B1(n_349),
.B2(n_375),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_464),
.B(n_475),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_423),
.B(n_380),
.C(n_381),
.Y(n_471)
);

CKINVDCx20_ASAP7_75t_R g472 ( 
.A(n_399),
.Y(n_472)
);

AND2x2_ASAP7_75t_L g490 ( 
.A(n_472),
.B(n_390),
.Y(n_490)
);

OAI21xp5_ASAP7_75t_L g474 ( 
.A1(n_421),
.A2(n_346),
.B(n_370),
.Y(n_474)
);

OAI21xp5_ASAP7_75t_L g501 ( 
.A1(n_474),
.A2(n_413),
.B(n_390),
.Y(n_501)
);

OAI22xp5_ASAP7_75t_L g531 ( 
.A1(n_476),
.A2(n_503),
.B1(n_444),
.B2(n_443),
.Y(n_531)
);

AOI22xp5_ASAP7_75t_SL g547 ( 
.A1(n_477),
.A2(n_454),
.B1(n_461),
.B2(n_469),
.Y(n_547)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_438),
.Y(n_478)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_478),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_479),
.B(n_482),
.C(n_483),
.Y(n_522)
);

CKINVDCx16_ASAP7_75t_R g481 ( 
.A(n_445),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_SL g552 ( 
.A(n_481),
.B(n_484),
.Y(n_552)
);

XOR2xp5_ASAP7_75t_L g482 ( 
.A(n_456),
.B(n_458),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_456),
.B(n_397),
.C(n_389),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_SL g484 ( 
.A(n_465),
.B(n_407),
.Y(n_484)
);

CKINVDCx20_ASAP7_75t_R g485 ( 
.A(n_448),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_485),
.B(n_499),
.Y(n_520)
);

XNOR2xp5_ASAP7_75t_L g486 ( 
.A(n_456),
.B(n_389),
.Y(n_486)
);

XOR2xp5_ASAP7_75t_L g518 ( 
.A(n_486),
.B(n_500),
.Y(n_518)
);

OAI22xp5_ASAP7_75t_SL g488 ( 
.A1(n_450),
.A2(n_435),
.B1(n_472),
.B2(n_433),
.Y(n_488)
);

AOI22xp5_ASAP7_75t_L g539 ( 
.A1(n_488),
.A2(n_514),
.B1(n_515),
.B2(n_449),
.Y(n_539)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_438),
.Y(n_489)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_489),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_490),
.Y(n_535)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_442),
.Y(n_492)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_492),
.Y(n_536)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_442),
.Y(n_493)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_493),
.Y(n_538)
);

BUFx6f_ASAP7_75t_L g494 ( 
.A(n_468),
.Y(n_494)
);

CKINVDCx20_ASAP7_75t_R g519 ( 
.A(n_494),
.Y(n_519)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_475),
.Y(n_495)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_495),
.Y(n_540)
);

AOI21xp5_ASAP7_75t_L g523 ( 
.A1(n_496),
.A2(n_501),
.B(n_509),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_SL g497 ( 
.A(n_462),
.B(n_430),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_497),
.B(n_505),
.Y(n_532)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_458),
.B(n_397),
.C(n_382),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g525 ( 
.A(n_498),
.B(n_506),
.C(n_446),
.Y(n_525)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_445),
.Y(n_499)
);

XNOR2xp5_ASAP7_75t_L g500 ( 
.A(n_459),
.B(n_431),
.Y(n_500)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_464),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_502),
.B(n_504),
.Y(n_530)
);

AOI22xp5_ASAP7_75t_SL g503 ( 
.A1(n_467),
.A2(n_429),
.B1(n_427),
.B2(n_400),
.Y(n_503)
);

CKINVDCx20_ASAP7_75t_R g504 ( 
.A(n_448),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_462),
.B(n_393),
.Y(n_505)
);

XOR2xp5_ASAP7_75t_L g506 ( 
.A(n_463),
.B(n_410),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_466),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_507),
.B(n_511),
.Y(n_541)
);

OAI21xp5_ASAP7_75t_L g509 ( 
.A1(n_446),
.A2(n_388),
.B(n_404),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_463),
.B(n_465),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g551 ( 
.A(n_510),
.B(n_440),
.Y(n_551)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_466),
.Y(n_511)
);

OAI22xp5_ASAP7_75t_SL g514 ( 
.A1(n_450),
.A2(n_406),
.B1(n_412),
.B2(n_425),
.Y(n_514)
);

OAI22xp33_ASAP7_75t_L g515 ( 
.A1(n_467),
.A2(n_414),
.B1(n_395),
.B2(n_422),
.Y(n_515)
);

CKINVDCx16_ASAP7_75t_R g516 ( 
.A(n_480),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_516),
.B(n_521),
.Y(n_578)
);

XNOR2xp5_ASAP7_75t_L g517 ( 
.A(n_482),
.B(n_457),
.Y(n_517)
);

XOR2xp5_ASAP7_75t_L g563 ( 
.A(n_517),
.B(n_528),
.Y(n_563)
);

CKINVDCx20_ASAP7_75t_R g521 ( 
.A(n_487),
.Y(n_521)
);

XNOR2xp5_ASAP7_75t_L g566 ( 
.A(n_525),
.B(n_506),
.Y(n_566)
);

OAI22xp5_ASAP7_75t_SL g526 ( 
.A1(n_476),
.A2(n_450),
.B1(n_435),
.B2(n_457),
.Y(n_526)
);

AOI22xp5_ASAP7_75t_L g556 ( 
.A1(n_526),
.A2(n_527),
.B1(n_537),
.B2(n_549),
.Y(n_556)
);

OAI22xp5_ASAP7_75t_SL g527 ( 
.A1(n_491),
.A2(n_433),
.B1(n_447),
.B2(n_453),
.Y(n_527)
);

XOR2xp5_ASAP7_75t_L g528 ( 
.A(n_486),
.B(n_471),
.Y(n_528)
);

XNOR2xp5_ASAP7_75t_SL g529 ( 
.A(n_483),
.B(n_459),
.Y(n_529)
);

XNOR2xp5_ASAP7_75t_SL g560 ( 
.A(n_529),
.B(n_528),
.Y(n_560)
);

OAI22xp5_ASAP7_75t_L g559 ( 
.A1(n_531),
.A2(n_533),
.B1(n_539),
.B2(n_542),
.Y(n_559)
);

OAI22xp5_ASAP7_75t_L g533 ( 
.A1(n_503),
.A2(n_460),
.B1(n_439),
.B2(n_470),
.Y(n_533)
);

OAI22xp5_ASAP7_75t_SL g537 ( 
.A1(n_491),
.A2(n_439),
.B1(n_434),
.B2(n_461),
.Y(n_537)
);

AOI22xp5_ASAP7_75t_L g542 ( 
.A1(n_488),
.A2(n_449),
.B1(n_436),
.B2(n_437),
.Y(n_542)
);

XOR2xp5_ASAP7_75t_L g543 ( 
.A(n_479),
.B(n_471),
.Y(n_543)
);

MAJIxp5_ASAP7_75t_L g562 ( 
.A(n_543),
.B(n_544),
.C(n_550),
.Y(n_562)
);

XOR2xp5_ASAP7_75t_L g544 ( 
.A(n_500),
.B(n_434),
.Y(n_544)
);

AOI22x1_ASAP7_75t_L g545 ( 
.A1(n_480),
.A2(n_469),
.B1(n_474),
.B2(n_455),
.Y(n_545)
);

HB1xp67_ASAP7_75t_L g564 ( 
.A(n_545),
.Y(n_564)
);

CKINVDCx20_ASAP7_75t_R g546 ( 
.A(n_480),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_546),
.B(n_514),
.Y(n_580)
);

OAI22xp5_ASAP7_75t_SL g582 ( 
.A1(n_547),
.A2(n_468),
.B1(n_451),
.B2(n_494),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_507),
.B(n_440),
.Y(n_548)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_548),
.Y(n_568)
);

OAI22xp5_ASAP7_75t_SL g549 ( 
.A1(n_495),
.A2(n_474),
.B1(n_454),
.B2(n_437),
.Y(n_549)
);

XOR2xp5_ASAP7_75t_L g550 ( 
.A(n_498),
.B(n_441),
.Y(n_550)
);

NAND3xp33_ASAP7_75t_L g570 ( 
.A(n_551),
.B(n_553),
.C(n_512),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_L g553 ( 
.A(n_511),
.B(n_473),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_513),
.B(n_469),
.Y(n_554)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_554),
.Y(n_581)
);

OAI22xp5_ASAP7_75t_L g555 ( 
.A1(n_502),
.A2(n_452),
.B1(n_473),
.B2(n_469),
.Y(n_555)
);

BUFx2_ASAP7_75t_L g577 ( 
.A(n_555),
.Y(n_577)
);

OAI21xp5_ASAP7_75t_SL g557 ( 
.A1(n_523),
.A2(n_508),
.B(n_509),
.Y(n_557)
);

AOI21xp5_ASAP7_75t_L g591 ( 
.A1(n_557),
.A2(n_565),
.B(n_575),
.Y(n_591)
);

AOI22xp5_ASAP7_75t_L g558 ( 
.A1(n_526),
.A2(n_508),
.B1(n_501),
.B2(n_490),
.Y(n_558)
);

OAI22xp5_ASAP7_75t_L g596 ( 
.A1(n_558),
.A2(n_567),
.B1(n_570),
.B2(n_573),
.Y(n_596)
);

XNOR2xp5_ASAP7_75t_L g595 ( 
.A(n_560),
.B(n_566),
.Y(n_595)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_524),
.Y(n_561)
);

INVx1_ASAP7_75t_SL g615 ( 
.A(n_561),
.Y(n_615)
);

AOI21xp5_ASAP7_75t_L g565 ( 
.A1(n_523),
.A2(n_490),
.B(n_496),
.Y(n_565)
);

AOI22xp5_ASAP7_75t_L g567 ( 
.A1(n_527),
.A2(n_512),
.B1(n_504),
.B2(n_485),
.Y(n_567)
);

XNOR2xp5_ASAP7_75t_L g569 ( 
.A(n_518),
.B(n_499),
.Y(n_569)
);

XNOR2xp5_ASAP7_75t_L g604 ( 
.A(n_569),
.B(n_585),
.Y(n_604)
);

MAJIxp5_ASAP7_75t_L g571 ( 
.A(n_543),
.B(n_478),
.C(n_493),
.Y(n_571)
);

MAJIxp5_ASAP7_75t_L g593 ( 
.A(n_571),
.B(n_572),
.C(n_576),
.Y(n_593)
);

MAJIxp5_ASAP7_75t_L g572 ( 
.A(n_522),
.B(n_492),
.C(n_489),
.Y(n_572)
);

CKINVDCx14_ASAP7_75t_R g573 ( 
.A(n_552),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_SL g574 ( 
.A(n_532),
.B(n_428),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_SL g592 ( 
.A(n_574),
.B(n_583),
.Y(n_592)
);

AOI21xp5_ASAP7_75t_L g575 ( 
.A1(n_546),
.A2(n_515),
.B(n_513),
.Y(n_575)
);

MAJIxp5_ASAP7_75t_L g576 ( 
.A(n_522),
.B(n_518),
.C(n_525),
.Y(n_576)
);

MAJIxp5_ASAP7_75t_L g579 ( 
.A(n_550),
.B(n_451),
.C(n_369),
.Y(n_579)
);

MAJIxp5_ASAP7_75t_L g594 ( 
.A(n_579),
.B(n_588),
.C(n_530),
.Y(n_594)
);

CKINVDCx20_ASAP7_75t_R g614 ( 
.A(n_580),
.Y(n_614)
);

AOI22xp5_ASAP7_75t_L g597 ( 
.A1(n_582),
.A2(n_539),
.B1(n_549),
.B2(n_542),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_SL g583 ( 
.A(n_521),
.B(n_426),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_541),
.B(n_424),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_SL g599 ( 
.A(n_584),
.B(n_586),
.Y(n_599)
);

XNOR2xp5_ASAP7_75t_L g585 ( 
.A(n_529),
.B(n_408),
.Y(n_585)
);

CKINVDCx16_ASAP7_75t_R g586 ( 
.A(n_548),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_541),
.Y(n_587)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_587),
.Y(n_611)
);

MAJIxp5_ASAP7_75t_L g588 ( 
.A(n_517),
.B(n_544),
.C(n_535),
.Y(n_588)
);

AOI22xp5_ASAP7_75t_L g589 ( 
.A1(n_554),
.A2(n_468),
.B1(n_354),
.B2(n_370),
.Y(n_589)
);

OAI22xp5_ASAP7_75t_L g606 ( 
.A1(n_589),
.A2(n_545),
.B1(n_519),
.B2(n_536),
.Y(n_606)
);

OAI21xp5_ASAP7_75t_L g590 ( 
.A1(n_535),
.A2(n_369),
.B(n_341),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_590),
.B(n_561),
.Y(n_613)
);

XNOR2xp5_ASAP7_75t_L g621 ( 
.A(n_594),
.B(n_607),
.Y(n_621)
);

INVxp33_ASAP7_75t_L g640 ( 
.A(n_597),
.Y(n_640)
);

HB1xp67_ASAP7_75t_L g598 ( 
.A(n_572),
.Y(n_598)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_598),
.Y(n_628)
);

MAJIxp5_ASAP7_75t_L g600 ( 
.A(n_563),
.B(n_540),
.C(n_520),
.Y(n_600)
);

MAJIxp5_ASAP7_75t_L g623 ( 
.A(n_600),
.B(n_605),
.C(n_608),
.Y(n_623)
);

AOI22xp5_ASAP7_75t_L g601 ( 
.A1(n_577),
.A2(n_530),
.B1(n_537),
.B2(n_540),
.Y(n_601)
);

AOI22xp5_ASAP7_75t_L g633 ( 
.A1(n_601),
.A2(n_606),
.B1(n_609),
.B2(n_610),
.Y(n_633)
);

HB1xp67_ASAP7_75t_L g602 ( 
.A(n_569),
.Y(n_602)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_602),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_L g603 ( 
.A(n_571),
.B(n_588),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_SL g620 ( 
.A(n_603),
.B(n_618),
.Y(n_620)
);

MAJIxp5_ASAP7_75t_L g605 ( 
.A(n_563),
.B(n_520),
.C(n_547),
.Y(n_605)
);

XNOR2xp5_ASAP7_75t_L g607 ( 
.A(n_576),
.B(n_545),
.Y(n_607)
);

MAJIxp5_ASAP7_75t_L g608 ( 
.A(n_562),
.B(n_538),
.C(n_536),
.Y(n_608)
);

OAI22xp5_ASAP7_75t_SL g609 ( 
.A1(n_577),
.A2(n_534),
.B1(n_524),
.B2(n_538),
.Y(n_609)
);

AOI22xp5_ASAP7_75t_L g610 ( 
.A1(n_559),
.A2(n_534),
.B1(n_519),
.B2(n_381),
.Y(n_610)
);

CKINVDCx16_ASAP7_75t_R g612 ( 
.A(n_578),
.Y(n_612)
);

NOR2xp33_ASAP7_75t_L g619 ( 
.A(n_612),
.B(n_568),
.Y(n_619)
);

INVx1_ASAP7_75t_SL g626 ( 
.A(n_613),
.Y(n_626)
);

AOI22xp5_ASAP7_75t_L g616 ( 
.A1(n_564),
.A2(n_341),
.B1(n_336),
.B2(n_322),
.Y(n_616)
);

AOI22xp5_ASAP7_75t_L g639 ( 
.A1(n_616),
.A2(n_615),
.B1(n_590),
.B2(n_582),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_567),
.B(n_322),
.Y(n_617)
);

CKINVDCx20_ASAP7_75t_R g622 ( 
.A(n_617),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g618 ( 
.A(n_579),
.B(n_336),
.Y(n_618)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_619),
.Y(n_648)
);

MAJIxp5_ASAP7_75t_L g624 ( 
.A(n_593),
.B(n_562),
.C(n_566),
.Y(n_624)
);

MAJIxp5_ASAP7_75t_L g659 ( 
.A(n_624),
.B(n_630),
.C(n_641),
.Y(n_659)
);

AOI21xp5_ASAP7_75t_SL g625 ( 
.A1(n_596),
.A2(n_557),
.B(n_581),
.Y(n_625)
);

OAI21xp5_ASAP7_75t_L g644 ( 
.A1(n_625),
.A2(n_601),
.B(n_617),
.Y(n_644)
);

XNOR2xp5_ASAP7_75t_L g627 ( 
.A(n_608),
.B(n_585),
.Y(n_627)
);

XNOR2xp5_ASAP7_75t_L g662 ( 
.A(n_627),
.B(n_629),
.Y(n_662)
);

XNOR2xp5_ASAP7_75t_L g629 ( 
.A(n_593),
.B(n_560),
.Y(n_629)
);

MAJIxp5_ASAP7_75t_L g630 ( 
.A(n_594),
.B(n_558),
.C(n_556),
.Y(n_630)
);

XOR2xp5_ASAP7_75t_L g631 ( 
.A(n_607),
.B(n_565),
.Y(n_631)
);

XNOR2xp5_ASAP7_75t_L g643 ( 
.A(n_631),
.B(n_636),
.Y(n_643)
);

OAI21xp5_ASAP7_75t_L g632 ( 
.A1(n_591),
.A2(n_556),
.B(n_575),
.Y(n_632)
);

AO21x1_ASAP7_75t_L g660 ( 
.A1(n_632),
.A2(n_642),
.B(n_595),
.Y(n_660)
);

OAI21xp5_ASAP7_75t_SL g635 ( 
.A1(n_591),
.A2(n_614),
.B(n_599),
.Y(n_635)
);

NOR2xp33_ASAP7_75t_SL g654 ( 
.A(n_635),
.B(n_638),
.Y(n_654)
);

XOR2xp5_ASAP7_75t_L g636 ( 
.A(n_600),
.B(n_605),
.Y(n_636)
);

HB1xp67_ASAP7_75t_L g637 ( 
.A(n_592),
.Y(n_637)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_637),
.Y(n_649)
);

CKINVDCx20_ASAP7_75t_R g638 ( 
.A(n_609),
.Y(n_638)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_639),
.Y(n_650)
);

XNOR2xp5_ASAP7_75t_SL g641 ( 
.A(n_595),
.B(n_589),
.Y(n_641)
);

NOR2xp67_ASAP7_75t_L g656 ( 
.A(n_641),
.B(n_604),
.Y(n_656)
);

OAI21xp5_ASAP7_75t_L g642 ( 
.A1(n_597),
.A2(n_287),
.B(n_252),
.Y(n_642)
);

OR2x2_ASAP7_75t_L g671 ( 
.A(n_644),
.B(n_658),
.Y(n_671)
);

OAI21xp5_ASAP7_75t_SL g645 ( 
.A1(n_625),
.A2(n_611),
.B(n_613),
.Y(n_645)
);

OAI21xp5_ASAP7_75t_SL g676 ( 
.A1(n_645),
.A2(n_3),
.B(n_4),
.Y(n_676)
);

NOR2xp33_ASAP7_75t_L g646 ( 
.A(n_620),
.B(n_611),
.Y(n_646)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_646),
.Y(n_665)
);

AND2x2_ASAP7_75t_L g647 ( 
.A(n_632),
.B(n_610),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_647),
.B(n_651),
.Y(n_670)
);

AND2x2_ASAP7_75t_L g651 ( 
.A(n_633),
.B(n_615),
.Y(n_651)
);

NOR2xp33_ASAP7_75t_L g652 ( 
.A(n_628),
.B(n_604),
.Y(n_652)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_652),
.Y(n_677)
);

INVxp67_ASAP7_75t_L g653 ( 
.A(n_634),
.Y(n_653)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_653),
.Y(n_678)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_626),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_655),
.B(n_657),
.Y(n_679)
);

OAI21xp5_ASAP7_75t_L g669 ( 
.A1(n_656),
.A2(n_627),
.B(n_629),
.Y(n_669)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_626),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_622),
.B(n_616),
.Y(n_658)
);

NOR2xp33_ASAP7_75t_L g672 ( 
.A(n_659),
.B(n_206),
.Y(n_672)
);

XOR2xp5_ASAP7_75t_L g664 ( 
.A(n_660),
.B(n_640),
.Y(n_664)
);

MAJIxp5_ASAP7_75t_L g661 ( 
.A(n_630),
.B(n_220),
.C(n_206),
.Y(n_661)
);

MAJIxp5_ASAP7_75t_L g663 ( 
.A(n_661),
.B(n_624),
.C(n_631),
.Y(n_663)
);

XNOR2xp5_ASAP7_75t_L g684 ( 
.A(n_663),
.B(n_664),
.Y(n_684)
);

OAI22xp5_ASAP7_75t_SL g666 ( 
.A1(n_650),
.A2(n_640),
.B1(n_639),
.B2(n_642),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_666),
.B(n_668),
.Y(n_687)
);

AOI21xp5_ASAP7_75t_L g667 ( 
.A1(n_654),
.A2(n_621),
.B(n_623),
.Y(n_667)
);

AOI21xp5_ASAP7_75t_L g680 ( 
.A1(n_667),
.A2(n_669),
.B(n_662),
.Y(n_680)
);

AOI22xp5_ASAP7_75t_L g668 ( 
.A1(n_651),
.A2(n_621),
.B1(n_636),
.B2(n_623),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_672),
.B(n_673),
.Y(n_689)
);

OAI22xp5_ASAP7_75t_SL g673 ( 
.A1(n_647),
.A2(n_220),
.B1(n_211),
.B2(n_5),
.Y(n_673)
);

NAND2x1p5_ASAP7_75t_L g674 ( 
.A(n_647),
.B(n_211),
.Y(n_674)
);

OAI21xp5_ASAP7_75t_L g683 ( 
.A1(n_674),
.A2(n_658),
.B(n_653),
.Y(n_683)
);

NOR2xp33_ASAP7_75t_L g675 ( 
.A(n_649),
.B(n_211),
.Y(n_675)
);

NOR2xp33_ASAP7_75t_SL g686 ( 
.A(n_675),
.B(n_651),
.Y(n_686)
);

AOI21xp5_ASAP7_75t_SL g682 ( 
.A1(n_676),
.A2(n_645),
.B(n_644),
.Y(n_682)
);

AOI21x1_ASAP7_75t_SL g697 ( 
.A1(n_680),
.A2(n_682),
.B(n_679),
.Y(n_697)
);

NOR2xp33_ASAP7_75t_L g681 ( 
.A(n_665),
.B(n_648),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_681),
.B(n_685),
.Y(n_695)
);

INVxp67_ASAP7_75t_L g698 ( 
.A(n_683),
.Y(n_698)
);

NOR2xp33_ASAP7_75t_L g685 ( 
.A(n_677),
.B(n_659),
.Y(n_685)
);

AOI22xp5_ASAP7_75t_L g701 ( 
.A1(n_686),
.A2(n_690),
.B1(n_691),
.B2(n_666),
.Y(n_701)
);

XOR2xp5_ASAP7_75t_L g688 ( 
.A(n_669),
.B(n_643),
.Y(n_688)
);

MAJIxp5_ASAP7_75t_L g694 ( 
.A(n_688),
.B(n_663),
.C(n_664),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_SL g690 ( 
.A(n_667),
.B(n_662),
.Y(n_690)
);

NOR2xp33_ASAP7_75t_L g691 ( 
.A(n_678),
.B(n_643),
.Y(n_691)
);

NOR2xp33_ASAP7_75t_SL g692 ( 
.A(n_668),
.B(n_660),
.Y(n_692)
);

AOI21xp5_ASAP7_75t_L g699 ( 
.A1(n_692),
.A2(n_671),
.B(n_670),
.Y(n_699)
);

AOI21x1_ASAP7_75t_L g693 ( 
.A1(n_687),
.A2(n_671),
.B(n_679),
.Y(n_693)
);

OAI21x1_ASAP7_75t_SL g704 ( 
.A1(n_693),
.A2(n_697),
.B(n_699),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_694),
.B(n_696),
.Y(n_706)
);

INVxp67_ASAP7_75t_L g696 ( 
.A(n_688),
.Y(n_696)
);

OAI21xp5_ASAP7_75t_SL g700 ( 
.A1(n_682),
.A2(n_670),
.B(n_674),
.Y(n_700)
);

AOI21xp5_ASAP7_75t_SL g703 ( 
.A1(n_700),
.A2(n_684),
.B(n_674),
.Y(n_703)
);

NAND3xp33_ASAP7_75t_L g702 ( 
.A(n_701),
.B(n_684),
.C(n_689),
.Y(n_702)
);

AOI21xp5_ASAP7_75t_L g708 ( 
.A1(n_702),
.A2(n_703),
.B(n_705),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_SL g705 ( 
.A(n_695),
.B(n_661),
.Y(n_705)
);

MAJIxp5_ASAP7_75t_L g707 ( 
.A(n_706),
.B(n_698),
.C(n_673),
.Y(n_707)
);

MAJIxp5_ASAP7_75t_L g710 ( 
.A(n_707),
.B(n_709),
.C(n_4),
.Y(n_710)
);

MAJIxp5_ASAP7_75t_L g709 ( 
.A(n_704),
.B(n_698),
.C(n_676),
.Y(n_709)
);

AOI21xp5_ASAP7_75t_L g712 ( 
.A1(n_710),
.A2(n_711),
.B(n_5),
.Y(n_712)
);

NOR2xp33_ASAP7_75t_SL g711 ( 
.A(n_708),
.B(n_4),
.Y(n_711)
);

OAI21xp5_ASAP7_75t_L g713 ( 
.A1(n_712),
.A2(n_5),
.B(n_6),
.Y(n_713)
);

NOR2xp33_ASAP7_75t_L g714 ( 
.A(n_713),
.B(n_5),
.Y(n_714)
);


endmodule