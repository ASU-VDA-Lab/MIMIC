module fake_netlist_5_2280_n_929 (n_137, n_168, n_164, n_191, n_91, n_82, n_122, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_189, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_173, n_25, n_53, n_160, n_188, n_190, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_55, n_99, n_2, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_929);

input n_137;
input n_168;
input n_164;
input n_191;
input n_91;
input n_82;
input n_122;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_173;
input n_25;
input n_53;
input n_160;
input n_188;
input n_190;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_929;

wire n_924;
wire n_676;
wire n_294;
wire n_431;
wire n_318;
wire n_380;
wire n_419;
wire n_653;
wire n_611;
wire n_444;
wire n_642;
wire n_469;
wire n_615;
wire n_851;
wire n_194;
wire n_316;
wire n_785;
wire n_389;
wire n_855;
wire n_843;
wire n_549;
wire n_684;
wire n_850;
wire n_418;
wire n_248;
wire n_315;
wire n_268;
wire n_523;
wire n_451;
wire n_532;
wire n_705;
wire n_619;
wire n_408;
wire n_865;
wire n_913;
wire n_678;
wire n_664;
wire n_376;
wire n_697;
wire n_503;
wire n_235;
wire n_226;
wire n_605;
wire n_776;
wire n_928;
wire n_667;
wire n_515;
wire n_790;
wire n_353;
wire n_351;
wire n_367;
wire n_643;
wire n_620;
wire n_916;
wire n_452;
wire n_885;
wire n_397;
wire n_493;
wire n_525;
wire n_880;
wire n_703;
wire n_698;
wire n_483;
wire n_544;
wire n_683;
wire n_780;
wire n_649;
wire n_552;
wire n_547;
wire n_721;
wire n_841;
wire n_564;
wire n_467;
wire n_802;
wire n_423;
wire n_840;
wire n_284;
wire n_501;
wire n_245;
wire n_823;
wire n_725;
wire n_280;
wire n_744;
wire n_590;
wire n_629;
wire n_672;
wire n_873;
wire n_378;
wire n_551;
wire n_762;
wire n_581;
wire n_688;
wire n_382;
wire n_554;
wire n_800;
wire n_898;
wire n_254;
wire n_690;
wire n_583;
wire n_718;
wire n_671;
wire n_819;
wire n_302;
wire n_265;
wire n_526;
wire n_915;
wire n_719;
wire n_293;
wire n_372;
wire n_443;
wire n_244;
wire n_677;
wire n_859;
wire n_864;
wire n_821;
wire n_198;
wire n_714;
wire n_447;
wire n_247;
wire n_314;
wire n_368;
wire n_433;
wire n_604;
wire n_321;
wire n_292;
wire n_909;
wire n_625;
wire n_854;
wire n_621;
wire n_753;
wire n_455;
wire n_674;
wire n_417;
wire n_612;
wire n_212;
wire n_385;
wire n_516;
wire n_498;
wire n_788;
wire n_507;
wire n_497;
wire n_689;
wire n_738;
wire n_912;
wire n_606;
wire n_559;
wire n_275;
wire n_640;
wire n_252;
wire n_624;
wire n_825;
wire n_295;
wire n_330;
wire n_877;
wire n_508;
wire n_739;
wire n_506;
wire n_737;
wire n_610;
wire n_692;
wire n_755;
wire n_509;
wire n_568;
wire n_373;
wire n_820;
wire n_757;
wire n_307;
wire n_633;
wire n_439;
wire n_530;
wire n_556;
wire n_209;
wire n_259;
wire n_448;
wire n_758;
wire n_668;
wire n_733;
wire n_375;
wire n_301;
wire n_828;
wire n_779;
wire n_576;
wire n_804;
wire n_867;
wire n_537;
wire n_902;
wire n_587;
wire n_659;
wire n_492;
wire n_792;
wire n_563;
wire n_756;
wire n_878;
wire n_524;
wire n_399;
wire n_341;
wire n_204;
wire n_394;
wire n_250;
wire n_579;
wire n_741;
wire n_548;
wire n_543;
wire n_260;
wire n_812;
wire n_842;
wire n_298;
wire n_650;
wire n_320;
wire n_694;
wire n_518;
wire n_505;
wire n_286;
wire n_883;
wire n_282;
wire n_752;
wire n_331;
wire n_906;
wire n_905;
wire n_406;
wire n_519;
wire n_470;
wire n_908;
wire n_782;
wire n_919;
wire n_325;
wire n_449;
wire n_862;
wire n_900;
wire n_724;
wire n_856;
wire n_546;
wire n_760;
wire n_658;
wire n_281;
wire n_918;
wire n_240;
wire n_381;
wire n_220;
wire n_291;
wire n_231;
wire n_257;
wire n_390;
wire n_731;
wire n_456;
wire n_371;
wire n_481;
wire n_535;
wire n_709;
wire n_540;
wire n_317;
wire n_618;
wire n_896;
wire n_323;
wire n_569;
wire n_769;
wire n_195;
wire n_356;
wire n_227;
wire n_592;
wire n_920;
wire n_894;
wire n_271;
wire n_831;
wire n_826;
wire n_335;
wire n_886;
wire n_654;
wire n_370;
wire n_234;
wire n_343;
wire n_379;
wire n_428;
wire n_308;
wire n_267;
wire n_514;
wire n_457;
wire n_570;
wire n_833;
wire n_297;
wire n_853;
wire n_603;
wire n_225;
wire n_377;
wire n_751;
wire n_484;
wire n_775;
wire n_219;
wire n_442;
wire n_814;
wire n_192;
wire n_636;
wire n_786;
wire n_600;
wire n_660;
wire n_223;
wire n_392;
wire n_655;
wire n_704;
wire n_787;
wire n_264;
wire n_669;
wire n_472;
wire n_750;
wire n_742;
wire n_454;
wire n_387;
wire n_771;
wire n_374;
wire n_276;
wire n_339;
wire n_882;
wire n_243;
wire n_398;
wire n_396;
wire n_635;
wire n_347;
wire n_763;
wire n_550;
wire n_522;
wire n_255;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_662;
wire n_459;
wire n_646;
wire n_211;
wire n_218;
wire n_400;
wire n_436;
wire n_290;
wire n_580;
wire n_221;
wire n_622;
wire n_723;
wire n_386;
wire n_578;
wire n_926;
wire n_287;
wire n_344;
wire n_848;
wire n_555;
wire n_783;
wire n_473;
wire n_422;
wire n_475;
wire n_777;
wire n_661;
wire n_682;
wire n_415;
wire n_485;
wire n_496;
wire n_355;
wire n_849;
wire n_486;
wire n_670;
wire n_816;
wire n_336;
wire n_584;
wire n_681;
wire n_591;
wire n_922;
wire n_521;
wire n_614;
wire n_663;
wire n_845;
wire n_337;
wire n_430;
wire n_313;
wire n_631;
wire n_673;
wire n_837;
wire n_528;
wire n_479;
wire n_510;
wire n_216;
wire n_680;
wire n_395;
wire n_432;
wire n_553;
wire n_727;
wire n_839;
wire n_901;
wire n_311;
wire n_813;
wire n_830;
wire n_773;
wire n_208;
wire n_743;
wire n_328;
wire n_214;
wire n_801;
wire n_299;
wire n_303;
wire n_369;
wire n_675;
wire n_888;
wire n_296;
wire n_613;
wire n_871;
wire n_241;
wire n_637;
wire n_357;
wire n_875;
wire n_598;
wire n_685;
wire n_608;
wire n_446;
wire n_445;
wire n_749;
wire n_829;
wire n_858;
wire n_923;
wire n_772;
wire n_691;
wire n_881;
wire n_717;
wire n_468;
wire n_499;
wire n_213;
wire n_342;
wire n_517;
wire n_482;
wire n_588;
wire n_361;
wire n_464;
wire n_789;
wire n_363;
wire n_402;
wire n_413;
wire n_734;
wire n_638;
wire n_700;
wire n_197;
wire n_796;
wire n_573;
wire n_866;
wire n_236;
wire n_388;
wire n_761;
wire n_249;
wire n_903;
wire n_740;
wire n_304;
wire n_329;
wire n_203;
wire n_274;
wire n_577;
wire n_384;
wire n_582;
wire n_460;
wire n_889;
wire n_277;
wire n_477;
wire n_338;
wire n_571;
wire n_461;
wire n_333;
wire n_693;
wire n_309;
wire n_512;
wire n_836;
wire n_462;
wire n_322;
wire n_567;
wire n_258;
wire n_652;
wire n_778;
wire n_306;
wire n_907;
wire n_722;
wire n_458;
wire n_288;
wire n_770;
wire n_844;
wire n_201;
wire n_263;
wire n_471;
wire n_609;
wire n_852;
wire n_224;
wire n_228;
wire n_283;
wire n_383;
wire n_711;
wire n_781;
wire n_834;
wire n_474;
wire n_765;
wire n_542;
wire n_463;
wire n_488;
wire n_595;
wire n_736;
wire n_502;
wire n_892;
wire n_893;
wire n_891;
wire n_239;
wire n_466;
wire n_420;
wire n_630;
wire n_489;
wire n_632;
wire n_699;
wire n_617;
wire n_310;
wire n_593;
wire n_504;
wire n_511;
wire n_748;
wire n_586;
wire n_846;
wire n_874;
wire n_465;
wire n_838;
wire n_358;
wire n_362;
wire n_876;
wire n_332;
wire n_273;
wire n_585;
wire n_349;
wire n_270;
wire n_616;
wire n_230;
wire n_601;
wire n_279;
wire n_917;
wire n_253;
wire n_261;
wire n_289;
wire n_745;
wire n_627;
wire n_767;
wire n_206;
wire n_217;
wire n_440;
wire n_726;
wire n_478;
wire n_793;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_648;
wire n_312;
wire n_476;
wire n_818;
wire n_429;
wire n_861;
wire n_534;
wire n_884;
wire n_899;
wire n_345;
wire n_210;
wire n_494;
wire n_641;
wire n_628;
wire n_365;
wire n_774;
wire n_729;
wire n_730;
wire n_911;
wire n_557;
wire n_354;
wire n_607;
wire n_575;
wire n_480;
wire n_647;
wire n_237;
wire n_425;
wire n_513;
wire n_407;
wire n_527;
wire n_679;
wire n_707;
wire n_710;
wire n_795;
wire n_695;
wire n_832;
wire n_857;
wire n_560;
wire n_656;
wire n_340;
wire n_207;
wire n_561;
wire n_346;
wire n_393;
wire n_229;
wire n_487;
wire n_495;
wire n_602;
wire n_665;
wire n_574;
wire n_437;
wire n_453;
wire n_403;
wire n_421;
wire n_879;
wire n_720;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_863;
wire n_910;
wire n_490;
wire n_805;
wire n_326;
wire n_794;
wire n_768;
wire n_921;
wire n_233;
wire n_404;
wire n_686;
wire n_205;
wire n_366;
wire n_572;
wire n_712;
wire n_847;
wire n_754;
wire n_815;
wire n_246;
wire n_596;
wire n_410;
wire n_558;
wire n_708;
wire n_269;
wire n_529;
wire n_735;
wire n_702;
wire n_285;
wire n_822;
wire n_412;
wire n_232;
wire n_327;
wire n_657;
wire n_644;
wire n_728;
wire n_895;
wire n_202;
wire n_266;
wire n_272;
wire n_491;
wire n_427;
wire n_791;
wire n_732;
wire n_193;
wire n_251;
wire n_352;
wire n_566;
wire n_426;
wire n_520;
wire n_565;
wire n_808;
wire n_409;
wire n_797;
wire n_887;
wire n_589;
wire n_716;
wire n_597;
wire n_500;
wire n_562;
wire n_300;
wire n_651;
wire n_435;
wire n_809;
wire n_870;
wire n_334;
wire n_599;
wire n_766;
wire n_811;
wire n_541;
wire n_807;
wire n_391;
wire n_701;
wire n_434;
wire n_645;
wire n_539;
wire n_835;
wire n_538;
wire n_666;
wire n_262;
wire n_803;
wire n_868;
wire n_238;
wire n_639;
wire n_799;
wire n_914;
wire n_687;
wire n_715;
wire n_411;
wire n_414;
wire n_319;
wire n_364;
wire n_927;
wire n_536;
wire n_531;
wire n_242;
wire n_817;
wire n_872;
wire n_360;
wire n_594;
wire n_764;
wire n_200;
wire n_890;
wire n_759;
wire n_222;
wire n_438;
wire n_806;
wire n_713;
wire n_904;
wire n_869;
wire n_324;
wire n_810;
wire n_634;
wire n_416;
wire n_199;
wire n_827;
wire n_401;
wire n_348;
wire n_626;
wire n_925;
wire n_424;
wire n_706;
wire n_746;
wire n_256;
wire n_305;
wire n_533;
wire n_747;
wire n_278;
wire n_784;

BUFx10_ASAP7_75t_L g192 ( 
.A(n_2),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_109),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_43),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_50),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_136),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_120),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g198 ( 
.A(n_142),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_188),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_41),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_133),
.Y(n_201)
);

HB1xp67_ASAP7_75t_L g202 ( 
.A(n_73),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_110),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_91),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_38),
.Y(n_205)
);

INVx2_ASAP7_75t_SL g206 ( 
.A(n_107),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_1),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_90),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_156),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_44),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_99),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_158),
.Y(n_212)
);

BUFx3_ASAP7_75t_L g213 ( 
.A(n_162),
.Y(n_213)
);

INVx4_ASAP7_75t_R g214 ( 
.A(n_119),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_29),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_85),
.Y(n_216)
);

BUFx3_ASAP7_75t_L g217 ( 
.A(n_111),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_145),
.Y(n_218)
);

HB1xp67_ASAP7_75t_L g219 ( 
.A(n_166),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_79),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_139),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_12),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_67),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_74),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_175),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_39),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_189),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_17),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_70),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_24),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_3),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_40),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_49),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_32),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_160),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_76),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_97),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_163),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_131),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_57),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_121),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_130),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_71),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_143),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_75),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_171),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_66),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_146),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_184),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_69),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_64),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_34),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_2),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_134),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_20),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_141),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_11),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_21),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_42),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_168),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_26),
.Y(n_261)
);

BUFx10_ASAP7_75t_L g262 ( 
.A(n_53),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_62),
.Y(n_263)
);

BUFx5_ASAP7_75t_L g264 ( 
.A(n_116),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_61),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_123),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_77),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_10),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_88),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_105),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_149),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_129),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_132),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_89),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_92),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_190),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_72),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_101),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_15),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_125),
.Y(n_280)
);

INVx2_ASAP7_75t_SL g281 ( 
.A(n_103),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_159),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_187),
.Y(n_283)
);

CKINVDCx16_ASAP7_75t_R g284 ( 
.A(n_36),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_95),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_257),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_268),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_207),
.Y(n_288)
);

BUFx2_ASAP7_75t_SL g289 ( 
.A(n_203),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_195),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_193),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_194),
.Y(n_292)
);

HB1xp67_ASAP7_75t_L g293 ( 
.A(n_222),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_196),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_201),
.Y(n_295)
);

HB1xp67_ASAP7_75t_L g296 ( 
.A(n_228),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_205),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_253),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_210),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_230),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_197),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_215),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_199),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_200),
.Y(n_304)
);

INVxp67_ASAP7_75t_SL g305 ( 
.A(n_202),
.Y(n_305)
);

INVxp67_ASAP7_75t_SL g306 ( 
.A(n_219),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_204),
.Y(n_307)
);

INVxp67_ASAP7_75t_SL g308 ( 
.A(n_213),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_220),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_226),
.B(n_0),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_231),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_235),
.B(n_0),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_234),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_237),
.Y(n_314)
);

INVxp67_ASAP7_75t_SL g315 ( 
.A(n_217),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_255),
.Y(n_316)
);

INVxp67_ASAP7_75t_L g317 ( 
.A(n_192),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_264),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_208),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_209),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_247),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_259),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_263),
.Y(n_323)
);

INVxp33_ASAP7_75t_SL g324 ( 
.A(n_258),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_212),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_279),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_272),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_252),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_274),
.Y(n_329)
);

INVxp67_ASAP7_75t_SL g330 ( 
.A(n_278),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_282),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_283),
.Y(n_332)
);

INVxp33_ASAP7_75t_SL g333 ( 
.A(n_216),
.Y(n_333)
);

NOR2xp67_ASAP7_75t_L g334 ( 
.A(n_211),
.B(n_1),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_265),
.Y(n_335)
);

HB1xp67_ASAP7_75t_L g336 ( 
.A(n_198),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_240),
.Y(n_337)
);

INVxp67_ASAP7_75t_L g338 ( 
.A(n_192),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_243),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_206),
.B(n_3),
.Y(n_340)
);

NOR2xp67_ASAP7_75t_L g341 ( 
.A(n_245),
.B(n_4),
.Y(n_341)
);

INVxp67_ASAP7_75t_SL g342 ( 
.A(n_281),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_270),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_221),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_239),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_223),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_262),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_262),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_264),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_224),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_345),
.Y(n_351)
);

AND2x2_ASAP7_75t_L g352 ( 
.A(n_308),
.B(n_284),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_291),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_318),
.Y(n_354)
);

BUFx6f_ASAP7_75t_L g355 ( 
.A(n_318),
.Y(n_355)
);

OA21x2_ASAP7_75t_L g356 ( 
.A1(n_349),
.A2(n_227),
.B(n_225),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_292),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_295),
.Y(n_358)
);

AND2x6_ASAP7_75t_L g359 ( 
.A(n_349),
.B(n_218),
.Y(n_359)
);

BUFx6f_ASAP7_75t_L g360 ( 
.A(n_337),
.Y(n_360)
);

AND2x2_ASAP7_75t_L g361 ( 
.A(n_315),
.B(n_330),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_286),
.Y(n_362)
);

NAND2xp33_ASAP7_75t_L g363 ( 
.A(n_297),
.B(n_218),
.Y(n_363)
);

BUFx6f_ASAP7_75t_L g364 ( 
.A(n_339),
.Y(n_364)
);

NAND2xp33_ASAP7_75t_SL g365 ( 
.A(n_347),
.B(n_348),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_299),
.Y(n_366)
);

BUFx6f_ASAP7_75t_L g367 ( 
.A(n_302),
.Y(n_367)
);

INVx3_ASAP7_75t_L g368 ( 
.A(n_309),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_313),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_314),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_321),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_322),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_323),
.Y(n_373)
);

OA21x2_ASAP7_75t_L g374 ( 
.A1(n_327),
.A2(n_232),
.B(n_229),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_329),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_324),
.B(n_233),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_290),
.B(n_238),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_331),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_332),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_287),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_342),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_334),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_341),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_340),
.Y(n_384)
);

NAND2xp33_ASAP7_75t_SL g385 ( 
.A(n_347),
.B(n_218),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_310),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_294),
.B(n_285),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_312),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_293),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_296),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_SL g391 ( 
.A(n_301),
.B(n_218),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_303),
.Y(n_392)
);

AND2x4_ASAP7_75t_L g393 ( 
.A(n_305),
.B(n_239),
.Y(n_393)
);

CKINVDCx16_ASAP7_75t_R g394 ( 
.A(n_328),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_306),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_304),
.Y(n_396)
);

INVxp67_ASAP7_75t_L g397 ( 
.A(n_336),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_SL g398 ( 
.A(n_307),
.B(n_236),
.Y(n_398)
);

BUFx3_ASAP7_75t_L g399 ( 
.A(n_319),
.Y(n_399)
);

HB1xp67_ASAP7_75t_L g400 ( 
.A(n_317),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_320),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_325),
.B(n_280),
.Y(n_402)
);

INVx1_ASAP7_75t_SL g403 ( 
.A(n_328),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_344),
.Y(n_404)
);

BUFx2_ASAP7_75t_L g405 ( 
.A(n_300),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_333),
.B(n_241),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_346),
.Y(n_407)
);

BUFx6f_ASAP7_75t_L g408 ( 
.A(n_355),
.Y(n_408)
);

AND2x4_ASAP7_75t_L g409 ( 
.A(n_393),
.B(n_350),
.Y(n_409)
);

AND2x2_ASAP7_75t_L g410 ( 
.A(n_352),
.B(n_289),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_354),
.B(n_264),
.Y(n_411)
);

OR2x2_ASAP7_75t_L g412 ( 
.A(n_352),
.B(n_338),
.Y(n_412)
);

INVxp67_ASAP7_75t_SL g413 ( 
.A(n_362),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_381),
.B(n_300),
.Y(n_414)
);

INVx4_ASAP7_75t_L g415 ( 
.A(n_355),
.Y(n_415)
);

AND2x2_ASAP7_75t_SL g416 ( 
.A(n_394),
.B(n_236),
.Y(n_416)
);

INVx6_ASAP7_75t_L g417 ( 
.A(n_393),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_395),
.B(n_311),
.Y(n_418)
);

INVx4_ASAP7_75t_L g419 ( 
.A(n_355),
.Y(n_419)
);

AND2x6_ASAP7_75t_L g420 ( 
.A(n_392),
.B(n_236),
.Y(n_420)
);

INVx4_ASAP7_75t_L g421 ( 
.A(n_355),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_353),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_357),
.Y(n_423)
);

INVx4_ASAP7_75t_L g424 ( 
.A(n_355),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_358),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_370),
.Y(n_426)
);

INVx3_ASAP7_75t_L g427 ( 
.A(n_367),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_371),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_SL g429 ( 
.A(n_393),
.B(n_236),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_372),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_378),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_388),
.B(n_386),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_379),
.Y(n_433)
);

INVxp67_ASAP7_75t_L g434 ( 
.A(n_400),
.Y(n_434)
);

AND2x4_ASAP7_75t_L g435 ( 
.A(n_392),
.B(n_407),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_362),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_367),
.Y(n_437)
);

OR2x2_ASAP7_75t_L g438 ( 
.A(n_389),
.B(n_242),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_360),
.Y(n_439)
);

BUFx4f_ASAP7_75t_L g440 ( 
.A(n_404),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_367),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_360),
.Y(n_442)
);

BUFx6f_ASAP7_75t_L g443 ( 
.A(n_367),
.Y(n_443)
);

INVx8_ASAP7_75t_L g444 ( 
.A(n_361),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_367),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_360),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_366),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_360),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_399),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_366),
.Y(n_450)
);

OR2x2_ASAP7_75t_L g451 ( 
.A(n_390),
.B(n_244),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_360),
.Y(n_452)
);

AND2x2_ASAP7_75t_L g453 ( 
.A(n_361),
.B(n_348),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_386),
.B(n_311),
.Y(n_454)
);

INVx1_ASAP7_75t_SL g455 ( 
.A(n_403),
.Y(n_455)
);

AND3x1_ASAP7_75t_L g456 ( 
.A(n_384),
.B(n_326),
.C(n_316),
.Y(n_456)
);

INVx4_ASAP7_75t_L g457 ( 
.A(n_364),
.Y(n_457)
);

BUFx3_ASAP7_75t_L g458 ( 
.A(n_399),
.Y(n_458)
);

AND2x4_ASAP7_75t_L g459 ( 
.A(n_407),
.B(n_404),
.Y(n_459)
);

INVx2_ASAP7_75t_SL g460 ( 
.A(n_391),
.Y(n_460)
);

HB1xp67_ASAP7_75t_L g461 ( 
.A(n_382),
.Y(n_461)
);

INVx4_ASAP7_75t_L g462 ( 
.A(n_364),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_369),
.Y(n_463)
);

BUFx2_ASAP7_75t_L g464 ( 
.A(n_397),
.Y(n_464)
);

AND2x4_ASAP7_75t_L g465 ( 
.A(n_396),
.B(n_246),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_SL g466 ( 
.A(n_391),
.B(n_267),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_364),
.Y(n_467)
);

INVx6_ASAP7_75t_L g468 ( 
.A(n_364),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_369),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_SL g470 ( 
.A(n_398),
.B(n_267),
.Y(n_470)
);

INVx4_ASAP7_75t_L g471 ( 
.A(n_364),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_373),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_373),
.Y(n_473)
);

INVx5_ASAP7_75t_L g474 ( 
.A(n_359),
.Y(n_474)
);

BUFx6f_ASAP7_75t_L g475 ( 
.A(n_354),
.Y(n_475)
);

BUFx3_ASAP7_75t_L g476 ( 
.A(n_368),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_375),
.Y(n_477)
);

AO22x2_ASAP7_75t_L g478 ( 
.A1(n_460),
.A2(n_398),
.B1(n_401),
.B2(n_383),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_436),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_422),
.Y(n_480)
);

NAND2xp33_ASAP7_75t_L g481 ( 
.A(n_444),
.B(n_377),
.Y(n_481)
);

AO22x2_ASAP7_75t_L g482 ( 
.A1(n_412),
.A2(n_385),
.B1(n_288),
.B2(n_298),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_432),
.B(n_406),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_423),
.Y(n_484)
);

AND2x2_ASAP7_75t_L g485 ( 
.A(n_454),
.B(n_376),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_475),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_425),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_432),
.B(n_417),
.Y(n_488)
);

AO22x2_ASAP7_75t_L g489 ( 
.A1(n_453),
.A2(n_385),
.B1(n_288),
.B2(n_298),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_426),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_417),
.B(n_387),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_428),
.Y(n_492)
);

AND2x2_ASAP7_75t_L g493 ( 
.A(n_454),
.B(n_335),
.Y(n_493)
);

AND2x4_ASAP7_75t_L g494 ( 
.A(n_476),
.B(n_380),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_417),
.B(n_402),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_430),
.Y(n_496)
);

INVxp67_ASAP7_75t_L g497 ( 
.A(n_418),
.Y(n_497)
);

AO22x2_ASAP7_75t_L g498 ( 
.A1(n_466),
.A2(n_365),
.B1(n_316),
.B2(n_326),
.Y(n_498)
);

AOI22xp5_ASAP7_75t_L g499 ( 
.A1(n_435),
.A2(n_374),
.B1(n_356),
.B2(n_343),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_431),
.Y(n_500)
);

OR2x6_ASAP7_75t_L g501 ( 
.A(n_458),
.B(n_405),
.Y(n_501)
);

AOI22xp5_ASAP7_75t_L g502 ( 
.A1(n_435),
.A2(n_374),
.B1(n_356),
.B2(n_343),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_413),
.B(n_356),
.Y(n_503)
);

AND2x2_ASAP7_75t_SL g504 ( 
.A(n_456),
.B(n_405),
.Y(n_504)
);

OR2x2_ASAP7_75t_SL g505 ( 
.A(n_438),
.B(n_365),
.Y(n_505)
);

OAI221xp5_ASAP7_75t_L g506 ( 
.A1(n_413),
.A2(n_375),
.B1(n_380),
.B2(n_368),
.C(n_351),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_444),
.B(n_433),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_447),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_450),
.Y(n_509)
);

AOI22xp5_ASAP7_75t_L g510 ( 
.A1(n_459),
.A2(n_374),
.B1(n_266),
.B2(n_248),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_434),
.B(n_414),
.Y(n_511)
);

AO22x2_ASAP7_75t_L g512 ( 
.A1(n_466),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_512)
);

BUFx3_ASAP7_75t_L g513 ( 
.A(n_459),
.Y(n_513)
);

INVxp67_ASAP7_75t_L g514 ( 
.A(n_418),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_463),
.Y(n_515)
);

OAI221xp5_ASAP7_75t_L g516 ( 
.A1(n_461),
.A2(n_368),
.B1(n_351),
.B2(n_249),
.C(n_277),
.Y(n_516)
);

INVxp67_ASAP7_75t_L g517 ( 
.A(n_464),
.Y(n_517)
);

AO22x2_ASAP7_75t_L g518 ( 
.A1(n_470),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_518)
);

AO22x2_ASAP7_75t_L g519 ( 
.A1(n_470),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_519)
);

NAND2x1p5_ASAP7_75t_L g520 ( 
.A(n_410),
.B(n_267),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_469),
.Y(n_521)
);

NAND2x1p5_ASAP7_75t_L g522 ( 
.A(n_409),
.B(n_267),
.Y(n_522)
);

INVx1_ASAP7_75t_SL g523 ( 
.A(n_455),
.Y(n_523)
);

OAI221xp5_ASAP7_75t_L g524 ( 
.A1(n_461),
.A2(n_261),
.B1(n_276),
.B2(n_275),
.C(n_273),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_475),
.Y(n_525)
);

CKINVDCx20_ASAP7_75t_R g526 ( 
.A(n_449),
.Y(n_526)
);

NAND3xp33_ASAP7_75t_L g527 ( 
.A(n_414),
.B(n_451),
.C(n_456),
.Y(n_527)
);

AND2x2_ASAP7_75t_L g528 ( 
.A(n_409),
.B(n_250),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_444),
.B(n_359),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_472),
.Y(n_530)
);

OR2x2_ASAP7_75t_L g531 ( 
.A(n_455),
.B(n_8),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_475),
.Y(n_532)
);

AOI22xp5_ASAP7_75t_L g533 ( 
.A1(n_440),
.A2(n_260),
.B1(n_256),
.B2(n_271),
.Y(n_533)
);

INVxp67_ASAP7_75t_L g534 ( 
.A(n_434),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_429),
.B(n_359),
.Y(n_535)
);

OAI22xp5_ASAP7_75t_SL g536 ( 
.A1(n_416),
.A2(n_251),
.B1(n_254),
.B2(n_269),
.Y(n_536)
);

NOR2xp67_ASAP7_75t_L g537 ( 
.A(n_465),
.B(n_25),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_473),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_477),
.Y(n_539)
);

AND2x4_ASAP7_75t_L g540 ( 
.A(n_465),
.B(n_239),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_429),
.B(n_359),
.Y(n_541)
);

INVx4_ASAP7_75t_L g542 ( 
.A(n_440),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_411),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_408),
.Y(n_544)
);

OAI221xp5_ASAP7_75t_L g545 ( 
.A1(n_411),
.A2(n_363),
.B1(n_214),
.B2(n_264),
.C(n_12),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_437),
.Y(n_546)
);

HAxp5_ASAP7_75t_SL g547 ( 
.A(n_441),
.B(n_9),
.CON(n_547),
.SN(n_547)
);

AO22x2_ASAP7_75t_L g548 ( 
.A1(n_445),
.A2(n_10),
.B1(n_11),
.B2(n_13),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_SL g549 ( 
.A(n_483),
.B(n_474),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_SL g550 ( 
.A(n_542),
.B(n_474),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_SL g551 ( 
.A(n_485),
.B(n_474),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_SL g552 ( 
.A(n_497),
.B(n_474),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_SL g553 ( 
.A(n_514),
.B(n_443),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_SL g554 ( 
.A(n_513),
.B(n_443),
.Y(n_554)
);

NAND2xp33_ASAP7_75t_SL g555 ( 
.A(n_536),
.B(n_443),
.Y(n_555)
);

AND2x4_ASAP7_75t_L g556 ( 
.A(n_494),
.B(n_480),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_SL g557 ( 
.A(n_511),
.B(n_408),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_488),
.B(n_427),
.Y(n_558)
);

AND2x4_ASAP7_75t_L g559 ( 
.A(n_494),
.B(n_484),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_SL g560 ( 
.A(n_523),
.B(n_408),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_SL g561 ( 
.A(n_507),
.B(n_427),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_543),
.B(n_439),
.Y(n_562)
);

AND2x4_ASAP7_75t_L g563 ( 
.A(n_487),
.B(n_442),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_SL g564 ( 
.A(n_527),
.B(n_446),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_SL g565 ( 
.A(n_534),
.B(n_448),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_491),
.B(n_452),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_SL g567 ( 
.A(n_540),
.B(n_467),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_SL g568 ( 
.A(n_540),
.B(n_457),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_SL g569 ( 
.A(n_517),
.B(n_457),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_SL g570 ( 
.A(n_537),
.B(n_471),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_SL g571 ( 
.A(n_495),
.B(n_471),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_SL g572 ( 
.A(n_490),
.B(n_462),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_SL g573 ( 
.A(n_492),
.B(n_462),
.Y(n_573)
);

AND2x2_ASAP7_75t_L g574 ( 
.A(n_493),
.B(n_468),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_SL g575 ( 
.A(n_496),
.B(n_415),
.Y(n_575)
);

NAND2xp33_ASAP7_75t_SL g576 ( 
.A(n_528),
.B(n_415),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_SL g577 ( 
.A(n_500),
.B(n_419),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_SL g578 ( 
.A(n_479),
.B(n_520),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_478),
.B(n_419),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_SL g580 ( 
.A(n_504),
.B(n_421),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_SL g581 ( 
.A(n_510),
.B(n_421),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_SL g582 ( 
.A(n_522),
.B(n_424),
.Y(n_582)
);

NAND2xp33_ASAP7_75t_SL g583 ( 
.A(n_526),
.B(n_424),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_SL g584 ( 
.A(n_508),
.B(n_264),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_SL g585 ( 
.A(n_509),
.B(n_264),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_SL g586 ( 
.A(n_515),
.B(n_420),
.Y(n_586)
);

NAND2xp33_ASAP7_75t_SL g587 ( 
.A(n_531),
.B(n_547),
.Y(n_587)
);

AND2x2_ASAP7_75t_L g588 ( 
.A(n_501),
.B(n_468),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_SL g589 ( 
.A(n_521),
.B(n_420),
.Y(n_589)
);

NAND2xp33_ASAP7_75t_SL g590 ( 
.A(n_529),
.B(n_420),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_SL g591 ( 
.A(n_530),
.B(n_420),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_SL g592 ( 
.A(n_538),
.B(n_468),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_SL g593 ( 
.A(n_533),
.B(n_27),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_SL g594 ( 
.A(n_499),
.B(n_28),
.Y(n_594)
);

NAND2xp33_ASAP7_75t_SL g595 ( 
.A(n_503),
.B(n_13),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_SL g596 ( 
.A(n_502),
.B(n_30),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_SL g597 ( 
.A(n_539),
.B(n_31),
.Y(n_597)
);

NAND2xp33_ASAP7_75t_SL g598 ( 
.A(n_535),
.B(n_541),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_478),
.B(n_359),
.Y(n_599)
);

XNOR2xp5_ASAP7_75t_SL g600 ( 
.A(n_482),
.B(n_14),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_SL g601 ( 
.A(n_486),
.B(n_33),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_SL g602 ( 
.A(n_525),
.B(n_35),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_532),
.B(n_359),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_SL g604 ( 
.A(n_546),
.B(n_37),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_SL g605 ( 
.A(n_544),
.B(n_45),
.Y(n_605)
);

NAND2xp33_ASAP7_75t_SL g606 ( 
.A(n_505),
.B(n_14),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_SL g607 ( 
.A(n_516),
.B(n_46),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_SL g608 ( 
.A(n_481),
.B(n_524),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_583),
.Y(n_609)
);

AO31x2_ASAP7_75t_L g610 ( 
.A1(n_579),
.A2(n_506),
.A3(n_545),
.B(n_519),
.Y(n_610)
);

AOI21xp5_ASAP7_75t_L g611 ( 
.A1(n_570),
.A2(n_363),
.B(n_501),
.Y(n_611)
);

AO31x2_ASAP7_75t_L g612 ( 
.A1(n_599),
.A2(n_519),
.A3(n_518),
.B(n_512),
.Y(n_612)
);

OAI21x1_ASAP7_75t_L g613 ( 
.A1(n_562),
.A2(n_512),
.B(n_518),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_566),
.B(n_558),
.Y(n_614)
);

OAI22xp5_ASAP7_75t_L g615 ( 
.A1(n_594),
.A2(n_548),
.B1(n_498),
.B2(n_482),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_SL g616 ( 
.A(n_556),
.B(n_489),
.Y(n_616)
);

HB1xp67_ASAP7_75t_L g617 ( 
.A(n_556),
.Y(n_617)
);

OA21x2_ASAP7_75t_L g618 ( 
.A1(n_564),
.A2(n_548),
.B(n_498),
.Y(n_618)
);

AO21x2_ASAP7_75t_L g619 ( 
.A1(n_596),
.A2(n_489),
.B(n_114),
.Y(n_619)
);

OAI22x1_ASAP7_75t_L g620 ( 
.A1(n_600),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_L g621 ( 
.A(n_587),
.B(n_16),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_L g622 ( 
.A(n_574),
.B(n_18),
.Y(n_622)
);

AOI21xp5_ASAP7_75t_L g623 ( 
.A1(n_571),
.A2(n_581),
.B(n_568),
.Y(n_623)
);

AND2x2_ASAP7_75t_L g624 ( 
.A(n_559),
.B(n_588),
.Y(n_624)
);

AND2x2_ASAP7_75t_L g625 ( 
.A(n_559),
.B(n_18),
.Y(n_625)
);

BUFx2_ASAP7_75t_L g626 ( 
.A(n_606),
.Y(n_626)
);

OAI21x1_ASAP7_75t_SL g627 ( 
.A1(n_603),
.A2(n_117),
.B(n_186),
.Y(n_627)
);

INVx2_ASAP7_75t_SL g628 ( 
.A(n_560),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_563),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_557),
.B(n_47),
.Y(n_630)
);

INVxp67_ASAP7_75t_SL g631 ( 
.A(n_563),
.Y(n_631)
);

OAI21x1_ASAP7_75t_L g632 ( 
.A1(n_561),
.A2(n_115),
.B(n_185),
.Y(n_632)
);

OAI21x1_ASAP7_75t_L g633 ( 
.A1(n_549),
.A2(n_113),
.B(n_183),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_608),
.B(n_48),
.Y(n_634)
);

BUFx2_ASAP7_75t_L g635 ( 
.A(n_555),
.Y(n_635)
);

OAI21x1_ASAP7_75t_L g636 ( 
.A1(n_551),
.A2(n_118),
.B(n_182),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_553),
.B(n_51),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_567),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_580),
.B(n_52),
.Y(n_639)
);

AOI21xp5_ASAP7_75t_L g640 ( 
.A1(n_598),
.A2(n_122),
.B(n_181),
.Y(n_640)
);

AOI21xp5_ASAP7_75t_L g641 ( 
.A1(n_582),
.A2(n_112),
.B(n_180),
.Y(n_641)
);

AO31x2_ASAP7_75t_L g642 ( 
.A1(n_595),
.A2(n_19),
.A3(n_20),
.B(n_21),
.Y(n_642)
);

OAI21xp5_ASAP7_75t_L g643 ( 
.A1(n_607),
.A2(n_124),
.B(n_179),
.Y(n_643)
);

OAI21xp33_ASAP7_75t_L g644 ( 
.A1(n_565),
.A2(n_19),
.B(n_22),
.Y(n_644)
);

OAI21xp5_ASAP7_75t_L g645 ( 
.A1(n_593),
.A2(n_584),
.B(n_585),
.Y(n_645)
);

BUFx2_ASAP7_75t_L g646 ( 
.A(n_576),
.Y(n_646)
);

OAI21x1_ASAP7_75t_L g647 ( 
.A1(n_575),
.A2(n_108),
.B(n_178),
.Y(n_647)
);

OAI21x1_ASAP7_75t_L g648 ( 
.A1(n_577),
.A2(n_106),
.B(n_177),
.Y(n_648)
);

OAI21x1_ASAP7_75t_L g649 ( 
.A1(n_572),
.A2(n_104),
.B(n_176),
.Y(n_649)
);

BUFx3_ASAP7_75t_L g650 ( 
.A(n_569),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_552),
.B(n_102),
.Y(n_651)
);

BUFx6f_ASAP7_75t_L g652 ( 
.A(n_554),
.Y(n_652)
);

AOI31xp67_ASAP7_75t_L g653 ( 
.A1(n_586),
.A2(n_126),
.A3(n_174),
.B(n_173),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_592),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_578),
.B(n_98),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_573),
.Y(n_656)
);

OAI21xp5_ASAP7_75t_L g657 ( 
.A1(n_590),
.A2(n_100),
.B(n_172),
.Y(n_657)
);

OAI21x1_ASAP7_75t_L g658 ( 
.A1(n_550),
.A2(n_96),
.B(n_170),
.Y(n_658)
);

AOI21xp5_ASAP7_75t_SL g659 ( 
.A1(n_604),
.A2(n_94),
.B(n_169),
.Y(n_659)
);

AOI22xp33_ASAP7_75t_L g660 ( 
.A1(n_621),
.A2(n_597),
.B1(n_605),
.B2(n_601),
.Y(n_660)
);

OR2x2_ASAP7_75t_L g661 ( 
.A(n_617),
.B(n_591),
.Y(n_661)
);

OR2x2_ASAP7_75t_L g662 ( 
.A(n_624),
.B(n_589),
.Y(n_662)
);

INVx3_ASAP7_75t_L g663 ( 
.A(n_636),
.Y(n_663)
);

AND2x4_ASAP7_75t_L g664 ( 
.A(n_629),
.B(n_602),
.Y(n_664)
);

AOI22xp5_ASAP7_75t_L g665 ( 
.A1(n_635),
.A2(n_22),
.B1(n_23),
.B2(n_24),
.Y(n_665)
);

AOI221xp5_ASAP7_75t_L g666 ( 
.A1(n_615),
.A2(n_23),
.B1(n_54),
.B2(n_55),
.C(n_56),
.Y(n_666)
);

AND2x6_ASAP7_75t_L g667 ( 
.A(n_634),
.B(n_58),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_654),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_638),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_653),
.Y(n_670)
);

OAI21x1_ASAP7_75t_L g671 ( 
.A1(n_632),
.A2(n_59),
.B(n_60),
.Y(n_671)
);

OAI22xp5_ASAP7_75t_L g672 ( 
.A1(n_631),
.A2(n_63),
.B1(n_65),
.B2(n_68),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_628),
.Y(n_673)
);

OAI21x1_ASAP7_75t_L g674 ( 
.A1(n_633),
.A2(n_623),
.B(n_647),
.Y(n_674)
);

AO31x2_ASAP7_75t_L g675 ( 
.A1(n_615),
.A2(n_78),
.A3(n_80),
.B(n_81),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_614),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_652),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_648),
.Y(n_678)
);

OA21x2_ASAP7_75t_L g679 ( 
.A1(n_657),
.A2(n_82),
.B(n_83),
.Y(n_679)
);

AO31x2_ASAP7_75t_L g680 ( 
.A1(n_634),
.A2(n_84),
.A3(n_86),
.B(n_87),
.Y(n_680)
);

INVx2_ASAP7_75t_SL g681 ( 
.A(n_652),
.Y(n_681)
);

OAI21x1_ASAP7_75t_L g682 ( 
.A1(n_649),
.A2(n_93),
.B(n_127),
.Y(n_682)
);

NOR2xp33_ASAP7_75t_L g683 ( 
.A(n_626),
.B(n_128),
.Y(n_683)
);

OA21x2_ASAP7_75t_L g684 ( 
.A1(n_657),
.A2(n_135),
.B(n_137),
.Y(n_684)
);

AOI22xp33_ASAP7_75t_L g685 ( 
.A1(n_644),
.A2(n_138),
.B1(n_140),
.B2(n_144),
.Y(n_685)
);

OR2x2_ASAP7_75t_L g686 ( 
.A(n_616),
.B(n_147),
.Y(n_686)
);

OAI21x1_ASAP7_75t_L g687 ( 
.A1(n_658),
.A2(n_148),
.B(n_150),
.Y(n_687)
);

OAI21x1_ASAP7_75t_L g688 ( 
.A1(n_640),
.A2(n_151),
.B(n_152),
.Y(n_688)
);

BUFx6f_ASAP7_75t_L g689 ( 
.A(n_652),
.Y(n_689)
);

NAND2x1p5_ASAP7_75t_L g690 ( 
.A(n_646),
.B(n_153),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_625),
.Y(n_691)
);

OAI21xp5_ASAP7_75t_L g692 ( 
.A1(n_630),
.A2(n_154),
.B(n_155),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_613),
.Y(n_693)
);

AND2x2_ASAP7_75t_L g694 ( 
.A(n_622),
.B(n_157),
.Y(n_694)
);

OAI21x1_ASAP7_75t_L g695 ( 
.A1(n_640),
.A2(n_161),
.B(n_164),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_655),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_656),
.Y(n_697)
);

OA21x2_ASAP7_75t_L g698 ( 
.A1(n_643),
.A2(n_165),
.B(n_167),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_610),
.Y(n_699)
);

BUFx2_ASAP7_75t_L g700 ( 
.A(n_609),
.Y(n_700)
);

OAI21x1_ASAP7_75t_L g701 ( 
.A1(n_674),
.A2(n_627),
.B(n_643),
.Y(n_701)
);

HB1xp67_ASAP7_75t_L g702 ( 
.A(n_691),
.Y(n_702)
);

OR2x2_ASAP7_75t_L g703 ( 
.A(n_699),
.B(n_612),
.Y(n_703)
);

AND2x2_ASAP7_75t_L g704 ( 
.A(n_676),
.B(n_612),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_693),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_676),
.Y(n_706)
);

HB1xp67_ASAP7_75t_L g707 ( 
.A(n_689),
.Y(n_707)
);

OAI22xp5_ASAP7_75t_L g708 ( 
.A1(n_696),
.A2(n_650),
.B1(n_639),
.B2(n_637),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_699),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_697),
.Y(n_710)
);

AND2x2_ASAP7_75t_L g711 ( 
.A(n_697),
.B(n_612),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_669),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_668),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_675),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_675),
.Y(n_715)
);

INVxp67_ASAP7_75t_L g716 ( 
.A(n_700),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_675),
.Y(n_717)
);

NAND2x1_ASAP7_75t_L g718 ( 
.A(n_663),
.B(n_659),
.Y(n_718)
);

BUFx10_ASAP7_75t_L g719 ( 
.A(n_683),
.Y(n_719)
);

NOR2xp33_ASAP7_75t_L g720 ( 
.A(n_683),
.B(n_639),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_675),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_661),
.Y(n_722)
);

BUFx2_ASAP7_75t_L g723 ( 
.A(n_689),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_677),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_673),
.Y(n_725)
);

HB1xp67_ASAP7_75t_L g726 ( 
.A(n_689),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_680),
.Y(n_727)
);

HB1xp67_ASAP7_75t_L g728 ( 
.A(n_689),
.Y(n_728)
);

INVxp67_ASAP7_75t_L g729 ( 
.A(n_681),
.Y(n_729)
);

AOI21x1_ASAP7_75t_L g730 ( 
.A1(n_670),
.A2(n_630),
.B(n_611),
.Y(n_730)
);

AND2x2_ASAP7_75t_L g731 ( 
.A(n_694),
.B(n_618),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_680),
.Y(n_732)
);

INVx3_ASAP7_75t_L g733 ( 
.A(n_687),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_678),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_688),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_680),
.Y(n_736)
);

AOI22xp33_ASAP7_75t_L g737 ( 
.A1(n_666),
.A2(n_619),
.B1(n_618),
.B2(n_620),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_688),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_680),
.Y(n_739)
);

CKINVDCx16_ASAP7_75t_R g740 ( 
.A(n_681),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_679),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_695),
.Y(n_742)
);

INVx3_ASAP7_75t_L g743 ( 
.A(n_687),
.Y(n_743)
);

AND2x2_ASAP7_75t_L g744 ( 
.A(n_690),
.B(n_619),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_679),
.Y(n_745)
);

HB1xp67_ASAP7_75t_L g746 ( 
.A(n_662),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_679),
.Y(n_747)
);

HB1xp67_ASAP7_75t_L g748 ( 
.A(n_664),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_664),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_695),
.Y(n_750)
);

NOR2xp33_ASAP7_75t_R g751 ( 
.A(n_740),
.B(n_686),
.Y(n_751)
);

NAND2xp33_ASAP7_75t_R g752 ( 
.A(n_720),
.B(n_684),
.Y(n_752)
);

INVxp33_ASAP7_75t_L g753 ( 
.A(n_746),
.Y(n_753)
);

NAND2xp33_ASAP7_75t_R g754 ( 
.A(n_744),
.B(n_684),
.Y(n_754)
);

NAND2xp33_ASAP7_75t_R g755 ( 
.A(n_744),
.B(n_684),
.Y(n_755)
);

BUFx3_ASAP7_75t_L g756 ( 
.A(n_723),
.Y(n_756)
);

AND2x4_ASAP7_75t_L g757 ( 
.A(n_723),
.B(n_664),
.Y(n_757)
);

AND2x4_ASAP7_75t_L g758 ( 
.A(n_749),
.B(n_748),
.Y(n_758)
);

AND2x4_ASAP7_75t_L g759 ( 
.A(n_716),
.B(n_651),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_722),
.B(n_665),
.Y(n_760)
);

NOR2xp33_ASAP7_75t_R g761 ( 
.A(n_719),
.B(n_667),
.Y(n_761)
);

NAND2xp33_ASAP7_75t_R g762 ( 
.A(n_731),
.B(n_698),
.Y(n_762)
);

BUFx3_ASAP7_75t_L g763 ( 
.A(n_725),
.Y(n_763)
);

NAND2xp33_ASAP7_75t_R g764 ( 
.A(n_731),
.B(n_698),
.Y(n_764)
);

NOR2xp33_ASAP7_75t_R g765 ( 
.A(n_719),
.B(n_667),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_713),
.Y(n_766)
);

NOR2xp33_ASAP7_75t_R g767 ( 
.A(n_719),
.B(n_667),
.Y(n_767)
);

NOR2xp33_ASAP7_75t_R g768 ( 
.A(n_707),
.B(n_667),
.Y(n_768)
);

NOR2xp33_ASAP7_75t_R g769 ( 
.A(n_726),
.B(n_667),
.Y(n_769)
);

CKINVDCx16_ASAP7_75t_R g770 ( 
.A(n_728),
.Y(n_770)
);

OR2x6_ASAP7_75t_L g771 ( 
.A(n_713),
.B(n_690),
.Y(n_771)
);

INVxp67_ASAP7_75t_L g772 ( 
.A(n_702),
.Y(n_772)
);

OR2x2_ASAP7_75t_L g773 ( 
.A(n_704),
.B(n_711),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_706),
.B(n_642),
.Y(n_774)
);

AND2x4_ASAP7_75t_L g775 ( 
.A(n_729),
.B(n_651),
.Y(n_775)
);

INVxp67_ASAP7_75t_L g776 ( 
.A(n_724),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_706),
.B(n_642),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_705),
.Y(n_778)
);

OR2x6_ASAP7_75t_L g779 ( 
.A(n_710),
.B(n_672),
.Y(n_779)
);

NAND2xp33_ASAP7_75t_R g780 ( 
.A(n_711),
.B(n_698),
.Y(n_780)
);

BUFx3_ASAP7_75t_L g781 ( 
.A(n_712),
.Y(n_781)
);

OR2x2_ASAP7_75t_L g782 ( 
.A(n_704),
.B(n_642),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_705),
.Y(n_783)
);

NAND2xp33_ASAP7_75t_R g784 ( 
.A(n_712),
.B(n_655),
.Y(n_784)
);

INVxp67_ASAP7_75t_L g785 ( 
.A(n_710),
.Y(n_785)
);

BUFx10_ASAP7_75t_L g786 ( 
.A(n_727),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_709),
.Y(n_787)
);

NOR2xp33_ASAP7_75t_R g788 ( 
.A(n_703),
.B(n_663),
.Y(n_788)
);

INVxp67_ASAP7_75t_L g789 ( 
.A(n_703),
.Y(n_789)
);

NOR2xp33_ASAP7_75t_L g790 ( 
.A(n_708),
.B(n_692),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_778),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_783),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_787),
.Y(n_793)
);

INVxp67_ASAP7_75t_SL g794 ( 
.A(n_772),
.Y(n_794)
);

HB1xp67_ASAP7_75t_L g795 ( 
.A(n_781),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_789),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_774),
.Y(n_797)
);

AND2x2_ASAP7_75t_L g798 ( 
.A(n_773),
.B(n_715),
.Y(n_798)
);

AND2x4_ASAP7_75t_L g799 ( 
.A(n_758),
.B(n_782),
.Y(n_799)
);

OR2x2_ASAP7_75t_L g800 ( 
.A(n_777),
.B(n_727),
.Y(n_800)
);

OR2x2_ASAP7_75t_L g801 ( 
.A(n_776),
.B(n_732),
.Y(n_801)
);

HB1xp67_ASAP7_75t_L g802 ( 
.A(n_763),
.Y(n_802)
);

AND2x2_ASAP7_75t_L g803 ( 
.A(n_766),
.B(n_721),
.Y(n_803)
);

AND2x2_ASAP7_75t_L g804 ( 
.A(n_785),
.B(n_721),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_786),
.Y(n_805)
);

AND2x2_ASAP7_75t_L g806 ( 
.A(n_758),
.B(n_715),
.Y(n_806)
);

NAND3xp33_ASAP7_75t_L g807 ( 
.A(n_790),
.B(n_752),
.C(n_737),
.Y(n_807)
);

OR2x2_ASAP7_75t_L g808 ( 
.A(n_770),
.B(n_736),
.Y(n_808)
);

AND2x2_ASAP7_75t_L g809 ( 
.A(n_757),
.B(n_717),
.Y(n_809)
);

HB1xp67_ASAP7_75t_L g810 ( 
.A(n_784),
.Y(n_810)
);

HB1xp67_ASAP7_75t_L g811 ( 
.A(n_788),
.Y(n_811)
);

BUFx2_ASAP7_75t_L g812 ( 
.A(n_756),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_757),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_779),
.Y(n_814)
);

AND2x2_ASAP7_75t_L g815 ( 
.A(n_753),
.B(n_717),
.Y(n_815)
);

AOI22xp33_ASAP7_75t_L g816 ( 
.A1(n_751),
.A2(n_759),
.B1(n_685),
.B2(n_771),
.Y(n_816)
);

AND2x4_ASAP7_75t_L g817 ( 
.A(n_805),
.B(n_736),
.Y(n_817)
);

INVx5_ASAP7_75t_L g818 ( 
.A(n_805),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_791),
.Y(n_819)
);

INVx4_ASAP7_75t_L g820 ( 
.A(n_812),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_794),
.B(n_760),
.Y(n_821)
);

INVxp67_ASAP7_75t_SL g822 ( 
.A(n_810),
.Y(n_822)
);

BUFx2_ASAP7_75t_L g823 ( 
.A(n_814),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_791),
.Y(n_824)
);

BUFx6f_ASAP7_75t_L g825 ( 
.A(n_814),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_793),
.Y(n_826)
);

AND2x2_ASAP7_75t_L g827 ( 
.A(n_798),
.B(n_799),
.Y(n_827)
);

OR2x2_ASAP7_75t_L g828 ( 
.A(n_800),
.B(n_732),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_793),
.Y(n_829)
);

AND2x2_ASAP7_75t_L g830 ( 
.A(n_798),
.B(n_714),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_792),
.Y(n_831)
);

NOR2x1_ASAP7_75t_L g832 ( 
.A(n_807),
.B(n_771),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_803),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_829),
.Y(n_834)
);

AND2x4_ASAP7_75t_L g835 ( 
.A(n_818),
.B(n_812),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_829),
.Y(n_836)
);

OR2x2_ASAP7_75t_L g837 ( 
.A(n_822),
.B(n_808),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_821),
.B(n_796),
.Y(n_838)
);

AND2x2_ASAP7_75t_L g839 ( 
.A(n_827),
.B(n_799),
.Y(n_839)
);

INVxp67_ASAP7_75t_SL g840 ( 
.A(n_828),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_827),
.B(n_815),
.Y(n_841)
);

INVxp67_ASAP7_75t_L g842 ( 
.A(n_823),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_823),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_831),
.B(n_815),
.Y(n_844)
);

AND2x2_ASAP7_75t_L g845 ( 
.A(n_820),
.B(n_799),
.Y(n_845)
);

CKINVDCx14_ASAP7_75t_R g846 ( 
.A(n_820),
.Y(n_846)
);

INVx2_ASAP7_75t_SL g847 ( 
.A(n_839),
.Y(n_847)
);

NOR2x1_ASAP7_75t_L g848 ( 
.A(n_835),
.B(n_820),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_838),
.B(n_802),
.Y(n_849)
);

NAND2xp33_ASAP7_75t_SL g850 ( 
.A(n_837),
.B(n_769),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_844),
.B(n_795),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_841),
.B(n_825),
.Y(n_852)
);

AOI22xp33_ASAP7_75t_L g853 ( 
.A1(n_850),
.A2(n_832),
.B1(n_816),
.B2(n_685),
.Y(n_853)
);

INVx1_ASAP7_75t_SL g854 ( 
.A(n_849),
.Y(n_854)
);

AND2x2_ASAP7_75t_L g855 ( 
.A(n_847),
.B(n_845),
.Y(n_855)
);

INVxp67_ASAP7_75t_L g856 ( 
.A(n_851),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_852),
.Y(n_857)
);

INVx1_ASAP7_75t_SL g858 ( 
.A(n_854),
.Y(n_858)
);

AOI21xp5_ASAP7_75t_L g859 ( 
.A1(n_856),
.A2(n_848),
.B(n_846),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_857),
.B(n_840),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_855),
.B(n_840),
.Y(n_861)
);

AND2x2_ASAP7_75t_L g862 ( 
.A(n_858),
.B(n_846),
.Y(n_862)
);

AND2x2_ASAP7_75t_L g863 ( 
.A(n_859),
.B(n_843),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_861),
.B(n_842),
.Y(n_864)
);

INVx2_ASAP7_75t_L g865 ( 
.A(n_862),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_864),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_863),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_864),
.Y(n_868)
);

NOR2xp33_ASAP7_75t_L g869 ( 
.A(n_865),
.B(n_860),
.Y(n_869)
);

NAND4xp25_ASAP7_75t_L g870 ( 
.A(n_865),
.B(n_853),
.C(n_775),
.D(n_835),
.Y(n_870)
);

NAND3xp33_ASAP7_75t_L g871 ( 
.A(n_867),
.B(n_868),
.C(n_866),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_865),
.B(n_842),
.Y(n_872)
);

AOI21xp5_ASAP7_75t_L g873 ( 
.A1(n_865),
.A2(n_853),
.B(n_811),
.Y(n_873)
);

NOR2xp33_ASAP7_75t_SL g874 ( 
.A(n_865),
.B(n_818),
.Y(n_874)
);

AOI221xp5_ASAP7_75t_L g875 ( 
.A1(n_867),
.A2(n_817),
.B1(n_825),
.B2(n_834),
.C(n_826),
.Y(n_875)
);

NAND4xp25_ASAP7_75t_L g876 ( 
.A(n_869),
.B(n_808),
.C(n_813),
.D(n_754),
.Y(n_876)
);

OAI22xp5_ASAP7_75t_L g877 ( 
.A1(n_873),
.A2(n_818),
.B1(n_825),
.B2(n_836),
.Y(n_877)
);

OAI211xp5_ASAP7_75t_SL g878 ( 
.A1(n_871),
.A2(n_660),
.B(n_641),
.C(n_813),
.Y(n_878)
);

AOI31xp33_ASAP7_75t_L g879 ( 
.A1(n_872),
.A2(n_755),
.A3(n_660),
.B(n_762),
.Y(n_879)
);

OAI211xp5_ASAP7_75t_SL g880 ( 
.A1(n_875),
.A2(n_819),
.B(n_824),
.C(n_797),
.Y(n_880)
);

NOR2xp33_ASAP7_75t_L g881 ( 
.A(n_870),
.B(n_825),
.Y(n_881)
);

OAI221xp5_ASAP7_75t_L g882 ( 
.A1(n_874),
.A2(n_818),
.B1(n_825),
.B2(n_764),
.C(n_780),
.Y(n_882)
);

NOR2xp33_ASAP7_75t_L g883 ( 
.A(n_869),
.B(n_818),
.Y(n_883)
);

AOI22xp5_ASAP7_75t_L g884 ( 
.A1(n_869),
.A2(n_817),
.B1(n_797),
.B2(n_809),
.Y(n_884)
);

NOR4xp75_ASAP7_75t_L g885 ( 
.A(n_877),
.B(n_718),
.C(n_830),
.D(n_645),
.Y(n_885)
);

INVx2_ASAP7_75t_SL g886 ( 
.A(n_883),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_881),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_884),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_878),
.Y(n_889)
);

NAND4xp75_ASAP7_75t_L g890 ( 
.A(n_880),
.B(n_645),
.C(n_804),
.D(n_714),
.Y(n_890)
);

HB1xp67_ASAP7_75t_L g891 ( 
.A(n_876),
.Y(n_891)
);

INVx1_ASAP7_75t_SL g892 ( 
.A(n_879),
.Y(n_892)
);

NOR3xp33_ASAP7_75t_SL g893 ( 
.A(n_887),
.B(n_882),
.C(n_739),
.Y(n_893)
);

NOR2xp33_ASAP7_75t_R g894 ( 
.A(n_886),
.B(n_191),
.Y(n_894)
);

NAND2xp33_ASAP7_75t_SL g895 ( 
.A(n_888),
.B(n_761),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_892),
.B(n_836),
.Y(n_896)
);

NOR3xp33_ASAP7_75t_SL g897 ( 
.A(n_889),
.B(n_739),
.C(n_765),
.Y(n_897)
);

NAND2xp33_ASAP7_75t_SL g898 ( 
.A(n_891),
.B(n_767),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_SL g899 ( 
.A(n_892),
.B(n_817),
.Y(n_899)
);

NOR3xp33_ASAP7_75t_SL g900 ( 
.A(n_890),
.B(n_768),
.C(n_747),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_885),
.B(n_831),
.Y(n_901)
);

NAND3xp33_ASAP7_75t_SL g902 ( 
.A(n_892),
.B(n_718),
.C(n_801),
.Y(n_902)
);

OR3x1_ASAP7_75t_L g903 ( 
.A(n_902),
.B(n_745),
.C(n_747),
.Y(n_903)
);

INVx1_ASAP7_75t_SL g904 ( 
.A(n_894),
.Y(n_904)
);

NAND3xp33_ASAP7_75t_L g905 ( 
.A(n_898),
.B(n_801),
.C(n_828),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_896),
.Y(n_906)
);

NAND4xp75_ASAP7_75t_L g907 ( 
.A(n_899),
.B(n_830),
.C(n_804),
.D(n_809),
.Y(n_907)
);

AOI22x1_ASAP7_75t_L g908 ( 
.A1(n_895),
.A2(n_800),
.B1(n_735),
.B2(n_750),
.Y(n_908)
);

NAND4xp25_ASAP7_75t_L g909 ( 
.A(n_901),
.B(n_806),
.C(n_803),
.D(n_750),
.Y(n_909)
);

AOI22xp5_ASAP7_75t_L g910 ( 
.A1(n_897),
.A2(n_806),
.B1(n_833),
.B2(n_779),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_893),
.Y(n_911)
);

NAND3xp33_ASAP7_75t_SL g912 ( 
.A(n_900),
.B(n_833),
.C(n_745),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_906),
.Y(n_913)
);

OA22x2_ASAP7_75t_L g914 ( 
.A1(n_911),
.A2(n_741),
.B1(n_682),
.B2(n_671),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_904),
.Y(n_915)
);

OAI22xp5_ASAP7_75t_SL g916 ( 
.A1(n_903),
.A2(n_741),
.B1(n_742),
.B2(n_738),
.Y(n_916)
);

INVx2_ASAP7_75t_SL g917 ( 
.A(n_908),
.Y(n_917)
);

HB1xp67_ASAP7_75t_L g918 ( 
.A(n_907),
.Y(n_918)
);

OAI21xp5_ASAP7_75t_L g919 ( 
.A1(n_918),
.A2(n_915),
.B(n_913),
.Y(n_919)
);

AOI22xp33_ASAP7_75t_L g920 ( 
.A1(n_917),
.A2(n_912),
.B1(n_909),
.B2(n_905),
.Y(n_920)
);

AOI22x1_ASAP7_75t_L g921 ( 
.A1(n_916),
.A2(n_910),
.B1(n_742),
.B2(n_738),
.Y(n_921)
);

AOI31xp33_ASAP7_75t_L g922 ( 
.A1(n_919),
.A2(n_914),
.A3(n_735),
.B(n_734),
.Y(n_922)
);

AOI22xp33_ASAP7_75t_L g923 ( 
.A1(n_920),
.A2(n_921),
.B1(n_733),
.B2(n_743),
.Y(n_923)
);

OAI22xp5_ASAP7_75t_L g924 ( 
.A1(n_920),
.A2(n_743),
.B1(n_733),
.B2(n_663),
.Y(n_924)
);

XOR2xp5_ASAP7_75t_L g925 ( 
.A(n_924),
.B(n_730),
.Y(n_925)
);

AOI22xp33_ASAP7_75t_L g926 ( 
.A1(n_925),
.A2(n_923),
.B1(n_922),
.B2(n_743),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_926),
.Y(n_927)
);

OAI221xp5_ASAP7_75t_R g928 ( 
.A1(n_927),
.A2(n_682),
.B1(n_671),
.B2(n_610),
.C(n_730),
.Y(n_928)
);

AOI211xp5_ASAP7_75t_L g929 ( 
.A1(n_928),
.A2(n_701),
.B(n_674),
.C(n_734),
.Y(n_929)
);


endmodule