module fake_netlist_6_939_n_3307 (n_52, n_591, n_435, n_1, n_91, n_793, n_326, n_801, n_256, n_853, n_440, n_587, n_695, n_507, n_909, n_580, n_762, n_881, n_875, n_209, n_367, n_465, n_680, n_741, n_760, n_590, n_625, n_63, n_661, n_223, n_278, n_341, n_362, n_148, n_226, n_828, n_161, n_22, n_208, n_462, n_68, n_607, n_671, n_726, n_316, n_419, n_28, n_304, n_212, n_700, n_50, n_694, n_7, n_740, n_578, n_703, n_144, n_365, n_125, n_168, n_384, n_297, n_595, n_627, n_524, n_342, n_77, n_820, n_783, n_106, n_725, n_358, n_160, n_751, n_449, n_131, n_749, n_798, n_188, n_310, n_509, n_186, n_245, n_0, n_368, n_575, n_677, n_805, n_396, n_495, n_815, n_350, n_78, n_84, n_585, n_732, n_568, n_392, n_840, n_442, n_480, n_142, n_874, n_724, n_143, n_382, n_673, n_180, n_62, n_628, n_883, n_557, n_823, n_349, n_643, n_233, n_617, n_698, n_898, n_845, n_255, n_807, n_739, n_284, n_400, n_140, n_337, n_865, n_893, n_214, n_485, n_67, n_15, n_443, n_246, n_892, n_768, n_38, n_471, n_289, n_421, n_781, n_424, n_789, n_615, n_59, n_181, n_182, n_238, n_573, n_769, n_202, n_320, n_108, n_639, n_676, n_327, n_794, n_727, n_894, n_369, n_597, n_685, n_280, n_287, n_832, n_353, n_610, n_555, n_389, n_814, n_415, n_830, n_65, n_230, n_605, n_461, n_873, n_141, n_383, n_826, n_669, n_200, n_447, n_176, n_872, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_517, n_718, n_747, n_852, n_667, n_71, n_74, n_229, n_542, n_847, n_644, n_682, n_851, n_621, n_305, n_72, n_721, n_750, n_532, n_742, n_173, n_535, n_691, n_250, n_372, n_468, n_544, n_901, n_111, n_504, n_314, n_378, n_413, n_377, n_791, n_35, n_183, n_510, n_837, n_836, n_79, n_863, n_375, n_601, n_338, n_522, n_466, n_704, n_748, n_506, n_56, n_763, n_360, n_603, n_119, n_235, n_536, n_895, n_866, n_622, n_147, n_191, n_340, n_710, n_387, n_452, n_616, n_658, n_744, n_39, n_344, n_73, n_581, n_428, n_761, n_785, n_746, n_609, n_765, n_432, n_641, n_822, n_693, n_101, n_167, n_631, n_174, n_127, n_516, n_153, n_720, n_525, n_758, n_842, n_611, n_156, n_491, n_878, n_145, n_42, n_133, n_656, n_772, n_96, n_8, n_843, n_797, n_666, n_371, n_795, n_770, n_567, n_899, n_189, n_738, n_405, n_213, n_538, n_294, n_302, n_499, n_380, n_838, n_129, n_705, n_647, n_197, n_11, n_137, n_17, n_343, n_844, n_448, n_886, n_20, n_494, n_539, n_493, n_397, n_155, n_109, n_614, n_529, n_445, n_425, n_684, n_122, n_888, n_45, n_454, n_34, n_218, n_638, n_70, n_234, n_910, n_37, n_486, n_911, n_381, n_82, n_27, n_236, n_653, n_887, n_752, n_908, n_112, n_172, n_713, n_648, n_657, n_576, n_472, n_270, n_239, n_126, n_414, n_97, n_563, n_58, n_782, n_490, n_803, n_290, n_220, n_809, n_118, n_224, n_48, n_25, n_93, n_839, n_80, n_734, n_708, n_196, n_402, n_352, n_668, n_478, n_626, n_574, n_779, n_9, n_800, n_460, n_107, n_907, n_854, n_6, n_417, n_14, n_446, n_498, n_662, n_89, n_374, n_659, n_709, n_870, n_366, n_904, n_777, n_407, n_913, n_450, n_103, n_808, n_867, n_272, n_526, n_185, n_712, n_348, n_711, n_579, n_69, n_376, n_390, n_473, n_293, n_31, n_334, n_559, n_53, n_370, n_44, n_458, n_232, n_650, n_16, n_163, n_717, n_46, n_330, n_771, n_470, n_475, n_298, n_18, n_492, n_281, n_258, n_551, n_154, n_699, n_456, n_564, n_98, n_260, n_265, n_313, n_451, n_624, n_824, n_279, n_686, n_796, n_252, n_757, n_228, n_565, n_594, n_719, n_356, n_577, n_166, n_184, n_552, n_619, n_885, n_216, n_455, n_896, n_83, n_521, n_363, n_572, n_912, n_395, n_813, n_592, n_745, n_654, n_323, n_829, n_606, n_393, n_818, n_411, n_503, n_716, n_152, n_623, n_92, n_884, n_599, n_513, n_855, n_776, n_321, n_645, n_331, n_105, n_227, n_132, n_868, n_570, n_731, n_859, n_406, n_483, n_735, n_102, n_204, n_482, n_755, n_474, n_527, n_261, n_608, n_620, n_420, n_683, n_630, n_312, n_394, n_32, n_66, n_130, n_519, n_541, n_512, n_164, n_292, n_100, n_121, n_307, n_469, n_433, n_500, n_23, n_792, n_880, n_476, n_714, n_2, n_291, n_219, n_543, n_889, n_357, n_150, n_264, n_263, n_589, n_860, n_481, n_788, n_819, n_821, n_325, n_767, n_804, n_329, n_464, n_600, n_831, n_802, n_561, n_33, n_477, n_549, n_533, n_408, n_806, n_864, n_879, n_61, n_237, n_584, n_244, n_399, n_76, n_243, n_124, n_548, n_905, n_94, n_282, n_436, n_833, n_116, n_211, n_523, n_117, n_175, n_322, n_707, n_345, n_409, n_231, n_354, n_689, n_40, n_799, n_505, n_240, n_756, n_139, n_319, n_41, n_134, n_547, n_537, n_273, n_558, n_810, n_635, n_95, n_787, n_311, n_10, n_403, n_723, n_253, n_634, n_583, n_596, n_123, n_136, n_546, n_562, n_249, n_201, n_386, n_764, n_556, n_159, n_157, n_162, n_692, n_733, n_754, n_115, n_487, n_550, n_128, n_241, n_30, n_275, n_553, n_43, n_652, n_849, n_560, n_753, n_642, n_276, n_569, n_441, n_221, n_811, n_882, n_444, n_586, n_423, n_146, n_737, n_318, n_303, n_511, n_715, n_467, n_306, n_21, n_193, n_269, n_359, n_346, n_88, n_3, n_416, n_530, n_277, n_520, n_418, n_113, n_618, n_790, n_582, n_4, n_199, n_138, n_266, n_296, n_861, n_674, n_857, n_871, n_775, n_571, n_268, n_271, n_404, n_651, n_439, n_158, n_217, n_49, n_210, n_299, n_518, n_206, n_679, n_5, n_453, n_612, n_633, n_665, n_902, n_333, n_588, n_215, n_178, n_247, n_225, n_308, n_309, n_914, n_759, n_355, n_426, n_317, n_149, n_632, n_702, n_431, n_90, n_347, n_812, n_24, n_459, n_54, n_502, n_328, n_672, n_534, n_488, n_429, n_373, n_87, n_195, n_285, n_497, n_780, n_773, n_675, n_903, n_85, n_99, n_257, n_730, n_655, n_13, n_706, n_786, n_670, n_203, n_286, n_254, n_207, n_834, n_242, n_835, n_19, n_47, n_690, n_29, n_850, n_75, n_401, n_324, n_743, n_766, n_816, n_335, n_430, n_463, n_545, n_489, n_877, n_205, n_604, n_848, n_120, n_251, n_301, n_274, n_636, n_825, n_728, n_681, n_729, n_110, n_151, n_876, n_774, n_412, n_640, n_81, n_660, n_36, n_26, n_55, n_267, n_438, n_339, n_784, n_315, n_434, n_515, n_64, n_288, n_427, n_479, n_496, n_598, n_422, n_696, n_906, n_688, n_722, n_862, n_135, n_165, n_351, n_869, n_437, n_259, n_177, n_540, n_593, n_514, n_646, n_528, n_391, n_457, n_687, n_697, n_364, n_890, n_637, n_295, n_385, n_701, n_817, n_629, n_388, n_190, n_858, n_262, n_484, n_613, n_736, n_187, n_897, n_900, n_846, n_501, n_841, n_531, n_827, n_60, n_361, n_508, n_663, n_856, n_379, n_170, n_778, n_332, n_891, n_336, n_12, n_398, n_410, n_566, n_554, n_602, n_194, n_664, n_171, n_678, n_192, n_57, n_169, n_51, n_649, n_283, n_3307);

input n_52;
input n_591;
input n_435;
input n_1;
input n_91;
input n_793;
input n_326;
input n_801;
input n_256;
input n_853;
input n_440;
input n_587;
input n_695;
input n_507;
input n_909;
input n_580;
input n_762;
input n_881;
input n_875;
input n_209;
input n_367;
input n_465;
input n_680;
input n_741;
input n_760;
input n_590;
input n_625;
input n_63;
input n_661;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_828;
input n_161;
input n_22;
input n_208;
input n_462;
input n_68;
input n_607;
input n_671;
input n_726;
input n_316;
input n_419;
input n_28;
input n_304;
input n_212;
input n_700;
input n_50;
input n_694;
input n_7;
input n_740;
input n_578;
input n_703;
input n_144;
input n_365;
input n_125;
input n_168;
input n_384;
input n_297;
input n_595;
input n_627;
input n_524;
input n_342;
input n_77;
input n_820;
input n_783;
input n_106;
input n_725;
input n_358;
input n_160;
input n_751;
input n_449;
input n_131;
input n_749;
input n_798;
input n_188;
input n_310;
input n_509;
input n_186;
input n_245;
input n_0;
input n_368;
input n_575;
input n_677;
input n_805;
input n_396;
input n_495;
input n_815;
input n_350;
input n_78;
input n_84;
input n_585;
input n_732;
input n_568;
input n_392;
input n_840;
input n_442;
input n_480;
input n_142;
input n_874;
input n_724;
input n_143;
input n_382;
input n_673;
input n_180;
input n_62;
input n_628;
input n_883;
input n_557;
input n_823;
input n_349;
input n_643;
input n_233;
input n_617;
input n_698;
input n_898;
input n_845;
input n_255;
input n_807;
input n_739;
input n_284;
input n_400;
input n_140;
input n_337;
input n_865;
input n_893;
input n_214;
input n_485;
input n_67;
input n_15;
input n_443;
input n_246;
input n_892;
input n_768;
input n_38;
input n_471;
input n_289;
input n_421;
input n_781;
input n_424;
input n_789;
input n_615;
input n_59;
input n_181;
input n_182;
input n_238;
input n_573;
input n_769;
input n_202;
input n_320;
input n_108;
input n_639;
input n_676;
input n_327;
input n_794;
input n_727;
input n_894;
input n_369;
input n_597;
input n_685;
input n_280;
input n_287;
input n_832;
input n_353;
input n_610;
input n_555;
input n_389;
input n_814;
input n_415;
input n_830;
input n_65;
input n_230;
input n_605;
input n_461;
input n_873;
input n_141;
input n_383;
input n_826;
input n_669;
input n_200;
input n_447;
input n_176;
input n_872;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_517;
input n_718;
input n_747;
input n_852;
input n_667;
input n_71;
input n_74;
input n_229;
input n_542;
input n_847;
input n_644;
input n_682;
input n_851;
input n_621;
input n_305;
input n_72;
input n_721;
input n_750;
input n_532;
input n_742;
input n_173;
input n_535;
input n_691;
input n_250;
input n_372;
input n_468;
input n_544;
input n_901;
input n_111;
input n_504;
input n_314;
input n_378;
input n_413;
input n_377;
input n_791;
input n_35;
input n_183;
input n_510;
input n_837;
input n_836;
input n_79;
input n_863;
input n_375;
input n_601;
input n_338;
input n_522;
input n_466;
input n_704;
input n_748;
input n_506;
input n_56;
input n_763;
input n_360;
input n_603;
input n_119;
input n_235;
input n_536;
input n_895;
input n_866;
input n_622;
input n_147;
input n_191;
input n_340;
input n_710;
input n_387;
input n_452;
input n_616;
input n_658;
input n_744;
input n_39;
input n_344;
input n_73;
input n_581;
input n_428;
input n_761;
input n_785;
input n_746;
input n_609;
input n_765;
input n_432;
input n_641;
input n_822;
input n_693;
input n_101;
input n_167;
input n_631;
input n_174;
input n_127;
input n_516;
input n_153;
input n_720;
input n_525;
input n_758;
input n_842;
input n_611;
input n_156;
input n_491;
input n_878;
input n_145;
input n_42;
input n_133;
input n_656;
input n_772;
input n_96;
input n_8;
input n_843;
input n_797;
input n_666;
input n_371;
input n_795;
input n_770;
input n_567;
input n_899;
input n_189;
input n_738;
input n_405;
input n_213;
input n_538;
input n_294;
input n_302;
input n_499;
input n_380;
input n_838;
input n_129;
input n_705;
input n_647;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_844;
input n_448;
input n_886;
input n_20;
input n_494;
input n_539;
input n_493;
input n_397;
input n_155;
input n_109;
input n_614;
input n_529;
input n_445;
input n_425;
input n_684;
input n_122;
input n_888;
input n_45;
input n_454;
input n_34;
input n_218;
input n_638;
input n_70;
input n_234;
input n_910;
input n_37;
input n_486;
input n_911;
input n_381;
input n_82;
input n_27;
input n_236;
input n_653;
input n_887;
input n_752;
input n_908;
input n_112;
input n_172;
input n_713;
input n_648;
input n_657;
input n_576;
input n_472;
input n_270;
input n_239;
input n_126;
input n_414;
input n_97;
input n_563;
input n_58;
input n_782;
input n_490;
input n_803;
input n_290;
input n_220;
input n_809;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_839;
input n_80;
input n_734;
input n_708;
input n_196;
input n_402;
input n_352;
input n_668;
input n_478;
input n_626;
input n_574;
input n_779;
input n_9;
input n_800;
input n_460;
input n_107;
input n_907;
input n_854;
input n_6;
input n_417;
input n_14;
input n_446;
input n_498;
input n_662;
input n_89;
input n_374;
input n_659;
input n_709;
input n_870;
input n_366;
input n_904;
input n_777;
input n_407;
input n_913;
input n_450;
input n_103;
input n_808;
input n_867;
input n_272;
input n_526;
input n_185;
input n_712;
input n_348;
input n_711;
input n_579;
input n_69;
input n_376;
input n_390;
input n_473;
input n_293;
input n_31;
input n_334;
input n_559;
input n_53;
input n_370;
input n_44;
input n_458;
input n_232;
input n_650;
input n_16;
input n_163;
input n_717;
input n_46;
input n_330;
input n_771;
input n_470;
input n_475;
input n_298;
input n_18;
input n_492;
input n_281;
input n_258;
input n_551;
input n_154;
input n_699;
input n_456;
input n_564;
input n_98;
input n_260;
input n_265;
input n_313;
input n_451;
input n_624;
input n_824;
input n_279;
input n_686;
input n_796;
input n_252;
input n_757;
input n_228;
input n_565;
input n_594;
input n_719;
input n_356;
input n_577;
input n_166;
input n_184;
input n_552;
input n_619;
input n_885;
input n_216;
input n_455;
input n_896;
input n_83;
input n_521;
input n_363;
input n_572;
input n_912;
input n_395;
input n_813;
input n_592;
input n_745;
input n_654;
input n_323;
input n_829;
input n_606;
input n_393;
input n_818;
input n_411;
input n_503;
input n_716;
input n_152;
input n_623;
input n_92;
input n_884;
input n_599;
input n_513;
input n_855;
input n_776;
input n_321;
input n_645;
input n_331;
input n_105;
input n_227;
input n_132;
input n_868;
input n_570;
input n_731;
input n_859;
input n_406;
input n_483;
input n_735;
input n_102;
input n_204;
input n_482;
input n_755;
input n_474;
input n_527;
input n_261;
input n_608;
input n_620;
input n_420;
input n_683;
input n_630;
input n_312;
input n_394;
input n_32;
input n_66;
input n_130;
input n_519;
input n_541;
input n_512;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_469;
input n_433;
input n_500;
input n_23;
input n_792;
input n_880;
input n_476;
input n_714;
input n_2;
input n_291;
input n_219;
input n_543;
input n_889;
input n_357;
input n_150;
input n_264;
input n_263;
input n_589;
input n_860;
input n_481;
input n_788;
input n_819;
input n_821;
input n_325;
input n_767;
input n_804;
input n_329;
input n_464;
input n_600;
input n_831;
input n_802;
input n_561;
input n_33;
input n_477;
input n_549;
input n_533;
input n_408;
input n_806;
input n_864;
input n_879;
input n_61;
input n_237;
input n_584;
input n_244;
input n_399;
input n_76;
input n_243;
input n_124;
input n_548;
input n_905;
input n_94;
input n_282;
input n_436;
input n_833;
input n_116;
input n_211;
input n_523;
input n_117;
input n_175;
input n_322;
input n_707;
input n_345;
input n_409;
input n_231;
input n_354;
input n_689;
input n_40;
input n_799;
input n_505;
input n_240;
input n_756;
input n_139;
input n_319;
input n_41;
input n_134;
input n_547;
input n_537;
input n_273;
input n_558;
input n_810;
input n_635;
input n_95;
input n_787;
input n_311;
input n_10;
input n_403;
input n_723;
input n_253;
input n_634;
input n_583;
input n_596;
input n_123;
input n_136;
input n_546;
input n_562;
input n_249;
input n_201;
input n_386;
input n_764;
input n_556;
input n_159;
input n_157;
input n_162;
input n_692;
input n_733;
input n_754;
input n_115;
input n_487;
input n_550;
input n_128;
input n_241;
input n_30;
input n_275;
input n_553;
input n_43;
input n_652;
input n_849;
input n_560;
input n_753;
input n_642;
input n_276;
input n_569;
input n_441;
input n_221;
input n_811;
input n_882;
input n_444;
input n_586;
input n_423;
input n_146;
input n_737;
input n_318;
input n_303;
input n_511;
input n_715;
input n_467;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_346;
input n_88;
input n_3;
input n_416;
input n_530;
input n_277;
input n_520;
input n_418;
input n_113;
input n_618;
input n_790;
input n_582;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_861;
input n_674;
input n_857;
input n_871;
input n_775;
input n_571;
input n_268;
input n_271;
input n_404;
input n_651;
input n_439;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_518;
input n_206;
input n_679;
input n_5;
input n_453;
input n_612;
input n_633;
input n_665;
input n_902;
input n_333;
input n_588;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_914;
input n_759;
input n_355;
input n_426;
input n_317;
input n_149;
input n_632;
input n_702;
input n_431;
input n_90;
input n_347;
input n_812;
input n_24;
input n_459;
input n_54;
input n_502;
input n_328;
input n_672;
input n_534;
input n_488;
input n_429;
input n_373;
input n_87;
input n_195;
input n_285;
input n_497;
input n_780;
input n_773;
input n_675;
input n_903;
input n_85;
input n_99;
input n_257;
input n_730;
input n_655;
input n_13;
input n_706;
input n_786;
input n_670;
input n_203;
input n_286;
input n_254;
input n_207;
input n_834;
input n_242;
input n_835;
input n_19;
input n_47;
input n_690;
input n_29;
input n_850;
input n_75;
input n_401;
input n_324;
input n_743;
input n_766;
input n_816;
input n_335;
input n_430;
input n_463;
input n_545;
input n_489;
input n_877;
input n_205;
input n_604;
input n_848;
input n_120;
input n_251;
input n_301;
input n_274;
input n_636;
input n_825;
input n_728;
input n_681;
input n_729;
input n_110;
input n_151;
input n_876;
input n_774;
input n_412;
input n_640;
input n_81;
input n_660;
input n_36;
input n_26;
input n_55;
input n_267;
input n_438;
input n_339;
input n_784;
input n_315;
input n_434;
input n_515;
input n_64;
input n_288;
input n_427;
input n_479;
input n_496;
input n_598;
input n_422;
input n_696;
input n_906;
input n_688;
input n_722;
input n_862;
input n_135;
input n_165;
input n_351;
input n_869;
input n_437;
input n_259;
input n_177;
input n_540;
input n_593;
input n_514;
input n_646;
input n_528;
input n_391;
input n_457;
input n_687;
input n_697;
input n_364;
input n_890;
input n_637;
input n_295;
input n_385;
input n_701;
input n_817;
input n_629;
input n_388;
input n_190;
input n_858;
input n_262;
input n_484;
input n_613;
input n_736;
input n_187;
input n_897;
input n_900;
input n_846;
input n_501;
input n_841;
input n_531;
input n_827;
input n_60;
input n_361;
input n_508;
input n_663;
input n_856;
input n_379;
input n_170;
input n_778;
input n_332;
input n_891;
input n_336;
input n_12;
input n_398;
input n_410;
input n_566;
input n_554;
input n_602;
input n_194;
input n_664;
input n_171;
input n_678;
input n_192;
input n_57;
input n_169;
input n_51;
input n_649;
input n_283;

output n_3307;

wire n_992;
wire n_2542;
wire n_1671;
wire n_2817;
wire n_1613;
wire n_1458;
wire n_1234;
wire n_2576;
wire n_3254;
wire n_1199;
wire n_1674;
wire n_1027;
wire n_1351;
wire n_3266;
wire n_1189;
wire n_3152;
wire n_1212;
wire n_2157;
wire n_2332;
wire n_1307;
wire n_3178;
wire n_2003;
wire n_1038;
wire n_1581;
wire n_1003;
wire n_1237;
wire n_1061;
wire n_2353;
wire n_2534;
wire n_3089;
wire n_3301;
wire n_1357;
wire n_1853;
wire n_2451;
wire n_1738;
wire n_2243;
wire n_1575;
wire n_1854;
wire n_2324;
wire n_3088;
wire n_1923;
wire n_3257;
wire n_1342;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_2260;
wire n_3222;
wire n_1708;
wire n_1151;
wire n_2977;
wire n_1739;
wire n_2051;
wire n_2317;
wire n_1380;
wire n_2359;
wire n_2847;
wire n_1402;
wire n_2557;
wire n_1688;
wire n_1691;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_2405;
wire n_1160;
wire n_2647;
wire n_1238;
wire n_1991;
wire n_2570;
wire n_2179;
wire n_2386;
wire n_2997;
wire n_1724;
wire n_1032;
wire n_2336;
wire n_1247;
wire n_1547;
wire n_2521;
wire n_3046;
wire n_2956;
wire n_1553;
wire n_1099;
wire n_2491;
wire n_1264;
wire n_1192;
wire n_1844;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_2211;
wire n_1370;
wire n_1786;
wire n_2382;
wire n_2672;
wire n_3030;
wire n_2291;
wire n_2299;
wire n_1371;
wire n_1285;
wire n_2886;
wire n_2974;
wire n_1985;
wire n_2989;
wire n_2838;
wire n_2184;
wire n_2982;
wire n_1803;
wire n_1172;
wire n_2509;
wire n_2513;
wire n_3282;
wire n_1590;
wire n_2645;
wire n_1532;
wire n_2313;
wire n_2628;
wire n_3071;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_2926;
wire n_1704;
wire n_1078;
wire n_1711;
wire n_2247;
wire n_3106;
wire n_1140;
wire n_2630;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_2344;
wire n_1579;
wire n_3275;
wire n_2365;
wire n_2470;
wire n_2321;
wire n_1263;
wire n_2019;
wire n_3031;
wire n_2074;
wire n_2447;
wire n_2919;
wire n_2129;
wire n_2340;
wire n_1261;
wire n_945;
wire n_2286;
wire n_1649;
wire n_2018;
wire n_2094;
wire n_3080;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_2356;
wire n_2399;
wire n_1422;
wire n_1772;
wire n_1232;
wire n_1572;
wire n_1874;
wire n_3165;
wire n_1119;
wire n_2865;
wire n_2825;
wire n_2013;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_2510;
wire n_1541;
wire n_1300;
wire n_2480;
wire n_2739;
wire n_3023;
wire n_3232;
wire n_1313;
wire n_2791;
wire n_3251;
wire n_1056;
wire n_2212;
wire n_3048;
wire n_1455;
wire n_2418;
wire n_2864;
wire n_1163;
wire n_2729;
wire n_3063;
wire n_1180;
wire n_2256;
wire n_2582;
wire n_943;
wire n_1798;
wire n_1550;
wire n_2703;
wire n_2786;
wire n_1591;
wire n_3122;
wire n_2806;
wire n_1344;
wire n_3261;
wire n_2730;
wire n_2495;
wire n_940;
wire n_1781;
wire n_1971;
wire n_2058;
wire n_2090;
wire n_2603;
wire n_2660;
wire n_3028;
wire n_2981;
wire n_3076;
wire n_2173;
wire n_2004;
wire n_1106;
wire n_1471;
wire n_953;
wire n_1094;
wire n_3077;
wire n_1345;
wire n_1820;
wire n_2873;
wire n_3107;
wire n_2880;
wire n_3225;
wire n_2394;
wire n_2108;
wire n_1421;
wire n_2836;
wire n_1936;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_2378;
wire n_1660;
wire n_1961;
wire n_3047;
wire n_1280;
wire n_2655;
wire n_1400;
wire n_2625;
wire n_3296;
wire n_2843;
wire n_1467;
wire n_3297;
wire n_976;
wire n_3067;
wire n_2155;
wire n_2686;
wire n_1445;
wire n_2364;
wire n_2551;
wire n_1526;
wire n_1560;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_2996;
wire n_2599;
wire n_2985;
wire n_1978;
wire n_2085;
wire n_917;
wire n_2370;
wire n_2612;
wire n_1446;
wire n_2591;
wire n_1815;
wire n_2214;
wire n_1658;
wire n_2593;
wire n_3269;
wire n_1230;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_2613;
wire n_1333;
wire n_2496;
wire n_2708;
wire n_1648;
wire n_3189;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_2725;
wire n_2277;
wire n_3164;
wire n_1558;
wire n_1732;
wire n_2300;
wire n_1986;
wire n_2397;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_2190;
wire n_2907;
wire n_2735;
wire n_1843;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_2778;
wire n_2850;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_1441;
wire n_1123;
wire n_1309;
wire n_2104;
wire n_1381;
wire n_2961;
wire n_1699;
wire n_916;
wire n_2093;
wire n_2633;
wire n_2207;
wire n_1970;
wire n_2770;
wire n_2101;
wire n_2696;
wire n_2059;
wire n_2198;
wire n_2669;
wire n_2925;
wire n_2073;
wire n_2273;
wire n_2546;
wire n_3272;
wire n_3193;
wire n_2522;
wire n_2792;
wire n_1328;
wire n_1957;
wire n_2917;
wire n_2616;
wire n_3118;
wire n_1907;
wire n_2529;
wire n_1162;
wire n_1530;
wire n_939;
wire n_1543;
wire n_2811;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_982;
wire n_2674;
wire n_2832;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_932;
wire n_2831;
wire n_2998;
wire n_1876;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_979;
wire n_1873;
wire n_1866;
wire n_1680;
wire n_993;
wire n_2692;
wire n_3248;
wire n_2031;
wire n_2130;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_2228;
wire n_1988;
wire n_2941;
wire n_1278;
wire n_2455;
wire n_2876;
wire n_2654;
wire n_3036;
wire n_2469;
wire n_1064;
wire n_3099;
wire n_1396;
wire n_2355;
wire n_966;
wire n_2908;
wire n_3168;
wire n_2751;
wire n_2764;
wire n_1663;
wire n_2895;
wire n_2009;
wire n_1793;
wire n_2922;
wire n_1233;
wire n_1289;
wire n_2714;
wire n_2245;
wire n_3092;
wire n_3055;
wire n_2068;
wire n_1107;
wire n_2866;
wire n_2457;
wire n_3294;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_2580;
wire n_2176;
wire n_2072;
wire n_1354;
wire n_2821;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_2459;
wire n_1111;
wire n_1713;
wire n_2971;
wire n_2678;
wire n_1251;
wire n_1265;
wire n_2711;
wire n_1726;
wire n_1950;
wire n_1563;
wire n_1912;
wire n_2434;
wire n_1982;
wire n_2878;
wire n_3012;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_2818;
wire n_2428;
wire n_3247;
wire n_3069;
wire n_922;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_2664;
wire n_1722;
wire n_1664;
wire n_2641;
wire n_3022;
wire n_3052;
wire n_1165;
wire n_2008;
wire n_2749;
wire n_3298;
wire n_2192;
wire n_3281;
wire n_2254;
wire n_2345;
wire n_1926;
wire n_1175;
wire n_3273;
wire n_1386;
wire n_2311;
wire n_1896;
wire n_2965;
wire n_1747;
wire n_3058;
wire n_1012;
wire n_2624;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_2350;
wire n_2804;
wire n_2453;
wire n_2193;
wire n_2676;
wire n_1655;
wire n_928;
wire n_1214;
wire n_1801;
wire n_1886;
wire n_2347;
wire n_2092;
wire n_1654;
wire n_1157;
wire n_1750;
wire n_2994;
wire n_1462;
wire n_3153;
wire n_1188;
wire n_1752;
wire n_1813;
wire n_2514;
wire n_2206;
wire n_2810;
wire n_2967;
wire n_2319;
wire n_2519;
wire n_2916;
wire n_1063;
wire n_1588;
wire n_2963;
wire n_2947;
wire n_2467;
wire n_2602;
wire n_2468;
wire n_3145;
wire n_1124;
wire n_1624;
wire n_2096;
wire n_2980;
wire n_1965;
wire n_2476;
wire n_3280;
wire n_1515;
wire n_961;
wire n_1317;
wire n_1082;
wire n_3227;
wire n_2733;
wire n_2824;
wire n_3289;
wire n_2377;
wire n_2178;
wire n_3271;
wire n_950;
wire n_2812;
wire n_2644;
wire n_2036;
wire n_2976;
wire n_2152;
wire n_1709;
wire n_3009;
wire n_2652;
wire n_2411;
wire n_2525;
wire n_1825;
wire n_2393;
wire n_1757;
wire n_1796;
wire n_2657;
wire n_1792;
wire n_2067;
wire n_2136;
wire n_2921;
wire n_2409;
wire n_2082;
wire n_2252;
wire n_1412;
wire n_2497;
wire n_2687;
wire n_3237;
wire n_949;
wire n_1630;
wire n_2887;
wire n_2075;
wire n_2194;
wire n_2972;
wire n_2619;
wire n_3139;
wire n_2763;
wire n_2762;
wire n_1987;
wire n_968;
wire n_1369;
wire n_2271;
wire n_1008;
wire n_3192;
wire n_1546;
wire n_2583;
wire n_2606;
wire n_2279;
wire n_1052;
wire n_1033;
wire n_2794;
wire n_1296;
wire n_2663;
wire n_1990;
wire n_2391;
wire n_2431;
wire n_3073;
wire n_2987;
wire n_2938;
wire n_2150;
wire n_1294;
wire n_2943;
wire n_1420;
wire n_2078;
wire n_1634;
wire n_3252;
wire n_2932;
wire n_1767;
wire n_3253;
wire n_1779;
wire n_1465;
wire n_3209;
wire n_2622;
wire n_1858;
wire n_1044;
wire n_2658;
wire n_2665;
wire n_2165;
wire n_2133;
wire n_1712;
wire n_3021;
wire n_1391;
wire n_1523;
wire n_2750;
wire n_2893;
wire n_2775;
wire n_1208;
wire n_2558;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_2954;
wire n_2728;
wire n_2349;
wire n_3128;
wire n_2684;
wire n_2712;
wire n_1072;
wire n_3146;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_1100;
wire n_1487;
wire n_2691;
wire n_2913;
wire n_1756;
wire n_3183;
wire n_1128;
wire n_2493;
wire n_2230;
wire n_2705;
wire n_1969;
wire n_2690;
wire n_1071;
wire n_1565;
wire n_1067;
wire n_1493;
wire n_2145;
wire n_1968;
wire n_1952;
wire n_2573;
wire n_2646;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_2535;
wire n_2631;
wire n_1364;
wire n_3078;
wire n_2436;
wire n_2870;
wire n_1249;
wire n_2706;
wire n_1293;
wire n_2693;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_3159;
wire n_1451;
wire n_963;
wire n_2767;
wire n_1839;
wire n_2341;
wire n_1765;
wire n_2707;
wire n_3240;
wire n_1514;
wire n_1863;
wire n_3037;
wire n_1646;
wire n_3293;
wire n_1714;
wire n_1139;
wire n_3179;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_2897;
wire n_2537;
wire n_2554;
wire n_996;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_1513;
wire n_2747;
wire n_3171;
wire n_1913;
wire n_2097;
wire n_2170;
wire n_1488;
wire n_2853;
wire n_1808;
wire n_3053;
wire n_948;
wire n_2517;
wire n_2713;
wire n_2148;
wire n_977;
wire n_2339;
wire n_1005;
wire n_1947;
wire n_2765;
wire n_2861;
wire n_3158;
wire n_1788;
wire n_1999;
wire n_2731;
wire n_2590;
wire n_2643;
wire n_3150;
wire n_3018;
wire n_1469;
wire n_2060;
wire n_2608;
wire n_1838;
wire n_2638;
wire n_1835;
wire n_1776;
wire n_1766;
wire n_1959;
wire n_3133;
wire n_2002;
wire n_2650;
wire n_2138;
wire n_1492;
wire n_987;
wire n_2414;
wire n_1340;
wire n_3014;
wire n_3166;
wire n_1771;
wire n_2316;
wire n_3104;
wire n_3148;
wire n_2262;
wire n_3229;
wire n_1707;
wire n_2239;
wire n_3082;
wire n_1432;
wire n_2208;
wire n_989;
wire n_2604;
wire n_2407;
wire n_1277;
wire n_2816;
wire n_2689;
wire n_2933;
wire n_1473;
wire n_2191;
wire n_1723;
wire n_2717;
wire n_1246;
wire n_1878;
wire n_2574;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_2842;
wire n_2675;
wire n_1426;
wire n_1004;
wire n_1176;
wire n_2134;
wire n_1529;
wire n_2335;
wire n_2473;
wire n_1022;
wire n_2069;
wire n_2307;
wire n_2362;
wire n_2539;
wire n_2698;
wire n_2667;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_3119;
wire n_2948;
wire n_1577;
wire n_2958;
wire n_2297;
wire n_1181;
wire n_2119;
wire n_1822;
wire n_2936;
wire n_947;
wire n_3224;
wire n_1117;
wire n_2489;
wire n_1448;
wire n_1087;
wire n_3173;
wire n_1992;
wire n_1049;
wire n_3223;
wire n_2771;
wire n_2445;
wire n_3020;
wire n_2057;
wire n_2103;
wire n_3140;
wire n_3185;
wire n_2605;
wire n_1666;
wire n_2772;
wire n_1505;
wire n_1717;
wire n_926;
wire n_1817;
wire n_2449;
wire n_927;
wire n_2610;
wire n_3129;
wire n_1849;
wire n_2848;
wire n_919;
wire n_2868;
wire n_1698;
wire n_2231;
wire n_929;
wire n_2520;
wire n_1228;
wire n_2857;
wire n_1568;
wire n_1490;
wire n_2372;
wire n_1299;
wire n_2896;
wire n_2718;
wire n_3019;
wire n_2639;
wire n_1183;
wire n_1436;
wire n_2898;
wire n_2251;
wire n_1384;
wire n_2494;
wire n_2959;
wire n_2501;
wire n_3203;
wire n_2238;
wire n_2368;
wire n_1070;
wire n_2403;
wire n_2837;
wire n_998;
wire n_3200;
wire n_1665;
wire n_3259;
wire n_2524;
wire n_3167;
wire n_1383;
wire n_2460;
wire n_1178;
wire n_2127;
wire n_1424;
wire n_2338;
wire n_1073;
wire n_1000;
wire n_1195;
wire n_3025;
wire n_2137;
wire n_1626;
wire n_3191;
wire n_1507;
wire n_2482;
wire n_2532;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_3006;
wire n_2481;
wire n_1857;
wire n_1519;
wire n_2144;
wire n_3056;
wire n_1284;
wire n_1604;
wire n_2296;
wire n_2424;
wire n_3201;
wire n_1142;
wire n_2849;
wire n_1475;
wire n_1774;
wire n_1048;
wire n_1398;
wire n_1201;
wire n_2354;
wire n_2682;
wire n_3032;
wire n_3103;
wire n_2589;
wire n_1395;
wire n_2110;
wire n_2199;
wire n_2661;
wire n_2877;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_931;
wire n_1021;
wire n_2442;
wire n_1207;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_3072;
wire n_3087;
wire n_2053;
wire n_2259;
wire n_2121;
wire n_2773;
wire n_2545;
wire n_2432;
wire n_2710;
wire n_1478;
wire n_1310;
wire n_3142;
wire n_2966;
wire n_2294;
wire n_1363;
wire n_2581;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_1314;
wire n_1837;
wire n_964;
wire n_2218;
wire n_2788;
wire n_3196;
wire n_2435;
wire n_954;
wire n_2504;
wire n_2797;
wire n_2623;
wire n_1110;
wire n_2213;
wire n_1410;
wire n_2389;
wire n_1440;
wire n_2132;
wire n_2892;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_2748;
wire n_1483;
wire n_1834;
wire n_2331;
wire n_1372;
wire n_2292;
wire n_2860;
wire n_2330;
wire n_1457;
wire n_1719;
wire n_1339;
wire n_1787;
wire n_2701;
wire n_2475;
wire n_2511;
wire n_1993;
wire n_2281;
wire n_1427;
wire n_2416;
wire n_2745;
wire n_2617;
wire n_2776;
wire n_1466;
wire n_1919;
wire n_1080;
wire n_1877;
wire n_3144;
wire n_3211;
wire n_3244;
wire n_1141;
wire n_1268;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_2323;
wire n_1893;
wire n_2784;
wire n_2209;
wire n_2301;
wire n_3287;
wire n_2387;
wire n_1755;
wire n_1602;
wire n_2421;
wire n_1136;
wire n_3270;
wire n_2618;
wire n_2025;
wire n_2357;
wire n_2846;
wire n_2464;
wire n_3265;
wire n_1125;
wire n_970;
wire n_3306;
wire n_2488;
wire n_2224;
wire n_1980;
wire n_995;
wire n_1159;
wire n_2329;
wire n_1092;
wire n_2237;
wire n_3026;
wire n_1060;
wire n_1951;
wire n_2250;
wire n_3090;
wire n_3033;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_2990;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_2115;
wire n_2410;
wire n_2552;
wire n_1053;
wire n_3302;
wire n_2374;
wire n_1681;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_2929;
wire n_2780;
wire n_3226;
wire n_2596;
wire n_2274;
wire n_3163;
wire n_1153;
wire n_1618;
wire n_1531;
wire n_2828;
wire n_1185;
wire n_2384;
wire n_1745;
wire n_3127;
wire n_2724;
wire n_1831;
wire n_2585;
wire n_2621;
wire n_1653;
wire n_2352;
wire n_1679;
wire n_1625;
wire n_2601;
wire n_2160;
wire n_1453;
wire n_2146;
wire n_2226;
wire n_2131;
wire n_2502;
wire n_2801;
wire n_2920;
wire n_1901;
wire n_920;
wire n_1374;
wire n_2556;
wire n_2648;
wire n_3212;
wire n_1315;
wire n_1647;
wire n_2575;
wire n_2754;
wire n_1224;
wire n_2783;
wire n_2306;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_3188;
wire n_1933;
wire n_2462;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_2889;
wire n_3243;
wire n_1617;
wire n_3260;
wire n_1470;
wire n_2550;
wire n_3093;
wire n_3175;
wire n_3214;
wire n_1243;
wire n_2732;
wire n_2928;
wire n_1096;
wire n_2249;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_2227;
wire n_2270;
wire n_2822;
wire n_1425;
wire n_3169;
wire n_3205;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_3284;
wire n_983;
wire n_3109;
wire n_2023;
wire n_2572;
wire n_2204;
wire n_1520;
wire n_2720;
wire n_3126;
wire n_2159;
wire n_1390;
wire n_2289;
wire n_1077;
wire n_1733;
wire n_2315;
wire n_1419;
wire n_2863;
wire n_3299;
wire n_2955;
wire n_2995;
wire n_1731;
wire n_2158;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_3051;
wire n_1437;
wire n_2135;
wire n_1645;
wire n_1832;
wire n_1687;
wire n_1439;
wire n_2328;
wire n_1323;
wire n_2859;
wire n_2202;
wire n_2049;
wire n_1331;
wire n_2627;
wire n_956;
wire n_960;
wire n_2276;
wire n_3234;
wire n_2803;
wire n_2100;
wire n_2993;
wire n_1668;
wire n_2777;
wire n_1134;
wire n_3016;
wire n_3004;
wire n_3202;
wire n_2830;
wire n_2781;
wire n_3220;
wire n_1129;
wire n_2829;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_2181;
wire n_1869;
wire n_2911;
wire n_1764;
wire n_1429;
wire n_2826;
wire n_1610;
wire n_3084;
wire n_1889;
wire n_2379;
wire n_2016;
wire n_1905;
wire n_2343;
wire n_1593;
wire n_1202;
wire n_1030;
wire n_1937;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_2942;
wire n_1079;
wire n_2515;
wire n_1744;
wire n_2139;
wire n_2142;
wire n_1551;
wire n_2448;
wire n_1103;
wire n_2875;
wire n_2555;
wire n_2219;
wire n_1203;
wire n_2851;
wire n_2327;
wire n_951;
wire n_2201;
wire n_952;
wire n_999;
wire n_1254;
wire n_2841;
wire n_2420;
wire n_2984;
wire n_994;
wire n_2263;
wire n_3291;
wire n_2304;
wire n_1508;
wire n_2487;
wire n_974;
wire n_2983;
wire n_2240;
wire n_2278;
wire n_2656;
wire n_2538;
wire n_2597;
wire n_2375;
wire n_3113;
wire n_3194;
wire n_3250;
wire n_1934;
wire n_3276;
wire n_1020;
wire n_1042;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_2756;
wire n_1871;
wire n_2924;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_2884;
wire n_1549;
wire n_1510;
wire n_3120;
wire n_1468;
wire n_2855;
wire n_1859;
wire n_2102;
wire n_2563;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_2156;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_2598;
wire n_1270;
wire n_2549;
wire n_1187;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_2153;
wire n_2544;
wire n_2381;
wire n_2052;
wire n_1847;
wire n_2302;
wire n_1667;
wire n_1206;
wire n_3230;
wire n_1037;
wire n_1397;
wire n_3268;
wire n_3236;
wire n_1279;
wire n_1115;
wire n_1499;
wire n_2755;
wire n_3141;
wire n_923;
wire n_1409;
wire n_1841;
wire n_2637;
wire n_2823;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_3112;
wire n_2819;
wire n_3195;
wire n_2526;
wire n_3041;
wire n_2423;
wire n_1057;
wire n_3277;
wire n_3108;
wire n_2548;
wire n_991;
wire n_2785;
wire n_1657;
wire n_1126;
wire n_2412;
wire n_1997;
wire n_2636;
wire n_3131;
wire n_2439;
wire n_1108;
wire n_1818;
wire n_2404;
wire n_1182;
wire n_1298;
wire n_2559;
wire n_2177;
wire n_2595;
wire n_2088;
wire n_1611;
wire n_2740;
wire n_1601;
wire n_3011;
wire n_1960;
wire n_2694;
wire n_2061;
wire n_1686;
wire n_2757;
wire n_2337;
wire n_2401;
wire n_1356;
wire n_1589;
wire n_3042;
wire n_3213;
wire n_2309;
wire n_2900;
wire n_2957;
wire n_2607;
wire n_1740;
wire n_2737;
wire n_1497;
wire n_2890;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_3228;
wire n_1320;
wire n_2716;
wire n_3249;
wire n_3081;
wire n_2452;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_2722;
wire n_1452;
wire n_2854;
wire n_3010;
wire n_2499;
wire n_3043;
wire n_1622;
wire n_1586;
wire n_2543;
wire n_2264;
wire n_1694;
wire n_1535;
wire n_3137;
wire n_2486;
wire n_3132;
wire n_2571;
wire n_3138;
wire n_1596;
wire n_3177;
wire n_1190;
wire n_1734;
wire n_3172;
wire n_2902;
wire n_3217;
wire n_1983;
wire n_1938;
wire n_2498;
wire n_2220;
wire n_2577;
wire n_1262;
wire n_2472;
wire n_1891;
wire n_2171;
wire n_1213;
wire n_3238;
wire n_2235;
wire n_2988;
wire n_3136;
wire n_1350;
wire n_1673;
wire n_2232;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_2392;
wire n_2894;
wire n_2790;
wire n_2037;
wire n_2808;
wire n_2298;
wire n_2326;
wire n_1539;
wire n_1043;
wire n_3040;
wire n_1797;
wire n_3279;
wire n_1608;
wire n_986;
wire n_2305;
wire n_2120;
wire n_1472;
wire n_2050;
wire n_2373;
wire n_2164;
wire n_2402;
wire n_2225;
wire n_1081;
wire n_1870;
wire n_2964;
wire n_1692;
wire n_1084;
wire n_1171;
wire n_2169;
wire n_2371;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_2187;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_3262;
wire n_2904;
wire n_2244;
wire n_3013;
wire n_2586;
wire n_1684;
wire n_921;
wire n_2446;
wire n_1346;
wire n_1642;
wire n_1352;
wire n_2789;
wire n_3105;
wire n_3210;
wire n_2872;
wire n_937;
wire n_2257;
wire n_1682;
wire n_2017;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_2272;
wire n_2699;
wire n_2200;
wire n_3029;
wire n_1046;
wire n_2560;
wire n_1940;
wire n_1979;
wire n_2760;
wire n_2704;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_2738;
wire n_1405;
wire n_972;
wire n_2376;
wire n_1406;
wire n_2766;
wire n_1332;
wire n_2670;
wire n_2700;
wire n_962;
wire n_1041;
wire n_2346;
wire n_3134;
wire n_1569;
wire n_936;
wire n_3045;
wire n_3115;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_3278;
wire n_2342;
wire n_2167;
wire n_2084;
wire n_2970;
wire n_2882;
wire n_2541;
wire n_2940;
wire n_2518;
wire n_2458;
wire n_1222;
wire n_1823;
wire n_2479;
wire n_3050;
wire n_2782;
wire n_1974;
wire n_2673;
wire n_2456;
wire n_1720;
wire n_2527;
wire n_934;
wire n_1637;
wire n_2635;
wire n_1407;
wire n_1795;
wire n_2768;
wire n_2871;
wire n_2688;
wire n_1341;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_2314;
wire n_942;
wire n_3003;
wire n_2798;
wire n_2852;
wire n_1524;
wire n_2229;
wire n_1964;
wire n_2288;
wire n_1920;
wire n_2753;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_3292;
wire n_1545;
wire n_2007;
wire n_3121;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_3184;
wire n_1544;
wire n_1485;
wire n_2258;
wire n_1640;
wire n_1846;
wire n_3245;
wire n_3075;
wire n_2406;
wire n_2390;
wire n_959;
wire n_2310;
wire n_2506;
wire n_2141;
wire n_2562;
wire n_2642;
wire n_1343;
wire n_1522;
wire n_2734;
wire n_1782;
wire n_2383;
wire n_2626;
wire n_1676;
wire n_1830;
wire n_2351;
wire n_1567;
wire n_1319;
wire n_2986;
wire n_1900;
wire n_3246;
wire n_1548;
wire n_3044;
wire n_2973;
wire n_1155;
wire n_2536;
wire n_2196;
wire n_2629;
wire n_1633;
wire n_2195;
wire n_3208;
wire n_2809;
wire n_3007;
wire n_2172;
wire n_2835;
wire n_1416;
wire n_1528;
wire n_2820;
wire n_2293;
wire n_1146;
wire n_2021;
wire n_2454;
wire n_2114;
wire n_3074;
wire n_3174;
wire n_1086;
wire n_1066;
wire n_3102;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_1282;
wire n_2561;
wire n_2567;
wire n_2322;
wire n_2154;
wire n_2727;
wire n_2962;
wire n_2939;
wire n_1906;
wire n_1484;
wire n_2992;
wire n_3305;
wire n_1321;
wire n_1241;
wire n_1672;
wire n_2533;
wire n_3157;
wire n_1758;
wire n_3221;
wire n_3267;
wire n_2283;
wire n_2869;
wire n_2422;
wire n_1925;
wire n_1914;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_2759;
wire n_2945;
wire n_3061;
wire n_2361;
wire n_1373;
wire n_1292;
wire n_2266;
wire n_2960;
wire n_3005;
wire n_2427;
wire n_3151;
wire n_1029;
wire n_1447;
wire n_2388;
wire n_2056;
wire n_2611;
wire n_2901;
wire n_3258;
wire n_1706;
wire n_1498;
wire n_3143;
wire n_2653;
wire n_2417;
wire n_3000;
wire n_1210;
wire n_1248;
wire n_1556;
wire n_2189;
wire n_2680;
wire n_2246;
wire n_1047;
wire n_3149;
wire n_1984;
wire n_2236;
wire n_1385;
wire n_3156;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_2834;
wire n_3207;
wire n_2668;
wire n_2441;
wire n_1257;
wire n_3008;
wire n_1751;
wire n_2840;
wire n_3197;
wire n_3242;
wire n_1375;
wire n_1941;
wire n_2128;
wire n_1045;
wire n_1794;
wire n_1650;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_2398;
wire n_1872;
wire n_3091;
wire n_2695;
wire n_3124;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_1949;
wire n_2888;
wire n_2671;
wire n_2761;
wire n_2885;
wire n_2793;
wire n_2715;
wire n_2923;
wire n_1804;
wire n_1727;
wire n_2508;
wire n_1019;
wire n_2054;
wire n_2845;
wire n_1337;
wire n_3097;
wire n_2062;
wire n_2041;
wire n_2975;
wire n_1477;
wire n_1360;
wire n_2839;
wire n_1860;
wire n_2856;
wire n_1904;
wire n_2874;
wire n_1200;
wire n_2070;
wire n_2588;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_2484;
wire n_2348;
wire n_2944;
wire n_2614;
wire n_2126;
wire n_1154;
wire n_1600;
wire n_1113;
wire n_2833;
wire n_2253;
wire n_2758;
wire n_2366;
wire n_1098;
wire n_2937;
wire n_1329;
wire n_2045;
wire n_2261;
wire n_2216;
wire n_2210;
wire n_3300;
wire n_2978;
wire n_2066;
wire n_1476;
wire n_2516;
wire n_1001;
wire n_1800;
wire n_2241;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_2903;
wire n_2827;
wire n_1177;
wire n_3216;
wire n_1150;
wire n_3190;
wire n_1562;
wire n_1690;
wire n_1191;
wire n_1826;
wire n_1023;
wire n_1882;
wire n_2951;
wire n_1118;
wire n_1076;
wire n_2949;
wire n_1807;
wire n_1007;
wire n_1929;
wire n_1378;
wire n_2369;
wire n_1592;
wire n_1759;
wire n_2719;
wire n_1814;
wire n_1631;
wire n_1377;
wire n_1879;
wire n_1542;
wire n_2587;
wire n_3199;
wire n_2931;
wire n_1678;
wire n_2569;
wire n_2400;
wire n_1716;
wire n_1256;
wire n_1953;
wire n_933;
wire n_3303;
wire n_978;
wire n_2752;
wire n_3135;
wire n_1976;
wire n_2905;
wire n_1291;
wire n_1217;
wire n_1824;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_1435;
wire n_969;
wire n_988;
wire n_2140;
wire n_3160;
wire n_1065;
wire n_2796;
wire n_3255;
wire n_2507;
wire n_1401;
wire n_2358;
wire n_1255;
wire n_1516;
wire n_1536;
wire n_2186;
wire n_2163;
wire n_2029;
wire n_2815;
wire n_1204;
wire n_3034;
wire n_1132;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_955;
wire n_1379;
wire n_2528;
wire n_2814;
wire n_2787;
wire n_1338;
wire n_1097;
wire n_2969;
wire n_2395;
wire n_935;
wire n_3027;
wire n_1554;
wire n_3231;
wire n_1130;
wire n_3083;
wire n_2979;
wire n_1810;
wire n_2953;
wire n_2380;
wire n_1120;
wire n_1583;
wire n_3049;
wire n_1730;
wire n_2295;
wire n_2746;
wire n_2946;
wire n_1643;
wire n_2020;
wire n_2500;
wire n_2269;
wire n_1729;
wire n_2290;
wire n_2048;
wire n_2005;
wire n_2565;
wire n_1389;
wire n_1105;
wire n_3117;
wire n_1461;
wire n_2076;
wire n_2736;
wire n_2883;
wire n_1408;
wire n_1196;
wire n_1598;
wire n_2935;
wire n_3015;
wire n_2175;
wire n_2182;
wire n_2910;
wire n_1283;
wire n_2385;
wire n_918;
wire n_1848;
wire n_1114;
wire n_1785;
wire n_1147;
wire n_1754;
wire n_2149;
wire n_3057;
wire n_3154;
wire n_2396;
wire n_1506;
wire n_2584;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_1227;
wire n_2485;
wire n_2450;
wire n_2284;
wire n_2566;
wire n_2287;
wire n_971;
wire n_2702;
wire n_3241;
wire n_946;
wire n_2906;
wire n_1303;
wire n_2769;
wire n_1205;
wire n_2492;
wire n_1258;
wire n_2438;
wire n_2914;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_2463;
wire n_2881;
wire n_1677;
wire n_1116;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_3064;
wire n_1780;
wire n_3100;
wire n_1689;
wire n_2180;
wire n_2858;
wire n_3062;
wire n_2679;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_3215;
wire n_2952;
wire n_1017;
wire n_3068;
wire n_2117;
wire n_2234;
wire n_2779;
wire n_2685;
wire n_1083;
wire n_1561;
wire n_2741;
wire n_3114;
wire n_930;
wire n_2275;
wire n_1112;
wire n_2465;
wire n_2620;
wire n_2081;
wire n_2168;
wire n_2568;
wire n_2022;
wire n_1945;
wire n_2203;
wire n_1721;
wire n_1656;
wire n_1460;
wire n_2112;
wire n_2255;
wire n_1464;
wire n_1737;
wire n_2430;
wire n_1414;
wire n_2649;
wire n_2721;
wire n_944;
wire n_2034;
wire n_1028;
wire n_2106;
wire n_2862;
wire n_2265;
wire n_2615;
wire n_2683;
wire n_1922;
wire n_2032;
wire n_2744;
wire n_1011;
wire n_2474;
wire n_1566;
wire n_1215;
wire n_2444;
wire n_2437;
wire n_2743;
wire n_1973;
wire n_3181;
wire n_2267;
wire n_3035;
wire n_990;
wire n_1500;
wire n_1537;
wire n_1821;
wire n_2205;
wire n_3204;
wire n_1104;
wire n_1058;
wire n_2312;
wire n_1122;
wire n_1253;
wire n_1266;
wire n_2242;
wire n_1509;
wire n_1693;
wire n_2934;
wire n_3290;
wire n_1109;
wire n_2222;
wire n_3256;
wire n_1276;
wire n_3176;
wire n_2015;
wire n_2118;
wire n_2111;
wire n_2466;
wire n_2915;
wire n_2530;
wire n_1148;
wire n_2188;
wire n_2505;
wire n_1989;
wire n_1161;
wire n_2609;
wire n_1085;
wire n_2802;
wire n_2999;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_1584;
wire n_2425;
wire n_924;
wire n_1582;
wire n_2318;
wire n_3286;
wire n_2408;
wire n_1149;
wire n_3170;
wire n_1184;
wire n_2483;
wire n_2950;
wire n_1972;
wire n_3060;
wire n_3304;
wire n_2592;
wire n_1525;
wire n_3098;
wire n_2594;
wire n_2666;
wire n_1585;
wire n_1851;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_2564;
wire n_1816;
wire n_2503;
wire n_2433;
wire n_1518;
wire n_1362;
wire n_1156;
wire n_3123;
wire n_2600;
wire n_984;
wire n_1829;
wire n_2035;
wire n_3024;
wire n_1450;
wire n_1638;
wire n_3038;
wire n_3086;
wire n_2033;
wire n_1789;
wire n_2531;
wire n_1770;
wire n_3285;
wire n_2523;
wire n_1218;
wire n_2413;
wire n_1482;
wire n_981;
wire n_1349;
wire n_1144;
wire n_2071;
wire n_3219;
wire n_2429;
wire n_3130;
wire n_985;
wire n_2233;
wire n_2440;
wire n_2723;
wire n_3233;
wire n_997;
wire n_1710;
wire n_2800;
wire n_2161;
wire n_1301;
wire n_2805;
wire n_980;
wire n_2681;
wire n_1306;
wire n_3264;
wire n_2010;
wire n_2282;
wire n_1651;
wire n_1198;
wire n_3096;
wire n_2360;
wire n_2047;
wire n_2651;
wire n_2095;
wire n_3239;
wire n_1609;
wire n_2174;
wire n_3161;
wire n_2799;
wire n_2334;
wire n_3295;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_3066;
wire n_1574;
wire n_2426;
wire n_2490;
wire n_2844;
wire n_3101;
wire n_2303;
wire n_1619;
wire n_2478;
wire n_1981;
wire n_2285;
wire n_1606;
wire n_1133;
wire n_1194;
wire n_2742;
wire n_2640;
wire n_1051;
wire n_1552;
wire n_2918;
wire n_3288;
wire n_1996;
wire n_2367;
wire n_2867;
wire n_3198;
wire n_1039;
wire n_1442;
wire n_2726;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_3125;
wire n_1158;
wire n_2909;
wire n_2248;
wire n_941;
wire n_975;
wire n_3206;
wire n_1031;
wire n_1305;
wire n_2363;
wire n_2578;
wire n_2662;
wire n_3147;
wire n_3116;
wire n_1753;
wire n_3095;
wire n_3180;
wire n_2795;
wire n_2471;
wire n_3187;
wire n_2540;
wire n_973;
wire n_2807;
wire n_1921;
wire n_3218;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_2217;
wire n_2197;
wire n_2065;
wire n_2879;
wire n_967;
wire n_2215;
wire n_2461;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_2968;
wire n_1170;
wire n_1629;
wire n_2221;
wire n_1260;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_2553;
wire n_1040;
wire n_915;
wire n_3059;
wire n_1166;
wire n_2038;
wire n_2891;
wire n_1131;
wire n_2634;
wire n_1761;
wire n_2709;
wire n_3155;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_3110;
wire n_1632;
wire n_1890;
wire n_3017;
wire n_1805;
wire n_2477;
wire n_1888;
wire n_1557;
wire n_2280;
wire n_1833;
wire n_1311;
wire n_1494;
wire n_2325;
wire n_1850;
wire n_1898;
wire n_2443;
wire n_2697;
wire n_3235;
wire n_2308;
wire n_2162;
wire n_1868;
wire n_2333;
wire n_2079;
wire n_3001;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_2512;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_2086;
wire n_2185;
wire n_2927;
wire n_1836;
wire n_2774;
wire n_3039;
wire n_1226;
wire n_3162;
wire n_1274;
wire n_1486;
wire n_2166;
wire n_3094;
wire n_2899;
wire n_3274;
wire n_3186;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_1958;
wire n_2077;
wire n_1059;
wire n_1197;
wire n_3065;
wire n_2632;
wire n_2579;
wire n_2105;
wire n_3079;
wire n_2098;
wire n_3085;
wire n_1423;
wire n_2813;
wire n_1935;
wire n_2027;
wire n_3070;
wire n_2223;
wire n_2091;
wire n_3263;
wire n_2991;
wire n_1915;
wire n_1621;
wire n_1748;
wire n_2547;
wire n_2415;
wire n_1449;
wire n_2912;
wire n_2659;
wire n_2930;
wire n_1025;
wire n_2419;
wire n_3111;
wire n_2116;
wire n_2320;
wire n_1885;
wire n_2677;
wire n_1013;
wire n_3182;
wire n_1259;
wire n_3054;
wire n_3283;
wire n_2183;
wire n_3002;
wire n_1538;
wire n_1742;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g915 ( 
.A(n_640),
.Y(n_915)
);

CKINVDCx5p33_ASAP7_75t_R g916 ( 
.A(n_856),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_894),
.Y(n_917)
);

BUFx3_ASAP7_75t_L g918 ( 
.A(n_343),
.Y(n_918)
);

CKINVDCx5p33_ASAP7_75t_R g919 ( 
.A(n_897),
.Y(n_919)
);

CKINVDCx5p33_ASAP7_75t_R g920 ( 
.A(n_475),
.Y(n_920)
);

CKINVDCx5p33_ASAP7_75t_R g921 ( 
.A(n_213),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_892),
.Y(n_922)
);

CKINVDCx5p33_ASAP7_75t_R g923 ( 
.A(n_568),
.Y(n_923)
);

CKINVDCx5p33_ASAP7_75t_R g924 ( 
.A(n_653),
.Y(n_924)
);

CKINVDCx20_ASAP7_75t_R g925 ( 
.A(n_794),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_723),
.Y(n_926)
);

CKINVDCx5p33_ASAP7_75t_R g927 ( 
.A(n_783),
.Y(n_927)
);

CKINVDCx5p33_ASAP7_75t_R g928 ( 
.A(n_492),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_730),
.Y(n_929)
);

CKINVDCx5p33_ASAP7_75t_R g930 ( 
.A(n_364),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_392),
.Y(n_931)
);

CKINVDCx5p33_ASAP7_75t_R g932 ( 
.A(n_843),
.Y(n_932)
);

CKINVDCx5p33_ASAP7_75t_R g933 ( 
.A(n_790),
.Y(n_933)
);

CKINVDCx5p33_ASAP7_75t_R g934 ( 
.A(n_699),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_860),
.Y(n_935)
);

CKINVDCx5p33_ASAP7_75t_R g936 ( 
.A(n_583),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_152),
.Y(n_937)
);

INVx2_ASAP7_75t_L g938 ( 
.A(n_765),
.Y(n_938)
);

BUFx6f_ASAP7_75t_L g939 ( 
.A(n_478),
.Y(n_939)
);

CKINVDCx5p33_ASAP7_75t_R g940 ( 
.A(n_775),
.Y(n_940)
);

BUFx6f_ASAP7_75t_L g941 ( 
.A(n_728),
.Y(n_941)
);

CKINVDCx5p33_ASAP7_75t_R g942 ( 
.A(n_23),
.Y(n_942)
);

CKINVDCx12_ASAP7_75t_R g943 ( 
.A(n_637),
.Y(n_943)
);

INVx2_ASAP7_75t_SL g944 ( 
.A(n_803),
.Y(n_944)
);

INVx2_ASAP7_75t_SL g945 ( 
.A(n_810),
.Y(n_945)
);

CKINVDCx5p33_ASAP7_75t_R g946 ( 
.A(n_625),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_508),
.Y(n_947)
);

CKINVDCx5p33_ASAP7_75t_R g948 ( 
.A(n_777),
.Y(n_948)
);

CKINVDCx20_ASAP7_75t_R g949 ( 
.A(n_908),
.Y(n_949)
);

CKINVDCx5p33_ASAP7_75t_R g950 ( 
.A(n_795),
.Y(n_950)
);

CKINVDCx5p33_ASAP7_75t_R g951 ( 
.A(n_757),
.Y(n_951)
);

CKINVDCx5p33_ASAP7_75t_R g952 ( 
.A(n_887),
.Y(n_952)
);

CKINVDCx5p33_ASAP7_75t_R g953 ( 
.A(n_913),
.Y(n_953)
);

CKINVDCx5p33_ASAP7_75t_R g954 ( 
.A(n_838),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_479),
.Y(n_955)
);

CKINVDCx5p33_ASAP7_75t_R g956 ( 
.A(n_39),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_798),
.Y(n_957)
);

INVx2_ASAP7_75t_SL g958 ( 
.A(n_842),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_114),
.Y(n_959)
);

CKINVDCx5p33_ASAP7_75t_R g960 ( 
.A(n_24),
.Y(n_960)
);

CKINVDCx5p33_ASAP7_75t_R g961 ( 
.A(n_793),
.Y(n_961)
);

CKINVDCx5p33_ASAP7_75t_R g962 ( 
.A(n_634),
.Y(n_962)
);

CKINVDCx5p33_ASAP7_75t_R g963 ( 
.A(n_812),
.Y(n_963)
);

CKINVDCx5p33_ASAP7_75t_R g964 ( 
.A(n_586),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_71),
.Y(n_965)
);

CKINVDCx5p33_ASAP7_75t_R g966 ( 
.A(n_181),
.Y(n_966)
);

CKINVDCx20_ASAP7_75t_R g967 ( 
.A(n_679),
.Y(n_967)
);

CKINVDCx5p33_ASAP7_75t_R g968 ( 
.A(n_203),
.Y(n_968)
);

CKINVDCx20_ASAP7_75t_R g969 ( 
.A(n_697),
.Y(n_969)
);

CKINVDCx5p33_ASAP7_75t_R g970 ( 
.A(n_739),
.Y(n_970)
);

CKINVDCx20_ASAP7_75t_R g971 ( 
.A(n_161),
.Y(n_971)
);

CKINVDCx5p33_ASAP7_75t_R g972 ( 
.A(n_379),
.Y(n_972)
);

CKINVDCx5p33_ASAP7_75t_R g973 ( 
.A(n_752),
.Y(n_973)
);

CKINVDCx20_ASAP7_75t_R g974 ( 
.A(n_449),
.Y(n_974)
);

INVx1_ASAP7_75t_SL g975 ( 
.A(n_901),
.Y(n_975)
);

CKINVDCx5p33_ASAP7_75t_R g976 ( 
.A(n_893),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_885),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_857),
.Y(n_978)
);

BUFx3_ASAP7_75t_L g979 ( 
.A(n_802),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_822),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_776),
.Y(n_981)
);

BUFx5_ASAP7_75t_L g982 ( 
.A(n_796),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_809),
.Y(n_983)
);

CKINVDCx5p33_ASAP7_75t_R g984 ( 
.A(n_787),
.Y(n_984)
);

CKINVDCx5p33_ASAP7_75t_R g985 ( 
.A(n_761),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_316),
.Y(n_986)
);

CKINVDCx5p33_ASAP7_75t_R g987 ( 
.A(n_419),
.Y(n_987)
);

INVx2_ASAP7_75t_SL g988 ( 
.A(n_789),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_759),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_346),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_767),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_468),
.Y(n_992)
);

CKINVDCx5p33_ASAP7_75t_R g993 ( 
.A(n_263),
.Y(n_993)
);

CKINVDCx5p33_ASAP7_75t_R g994 ( 
.A(n_294),
.Y(n_994)
);

CKINVDCx5p33_ASAP7_75t_R g995 ( 
.A(n_154),
.Y(n_995)
);

CKINVDCx5p33_ASAP7_75t_R g996 ( 
.A(n_826),
.Y(n_996)
);

CKINVDCx5p33_ASAP7_75t_R g997 ( 
.A(n_876),
.Y(n_997)
);

CKINVDCx5p33_ASAP7_75t_R g998 ( 
.A(n_313),
.Y(n_998)
);

CKINVDCx5p33_ASAP7_75t_R g999 ( 
.A(n_855),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_153),
.Y(n_1000)
);

BUFx10_ASAP7_75t_L g1001 ( 
.A(n_907),
.Y(n_1001)
);

BUFx3_ASAP7_75t_L g1002 ( 
.A(n_59),
.Y(n_1002)
);

CKINVDCx5p33_ASAP7_75t_R g1003 ( 
.A(n_365),
.Y(n_1003)
);

CKINVDCx5p33_ASAP7_75t_R g1004 ( 
.A(n_274),
.Y(n_1004)
);

INVx2_ASAP7_75t_SL g1005 ( 
.A(n_483),
.Y(n_1005)
);

CKINVDCx5p33_ASAP7_75t_R g1006 ( 
.A(n_319),
.Y(n_1006)
);

INVx2_ASAP7_75t_L g1007 ( 
.A(n_845),
.Y(n_1007)
);

CKINVDCx5p33_ASAP7_75t_R g1008 ( 
.A(n_872),
.Y(n_1008)
);

BUFx6f_ASAP7_75t_L g1009 ( 
.A(n_881),
.Y(n_1009)
);

CKINVDCx5p33_ASAP7_75t_R g1010 ( 
.A(n_824),
.Y(n_1010)
);

INVxp67_ASAP7_75t_L g1011 ( 
.A(n_766),
.Y(n_1011)
);

CKINVDCx5p33_ASAP7_75t_R g1012 ( 
.A(n_424),
.Y(n_1012)
);

BUFx2_ASAP7_75t_L g1013 ( 
.A(n_813),
.Y(n_1013)
);

CKINVDCx5p33_ASAP7_75t_R g1014 ( 
.A(n_423),
.Y(n_1014)
);

BUFx3_ASAP7_75t_L g1015 ( 
.A(n_517),
.Y(n_1015)
);

CKINVDCx5p33_ASAP7_75t_R g1016 ( 
.A(n_779),
.Y(n_1016)
);

CKINVDCx5p33_ASAP7_75t_R g1017 ( 
.A(n_518),
.Y(n_1017)
);

BUFx8_ASAP7_75t_SL g1018 ( 
.A(n_764),
.Y(n_1018)
);

CKINVDCx5p33_ASAP7_75t_R g1019 ( 
.A(n_864),
.Y(n_1019)
);

INVxp67_ASAP7_75t_SL g1020 ( 
.A(n_199),
.Y(n_1020)
);

CKINVDCx5p33_ASAP7_75t_R g1021 ( 
.A(n_874),
.Y(n_1021)
);

CKINVDCx5p33_ASAP7_75t_R g1022 ( 
.A(n_904),
.Y(n_1022)
);

CKINVDCx5p33_ASAP7_75t_R g1023 ( 
.A(n_819),
.Y(n_1023)
);

CKINVDCx5p33_ASAP7_75t_R g1024 ( 
.A(n_556),
.Y(n_1024)
);

CKINVDCx5p33_ASAP7_75t_R g1025 ( 
.A(n_890),
.Y(n_1025)
);

INVxp67_ASAP7_75t_L g1026 ( 
.A(n_639),
.Y(n_1026)
);

CKINVDCx5p33_ASAP7_75t_R g1027 ( 
.A(n_624),
.Y(n_1027)
);

CKINVDCx20_ASAP7_75t_R g1028 ( 
.A(n_188),
.Y(n_1028)
);

CKINVDCx5p33_ASAP7_75t_R g1029 ( 
.A(n_623),
.Y(n_1029)
);

CKINVDCx5p33_ASAP7_75t_R g1030 ( 
.A(n_171),
.Y(n_1030)
);

CKINVDCx5p33_ASAP7_75t_R g1031 ( 
.A(n_769),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_891),
.Y(n_1032)
);

CKINVDCx5p33_ASAP7_75t_R g1033 ( 
.A(n_902),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_870),
.Y(n_1034)
);

CKINVDCx5p33_ASAP7_75t_R g1035 ( 
.A(n_286),
.Y(n_1035)
);

CKINVDCx5p33_ASAP7_75t_R g1036 ( 
.A(n_841),
.Y(n_1036)
);

INVx1_ASAP7_75t_SL g1037 ( 
.A(n_849),
.Y(n_1037)
);

CKINVDCx5p33_ASAP7_75t_R g1038 ( 
.A(n_205),
.Y(n_1038)
);

CKINVDCx5p33_ASAP7_75t_R g1039 ( 
.A(n_69),
.Y(n_1039)
);

CKINVDCx20_ASAP7_75t_R g1040 ( 
.A(n_259),
.Y(n_1040)
);

CKINVDCx5p33_ASAP7_75t_R g1041 ( 
.A(n_261),
.Y(n_1041)
);

CKINVDCx5p33_ASAP7_75t_R g1042 ( 
.A(n_792),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_176),
.Y(n_1043)
);

CKINVDCx5p33_ASAP7_75t_R g1044 ( 
.A(n_98),
.Y(n_1044)
);

CKINVDCx5p33_ASAP7_75t_R g1045 ( 
.A(n_116),
.Y(n_1045)
);

CKINVDCx5p33_ASAP7_75t_R g1046 ( 
.A(n_760),
.Y(n_1046)
);

CKINVDCx5p33_ASAP7_75t_R g1047 ( 
.A(n_521),
.Y(n_1047)
);

CKINVDCx5p33_ASAP7_75t_R g1048 ( 
.A(n_415),
.Y(n_1048)
);

CKINVDCx5p33_ASAP7_75t_R g1049 ( 
.A(n_350),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_563),
.Y(n_1050)
);

BUFx3_ASAP7_75t_L g1051 ( 
.A(n_436),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_633),
.Y(n_1052)
);

INVx1_ASAP7_75t_SL g1053 ( 
.A(n_246),
.Y(n_1053)
);

CKINVDCx5p33_ASAP7_75t_R g1054 ( 
.A(n_818),
.Y(n_1054)
);

INVx2_ASAP7_75t_L g1055 ( 
.A(n_905),
.Y(n_1055)
);

CKINVDCx5p33_ASAP7_75t_R g1056 ( 
.A(n_669),
.Y(n_1056)
);

CKINVDCx20_ASAP7_75t_R g1057 ( 
.A(n_117),
.Y(n_1057)
);

BUFx2_ASAP7_75t_L g1058 ( 
.A(n_846),
.Y(n_1058)
);

CKINVDCx5p33_ASAP7_75t_R g1059 ( 
.A(n_800),
.Y(n_1059)
);

INVx2_ASAP7_75t_SL g1060 ( 
.A(n_677),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_861),
.Y(n_1061)
);

CKINVDCx5p33_ASAP7_75t_R g1062 ( 
.A(n_797),
.Y(n_1062)
);

CKINVDCx5p33_ASAP7_75t_R g1063 ( 
.A(n_104),
.Y(n_1063)
);

CKINVDCx5p33_ASAP7_75t_R g1064 ( 
.A(n_368),
.Y(n_1064)
);

BUFx3_ASAP7_75t_L g1065 ( 
.A(n_119),
.Y(n_1065)
);

CKINVDCx5p33_ASAP7_75t_R g1066 ( 
.A(n_869),
.Y(n_1066)
);

CKINVDCx5p33_ASAP7_75t_R g1067 ( 
.A(n_361),
.Y(n_1067)
);

CKINVDCx5p33_ASAP7_75t_R g1068 ( 
.A(n_840),
.Y(n_1068)
);

CKINVDCx5p33_ASAP7_75t_R g1069 ( 
.A(n_820),
.Y(n_1069)
);

CKINVDCx5p33_ASAP7_75t_R g1070 ( 
.A(n_879),
.Y(n_1070)
);

CKINVDCx5p33_ASAP7_75t_R g1071 ( 
.A(n_873),
.Y(n_1071)
);

CKINVDCx5p33_ASAP7_75t_R g1072 ( 
.A(n_863),
.Y(n_1072)
);

CKINVDCx5p33_ASAP7_75t_R g1073 ( 
.A(n_770),
.Y(n_1073)
);

BUFx2_ASAP7_75t_SL g1074 ( 
.A(n_118),
.Y(n_1074)
);

INVx2_ASAP7_75t_L g1075 ( 
.A(n_829),
.Y(n_1075)
);

CKINVDCx5p33_ASAP7_75t_R g1076 ( 
.A(n_774),
.Y(n_1076)
);

BUFx6f_ASAP7_75t_L g1077 ( 
.A(n_200),
.Y(n_1077)
);

BUFx8_ASAP7_75t_SL g1078 ( 
.A(n_834),
.Y(n_1078)
);

CKINVDCx5p33_ASAP7_75t_R g1079 ( 
.A(n_763),
.Y(n_1079)
);

CKINVDCx5p33_ASAP7_75t_R g1080 ( 
.A(n_896),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_710),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_806),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_731),
.Y(n_1083)
);

INVx2_ASAP7_75t_L g1084 ( 
.A(n_836),
.Y(n_1084)
);

CKINVDCx5p33_ASAP7_75t_R g1085 ( 
.A(n_456),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_835),
.Y(n_1086)
);

INVx2_ASAP7_75t_SL g1087 ( 
.A(n_853),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_498),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_276),
.Y(n_1089)
);

CKINVDCx5p33_ASAP7_75t_R g1090 ( 
.A(n_663),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_295),
.Y(n_1091)
);

CKINVDCx5p33_ASAP7_75t_R g1092 ( 
.A(n_424),
.Y(n_1092)
);

BUFx6f_ASAP7_75t_L g1093 ( 
.A(n_744),
.Y(n_1093)
);

CKINVDCx5p33_ASAP7_75t_R g1094 ( 
.A(n_40),
.Y(n_1094)
);

CKINVDCx5p33_ASAP7_75t_R g1095 ( 
.A(n_815),
.Y(n_1095)
);

CKINVDCx5p33_ASAP7_75t_R g1096 ( 
.A(n_634),
.Y(n_1096)
);

CKINVDCx5p33_ASAP7_75t_R g1097 ( 
.A(n_871),
.Y(n_1097)
);

CKINVDCx16_ASAP7_75t_R g1098 ( 
.A(n_642),
.Y(n_1098)
);

BUFx5_ASAP7_75t_L g1099 ( 
.A(n_771),
.Y(n_1099)
);

CKINVDCx5p33_ASAP7_75t_R g1100 ( 
.A(n_823),
.Y(n_1100)
);

CKINVDCx5p33_ASAP7_75t_R g1101 ( 
.A(n_581),
.Y(n_1101)
);

CKINVDCx5p33_ASAP7_75t_R g1102 ( 
.A(n_490),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_828),
.Y(n_1103)
);

CKINVDCx5p33_ASAP7_75t_R g1104 ( 
.A(n_471),
.Y(n_1104)
);

CKINVDCx20_ASAP7_75t_R g1105 ( 
.A(n_626),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_886),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_900),
.Y(n_1107)
);

CKINVDCx5p33_ASAP7_75t_R g1108 ( 
.A(n_635),
.Y(n_1108)
);

CKINVDCx5p33_ASAP7_75t_R g1109 ( 
.A(n_158),
.Y(n_1109)
);

CKINVDCx5p33_ASAP7_75t_R g1110 ( 
.A(n_289),
.Y(n_1110)
);

INVx2_ASAP7_75t_SL g1111 ( 
.A(n_630),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_868),
.Y(n_1112)
);

CKINVDCx5p33_ASAP7_75t_R g1113 ( 
.A(n_883),
.Y(n_1113)
);

CKINVDCx5p33_ASAP7_75t_R g1114 ( 
.A(n_39),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_727),
.Y(n_1115)
);

CKINVDCx5p33_ASAP7_75t_R g1116 ( 
.A(n_203),
.Y(n_1116)
);

BUFx5_ASAP7_75t_L g1117 ( 
.A(n_854),
.Y(n_1117)
);

BUFx10_ASAP7_75t_L g1118 ( 
.A(n_307),
.Y(n_1118)
);

CKINVDCx5p33_ASAP7_75t_R g1119 ( 
.A(n_281),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_647),
.Y(n_1120)
);

CKINVDCx20_ASAP7_75t_R g1121 ( 
.A(n_564),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_218),
.Y(n_1122)
);

CKINVDCx5p33_ASAP7_75t_R g1123 ( 
.A(n_305),
.Y(n_1123)
);

CKINVDCx5p33_ASAP7_75t_R g1124 ( 
.A(n_756),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_831),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_163),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_707),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_244),
.Y(n_1128)
);

CKINVDCx5p33_ASAP7_75t_R g1129 ( 
.A(n_518),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_825),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_67),
.Y(n_1131)
);

BUFx3_ASAP7_75t_L g1132 ( 
.A(n_460),
.Y(n_1132)
);

CKINVDCx5p33_ASAP7_75t_R g1133 ( 
.A(n_395),
.Y(n_1133)
);

CKINVDCx5p33_ASAP7_75t_R g1134 ( 
.A(n_599),
.Y(n_1134)
);

CKINVDCx5p33_ASAP7_75t_R g1135 ( 
.A(n_430),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_808),
.Y(n_1136)
);

CKINVDCx5p33_ASAP7_75t_R g1137 ( 
.A(n_76),
.Y(n_1137)
);

CKINVDCx5p33_ASAP7_75t_R g1138 ( 
.A(n_844),
.Y(n_1138)
);

CKINVDCx5p33_ASAP7_75t_R g1139 ( 
.A(n_882),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_617),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_158),
.Y(n_1141)
);

INVx1_ASAP7_75t_SL g1142 ( 
.A(n_267),
.Y(n_1142)
);

CKINVDCx5p33_ASAP7_75t_R g1143 ( 
.A(n_814),
.Y(n_1143)
);

CKINVDCx5p33_ASAP7_75t_R g1144 ( 
.A(n_490),
.Y(n_1144)
);

INVx2_ASAP7_75t_L g1145 ( 
.A(n_762),
.Y(n_1145)
);

CKINVDCx5p33_ASAP7_75t_R g1146 ( 
.A(n_426),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_608),
.Y(n_1147)
);

CKINVDCx20_ASAP7_75t_R g1148 ( 
.A(n_805),
.Y(n_1148)
);

CKINVDCx5p33_ASAP7_75t_R g1149 ( 
.A(n_6),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_571),
.Y(n_1150)
);

CKINVDCx5p33_ASAP7_75t_R g1151 ( 
.A(n_827),
.Y(n_1151)
);

BUFx3_ASAP7_75t_L g1152 ( 
.A(n_743),
.Y(n_1152)
);

CKINVDCx16_ASAP7_75t_R g1153 ( 
.A(n_472),
.Y(n_1153)
);

INVx1_ASAP7_75t_SL g1154 ( 
.A(n_135),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_458),
.Y(n_1155)
);

CKINVDCx5p33_ASAP7_75t_R g1156 ( 
.A(n_628),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_116),
.Y(n_1157)
);

INVx2_ASAP7_75t_L g1158 ( 
.A(n_638),
.Y(n_1158)
);

BUFx10_ASAP7_75t_L g1159 ( 
.A(n_583),
.Y(n_1159)
);

CKINVDCx5p33_ASAP7_75t_R g1160 ( 
.A(n_592),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_541),
.Y(n_1161)
);

CKINVDCx5p33_ASAP7_75t_R g1162 ( 
.A(n_702),
.Y(n_1162)
);

CKINVDCx20_ASAP7_75t_R g1163 ( 
.A(n_632),
.Y(n_1163)
);

CKINVDCx5p33_ASAP7_75t_R g1164 ( 
.A(n_867),
.Y(n_1164)
);

CKINVDCx5p33_ASAP7_75t_R g1165 ( 
.A(n_629),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_459),
.Y(n_1166)
);

CKINVDCx5p33_ASAP7_75t_R g1167 ( 
.A(n_548),
.Y(n_1167)
);

INVxp67_ASAP7_75t_L g1168 ( 
.A(n_865),
.Y(n_1168)
);

CKINVDCx5p33_ASAP7_75t_R g1169 ( 
.A(n_866),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_875),
.Y(n_1170)
);

INVx1_ASAP7_75t_SL g1171 ( 
.A(n_592),
.Y(n_1171)
);

CKINVDCx5p33_ASAP7_75t_R g1172 ( 
.A(n_258),
.Y(n_1172)
);

INVx2_ASAP7_75t_L g1173 ( 
.A(n_295),
.Y(n_1173)
);

CKINVDCx5p33_ASAP7_75t_R g1174 ( 
.A(n_282),
.Y(n_1174)
);

HB1xp67_ASAP7_75t_L g1175 ( 
.A(n_343),
.Y(n_1175)
);

INVx2_ASAP7_75t_L g1176 ( 
.A(n_75),
.Y(n_1176)
);

CKINVDCx5p33_ASAP7_75t_R g1177 ( 
.A(n_785),
.Y(n_1177)
);

CKINVDCx5p33_ASAP7_75t_R g1178 ( 
.A(n_833),
.Y(n_1178)
);

BUFx6f_ASAP7_75t_L g1179 ( 
.A(n_593),
.Y(n_1179)
);

CKINVDCx5p33_ASAP7_75t_R g1180 ( 
.A(n_791),
.Y(n_1180)
);

CKINVDCx5p33_ASAP7_75t_R g1181 ( 
.A(n_898),
.Y(n_1181)
);

CKINVDCx5p33_ASAP7_75t_R g1182 ( 
.A(n_817),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_772),
.Y(n_1183)
);

CKINVDCx5p33_ASAP7_75t_R g1184 ( 
.A(n_375),
.Y(n_1184)
);

CKINVDCx5p33_ASAP7_75t_R g1185 ( 
.A(n_557),
.Y(n_1185)
);

INVx1_ASAP7_75t_SL g1186 ( 
.A(n_326),
.Y(n_1186)
);

CKINVDCx5p33_ASAP7_75t_R g1187 ( 
.A(n_906),
.Y(n_1187)
);

CKINVDCx5p33_ASAP7_75t_R g1188 ( 
.A(n_830),
.Y(n_1188)
);

CKINVDCx5p33_ASAP7_75t_R g1189 ( 
.A(n_895),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_851),
.Y(n_1190)
);

BUFx6f_ASAP7_75t_L g1191 ( 
.A(n_850),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_862),
.Y(n_1192)
);

BUFx10_ASAP7_75t_L g1193 ( 
.A(n_636),
.Y(n_1193)
);

CKINVDCx5p33_ASAP7_75t_R g1194 ( 
.A(n_222),
.Y(n_1194)
);

CKINVDCx5p33_ASAP7_75t_R g1195 ( 
.A(n_84),
.Y(n_1195)
);

BUFx5_ASAP7_75t_L g1196 ( 
.A(n_108),
.Y(n_1196)
);

INVx2_ASAP7_75t_SL g1197 ( 
.A(n_40),
.Y(n_1197)
);

CKINVDCx5p33_ASAP7_75t_R g1198 ( 
.A(n_816),
.Y(n_1198)
);

CKINVDCx20_ASAP7_75t_R g1199 ( 
.A(n_422),
.Y(n_1199)
);

CKINVDCx5p33_ASAP7_75t_R g1200 ( 
.A(n_631),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_9),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_878),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_804),
.Y(n_1203)
);

CKINVDCx5p33_ASAP7_75t_R g1204 ( 
.A(n_525),
.Y(n_1204)
);

CKINVDCx5p33_ASAP7_75t_R g1205 ( 
.A(n_859),
.Y(n_1205)
);

CKINVDCx20_ASAP7_75t_R g1206 ( 
.A(n_52),
.Y(n_1206)
);

CKINVDCx20_ASAP7_75t_R g1207 ( 
.A(n_89),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_271),
.Y(n_1208)
);

CKINVDCx5p33_ASAP7_75t_R g1209 ( 
.A(n_627),
.Y(n_1209)
);

INVx2_ASAP7_75t_SL g1210 ( 
.A(n_837),
.Y(n_1210)
);

CKINVDCx14_ASAP7_75t_R g1211 ( 
.A(n_347),
.Y(n_1211)
);

BUFx3_ASAP7_75t_L g1212 ( 
.A(n_562),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_801),
.Y(n_1213)
);

INVx1_ASAP7_75t_SL g1214 ( 
.A(n_848),
.Y(n_1214)
);

CKINVDCx5p33_ASAP7_75t_R g1215 ( 
.A(n_720),
.Y(n_1215)
);

CKINVDCx5p33_ASAP7_75t_R g1216 ( 
.A(n_546),
.Y(n_1216)
);

CKINVDCx5p33_ASAP7_75t_R g1217 ( 
.A(n_847),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_821),
.Y(n_1218)
);

CKINVDCx20_ASAP7_75t_R g1219 ( 
.A(n_788),
.Y(n_1219)
);

CKINVDCx5p33_ASAP7_75t_R g1220 ( 
.A(n_401),
.Y(n_1220)
);

CKINVDCx5p33_ASAP7_75t_R g1221 ( 
.A(n_688),
.Y(n_1221)
);

CKINVDCx20_ASAP7_75t_R g1222 ( 
.A(n_889),
.Y(n_1222)
);

CKINVDCx5p33_ASAP7_75t_R g1223 ( 
.A(n_888),
.Y(n_1223)
);

CKINVDCx5p33_ASAP7_75t_R g1224 ( 
.A(n_234),
.Y(n_1224)
);

CKINVDCx5p33_ASAP7_75t_R g1225 ( 
.A(n_449),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_347),
.Y(n_1226)
);

CKINVDCx5p33_ASAP7_75t_R g1227 ( 
.A(n_441),
.Y(n_1227)
);

INVx1_ASAP7_75t_SL g1228 ( 
.A(n_832),
.Y(n_1228)
);

CKINVDCx5p33_ASAP7_75t_R g1229 ( 
.A(n_45),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_504),
.Y(n_1230)
);

CKINVDCx5p33_ASAP7_75t_R g1231 ( 
.A(n_635),
.Y(n_1231)
);

CKINVDCx5p33_ASAP7_75t_R g1232 ( 
.A(n_44),
.Y(n_1232)
);

CKINVDCx5p33_ASAP7_75t_R g1233 ( 
.A(n_31),
.Y(n_1233)
);

CKINVDCx5p33_ASAP7_75t_R g1234 ( 
.A(n_773),
.Y(n_1234)
);

CKINVDCx5p33_ASAP7_75t_R g1235 ( 
.A(n_271),
.Y(n_1235)
);

CKINVDCx5p33_ASAP7_75t_R g1236 ( 
.A(n_214),
.Y(n_1236)
);

BUFx10_ASAP7_75t_L g1237 ( 
.A(n_877),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_339),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_914),
.Y(n_1239)
);

INVxp67_ASAP7_75t_L g1240 ( 
.A(n_63),
.Y(n_1240)
);

INVx2_ASAP7_75t_SL g1241 ( 
.A(n_289),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_55),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1),
.Y(n_1243)
);

INVx2_ASAP7_75t_SL g1244 ( 
.A(n_177),
.Y(n_1244)
);

INVx1_ASAP7_75t_SL g1245 ( 
.A(n_782),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_408),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_768),
.Y(n_1247)
);

CKINVDCx5p33_ASAP7_75t_R g1248 ( 
.A(n_807),
.Y(n_1248)
);

BUFx3_ASAP7_75t_L g1249 ( 
.A(n_46),
.Y(n_1249)
);

BUFx10_ASAP7_75t_L g1250 ( 
.A(n_304),
.Y(n_1250)
);

HB1xp67_ASAP7_75t_L g1251 ( 
.A(n_514),
.Y(n_1251)
);

CKINVDCx5p33_ASAP7_75t_R g1252 ( 
.A(n_780),
.Y(n_1252)
);

CKINVDCx5p33_ASAP7_75t_R g1253 ( 
.A(n_67),
.Y(n_1253)
);

CKINVDCx5p33_ASAP7_75t_R g1254 ( 
.A(n_903),
.Y(n_1254)
);

CKINVDCx5p33_ASAP7_75t_R g1255 ( 
.A(n_79),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_839),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_784),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_13),
.Y(n_1258)
);

CKINVDCx5p33_ASAP7_75t_R g1259 ( 
.A(n_407),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_578),
.Y(n_1260)
);

CKINVDCx5p33_ASAP7_75t_R g1261 ( 
.A(n_899),
.Y(n_1261)
);

BUFx2_ASAP7_75t_L g1262 ( 
.A(n_24),
.Y(n_1262)
);

CKINVDCx5p33_ASAP7_75t_R g1263 ( 
.A(n_811),
.Y(n_1263)
);

CKINVDCx20_ASAP7_75t_R g1264 ( 
.A(n_488),
.Y(n_1264)
);

CKINVDCx5p33_ASAP7_75t_R g1265 ( 
.A(n_781),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_293),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_799),
.Y(n_1267)
);

CKINVDCx5p33_ASAP7_75t_R g1268 ( 
.A(n_880),
.Y(n_1268)
);

CKINVDCx5p33_ASAP7_75t_R g1269 ( 
.A(n_325),
.Y(n_1269)
);

CKINVDCx5p33_ASAP7_75t_R g1270 ( 
.A(n_182),
.Y(n_1270)
);

HB1xp67_ASAP7_75t_L g1271 ( 
.A(n_740),
.Y(n_1271)
);

HB1xp67_ASAP7_75t_L g1272 ( 
.A(n_786),
.Y(n_1272)
);

BUFx2_ASAP7_75t_L g1273 ( 
.A(n_852),
.Y(n_1273)
);

CKINVDCx5p33_ASAP7_75t_R g1274 ( 
.A(n_220),
.Y(n_1274)
);

CKINVDCx5p33_ASAP7_75t_R g1275 ( 
.A(n_884),
.Y(n_1275)
);

CKINVDCx20_ASAP7_75t_R g1276 ( 
.A(n_858),
.Y(n_1276)
);

BUFx6f_ASAP7_75t_L g1277 ( 
.A(n_34),
.Y(n_1277)
);

CKINVDCx5p33_ASAP7_75t_R g1278 ( 
.A(n_186),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_360),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_148),
.Y(n_1280)
);

CKINVDCx5p33_ASAP7_75t_R g1281 ( 
.A(n_619),
.Y(n_1281)
);

CKINVDCx20_ASAP7_75t_R g1282 ( 
.A(n_304),
.Y(n_1282)
);

CKINVDCx5p33_ASAP7_75t_R g1283 ( 
.A(n_778),
.Y(n_1283)
);

CKINVDCx20_ASAP7_75t_R g1284 ( 
.A(n_925),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1196),
.Y(n_1285)
);

CKINVDCx20_ASAP7_75t_R g1286 ( 
.A(n_949),
.Y(n_1286)
);

BUFx10_ASAP7_75t_L g1287 ( 
.A(n_1175),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1196),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1196),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1196),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1196),
.Y(n_1291)
);

CKINVDCx5p33_ASAP7_75t_R g1292 ( 
.A(n_1018),
.Y(n_1292)
);

CKINVDCx5p33_ASAP7_75t_R g1293 ( 
.A(n_1078),
.Y(n_1293)
);

CKINVDCx5p33_ASAP7_75t_R g1294 ( 
.A(n_916),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_939),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_939),
.Y(n_1296)
);

CKINVDCx5p33_ASAP7_75t_R g1297 ( 
.A(n_919),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_939),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1077),
.Y(n_1299)
);

CKINVDCx5p33_ASAP7_75t_R g1300 ( 
.A(n_924),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1077),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1077),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1179),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1179),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1179),
.Y(n_1305)
);

INVxp67_ASAP7_75t_L g1306 ( 
.A(n_1262),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1277),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1277),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1277),
.Y(n_1309)
);

INVx2_ASAP7_75t_L g1310 ( 
.A(n_982),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_918),
.Y(n_1311)
);

INVxp67_ASAP7_75t_L g1312 ( 
.A(n_1251),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1002),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1015),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1051),
.Y(n_1315)
);

HB1xp67_ASAP7_75t_L g1316 ( 
.A(n_943),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1065),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1132),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1212),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1249),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_931),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_937),
.Y(n_1322)
);

INVx1_ASAP7_75t_SL g1323 ( 
.A(n_971),
.Y(n_1323)
);

CKINVDCx14_ASAP7_75t_R g1324 ( 
.A(n_1211),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_947),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_955),
.Y(n_1326)
);

INVxp67_ASAP7_75t_SL g1327 ( 
.A(n_1271),
.Y(n_1327)
);

CKINVDCx16_ASAP7_75t_R g1328 ( 
.A(n_1153),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_959),
.Y(n_1329)
);

INVx2_ASAP7_75t_L g1330 ( 
.A(n_982),
.Y(n_1330)
);

CKINVDCx20_ASAP7_75t_R g1331 ( 
.A(n_967),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_965),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_986),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_990),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_992),
.Y(n_1335)
);

INVxp33_ASAP7_75t_SL g1336 ( 
.A(n_915),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1000),
.Y(n_1337)
);

CKINVDCx5p33_ASAP7_75t_R g1338 ( 
.A(n_927),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1043),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1050),
.Y(n_1340)
);

CKINVDCx20_ASAP7_75t_R g1341 ( 
.A(n_969),
.Y(n_1341)
);

INVx1_ASAP7_75t_SL g1342 ( 
.A(n_974),
.Y(n_1342)
);

CKINVDCx5p33_ASAP7_75t_R g1343 ( 
.A(n_932),
.Y(n_1343)
);

CKINVDCx20_ASAP7_75t_R g1344 ( 
.A(n_1148),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1052),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1088),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1089),
.Y(n_1347)
);

CKINVDCx20_ASAP7_75t_R g1348 ( 
.A(n_1219),
.Y(n_1348)
);

BUFx2_ASAP7_75t_L g1349 ( 
.A(n_920),
.Y(n_1349)
);

INVx2_ASAP7_75t_L g1350 ( 
.A(n_982),
.Y(n_1350)
);

CKINVDCx16_ASAP7_75t_R g1351 ( 
.A(n_1098),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1091),
.Y(n_1352)
);

AND2x4_ASAP7_75t_L g1353 ( 
.A(n_1349),
.B(n_1273),
.Y(n_1353)
);

INVx3_ASAP7_75t_L g1354 ( 
.A(n_1295),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1296),
.Y(n_1355)
);

INVx2_ASAP7_75t_L g1356 ( 
.A(n_1298),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_L g1357 ( 
.A(n_1294),
.B(n_1297),
.Y(n_1357)
);

AND2x4_ASAP7_75t_L g1358 ( 
.A(n_1327),
.B(n_1013),
.Y(n_1358)
);

BUFx6f_ASAP7_75t_L g1359 ( 
.A(n_1299),
.Y(n_1359)
);

INVx2_ASAP7_75t_L g1360 ( 
.A(n_1301),
.Y(n_1360)
);

AND2x2_ASAP7_75t_L g1361 ( 
.A(n_1324),
.B(n_1058),
.Y(n_1361)
);

BUFx6f_ASAP7_75t_L g1362 ( 
.A(n_1302),
.Y(n_1362)
);

INVx2_ASAP7_75t_L g1363 ( 
.A(n_1303),
.Y(n_1363)
);

INVx2_ASAP7_75t_L g1364 ( 
.A(n_1304),
.Y(n_1364)
);

INVx2_ASAP7_75t_L g1365 ( 
.A(n_1305),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_SL g1366 ( 
.A(n_1351),
.B(n_1001),
.Y(n_1366)
);

BUFx6f_ASAP7_75t_L g1367 ( 
.A(n_1307),
.Y(n_1367)
);

INVx2_ASAP7_75t_L g1368 ( 
.A(n_1308),
.Y(n_1368)
);

CKINVDCx20_ASAP7_75t_R g1369 ( 
.A(n_1284),
.Y(n_1369)
);

BUFx6f_ASAP7_75t_L g1370 ( 
.A(n_1309),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1285),
.Y(n_1371)
);

INVx2_ASAP7_75t_L g1372 ( 
.A(n_1288),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1289),
.Y(n_1373)
);

AND2x4_ASAP7_75t_L g1374 ( 
.A(n_1306),
.B(n_1272),
.Y(n_1374)
);

INVx4_ASAP7_75t_L g1375 ( 
.A(n_1300),
.Y(n_1375)
);

BUFx6f_ASAP7_75t_L g1376 ( 
.A(n_1321),
.Y(n_1376)
);

AND2x4_ASAP7_75t_L g1377 ( 
.A(n_1312),
.B(n_979),
.Y(n_1377)
);

AND2x2_ASAP7_75t_SL g1378 ( 
.A(n_1328),
.B(n_1158),
.Y(n_1378)
);

AND2x4_ASAP7_75t_L g1379 ( 
.A(n_1316),
.B(n_1152),
.Y(n_1379)
);

AND2x6_ASAP7_75t_L g1380 ( 
.A(n_1311),
.B(n_1053),
.Y(n_1380)
);

INVx2_ASAP7_75t_L g1381 ( 
.A(n_1290),
.Y(n_1381)
);

INVx3_ASAP7_75t_L g1382 ( 
.A(n_1313),
.Y(n_1382)
);

INVx2_ASAP7_75t_L g1383 ( 
.A(n_1291),
.Y(n_1383)
);

HB1xp67_ASAP7_75t_L g1384 ( 
.A(n_1323),
.Y(n_1384)
);

BUFx6f_ASAP7_75t_L g1385 ( 
.A(n_1322),
.Y(n_1385)
);

AND2x4_ASAP7_75t_L g1386 ( 
.A(n_1338),
.B(n_1011),
.Y(n_1386)
);

INVx3_ASAP7_75t_L g1387 ( 
.A(n_1314),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1325),
.Y(n_1388)
);

BUFx6f_ASAP7_75t_L g1389 ( 
.A(n_1326),
.Y(n_1389)
);

CKINVDCx20_ASAP7_75t_R g1390 ( 
.A(n_1286),
.Y(n_1390)
);

INVx2_ASAP7_75t_L g1391 ( 
.A(n_1329),
.Y(n_1391)
);

BUFx6f_ASAP7_75t_L g1392 ( 
.A(n_1332),
.Y(n_1392)
);

INVx2_ASAP7_75t_L g1393 ( 
.A(n_1333),
.Y(n_1393)
);

AND2x4_ASAP7_75t_L g1394 ( 
.A(n_1343),
.B(n_1168),
.Y(n_1394)
);

INVxp67_ASAP7_75t_L g1395 ( 
.A(n_1342),
.Y(n_1395)
);

NAND2xp5_ASAP7_75t_L g1396 ( 
.A(n_1315),
.B(n_944),
.Y(n_1396)
);

NOR2xp33_ASAP7_75t_L g1397 ( 
.A(n_1336),
.B(n_975),
.Y(n_1397)
);

AOI22xp5_ASAP7_75t_L g1398 ( 
.A1(n_1292),
.A2(n_1222),
.B1(n_1276),
.B2(n_1020),
.Y(n_1398)
);

INVx2_ASAP7_75t_L g1399 ( 
.A(n_1334),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_SL g1400 ( 
.A(n_1293),
.B(n_1001),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1335),
.Y(n_1401)
);

INVx2_ASAP7_75t_L g1402 ( 
.A(n_1359),
.Y(n_1402)
);

CKINVDCx5p33_ASAP7_75t_R g1403 ( 
.A(n_1369),
.Y(n_1403)
);

NOR2xp33_ASAP7_75t_R g1404 ( 
.A(n_1390),
.B(n_1331),
.Y(n_1404)
);

BUFx2_ASAP7_75t_L g1405 ( 
.A(n_1395),
.Y(n_1405)
);

CKINVDCx5p33_ASAP7_75t_R g1406 ( 
.A(n_1375),
.Y(n_1406)
);

CKINVDCx5p33_ASAP7_75t_R g1407 ( 
.A(n_1384),
.Y(n_1407)
);

INVx2_ASAP7_75t_L g1408 ( 
.A(n_1359),
.Y(n_1408)
);

CKINVDCx5p33_ASAP7_75t_R g1409 ( 
.A(n_1357),
.Y(n_1409)
);

BUFx6f_ASAP7_75t_L g1410 ( 
.A(n_1376),
.Y(n_1410)
);

CKINVDCx5p33_ASAP7_75t_R g1411 ( 
.A(n_1397),
.Y(n_1411)
);

CKINVDCx5p33_ASAP7_75t_R g1412 ( 
.A(n_1398),
.Y(n_1412)
);

CKINVDCx5p33_ASAP7_75t_R g1413 ( 
.A(n_1386),
.Y(n_1413)
);

CKINVDCx5p33_ASAP7_75t_R g1414 ( 
.A(n_1394),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_L g1415 ( 
.A(n_1371),
.B(n_1373),
.Y(n_1415)
);

CKINVDCx20_ASAP7_75t_R g1416 ( 
.A(n_1400),
.Y(n_1416)
);

CKINVDCx20_ASAP7_75t_R g1417 ( 
.A(n_1366),
.Y(n_1417)
);

BUFx3_ASAP7_75t_L g1418 ( 
.A(n_1389),
.Y(n_1418)
);

NAND2xp33_ASAP7_75t_R g1419 ( 
.A(n_1353),
.B(n_921),
.Y(n_1419)
);

CKINVDCx20_ASAP7_75t_R g1420 ( 
.A(n_1361),
.Y(n_1420)
);

NOR2xp33_ASAP7_75t_R g1421 ( 
.A(n_1378),
.B(n_1341),
.Y(n_1421)
);

CKINVDCx5p33_ASAP7_75t_R g1422 ( 
.A(n_1377),
.Y(n_1422)
);

INVx8_ASAP7_75t_L g1423 ( 
.A(n_1379),
.Y(n_1423)
);

CKINVDCx16_ASAP7_75t_R g1424 ( 
.A(n_1358),
.Y(n_1424)
);

INVx2_ASAP7_75t_L g1425 ( 
.A(n_1362),
.Y(n_1425)
);

OA21x2_ASAP7_75t_L g1426 ( 
.A1(n_1372),
.A2(n_1330),
.B(n_1310),
.Y(n_1426)
);

INVx2_ASAP7_75t_L g1427 ( 
.A(n_1362),
.Y(n_1427)
);

NOR2xp33_ASAP7_75t_R g1428 ( 
.A(n_1382),
.B(n_1344),
.Y(n_1428)
);

CKINVDCx5p33_ASAP7_75t_R g1429 ( 
.A(n_1380),
.Y(n_1429)
);

AOI21x1_ASAP7_75t_L g1430 ( 
.A1(n_1381),
.A2(n_1350),
.B(n_922),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1388),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1401),
.Y(n_1432)
);

INVx2_ASAP7_75t_L g1433 ( 
.A(n_1367),
.Y(n_1433)
);

BUFx10_ASAP7_75t_L g1434 ( 
.A(n_1374),
.Y(n_1434)
);

CKINVDCx5p33_ASAP7_75t_R g1435 ( 
.A(n_1380),
.Y(n_1435)
);

NOR2xp67_ASAP7_75t_L g1436 ( 
.A(n_1387),
.B(n_1320),
.Y(n_1436)
);

CKINVDCx5p33_ASAP7_75t_R g1437 ( 
.A(n_1392),
.Y(n_1437)
);

CKINVDCx5p33_ASAP7_75t_R g1438 ( 
.A(n_1376),
.Y(n_1438)
);

OAI22xp33_ASAP7_75t_SL g1439 ( 
.A1(n_1396),
.A2(n_1005),
.B1(n_1197),
.B2(n_1111),
.Y(n_1439)
);

CKINVDCx5p33_ASAP7_75t_R g1440 ( 
.A(n_1385),
.Y(n_1440)
);

CKINVDCx5p33_ASAP7_75t_R g1441 ( 
.A(n_1385),
.Y(n_1441)
);

CKINVDCx5p33_ASAP7_75t_R g1442 ( 
.A(n_1367),
.Y(n_1442)
);

NOR2xp33_ASAP7_75t_L g1443 ( 
.A(n_1383),
.B(n_1287),
.Y(n_1443)
);

BUFx6f_ASAP7_75t_L g1444 ( 
.A(n_1370),
.Y(n_1444)
);

CKINVDCx5p33_ASAP7_75t_R g1445 ( 
.A(n_1370),
.Y(n_1445)
);

BUFx3_ASAP7_75t_L g1446 ( 
.A(n_1391),
.Y(n_1446)
);

NOR2xp67_ASAP7_75t_L g1447 ( 
.A(n_1354),
.B(n_1317),
.Y(n_1447)
);

INVx2_ASAP7_75t_L g1448 ( 
.A(n_1356),
.Y(n_1448)
);

CKINVDCx5p33_ASAP7_75t_R g1449 ( 
.A(n_1393),
.Y(n_1449)
);

AND2x2_ASAP7_75t_L g1450 ( 
.A(n_1399),
.B(n_1287),
.Y(n_1450)
);

BUFx6f_ASAP7_75t_L g1451 ( 
.A(n_1360),
.Y(n_1451)
);

INVxp67_ASAP7_75t_L g1452 ( 
.A(n_1355),
.Y(n_1452)
);

HB1xp67_ASAP7_75t_L g1453 ( 
.A(n_1363),
.Y(n_1453)
);

INVx4_ASAP7_75t_L g1454 ( 
.A(n_1364),
.Y(n_1454)
);

INVx2_ASAP7_75t_L g1455 ( 
.A(n_1365),
.Y(n_1455)
);

INVx2_ASAP7_75t_L g1456 ( 
.A(n_1368),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1388),
.Y(n_1457)
);

INVx2_ASAP7_75t_L g1458 ( 
.A(n_1359),
.Y(n_1458)
);

AND2x2_ASAP7_75t_L g1459 ( 
.A(n_1395),
.B(n_1318),
.Y(n_1459)
);

CKINVDCx5p33_ASAP7_75t_R g1460 ( 
.A(n_1369),
.Y(n_1460)
);

INVx2_ASAP7_75t_SL g1461 ( 
.A(n_1384),
.Y(n_1461)
);

CKINVDCx5p33_ASAP7_75t_R g1462 ( 
.A(n_1369),
.Y(n_1462)
);

OR2x2_ASAP7_75t_L g1463 ( 
.A(n_1395),
.B(n_1319),
.Y(n_1463)
);

CKINVDCx5p33_ASAP7_75t_R g1464 ( 
.A(n_1369),
.Y(n_1464)
);

CKINVDCx20_ASAP7_75t_R g1465 ( 
.A(n_1369),
.Y(n_1465)
);

AND2x2_ASAP7_75t_L g1466 ( 
.A(n_1395),
.B(n_1352),
.Y(n_1466)
);

CKINVDCx20_ASAP7_75t_R g1467 ( 
.A(n_1369),
.Y(n_1467)
);

NOR2xp33_ASAP7_75t_R g1468 ( 
.A(n_1369),
.B(n_1348),
.Y(n_1468)
);

CKINVDCx5p33_ASAP7_75t_R g1469 ( 
.A(n_1369),
.Y(n_1469)
);

NOR2xp67_ASAP7_75t_L g1470 ( 
.A(n_1395),
.B(n_933),
.Y(n_1470)
);

CKINVDCx5p33_ASAP7_75t_R g1471 ( 
.A(n_1369),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1388),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1388),
.Y(n_1473)
);

INVx2_ASAP7_75t_L g1474 ( 
.A(n_1448),
.Y(n_1474)
);

INVx3_ASAP7_75t_L g1475 ( 
.A(n_1410),
.Y(n_1475)
);

AND2x2_ASAP7_75t_L g1476 ( 
.A(n_1466),
.B(n_1337),
.Y(n_1476)
);

BUFx6f_ASAP7_75t_L g1477 ( 
.A(n_1410),
.Y(n_1477)
);

NAND2xp5_ASAP7_75t_L g1478 ( 
.A(n_1409),
.B(n_945),
.Y(n_1478)
);

NOR2xp33_ASAP7_75t_L g1479 ( 
.A(n_1411),
.B(n_1037),
.Y(n_1479)
);

NAND3xp33_ASAP7_75t_L g1480 ( 
.A(n_1459),
.B(n_928),
.C(n_923),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_L g1481 ( 
.A(n_1415),
.B(n_958),
.Y(n_1481)
);

AOI22xp5_ASAP7_75t_L g1482 ( 
.A1(n_1473),
.A2(n_1431),
.B1(n_1457),
.B2(n_1432),
.Y(n_1482)
);

OR2x6_ASAP7_75t_L g1483 ( 
.A(n_1461),
.B(n_1074),
.Y(n_1483)
);

NOR2xp33_ASAP7_75t_L g1484 ( 
.A(n_1405),
.B(n_1214),
.Y(n_1484)
);

INVx3_ASAP7_75t_L g1485 ( 
.A(n_1418),
.Y(n_1485)
);

OR2x2_ASAP7_75t_L g1486 ( 
.A(n_1463),
.B(n_1142),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1453),
.Y(n_1487)
);

NOR2xp33_ASAP7_75t_L g1488 ( 
.A(n_1449),
.B(n_1228),
.Y(n_1488)
);

AND2x4_ASAP7_75t_L g1489 ( 
.A(n_1402),
.B(n_1339),
.Y(n_1489)
);

INVx2_ASAP7_75t_L g1490 ( 
.A(n_1455),
.Y(n_1490)
);

INVx2_ASAP7_75t_SL g1491 ( 
.A(n_1407),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_L g1492 ( 
.A(n_1472),
.B(n_988),
.Y(n_1492)
);

NOR2xp33_ASAP7_75t_L g1493 ( 
.A(n_1406),
.B(n_1245),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1446),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1456),
.Y(n_1495)
);

AO22x1_ASAP7_75t_L g1496 ( 
.A1(n_1412),
.A2(n_1154),
.B1(n_1186),
.B2(n_1171),
.Y(n_1496)
);

BUFx6f_ASAP7_75t_L g1497 ( 
.A(n_1444),
.Y(n_1497)
);

INVx1_ASAP7_75t_SL g1498 ( 
.A(n_1428),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1452),
.Y(n_1499)
);

INVx2_ASAP7_75t_L g1500 ( 
.A(n_1426),
.Y(n_1500)
);

INVx2_ASAP7_75t_L g1501 ( 
.A(n_1426),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_L g1502 ( 
.A(n_1470),
.B(n_1060),
.Y(n_1502)
);

BUFx4_ASAP7_75t_L g1503 ( 
.A(n_1404),
.Y(n_1503)
);

BUFx6f_ASAP7_75t_L g1504 ( 
.A(n_1444),
.Y(n_1504)
);

BUFx2_ASAP7_75t_L g1505 ( 
.A(n_1468),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1408),
.Y(n_1506)
);

INVx2_ASAP7_75t_L g1507 ( 
.A(n_1451),
.Y(n_1507)
);

AOI22xp33_ASAP7_75t_L g1508 ( 
.A1(n_1439),
.A2(n_1007),
.B1(n_1055),
.B2(n_938),
.Y(n_1508)
);

BUFx3_ASAP7_75t_L g1509 ( 
.A(n_1437),
.Y(n_1509)
);

AND2x2_ASAP7_75t_L g1510 ( 
.A(n_1450),
.B(n_1438),
.Y(n_1510)
);

AND2x2_ASAP7_75t_SL g1511 ( 
.A(n_1424),
.B(n_1443),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1425),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1427),
.Y(n_1513)
);

HB1xp67_ASAP7_75t_L g1514 ( 
.A(n_1440),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1433),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1458),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1447),
.Y(n_1517)
);

INVx2_ASAP7_75t_L g1518 ( 
.A(n_1451),
.Y(n_1518)
);

AND2x2_ASAP7_75t_L g1519 ( 
.A(n_1441),
.B(n_1442),
.Y(n_1519)
);

CKINVDCx5p33_ASAP7_75t_R g1520 ( 
.A(n_1403),
.Y(n_1520)
);

INVxp67_ASAP7_75t_SL g1521 ( 
.A(n_1436),
.Y(n_1521)
);

BUFx3_ASAP7_75t_L g1522 ( 
.A(n_1465),
.Y(n_1522)
);

INVx4_ASAP7_75t_L g1523 ( 
.A(n_1445),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_SL g1524 ( 
.A(n_1429),
.B(n_1283),
.Y(n_1524)
);

BUFx2_ASAP7_75t_L g1525 ( 
.A(n_1421),
.Y(n_1525)
);

BUFx3_ASAP7_75t_L g1526 ( 
.A(n_1467),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1430),
.Y(n_1527)
);

BUFx6f_ASAP7_75t_L g1528 ( 
.A(n_1423),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1454),
.Y(n_1529)
);

INVx4_ASAP7_75t_L g1530 ( 
.A(n_1423),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_SL g1531 ( 
.A(n_1435),
.B(n_934),
.Y(n_1531)
);

AOI22xp5_ASAP7_75t_L g1532 ( 
.A1(n_1419),
.A2(n_948),
.B1(n_950),
.B2(n_940),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1422),
.Y(n_1533)
);

AOI22xp33_ASAP7_75t_L g1534 ( 
.A1(n_1420),
.A2(n_1084),
.B1(n_1145),
.B2(n_1075),
.Y(n_1534)
);

INVx3_ASAP7_75t_L g1535 ( 
.A(n_1434),
.Y(n_1535)
);

NAND3xp33_ASAP7_75t_L g1536 ( 
.A(n_1413),
.B(n_936),
.C(n_930),
.Y(n_1536)
);

NOR2xp33_ASAP7_75t_L g1537 ( 
.A(n_1414),
.B(n_1416),
.Y(n_1537)
);

INVx3_ASAP7_75t_L g1538 ( 
.A(n_1460),
.Y(n_1538)
);

CKINVDCx5p33_ASAP7_75t_R g1539 ( 
.A(n_1462),
.Y(n_1539)
);

NOR2xp33_ASAP7_75t_SL g1540 ( 
.A(n_1417),
.B(n_1028),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1464),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1469),
.Y(n_1542)
);

NOR2xp33_ASAP7_75t_L g1543 ( 
.A(n_1471),
.B(n_942),
.Y(n_1543)
);

AND2x4_ASAP7_75t_L g1544 ( 
.A(n_1418),
.B(n_1340),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_L g1545 ( 
.A(n_1409),
.B(n_1087),
.Y(n_1545)
);

NOR2xp33_ASAP7_75t_L g1546 ( 
.A(n_1411),
.B(n_946),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1466),
.B(n_1345),
.Y(n_1547)
);

NOR2x1p5_ASAP7_75t_L g1548 ( 
.A(n_1429),
.B(n_1274),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_L g1549 ( 
.A(n_1409),
.B(n_1210),
.Y(n_1549)
);

INVx3_ASAP7_75t_L g1550 ( 
.A(n_1410),
.Y(n_1550)
);

OR2x6_ASAP7_75t_L g1551 ( 
.A(n_1461),
.B(n_1241),
.Y(n_1551)
);

INVx1_ASAP7_75t_SL g1552 ( 
.A(n_1405),
.Y(n_1552)
);

INVxp67_ASAP7_75t_SL g1553 ( 
.A(n_1410),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_SL g1554 ( 
.A(n_1409),
.B(n_951),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_SL g1555 ( 
.A(n_1409),
.B(n_952),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1409),
.B(n_917),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1453),
.Y(n_1557)
);

OR2x6_ASAP7_75t_L g1558 ( 
.A(n_1461),
.B(n_1244),
.Y(n_1558)
);

NAND3xp33_ASAP7_75t_L g1559 ( 
.A(n_1411),
.B(n_960),
.C(n_956),
.Y(n_1559)
);

INVxp67_ASAP7_75t_SL g1560 ( 
.A(n_1410),
.Y(n_1560)
);

BUFx2_ASAP7_75t_L g1561 ( 
.A(n_1405),
.Y(n_1561)
);

BUFx3_ASAP7_75t_L g1562 ( 
.A(n_1418),
.Y(n_1562)
);

BUFx2_ASAP7_75t_L g1563 ( 
.A(n_1405),
.Y(n_1563)
);

AND2x6_ASAP7_75t_L g1564 ( 
.A(n_1466),
.B(n_926),
.Y(n_1564)
);

AOI22xp33_ASAP7_75t_L g1565 ( 
.A1(n_1431),
.A2(n_935),
.B1(n_957),
.B2(n_929),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1453),
.Y(n_1566)
);

INVx2_ASAP7_75t_L g1567 ( 
.A(n_1448),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1466),
.B(n_1346),
.Y(n_1568)
);

NOR2xp33_ASAP7_75t_L g1569 ( 
.A(n_1411),
.B(n_962),
.Y(n_1569)
);

CKINVDCx5p33_ASAP7_75t_R g1570 ( 
.A(n_1404),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1453),
.Y(n_1571)
);

NAND2xp5_ASAP7_75t_L g1572 ( 
.A(n_1409),
.B(n_977),
.Y(n_1572)
);

INVx2_ASAP7_75t_L g1573 ( 
.A(n_1448),
.Y(n_1573)
);

INVx2_ASAP7_75t_L g1574 ( 
.A(n_1448),
.Y(n_1574)
);

CKINVDCx16_ASAP7_75t_R g1575 ( 
.A(n_1404),
.Y(n_1575)
);

NOR2xp33_ASAP7_75t_L g1576 ( 
.A(n_1411),
.B(n_964),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1453),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1453),
.Y(n_1578)
);

INVx6_ASAP7_75t_L g1579 ( 
.A(n_1434),
.Y(n_1579)
);

INVx2_ASAP7_75t_L g1580 ( 
.A(n_1448),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_L g1581 ( 
.A(n_1409),
.B(n_978),
.Y(n_1581)
);

NOR2xp33_ASAP7_75t_L g1582 ( 
.A(n_1411),
.B(n_966),
.Y(n_1582)
);

BUFx6f_ASAP7_75t_L g1583 ( 
.A(n_1410),
.Y(n_1583)
);

BUFx10_ASAP7_75t_L g1584 ( 
.A(n_1407),
.Y(n_1584)
);

BUFx4f_ASAP7_75t_L g1585 ( 
.A(n_1405),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1453),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1466),
.B(n_1347),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1453),
.Y(n_1588)
);

INVx2_ASAP7_75t_L g1589 ( 
.A(n_1448),
.Y(n_1589)
);

OR2x2_ASAP7_75t_L g1590 ( 
.A(n_1405),
.B(n_1026),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_SL g1591 ( 
.A(n_1478),
.B(n_1545),
.Y(n_1591)
);

INVx2_ASAP7_75t_L g1592 ( 
.A(n_1500),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1489),
.Y(n_1593)
);

AOI22xp33_ASAP7_75t_L g1594 ( 
.A1(n_1479),
.A2(n_980),
.B1(n_983),
.B2(n_981),
.Y(n_1594)
);

AND2x4_ASAP7_75t_SL g1595 ( 
.A(n_1584),
.B(n_1237),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_L g1596 ( 
.A(n_1488),
.B(n_989),
.Y(n_1596)
);

AND2x4_ASAP7_75t_SL g1597 ( 
.A(n_1528),
.B(n_1237),
.Y(n_1597)
);

NOR2xp33_ASAP7_75t_L g1598 ( 
.A(n_1546),
.B(n_1040),
.Y(n_1598)
);

INVx6_ASAP7_75t_L g1599 ( 
.A(n_1579),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1495),
.Y(n_1600)
);

INVx2_ASAP7_75t_L g1601 ( 
.A(n_1501),
.Y(n_1601)
);

AOI22xp5_ASAP7_75t_L g1602 ( 
.A1(n_1493),
.A2(n_1032),
.B1(n_1034),
.B2(n_991),
.Y(n_1602)
);

INVx2_ASAP7_75t_SL g1603 ( 
.A(n_1585),
.Y(n_1603)
);

AOI21xp5_ASAP7_75t_L g1604 ( 
.A1(n_1521),
.A2(n_1081),
.B(n_1061),
.Y(n_1604)
);

AND2x2_ASAP7_75t_L g1605 ( 
.A(n_1510),
.B(n_1476),
.Y(n_1605)
);

OAI221xp5_ASAP7_75t_L g1606 ( 
.A1(n_1534),
.A2(n_1240),
.B1(n_1128),
.B2(n_1131),
.C(n_1126),
.Y(n_1606)
);

NAND3xp33_ASAP7_75t_L g1607 ( 
.A(n_1569),
.B(n_972),
.C(n_968),
.Y(n_1607)
);

AND2x4_ASAP7_75t_L g1608 ( 
.A(n_1528),
.B(n_1122),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_SL g1609 ( 
.A(n_1549),
.B(n_953),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_L g1610 ( 
.A(n_1547),
.B(n_1082),
.Y(n_1610)
);

NAND2xp33_ASAP7_75t_L g1611 ( 
.A(n_1564),
.B(n_982),
.Y(n_1611)
);

A2O1A1Ixp33_ASAP7_75t_L g1612 ( 
.A1(n_1484),
.A2(n_1086),
.B(n_1103),
.C(n_1083),
.Y(n_1612)
);

A2O1A1Ixp33_ASAP7_75t_L g1613 ( 
.A1(n_1556),
.A2(n_1107),
.B(n_1112),
.C(n_1106),
.Y(n_1613)
);

INVx2_ASAP7_75t_L g1614 ( 
.A(n_1474),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1490),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_L g1616 ( 
.A(n_1568),
.B(n_1115),
.Y(n_1616)
);

AND2x4_ASAP7_75t_L g1617 ( 
.A(n_1530),
.B(n_1140),
.Y(n_1617)
);

OR2x2_ASAP7_75t_L g1618 ( 
.A(n_1552),
.B(n_1269),
.Y(n_1618)
);

INVx2_ASAP7_75t_L g1619 ( 
.A(n_1567),
.Y(n_1619)
);

INVx3_ASAP7_75t_L g1620 ( 
.A(n_1477),
.Y(n_1620)
);

INVx2_ASAP7_75t_L g1621 ( 
.A(n_1573),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1574),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1580),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1589),
.Y(n_1624)
);

INVxp67_ASAP7_75t_SL g1625 ( 
.A(n_1477),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_L g1626 ( 
.A(n_1587),
.B(n_1120),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_SL g1627 ( 
.A(n_1572),
.B(n_954),
.Y(n_1627)
);

OAI22xp5_ASAP7_75t_SL g1628 ( 
.A1(n_1511),
.A2(n_1057),
.B1(n_1121),
.B2(n_1105),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_L g1629 ( 
.A(n_1581),
.B(n_1125),
.Y(n_1629)
);

BUFx6f_ASAP7_75t_L g1630 ( 
.A(n_1497),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1482),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_L g1632 ( 
.A(n_1576),
.B(n_1127),
.Y(n_1632)
);

INVx3_ASAP7_75t_L g1633 ( 
.A(n_1497),
.Y(n_1633)
);

INVx2_ASAP7_75t_L g1634 ( 
.A(n_1494),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_L g1635 ( 
.A(n_1582),
.B(n_1481),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_L g1636 ( 
.A(n_1499),
.B(n_1130),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_SL g1637 ( 
.A(n_1561),
.B(n_961),
.Y(n_1637)
);

BUFx2_ASAP7_75t_L g1638 ( 
.A(n_1563),
.Y(n_1638)
);

INVxp67_ASAP7_75t_L g1639 ( 
.A(n_1486),
.Y(n_1639)
);

INVx2_ASAP7_75t_L g1640 ( 
.A(n_1506),
.Y(n_1640)
);

INVx5_ASAP7_75t_L g1641 ( 
.A(n_1504),
.Y(n_1641)
);

NAND2xp5_ASAP7_75t_SL g1642 ( 
.A(n_1519),
.B(n_963),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_L g1643 ( 
.A(n_1564),
.B(n_1136),
.Y(n_1643)
);

OR2x2_ASAP7_75t_L g1644 ( 
.A(n_1590),
.B(n_1270),
.Y(n_1644)
);

AND2x6_ASAP7_75t_L g1645 ( 
.A(n_1509),
.B(n_1170),
.Y(n_1645)
);

NOR2xp33_ASAP7_75t_SL g1646 ( 
.A(n_1520),
.B(n_1163),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_SL g1647 ( 
.A(n_1491),
.B(n_1498),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1512),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_SL g1649 ( 
.A(n_1523),
.B(n_970),
.Y(n_1649)
);

OR2x6_ASAP7_75t_L g1650 ( 
.A(n_1522),
.B(n_1526),
.Y(n_1650)
);

AOI22xp33_ASAP7_75t_L g1651 ( 
.A1(n_1564),
.A2(n_1190),
.B1(n_1192),
.B2(n_1183),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_L g1652 ( 
.A(n_1517),
.B(n_1202),
.Y(n_1652)
);

INVx3_ASAP7_75t_L g1653 ( 
.A(n_1504),
.Y(n_1653)
);

INVx2_ASAP7_75t_L g1654 ( 
.A(n_1513),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1515),
.Y(n_1655)
);

INVxp67_ASAP7_75t_L g1656 ( 
.A(n_1514),
.Y(n_1656)
);

AND2x2_ASAP7_75t_L g1657 ( 
.A(n_1487),
.B(n_1118),
.Y(n_1657)
);

BUFx6f_ASAP7_75t_SL g1658 ( 
.A(n_1483),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_L g1659 ( 
.A(n_1502),
.B(n_1203),
.Y(n_1659)
);

HB1xp67_ASAP7_75t_L g1660 ( 
.A(n_1583),
.Y(n_1660)
);

INVx2_ASAP7_75t_L g1661 ( 
.A(n_1516),
.Y(n_1661)
);

OR2x6_ASAP7_75t_L g1662 ( 
.A(n_1538),
.B(n_1141),
.Y(n_1662)
);

NOR3xp33_ASAP7_75t_L g1663 ( 
.A(n_1543),
.B(n_993),
.C(n_987),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_L g1664 ( 
.A(n_1492),
.B(n_1213),
.Y(n_1664)
);

INVx2_ASAP7_75t_L g1665 ( 
.A(n_1527),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_SL g1666 ( 
.A(n_1559),
.B(n_973),
.Y(n_1666)
);

NOR2xp33_ASAP7_75t_L g1667 ( 
.A(n_1554),
.B(n_1199),
.Y(n_1667)
);

NOR2xp33_ASAP7_75t_L g1668 ( 
.A(n_1555),
.B(n_1540),
.Y(n_1668)
);

INVx2_ASAP7_75t_L g1669 ( 
.A(n_1507),
.Y(n_1669)
);

NAND2xp33_ASAP7_75t_L g1670 ( 
.A(n_1583),
.B(n_1099),
.Y(n_1670)
);

NAND2xp5_ASAP7_75t_SL g1671 ( 
.A(n_1575),
.B(n_976),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1529),
.B(n_1218),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_L g1673 ( 
.A(n_1532),
.B(n_1239),
.Y(n_1673)
);

INVx2_ASAP7_75t_L g1674 ( 
.A(n_1518),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_L g1675 ( 
.A(n_1557),
.B(n_1247),
.Y(n_1675)
);

NOR2xp33_ASAP7_75t_L g1676 ( 
.A(n_1570),
.B(n_1505),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1566),
.Y(n_1677)
);

INVx4_ASAP7_75t_L g1678 ( 
.A(n_1539),
.Y(n_1678)
);

BUFx8_ASAP7_75t_L g1679 ( 
.A(n_1541),
.Y(n_1679)
);

NOR3xp33_ASAP7_75t_L g1680 ( 
.A(n_1537),
.B(n_995),
.C(n_994),
.Y(n_1680)
);

NOR2xp33_ASAP7_75t_SL g1681 ( 
.A(n_1525),
.B(n_1206),
.Y(n_1681)
);

NAND2xp5_ASAP7_75t_L g1682 ( 
.A(n_1571),
.B(n_1256),
.Y(n_1682)
);

NOR2xp33_ASAP7_75t_L g1683 ( 
.A(n_1577),
.B(n_1207),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1578),
.B(n_1257),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_L g1685 ( 
.A(n_1586),
.B(n_1267),
.Y(n_1685)
);

NAND2xp5_ASAP7_75t_L g1686 ( 
.A(n_1588),
.B(n_984),
.Y(n_1686)
);

INVx2_ASAP7_75t_L g1687 ( 
.A(n_1475),
.Y(n_1687)
);

NOR2xp33_ASAP7_75t_L g1688 ( 
.A(n_1542),
.B(n_1264),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_L g1689 ( 
.A(n_1553),
.B(n_1560),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1544),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_L g1691 ( 
.A(n_1565),
.B(n_985),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_SL g1692 ( 
.A(n_1480),
.B(n_996),
.Y(n_1692)
);

OR2x6_ASAP7_75t_L g1693 ( 
.A(n_1535),
.B(n_1147),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1550),
.Y(n_1694)
);

INVx4_ASAP7_75t_L g1695 ( 
.A(n_1485),
.Y(n_1695)
);

NAND2xp5_ASAP7_75t_SL g1696 ( 
.A(n_1536),
.B(n_997),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_SL g1697 ( 
.A(n_1533),
.B(n_999),
.Y(n_1697)
);

BUFx5_ASAP7_75t_L g1698 ( 
.A(n_1562),
.Y(n_1698)
);

INVx2_ASAP7_75t_L g1699 ( 
.A(n_1483),
.Y(n_1699)
);

NOR2xp33_ASAP7_75t_L g1700 ( 
.A(n_1524),
.B(n_1282),
.Y(n_1700)
);

OR2x6_ASAP7_75t_L g1701 ( 
.A(n_1551),
.B(n_1150),
.Y(n_1701)
);

AND2x2_ASAP7_75t_L g1702 ( 
.A(n_1551),
.B(n_1118),
.Y(n_1702)
);

NOR2xp33_ASAP7_75t_L g1703 ( 
.A(n_1531),
.B(n_998),
.Y(n_1703)
);

NAND2xp5_ASAP7_75t_L g1704 ( 
.A(n_1508),
.B(n_1008),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1558),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1558),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1496),
.B(n_1548),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_SL g1708 ( 
.A(n_1503),
.B(n_1010),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1489),
.Y(n_1709)
);

NOR2xp33_ASAP7_75t_L g1710 ( 
.A(n_1479),
.B(n_1003),
.Y(n_1710)
);

HB1xp67_ASAP7_75t_L g1711 ( 
.A(n_1561),
.Y(n_1711)
);

NAND2xp5_ASAP7_75t_L g1712 ( 
.A(n_1479),
.B(n_1016),
.Y(n_1712)
);

AOI22xp33_ASAP7_75t_L g1713 ( 
.A1(n_1479),
.A2(n_982),
.B1(n_1117),
.B2(n_1099),
.Y(n_1713)
);

AND2x2_ASAP7_75t_L g1714 ( 
.A(n_1479),
.B(n_1159),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_1479),
.B(n_1019),
.Y(n_1715)
);

INVx8_ASAP7_75t_L g1716 ( 
.A(n_1528),
.Y(n_1716)
);

NOR2xp33_ASAP7_75t_L g1717 ( 
.A(n_1479),
.B(n_1004),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1489),
.Y(n_1718)
);

INVx4_ASAP7_75t_L g1719 ( 
.A(n_1528),
.Y(n_1719)
);

INVx2_ASAP7_75t_L g1720 ( 
.A(n_1500),
.Y(n_1720)
);

INVx2_ASAP7_75t_L g1721 ( 
.A(n_1500),
.Y(n_1721)
);

INVxp67_ASAP7_75t_L g1722 ( 
.A(n_1561),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_L g1723 ( 
.A(n_1479),
.B(n_1021),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1489),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_L g1725 ( 
.A(n_1479),
.B(n_1022),
.Y(n_1725)
);

AOI21xp5_ASAP7_75t_L g1726 ( 
.A1(n_1500),
.A2(n_1009),
.B(n_941),
.Y(n_1726)
);

NAND2xp5_ASAP7_75t_L g1727 ( 
.A(n_1479),
.B(n_1023),
.Y(n_1727)
);

AND2x2_ASAP7_75t_L g1728 ( 
.A(n_1479),
.B(n_1159),
.Y(n_1728)
);

CKINVDCx5p33_ASAP7_75t_R g1729 ( 
.A(n_1520),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_L g1730 ( 
.A(n_1479),
.B(n_1025),
.Y(n_1730)
);

OR2x6_ASAP7_75t_L g1731 ( 
.A(n_1509),
.B(n_1155),
.Y(n_1731)
);

AND2x2_ASAP7_75t_L g1732 ( 
.A(n_1479),
.B(n_1193),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1489),
.Y(n_1733)
);

NOR2xp33_ASAP7_75t_L g1734 ( 
.A(n_1479),
.B(n_1006),
.Y(n_1734)
);

NAND2xp5_ASAP7_75t_SL g1735 ( 
.A(n_1478),
.B(n_1031),
.Y(n_1735)
);

AND2x2_ASAP7_75t_L g1736 ( 
.A(n_1479),
.B(n_1193),
.Y(n_1736)
);

NOR2xp33_ASAP7_75t_SL g1737 ( 
.A(n_1552),
.B(n_1250),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1489),
.Y(n_1738)
);

NOR2x1_ASAP7_75t_L g1739 ( 
.A(n_1523),
.B(n_1157),
.Y(n_1739)
);

NOR2xp33_ASAP7_75t_L g1740 ( 
.A(n_1479),
.B(n_1012),
.Y(n_1740)
);

AND2x4_ASAP7_75t_L g1741 ( 
.A(n_1528),
.B(n_1161),
.Y(n_1741)
);

NAND2xp5_ASAP7_75t_L g1742 ( 
.A(n_1479),
.B(n_1033),
.Y(n_1742)
);

NAND2xp5_ASAP7_75t_L g1743 ( 
.A(n_1479),
.B(n_1036),
.Y(n_1743)
);

AND2x2_ASAP7_75t_L g1744 ( 
.A(n_1479),
.B(n_1250),
.Y(n_1744)
);

INVx2_ASAP7_75t_L g1745 ( 
.A(n_1500),
.Y(n_1745)
);

NOR2xp33_ASAP7_75t_L g1746 ( 
.A(n_1479),
.B(n_1014),
.Y(n_1746)
);

INVx2_ASAP7_75t_L g1747 ( 
.A(n_1500),
.Y(n_1747)
);

NAND2xp5_ASAP7_75t_L g1748 ( 
.A(n_1479),
.B(n_1042),
.Y(n_1748)
);

INVx2_ASAP7_75t_L g1749 ( 
.A(n_1500),
.Y(n_1749)
);

BUFx5_ASAP7_75t_L g1750 ( 
.A(n_1527),
.Y(n_1750)
);

AND2x6_ASAP7_75t_SL g1751 ( 
.A(n_1537),
.B(n_1166),
.Y(n_1751)
);

OAI21xp33_ASAP7_75t_L g1752 ( 
.A1(n_1710),
.A2(n_1024),
.B(n_1017),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1600),
.Y(n_1753)
);

INVx1_ASAP7_75t_SL g1754 ( 
.A(n_1638),
.Y(n_1754)
);

AOI21x1_ASAP7_75t_L g1755 ( 
.A1(n_1726),
.A2(n_1208),
.B(n_1201),
.Y(n_1755)
);

AOI21xp5_ASAP7_75t_L g1756 ( 
.A1(n_1591),
.A2(n_1009),
.B(n_941),
.Y(n_1756)
);

NAND2xp5_ASAP7_75t_L g1757 ( 
.A(n_1635),
.B(n_1046),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1665),
.Y(n_1758)
);

AOI21xp5_ASAP7_75t_L g1759 ( 
.A1(n_1592),
.A2(n_1009),
.B(n_941),
.Y(n_1759)
);

AOI21xp5_ASAP7_75t_L g1760 ( 
.A1(n_1601),
.A2(n_1191),
.B(n_1093),
.Y(n_1760)
);

INVx2_ASAP7_75t_L g1761 ( 
.A(n_1720),
.Y(n_1761)
);

INVx2_ASAP7_75t_L g1762 ( 
.A(n_1721),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1648),
.Y(n_1763)
);

NAND2xp5_ASAP7_75t_SL g1764 ( 
.A(n_1605),
.B(n_1054),
.Y(n_1764)
);

INVx4_ASAP7_75t_L g1765 ( 
.A(n_1641),
.Y(n_1765)
);

CKINVDCx5p33_ASAP7_75t_R g1766 ( 
.A(n_1729),
.Y(n_1766)
);

INVx2_ASAP7_75t_L g1767 ( 
.A(n_1745),
.Y(n_1767)
);

NAND2xp5_ASAP7_75t_SL g1768 ( 
.A(n_1668),
.B(n_1056),
.Y(n_1768)
);

NAND2xp5_ASAP7_75t_SL g1769 ( 
.A(n_1646),
.B(n_1059),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_SL g1770 ( 
.A(n_1631),
.B(n_1062),
.Y(n_1770)
);

INVxp67_ASAP7_75t_L g1771 ( 
.A(n_1711),
.Y(n_1771)
);

NAND2xp5_ASAP7_75t_L g1772 ( 
.A(n_1717),
.B(n_1066),
.Y(n_1772)
);

AOI21xp5_ASAP7_75t_L g1773 ( 
.A1(n_1747),
.A2(n_1191),
.B(n_1093),
.Y(n_1773)
);

AOI21xp5_ASAP7_75t_L g1774 ( 
.A1(n_1749),
.A2(n_1191),
.B(n_1093),
.Y(n_1774)
);

OAI21xp5_ASAP7_75t_L g1775 ( 
.A1(n_1673),
.A2(n_1069),
.B(n_1068),
.Y(n_1775)
);

NOR2xp33_ASAP7_75t_L g1776 ( 
.A(n_1598),
.B(n_1734),
.Y(n_1776)
);

AOI21xp5_ASAP7_75t_L g1777 ( 
.A1(n_1610),
.A2(n_1261),
.B(n_1254),
.Y(n_1777)
);

NAND2xp5_ASAP7_75t_L g1778 ( 
.A(n_1740),
.B(n_1070),
.Y(n_1778)
);

NAND2xp5_ASAP7_75t_SL g1779 ( 
.A(n_1639),
.B(n_1071),
.Y(n_1779)
);

NAND2xp5_ASAP7_75t_SL g1780 ( 
.A(n_1681),
.B(n_1072),
.Y(n_1780)
);

NAND2xp5_ASAP7_75t_L g1781 ( 
.A(n_1746),
.B(n_1073),
.Y(n_1781)
);

AOI21xp5_ASAP7_75t_L g1782 ( 
.A1(n_1616),
.A2(n_1265),
.B(n_1263),
.Y(n_1782)
);

AOI21xp5_ASAP7_75t_L g1783 ( 
.A1(n_1626),
.A2(n_1611),
.B(n_1689),
.Y(n_1783)
);

AOI21xp5_ASAP7_75t_L g1784 ( 
.A1(n_1712),
.A2(n_1748),
.B(n_1743),
.Y(n_1784)
);

NAND2xp5_ASAP7_75t_L g1785 ( 
.A(n_1596),
.B(n_1076),
.Y(n_1785)
);

AOI21xp5_ASAP7_75t_L g1786 ( 
.A1(n_1715),
.A2(n_1275),
.B(n_1268),
.Y(n_1786)
);

INVx2_ASAP7_75t_L g1787 ( 
.A(n_1750),
.Y(n_1787)
);

NOR2x1_ASAP7_75t_L g1788 ( 
.A(n_1678),
.B(n_1226),
.Y(n_1788)
);

INVx2_ASAP7_75t_L g1789 ( 
.A(n_1750),
.Y(n_1789)
);

INVx2_ASAP7_75t_L g1790 ( 
.A(n_1750),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1655),
.Y(n_1791)
);

INVxp67_ASAP7_75t_L g1792 ( 
.A(n_1618),
.Y(n_1792)
);

AOI21xp5_ASAP7_75t_L g1793 ( 
.A1(n_1723),
.A2(n_1080),
.B(n_1079),
.Y(n_1793)
);

NAND2xp5_ASAP7_75t_L g1794 ( 
.A(n_1725),
.B(n_1090),
.Y(n_1794)
);

AOI21xp5_ASAP7_75t_L g1795 ( 
.A1(n_1727),
.A2(n_1097),
.B(n_1095),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1615),
.Y(n_1796)
);

AOI21xp5_ASAP7_75t_L g1797 ( 
.A1(n_1730),
.A2(n_1252),
.B(n_1248),
.Y(n_1797)
);

AO21x1_ASAP7_75t_L g1798 ( 
.A1(n_1632),
.A2(n_1238),
.B(n_1230),
.Y(n_1798)
);

INVx2_ASAP7_75t_L g1799 ( 
.A(n_1750),
.Y(n_1799)
);

NAND2x1_ASAP7_75t_L g1800 ( 
.A(n_1614),
.B(n_1242),
.Y(n_1800)
);

NAND2xp5_ASAP7_75t_L g1801 ( 
.A(n_1742),
.B(n_1100),
.Y(n_1801)
);

AOI22xp5_ASAP7_75t_L g1802 ( 
.A1(n_1667),
.A2(n_1113),
.B1(n_1138),
.B2(n_1124),
.Y(n_1802)
);

NAND2xp5_ASAP7_75t_L g1803 ( 
.A(n_1714),
.B(n_1139),
.Y(n_1803)
);

AOI21xp5_ASAP7_75t_L g1804 ( 
.A1(n_1672),
.A2(n_1151),
.B(n_1143),
.Y(n_1804)
);

INVx2_ASAP7_75t_L g1805 ( 
.A(n_1619),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1622),
.Y(n_1806)
);

NAND2xp5_ASAP7_75t_L g1807 ( 
.A(n_1728),
.B(n_1162),
.Y(n_1807)
);

OAI21xp5_ASAP7_75t_L g1808 ( 
.A1(n_1629),
.A2(n_1169),
.B(n_1164),
.Y(n_1808)
);

AOI21xp5_ASAP7_75t_L g1809 ( 
.A1(n_1609),
.A2(n_1735),
.B(n_1627),
.Y(n_1809)
);

INVx2_ASAP7_75t_L g1810 ( 
.A(n_1621),
.Y(n_1810)
);

OAI22xp5_ASAP7_75t_L g1811 ( 
.A1(n_1695),
.A2(n_1178),
.B1(n_1180),
.B2(n_1177),
.Y(n_1811)
);

INVxp67_ASAP7_75t_L g1812 ( 
.A(n_1660),
.Y(n_1812)
);

NAND2xp5_ASAP7_75t_L g1813 ( 
.A(n_1732),
.B(n_1181),
.Y(n_1813)
);

AND2x4_ASAP7_75t_L g1814 ( 
.A(n_1719),
.B(n_1243),
.Y(n_1814)
);

AO22x1_ASAP7_75t_L g1815 ( 
.A1(n_1736),
.A2(n_1744),
.B1(n_1700),
.B2(n_1688),
.Y(n_1815)
);

NOR2xp33_ASAP7_75t_L g1816 ( 
.A(n_1722),
.B(n_1027),
.Y(n_1816)
);

OAI21xp5_ASAP7_75t_L g1817 ( 
.A1(n_1652),
.A2(n_1187),
.B(n_1182),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1623),
.Y(n_1818)
);

O2A1O1Ixp33_ASAP7_75t_L g1819 ( 
.A1(n_1612),
.A2(n_1258),
.B(n_1260),
.C(n_1246),
.Y(n_1819)
);

AOI21x1_ASAP7_75t_L g1820 ( 
.A1(n_1659),
.A2(n_1279),
.B(n_1266),
.Y(n_1820)
);

NAND2xp5_ASAP7_75t_L g1821 ( 
.A(n_1624),
.B(n_1188),
.Y(n_1821)
);

AOI22xp33_ASAP7_75t_L g1822 ( 
.A1(n_1594),
.A2(n_1117),
.B1(n_1099),
.B2(n_1189),
.Y(n_1822)
);

AOI21xp5_ASAP7_75t_L g1823 ( 
.A1(n_1697),
.A2(n_1205),
.B(n_1198),
.Y(n_1823)
);

AND2x2_ASAP7_75t_SL g1824 ( 
.A(n_1597),
.B(n_1173),
.Y(n_1824)
);

AOI21xp5_ASAP7_75t_L g1825 ( 
.A1(n_1704),
.A2(n_1234),
.B(n_1217),
.Y(n_1825)
);

AO22x1_ASAP7_75t_L g1826 ( 
.A1(n_1683),
.A2(n_1030),
.B1(n_1035),
.B2(n_1029),
.Y(n_1826)
);

OAI22xp5_ASAP7_75t_L g1827 ( 
.A1(n_1634),
.A2(n_1221),
.B1(n_1223),
.B2(n_1215),
.Y(n_1827)
);

AOI21x1_ASAP7_75t_L g1828 ( 
.A1(n_1664),
.A2(n_1280),
.B(n_1176),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1677),
.Y(n_1829)
);

NAND2xp5_ASAP7_75t_L g1830 ( 
.A(n_1636),
.B(n_1038),
.Y(n_1830)
);

NAND2xp5_ASAP7_75t_L g1831 ( 
.A(n_1703),
.B(n_1039),
.Y(n_1831)
);

AOI21xp5_ASAP7_75t_L g1832 ( 
.A1(n_1643),
.A2(n_643),
.B(n_641),
.Y(n_1832)
);

AOI22xp5_ASAP7_75t_L g1833 ( 
.A1(n_1607),
.A2(n_1117),
.B1(n_1099),
.B2(n_1044),
.Y(n_1833)
);

NAND2xp5_ASAP7_75t_L g1834 ( 
.A(n_1640),
.B(n_1041),
.Y(n_1834)
);

AND2x2_ASAP7_75t_L g1835 ( 
.A(n_1657),
.B(n_1045),
.Y(n_1835)
);

BUFx2_ASAP7_75t_L g1836 ( 
.A(n_1630),
.Y(n_1836)
);

AOI22xp33_ASAP7_75t_L g1837 ( 
.A1(n_1663),
.A2(n_1117),
.B1(n_1099),
.B2(n_1048),
.Y(n_1837)
);

NOR2xp33_ASAP7_75t_L g1838 ( 
.A(n_1676),
.B(n_1656),
.Y(n_1838)
);

AND2x4_ASAP7_75t_L g1839 ( 
.A(n_1641),
.B(n_644),
.Y(n_1839)
);

AOI22xp33_ASAP7_75t_L g1840 ( 
.A1(n_1713),
.A2(n_1117),
.B1(n_1049),
.B2(n_1063),
.Y(n_1840)
);

NAND2xp5_ASAP7_75t_L g1841 ( 
.A(n_1654),
.B(n_1047),
.Y(n_1841)
);

AOI21xp5_ASAP7_75t_L g1842 ( 
.A1(n_1686),
.A2(n_646),
.B(n_645),
.Y(n_1842)
);

NAND2xp5_ASAP7_75t_L g1843 ( 
.A(n_1661),
.B(n_1064),
.Y(n_1843)
);

NAND2xp5_ASAP7_75t_L g1844 ( 
.A(n_1602),
.B(n_1067),
.Y(n_1844)
);

INVx2_ASAP7_75t_L g1845 ( 
.A(n_1669),
.Y(n_1845)
);

O2A1O1Ixp33_ASAP7_75t_L g1846 ( 
.A1(n_1707),
.A2(n_1092),
.B(n_1094),
.C(n_1085),
.Y(n_1846)
);

AOI21xp5_ASAP7_75t_L g1847 ( 
.A1(n_1642),
.A2(n_649),
.B(n_648),
.Y(n_1847)
);

NAND2xp5_ASAP7_75t_L g1848 ( 
.A(n_1675),
.B(n_1096),
.Y(n_1848)
);

AOI21xp5_ASAP7_75t_L g1849 ( 
.A1(n_1692),
.A2(n_651),
.B(n_650),
.Y(n_1849)
);

NAND2xp5_ASAP7_75t_L g1850 ( 
.A(n_1682),
.B(n_1101),
.Y(n_1850)
);

NOR2xp33_ASAP7_75t_L g1851 ( 
.A(n_1628),
.B(n_1102),
.Y(n_1851)
);

AOI21xp5_ASAP7_75t_L g1852 ( 
.A1(n_1666),
.A2(n_654),
.B(n_652),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1674),
.Y(n_1853)
);

INVxp67_ASAP7_75t_L g1854 ( 
.A(n_1630),
.Y(n_1854)
);

OAI21xp5_ASAP7_75t_L g1855 ( 
.A1(n_1604),
.A2(n_1108),
.B(n_1104),
.Y(n_1855)
);

AOI21x1_ASAP7_75t_L g1856 ( 
.A1(n_1696),
.A2(n_656),
.B(n_655),
.Y(n_1856)
);

INVx2_ASAP7_75t_L g1857 ( 
.A(n_1687),
.Y(n_1857)
);

O2A1O1Ixp33_ASAP7_75t_L g1858 ( 
.A1(n_1613),
.A2(n_1110),
.B(n_1114),
.C(n_1109),
.Y(n_1858)
);

AOI21xp5_ASAP7_75t_L g1859 ( 
.A1(n_1691),
.A2(n_658),
.B(n_657),
.Y(n_1859)
);

INVx2_ASAP7_75t_L g1860 ( 
.A(n_1694),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1684),
.Y(n_1861)
);

AOI21xp5_ASAP7_75t_L g1862 ( 
.A1(n_1685),
.A2(n_660),
.B(n_659),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1593),
.Y(n_1863)
);

INVx2_ASAP7_75t_L g1864 ( 
.A(n_1709),
.Y(n_1864)
);

HB1xp67_ASAP7_75t_L g1865 ( 
.A(n_1620),
.Y(n_1865)
);

AOI21xp5_ASAP7_75t_L g1866 ( 
.A1(n_1649),
.A2(n_662),
.B(n_661),
.Y(n_1866)
);

NAND2xp5_ASAP7_75t_L g1867 ( 
.A(n_1698),
.B(n_1116),
.Y(n_1867)
);

NAND2xp5_ASAP7_75t_L g1868 ( 
.A(n_1698),
.B(n_1119),
.Y(n_1868)
);

AOI21xp5_ASAP7_75t_L g1869 ( 
.A1(n_1637),
.A2(n_665),
.B(n_664),
.Y(n_1869)
);

AOI21xp5_ASAP7_75t_L g1870 ( 
.A1(n_1783),
.A2(n_1647),
.B(n_1651),
.Y(n_1870)
);

AOI21xp5_ASAP7_75t_L g1871 ( 
.A1(n_1784),
.A2(n_1670),
.B(n_1718),
.Y(n_1871)
);

INVx2_ASAP7_75t_L g1872 ( 
.A(n_1753),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1829),
.Y(n_1873)
);

NOR2xp33_ASAP7_75t_L g1874 ( 
.A(n_1776),
.B(n_1644),
.Y(n_1874)
);

OAI21xp33_ASAP7_75t_SL g1875 ( 
.A1(n_1861),
.A2(n_1758),
.B(n_1770),
.Y(n_1875)
);

INVx2_ASAP7_75t_L g1876 ( 
.A(n_1763),
.Y(n_1876)
);

O2A1O1Ixp5_ASAP7_75t_L g1877 ( 
.A1(n_1815),
.A2(n_1671),
.B(n_1708),
.C(n_1699),
.Y(n_1877)
);

NAND2xp5_ASAP7_75t_L g1878 ( 
.A(n_1757),
.B(n_1698),
.Y(n_1878)
);

A2O1A1Ixp33_ASAP7_75t_SL g1879 ( 
.A1(n_1838),
.A2(n_1680),
.B(n_1706),
.C(n_1705),
.Y(n_1879)
);

NAND3xp33_ASAP7_75t_SL g1880 ( 
.A(n_1831),
.B(n_1737),
.C(n_1606),
.Y(n_1880)
);

HB1xp67_ASAP7_75t_L g1881 ( 
.A(n_1754),
.Y(n_1881)
);

AOI21xp5_ASAP7_75t_L g1882 ( 
.A1(n_1809),
.A2(n_1778),
.B(n_1772),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1791),
.Y(n_1883)
);

OAI22x1_ASAP7_75t_L g1884 ( 
.A1(n_1851),
.A2(n_1608),
.B1(n_1741),
.B2(n_1739),
.Y(n_1884)
);

O2A1O1Ixp33_ASAP7_75t_L g1885 ( 
.A1(n_1752),
.A2(n_1662),
.B(n_1702),
.C(n_1731),
.Y(n_1885)
);

NAND2xp5_ASAP7_75t_SL g1886 ( 
.A(n_1792),
.B(n_1698),
.Y(n_1886)
);

CKINVDCx8_ASAP7_75t_R g1887 ( 
.A(n_1766),
.Y(n_1887)
);

INVxp67_ASAP7_75t_L g1888 ( 
.A(n_1836),
.Y(n_1888)
);

NAND2xp5_ASAP7_75t_L g1889 ( 
.A(n_1781),
.B(n_1645),
.Y(n_1889)
);

O2A1O1Ixp33_ASAP7_75t_L g1890 ( 
.A1(n_1803),
.A2(n_1662),
.B(n_1731),
.C(n_1701),
.Y(n_1890)
);

AOI21xp5_ASAP7_75t_L g1891 ( 
.A1(n_1794),
.A2(n_1733),
.B(n_1724),
.Y(n_1891)
);

A2O1A1Ixp33_ASAP7_75t_L g1892 ( 
.A1(n_1858),
.A2(n_1846),
.B(n_1775),
.C(n_1855),
.Y(n_1892)
);

NAND3xp33_ASAP7_75t_L g1893 ( 
.A(n_1802),
.B(n_1679),
.C(n_1690),
.Y(n_1893)
);

AOI21xp5_ASAP7_75t_L g1894 ( 
.A1(n_1801),
.A2(n_1785),
.B(n_1787),
.Y(n_1894)
);

OR2x2_ASAP7_75t_L g1895 ( 
.A(n_1771),
.B(n_1650),
.Y(n_1895)
);

NOR2xp33_ASAP7_75t_L g1896 ( 
.A(n_1807),
.B(n_1603),
.Y(n_1896)
);

INVx1_ASAP7_75t_L g1897 ( 
.A(n_1761),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_1762),
.Y(n_1898)
);

NAND2xp5_ASAP7_75t_L g1899 ( 
.A(n_1830),
.B(n_1645),
.Y(n_1899)
);

AOI21xp5_ASAP7_75t_L g1900 ( 
.A1(n_1789),
.A2(n_1799),
.B(n_1790),
.Y(n_1900)
);

NOR2xp33_ASAP7_75t_L g1901 ( 
.A(n_1813),
.B(n_1650),
.Y(n_1901)
);

BUFx3_ASAP7_75t_L g1902 ( 
.A(n_1765),
.Y(n_1902)
);

O2A1O1Ixp33_ASAP7_75t_L g1903 ( 
.A1(n_1844),
.A2(n_1701),
.B(n_1738),
.C(n_1693),
.Y(n_1903)
);

INVx2_ASAP7_75t_L g1904 ( 
.A(n_1767),
.Y(n_1904)
);

NAND2xp5_ASAP7_75t_L g1905 ( 
.A(n_1848),
.B(n_1645),
.Y(n_1905)
);

CKINVDCx20_ASAP7_75t_R g1906 ( 
.A(n_1765),
.Y(n_1906)
);

NAND2xp5_ASAP7_75t_L g1907 ( 
.A(n_1850),
.B(n_1625),
.Y(n_1907)
);

NOR3xp33_ASAP7_75t_SL g1908 ( 
.A(n_1780),
.B(n_1129),
.C(n_1123),
.Y(n_1908)
);

INVx1_ASAP7_75t_L g1909 ( 
.A(n_1796),
.Y(n_1909)
);

OR2x2_ASAP7_75t_L g1910 ( 
.A(n_1834),
.B(n_1841),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1806),
.Y(n_1911)
);

OAI21xp33_ASAP7_75t_L g1912 ( 
.A1(n_1816),
.A2(n_1595),
.B(n_1693),
.Y(n_1912)
);

NAND2xp5_ASAP7_75t_L g1913 ( 
.A(n_1818),
.B(n_1843),
.Y(n_1913)
);

BUFx6f_ASAP7_75t_L g1914 ( 
.A(n_1839),
.Y(n_1914)
);

AOI21xp5_ASAP7_75t_L g1915 ( 
.A1(n_1859),
.A2(n_1617),
.B(n_1716),
.Y(n_1915)
);

AND2x2_ASAP7_75t_L g1916 ( 
.A(n_1835),
.B(n_1633),
.Y(n_1916)
);

BUFx3_ASAP7_75t_L g1917 ( 
.A(n_1865),
.Y(n_1917)
);

BUFx2_ASAP7_75t_L g1918 ( 
.A(n_1854),
.Y(n_1918)
);

A2O1A1Ixp33_ASAP7_75t_L g1919 ( 
.A1(n_1808),
.A2(n_1716),
.B(n_1653),
.C(n_1134),
.Y(n_1919)
);

NAND2xp5_ASAP7_75t_L g1920 ( 
.A(n_1805),
.B(n_1751),
.Y(n_1920)
);

O2A1O1Ixp33_ASAP7_75t_L g1921 ( 
.A1(n_1768),
.A2(n_1764),
.B(n_1769),
.C(n_1819),
.Y(n_1921)
);

OAI22xp5_ASAP7_75t_L g1922 ( 
.A1(n_1853),
.A2(n_1658),
.B1(n_1135),
.B2(n_1137),
.Y(n_1922)
);

CKINVDCx5p33_ASAP7_75t_R g1923 ( 
.A(n_1812),
.Y(n_1923)
);

OR2x4_ASAP7_75t_L g1924 ( 
.A(n_1863),
.B(n_1599),
.Y(n_1924)
);

HB1xp67_ASAP7_75t_L g1925 ( 
.A(n_1864),
.Y(n_1925)
);

O2A1O1Ixp33_ASAP7_75t_L g1926 ( 
.A1(n_1779),
.A2(n_1144),
.B(n_1146),
.C(n_1133),
.Y(n_1926)
);

AOI21xp5_ASAP7_75t_L g1927 ( 
.A1(n_1842),
.A2(n_667),
.B(n_666),
.Y(n_1927)
);

AOI21x1_ASAP7_75t_L g1928 ( 
.A1(n_1755),
.A2(n_670),
.B(n_668),
.Y(n_1928)
);

AOI21xp5_ASAP7_75t_L g1929 ( 
.A1(n_1849),
.A2(n_672),
.B(n_671),
.Y(n_1929)
);

AND2x4_ASAP7_75t_L g1930 ( 
.A(n_1857),
.B(n_673),
.Y(n_1930)
);

NAND2xp5_ASAP7_75t_L g1931 ( 
.A(n_1810),
.B(n_1149),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_1845),
.Y(n_1932)
);

OAI22xp5_ASAP7_75t_L g1933 ( 
.A1(n_1867),
.A2(n_1160),
.B1(n_1165),
.B2(n_1156),
.Y(n_1933)
);

O2A1O1Ixp33_ASAP7_75t_SL g1934 ( 
.A1(n_1847),
.A2(n_675),
.B(n_676),
.C(n_674),
.Y(n_1934)
);

O2A1O1Ixp5_ASAP7_75t_L g1935 ( 
.A1(n_1798),
.A2(n_1756),
.B(n_1817),
.C(n_1856),
.Y(n_1935)
);

INVx1_ASAP7_75t_L g1936 ( 
.A(n_1860),
.Y(n_1936)
);

INVx3_ASAP7_75t_L g1937 ( 
.A(n_1839),
.Y(n_1937)
);

OR2x2_ASAP7_75t_L g1938 ( 
.A(n_1868),
.B(n_1167),
.Y(n_1938)
);

O2A1O1Ixp33_ASAP7_75t_L g1939 ( 
.A1(n_1800),
.A2(n_1174),
.B(n_1184),
.C(n_1172),
.Y(n_1939)
);

O2A1O1Ixp5_ASAP7_75t_L g1940 ( 
.A1(n_1820),
.A2(n_2),
.B(n_0),
.C(n_1),
.Y(n_1940)
);

AOI21xp5_ASAP7_75t_L g1941 ( 
.A1(n_1852),
.A2(n_680),
.B(n_678),
.Y(n_1941)
);

AO21x1_ASAP7_75t_L g1942 ( 
.A1(n_1869),
.A2(n_3),
.B(n_2),
.Y(n_1942)
);

INVx1_ASAP7_75t_L g1943 ( 
.A(n_1828),
.Y(n_1943)
);

OR2x6_ASAP7_75t_L g1944 ( 
.A(n_1814),
.B(n_681),
.Y(n_1944)
);

INVx2_ASAP7_75t_L g1945 ( 
.A(n_1821),
.Y(n_1945)
);

CKINVDCx6p67_ASAP7_75t_R g1946 ( 
.A(n_1824),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1833),
.Y(n_1947)
);

CKINVDCx11_ASAP7_75t_R g1948 ( 
.A(n_1814),
.Y(n_1948)
);

BUFx6f_ASAP7_75t_L g1949 ( 
.A(n_1788),
.Y(n_1949)
);

AOI22x1_ASAP7_75t_L g1950 ( 
.A1(n_1825),
.A2(n_1194),
.B1(n_1195),
.B2(n_1185),
.Y(n_1950)
);

BUFx2_ASAP7_75t_L g1951 ( 
.A(n_1811),
.Y(n_1951)
);

NAND2xp5_ASAP7_75t_SL g1952 ( 
.A(n_1827),
.B(n_1200),
.Y(n_1952)
);

AOI22xp5_ASAP7_75t_L g1953 ( 
.A1(n_1826),
.A2(n_1209),
.B1(n_1216),
.B2(n_1204),
.Y(n_1953)
);

INVx1_ASAP7_75t_L g1954 ( 
.A(n_1759),
.Y(n_1954)
);

NAND2xp5_ASAP7_75t_SL g1955 ( 
.A(n_1786),
.B(n_1220),
.Y(n_1955)
);

CKINVDCx20_ASAP7_75t_R g1956 ( 
.A(n_1866),
.Y(n_1956)
);

NAND2xp5_ASAP7_75t_SL g1957 ( 
.A(n_1793),
.B(n_1224),
.Y(n_1957)
);

NOR2xp33_ASAP7_75t_L g1958 ( 
.A(n_1795),
.B(n_1225),
.Y(n_1958)
);

NAND2xp5_ASAP7_75t_L g1959 ( 
.A(n_1797),
.B(n_1227),
.Y(n_1959)
);

HB1xp67_ASAP7_75t_L g1960 ( 
.A(n_1777),
.Y(n_1960)
);

BUFx2_ASAP7_75t_L g1961 ( 
.A(n_1837),
.Y(n_1961)
);

OR2x6_ASAP7_75t_L g1962 ( 
.A(n_1832),
.B(n_682),
.Y(n_1962)
);

NAND2xp5_ASAP7_75t_L g1963 ( 
.A(n_1782),
.B(n_1804),
.Y(n_1963)
);

OR2x6_ASAP7_75t_SL g1964 ( 
.A(n_1840),
.B(n_1229),
.Y(n_1964)
);

NAND2xp5_ASAP7_75t_L g1965 ( 
.A(n_1823),
.B(n_1231),
.Y(n_1965)
);

AOI21x1_ASAP7_75t_L g1966 ( 
.A1(n_1760),
.A2(n_684),
.B(n_683),
.Y(n_1966)
);

INVx6_ASAP7_75t_L g1967 ( 
.A(n_1862),
.Y(n_1967)
);

AOI22xp33_ASAP7_75t_L g1968 ( 
.A1(n_1822),
.A2(n_1233),
.B1(n_1235),
.B2(n_1232),
.Y(n_1968)
);

NAND2xp5_ASAP7_75t_SL g1969 ( 
.A(n_1773),
.B(n_1236),
.Y(n_1969)
);

O2A1O1Ixp33_ASAP7_75t_SL g1970 ( 
.A1(n_1774),
.A2(n_686),
.B(n_687),
.C(n_685),
.Y(n_1970)
);

CKINVDCx11_ASAP7_75t_R g1971 ( 
.A(n_1754),
.Y(n_1971)
);

NAND2xp5_ASAP7_75t_L g1972 ( 
.A(n_1776),
.B(n_1253),
.Y(n_1972)
);

O2A1O1Ixp33_ASAP7_75t_L g1973 ( 
.A1(n_1776),
.A2(n_1259),
.B(n_1278),
.C(n_1255),
.Y(n_1973)
);

O2A1O1Ixp33_ASAP7_75t_L g1974 ( 
.A1(n_1776),
.A2(n_1281),
.B(n_4),
.C(n_0),
.Y(n_1974)
);

O2A1O1Ixp33_ASAP7_75t_L g1975 ( 
.A1(n_1776),
.A2(n_5),
.B(n_3),
.C(n_4),
.Y(n_1975)
);

AND3x1_ASAP7_75t_SL g1976 ( 
.A(n_1829),
.B(n_5),
.C(n_6),
.Y(n_1976)
);

AOI22xp33_ASAP7_75t_L g1977 ( 
.A1(n_1776),
.A2(n_9),
.B1(n_7),
.B2(n_8),
.Y(n_1977)
);

AOI22xp33_ASAP7_75t_SL g1978 ( 
.A1(n_1776),
.A2(n_10),
.B1(n_7),
.B2(n_8),
.Y(n_1978)
);

AND2x4_ASAP7_75t_L g1979 ( 
.A(n_1765),
.B(n_689),
.Y(n_1979)
);

NAND2xp5_ASAP7_75t_L g1980 ( 
.A(n_1776),
.B(n_10),
.Y(n_1980)
);

NOR2xp33_ASAP7_75t_L g1981 ( 
.A(n_1776),
.B(n_11),
.Y(n_1981)
);

AOI22xp5_ASAP7_75t_L g1982 ( 
.A1(n_1776),
.A2(n_13),
.B1(n_11),
.B2(n_12),
.Y(n_1982)
);

AOI222xp33_ASAP7_75t_L g1983 ( 
.A1(n_1776),
.A2(n_15),
.B1(n_17),
.B2(n_12),
.C1(n_14),
.C2(n_16),
.Y(n_1983)
);

A2O1A1Ixp33_ASAP7_75t_L g1984 ( 
.A1(n_1776),
.A2(n_16),
.B(n_14),
.C(n_15),
.Y(n_1984)
);

NAND2xp5_ASAP7_75t_L g1985 ( 
.A(n_1776),
.B(n_17),
.Y(n_1985)
);

CKINVDCx5p33_ASAP7_75t_R g1986 ( 
.A(n_1766),
.Y(n_1986)
);

NOR2xp33_ASAP7_75t_L g1987 ( 
.A(n_1776),
.B(n_18),
.Y(n_1987)
);

AND2x2_ASAP7_75t_L g1988 ( 
.A(n_1835),
.B(n_18),
.Y(n_1988)
);

OAI21xp33_ASAP7_75t_SL g1989 ( 
.A1(n_1776),
.A2(n_19),
.B(n_20),
.Y(n_1989)
);

OAI22xp5_ASAP7_75t_L g1990 ( 
.A1(n_1776),
.A2(n_21),
.B1(n_19),
.B2(n_20),
.Y(n_1990)
);

INVx5_ASAP7_75t_L g1991 ( 
.A(n_1765),
.Y(n_1991)
);

INVx3_ASAP7_75t_L g1992 ( 
.A(n_1765),
.Y(n_1992)
);

NOR3xp33_ASAP7_75t_SL g1993 ( 
.A(n_1776),
.B(n_21),
.C(n_22),
.Y(n_1993)
);

NOR2xp33_ASAP7_75t_L g1994 ( 
.A(n_1776),
.B(n_22),
.Y(n_1994)
);

NOR2xp33_ASAP7_75t_R g1995 ( 
.A(n_1766),
.B(n_690),
.Y(n_1995)
);

NAND2xp5_ASAP7_75t_L g1996 ( 
.A(n_1776),
.B(n_23),
.Y(n_1996)
);

INVx1_ASAP7_75t_L g1997 ( 
.A(n_1829),
.Y(n_1997)
);

OAI21xp5_ASAP7_75t_L g1998 ( 
.A1(n_1776),
.A2(n_692),
.B(n_691),
.Y(n_1998)
);

NOR2xp33_ASAP7_75t_L g1999 ( 
.A(n_1776),
.B(n_25),
.Y(n_1999)
);

AOI22xp5_ASAP7_75t_L g2000 ( 
.A1(n_1874),
.A2(n_27),
.B1(n_25),
.B2(n_26),
.Y(n_2000)
);

NAND2xp5_ASAP7_75t_L g2001 ( 
.A(n_1945),
.B(n_26),
.Y(n_2001)
);

CKINVDCx5p33_ASAP7_75t_R g2002 ( 
.A(n_1986),
.Y(n_2002)
);

NAND2xp5_ASAP7_75t_L g2003 ( 
.A(n_1972),
.B(n_27),
.Y(n_2003)
);

OA21x2_ASAP7_75t_L g2004 ( 
.A1(n_1943),
.A2(n_694),
.B(n_693),
.Y(n_2004)
);

NAND2xp5_ASAP7_75t_SL g2005 ( 
.A(n_1981),
.B(n_28),
.Y(n_2005)
);

OA21x2_ASAP7_75t_L g2006 ( 
.A1(n_1935),
.A2(n_696),
.B(n_695),
.Y(n_2006)
);

INVx2_ASAP7_75t_L g2007 ( 
.A(n_1872),
.Y(n_2007)
);

NAND2x1p5_ASAP7_75t_L g2008 ( 
.A(n_1991),
.B(n_698),
.Y(n_2008)
);

NAND2xp5_ASAP7_75t_L g2009 ( 
.A(n_1910),
.B(n_28),
.Y(n_2009)
);

AOI22xp5_ASAP7_75t_L g2010 ( 
.A1(n_1987),
.A2(n_31),
.B1(n_29),
.B2(n_30),
.Y(n_2010)
);

OAI21x1_ASAP7_75t_L g2011 ( 
.A1(n_1882),
.A2(n_701),
.B(n_700),
.Y(n_2011)
);

INVx5_ASAP7_75t_L g2012 ( 
.A(n_1914),
.Y(n_2012)
);

AOI21xp5_ASAP7_75t_L g2013 ( 
.A1(n_1894),
.A2(n_1870),
.B(n_1963),
.Y(n_2013)
);

BUFx6f_ASAP7_75t_L g2014 ( 
.A(n_1971),
.Y(n_2014)
);

OAI21x1_ASAP7_75t_L g2015 ( 
.A1(n_1871),
.A2(n_704),
.B(n_703),
.Y(n_2015)
);

AO32x2_ASAP7_75t_L g2016 ( 
.A1(n_1990),
.A2(n_32),
.A3(n_29),
.B1(n_30),
.B2(n_33),
.Y(n_2016)
);

NAND2xp5_ASAP7_75t_L g2017 ( 
.A(n_1994),
.B(n_32),
.Y(n_2017)
);

INVx1_ASAP7_75t_L g2018 ( 
.A(n_1876),
.Y(n_2018)
);

BUFx8_ASAP7_75t_L g2019 ( 
.A(n_1918),
.Y(n_2019)
);

INVx2_ASAP7_75t_L g2020 ( 
.A(n_1904),
.Y(n_2020)
);

OA21x2_ASAP7_75t_L g2021 ( 
.A1(n_1878),
.A2(n_706),
.B(n_705),
.Y(n_2021)
);

CKINVDCx5p33_ASAP7_75t_R g2022 ( 
.A(n_1887),
.Y(n_2022)
);

NOR4xp25_ASAP7_75t_L g2023 ( 
.A(n_1974),
.B(n_1975),
.C(n_1984),
.D(n_1999),
.Y(n_2023)
);

AOI221xp5_ASAP7_75t_SL g2024 ( 
.A1(n_1980),
.A2(n_35),
.B1(n_33),
.B2(n_34),
.C(n_36),
.Y(n_2024)
);

BUFx8_ASAP7_75t_L g2025 ( 
.A(n_1949),
.Y(n_2025)
);

AOI21x1_ASAP7_75t_L g2026 ( 
.A1(n_1960),
.A2(n_709),
.B(n_708),
.Y(n_2026)
);

AOI21x1_ASAP7_75t_L g2027 ( 
.A1(n_1889),
.A2(n_712),
.B(n_711),
.Y(n_2027)
);

NAND2xp5_ASAP7_75t_L g2028 ( 
.A(n_1907),
.B(n_35),
.Y(n_2028)
);

AOI21xp5_ASAP7_75t_L g2029 ( 
.A1(n_1892),
.A2(n_910),
.B(n_909),
.Y(n_2029)
);

OAI21xp5_ASAP7_75t_SL g2030 ( 
.A1(n_1885),
.A2(n_38),
.B(n_37),
.Y(n_2030)
);

NOR2xp33_ASAP7_75t_L g2031 ( 
.A(n_1923),
.B(n_713),
.Y(n_2031)
);

AO32x2_ASAP7_75t_L g2032 ( 
.A1(n_1933),
.A2(n_38),
.A3(n_36),
.B1(n_37),
.B2(n_41),
.Y(n_2032)
);

NAND2xp5_ASAP7_75t_L g2033 ( 
.A(n_1913),
.B(n_41),
.Y(n_2033)
);

NAND2xp5_ASAP7_75t_L g2034 ( 
.A(n_1896),
.B(n_42),
.Y(n_2034)
);

AO21x2_ASAP7_75t_L g2035 ( 
.A1(n_1954),
.A2(n_715),
.B(n_714),
.Y(n_2035)
);

AOI21xp5_ASAP7_75t_SL g2036 ( 
.A1(n_1998),
.A2(n_717),
.B(n_716),
.Y(n_2036)
);

INVx1_ASAP7_75t_L g2037 ( 
.A(n_1873),
.Y(n_2037)
);

NAND2xp5_ASAP7_75t_SL g2038 ( 
.A(n_1985),
.B(n_1996),
.Y(n_2038)
);

INVx1_ASAP7_75t_L g2039 ( 
.A(n_1883),
.Y(n_2039)
);

OAI21x1_ASAP7_75t_L g2040 ( 
.A1(n_1900),
.A2(n_719),
.B(n_718),
.Y(n_2040)
);

INVx1_ASAP7_75t_SL g2041 ( 
.A(n_1881),
.Y(n_2041)
);

AO31x2_ASAP7_75t_L g2042 ( 
.A1(n_1942),
.A2(n_1947),
.A3(n_1927),
.B(n_1919),
.Y(n_2042)
);

AND2x2_ASAP7_75t_L g2043 ( 
.A(n_1988),
.B(n_42),
.Y(n_2043)
);

NAND3xp33_ASAP7_75t_L g2044 ( 
.A(n_1983),
.B(n_43),
.C(n_44),
.Y(n_2044)
);

INVx8_ASAP7_75t_L g2045 ( 
.A(n_1991),
.Y(n_2045)
);

OAI21xp5_ASAP7_75t_SL g2046 ( 
.A1(n_1982),
.A2(n_1880),
.B(n_1978),
.Y(n_2046)
);

AND2x2_ASAP7_75t_L g2047 ( 
.A(n_1916),
.B(n_43),
.Y(n_2047)
);

BUFx6f_ASAP7_75t_L g2048 ( 
.A(n_1902),
.Y(n_2048)
);

O2A1O1Ixp5_ASAP7_75t_L g2049 ( 
.A1(n_1877),
.A2(n_47),
.B(n_45),
.C(n_46),
.Y(n_2049)
);

AO31x2_ASAP7_75t_L g2050 ( 
.A1(n_1929),
.A2(n_722),
.A3(n_724),
.B(n_721),
.Y(n_2050)
);

INVxp67_ASAP7_75t_L g2051 ( 
.A(n_1917),
.Y(n_2051)
);

BUFx6f_ASAP7_75t_L g2052 ( 
.A(n_1991),
.Y(n_2052)
);

INVx2_ASAP7_75t_L g2053 ( 
.A(n_1997),
.Y(n_2053)
);

OAI22xp5_ASAP7_75t_L g2054 ( 
.A1(n_1937),
.A2(n_49),
.B1(n_47),
.B2(n_48),
.Y(n_2054)
);

INVx1_ASAP7_75t_L g2055 ( 
.A(n_1909),
.Y(n_2055)
);

AOI221xp5_ASAP7_75t_SL g2056 ( 
.A1(n_1973),
.A2(n_50),
.B1(n_48),
.B2(n_49),
.C(n_51),
.Y(n_2056)
);

A2O1A1Ixp33_ASAP7_75t_L g2057 ( 
.A1(n_1958),
.A2(n_52),
.B(n_50),
.C(n_51),
.Y(n_2057)
);

OAI21x1_ASAP7_75t_L g2058 ( 
.A1(n_1928),
.A2(n_726),
.B(n_725),
.Y(n_2058)
);

BUFx6f_ASAP7_75t_L g2059 ( 
.A(n_1914),
.Y(n_2059)
);

OAI21xp5_ASAP7_75t_L g2060 ( 
.A1(n_1875),
.A2(n_53),
.B(n_54),
.Y(n_2060)
);

CKINVDCx5p33_ASAP7_75t_R g2061 ( 
.A(n_1906),
.Y(n_2061)
);

NAND2xp5_ASAP7_75t_L g2062 ( 
.A(n_1925),
.B(n_53),
.Y(n_2062)
);

OAI21x1_ASAP7_75t_L g2063 ( 
.A1(n_1966),
.A2(n_732),
.B(n_729),
.Y(n_2063)
);

NAND2xp5_ASAP7_75t_SL g2064 ( 
.A(n_1912),
.B(n_54),
.Y(n_2064)
);

NAND2xp5_ASAP7_75t_L g2065 ( 
.A(n_1901),
.B(n_55),
.Y(n_2065)
);

AOI21xp5_ASAP7_75t_L g2066 ( 
.A1(n_1891),
.A2(n_912),
.B(n_911),
.Y(n_2066)
);

NAND2xp5_ASAP7_75t_L g2067 ( 
.A(n_1899),
.B(n_56),
.Y(n_2067)
);

INVx1_ASAP7_75t_L g2068 ( 
.A(n_1911),
.Y(n_2068)
);

BUFx2_ASAP7_75t_L g2069 ( 
.A(n_1888),
.Y(n_2069)
);

NAND3xp33_ASAP7_75t_L g2070 ( 
.A(n_1993),
.B(n_56),
.C(n_57),
.Y(n_2070)
);

NOR2xp67_ASAP7_75t_SL g2071 ( 
.A(n_1893),
.B(n_57),
.Y(n_2071)
);

A2O1A1Ixp33_ASAP7_75t_L g2072 ( 
.A1(n_1921),
.A2(n_60),
.B(n_58),
.C(n_59),
.Y(n_2072)
);

NAND2xp5_ASAP7_75t_L g2073 ( 
.A(n_1905),
.B(n_58),
.Y(n_2073)
);

INVx1_ASAP7_75t_L g2074 ( 
.A(n_1936),
.Y(n_2074)
);

CKINVDCx5p33_ASAP7_75t_R g2075 ( 
.A(n_1995),
.Y(n_2075)
);

OAI21x1_ASAP7_75t_SL g2076 ( 
.A1(n_1915),
.A2(n_60),
.B(n_61),
.Y(n_2076)
);

NAND2xp5_ASAP7_75t_L g2077 ( 
.A(n_1951),
.B(n_61),
.Y(n_2077)
);

INVx1_ASAP7_75t_L g2078 ( 
.A(n_1897),
.Y(n_2078)
);

AND2x2_ASAP7_75t_L g2079 ( 
.A(n_1964),
.B(n_62),
.Y(n_2079)
);

OAI21xp5_ASAP7_75t_L g2080 ( 
.A1(n_1959),
.A2(n_1938),
.B(n_1961),
.Y(n_2080)
);

INVx1_ASAP7_75t_L g2081 ( 
.A(n_1898),
.Y(n_2081)
);

INVx1_ASAP7_75t_L g2082 ( 
.A(n_1932),
.Y(n_2082)
);

AO21x1_ASAP7_75t_L g2083 ( 
.A1(n_2060),
.A2(n_2030),
.B(n_2046),
.Y(n_2083)
);

AND2x4_ASAP7_75t_L g2084 ( 
.A(n_2012),
.B(n_1895),
.Y(n_2084)
);

OA21x2_ASAP7_75t_L g2085 ( 
.A1(n_2049),
.A2(n_1940),
.B(n_1941),
.Y(n_2085)
);

OAI21xp5_ASAP7_75t_L g2086 ( 
.A1(n_2023),
.A2(n_2080),
.B(n_2038),
.Y(n_2086)
);

INVx1_ASAP7_75t_L g2087 ( 
.A(n_2037),
.Y(n_2087)
);

INVx2_ASAP7_75t_L g2088 ( 
.A(n_2007),
.Y(n_2088)
);

OAI21x1_ASAP7_75t_L g2089 ( 
.A1(n_2013),
.A2(n_1969),
.B(n_1886),
.Y(n_2089)
);

AOI22xp33_ASAP7_75t_L g2090 ( 
.A1(n_2044),
.A2(n_1977),
.B1(n_1956),
.B2(n_1884),
.Y(n_2090)
);

INVx1_ASAP7_75t_L g2091 ( 
.A(n_2039),
.Y(n_2091)
);

INVx1_ASAP7_75t_L g2092 ( 
.A(n_2055),
.Y(n_2092)
);

BUFx6f_ASAP7_75t_L g2093 ( 
.A(n_2048),
.Y(n_2093)
);

AOI21xp5_ASAP7_75t_L g2094 ( 
.A1(n_2036),
.A2(n_1962),
.B(n_1934),
.Y(n_2094)
);

AO21x2_ASAP7_75t_L g2095 ( 
.A1(n_2029),
.A2(n_1957),
.B(n_1955),
.Y(n_2095)
);

AND2x2_ASAP7_75t_L g2096 ( 
.A(n_2047),
.B(n_1908),
.Y(n_2096)
);

HB1xp67_ASAP7_75t_L g2097 ( 
.A(n_2041),
.Y(n_2097)
);

INVx1_ASAP7_75t_L g2098 ( 
.A(n_2068),
.Y(n_2098)
);

OAI21x1_ASAP7_75t_L g2099 ( 
.A1(n_2011),
.A2(n_1965),
.B(n_1903),
.Y(n_2099)
);

INVx2_ASAP7_75t_L g2100 ( 
.A(n_2053),
.Y(n_2100)
);

NAND2x1p5_ASAP7_75t_L g2101 ( 
.A(n_2012),
.B(n_1992),
.Y(n_2101)
);

INVx2_ASAP7_75t_L g2102 ( 
.A(n_2020),
.Y(n_2102)
);

AOI21x1_ASAP7_75t_L g2103 ( 
.A1(n_2026),
.A2(n_1962),
.B(n_1952),
.Y(n_2103)
);

OR2x2_ASAP7_75t_L g2104 ( 
.A(n_2009),
.B(n_1920),
.Y(n_2104)
);

OAI21xp5_ASAP7_75t_L g2105 ( 
.A1(n_2072),
.A2(n_1926),
.B(n_1890),
.Y(n_2105)
);

NAND2xp5_ASAP7_75t_L g2106 ( 
.A(n_2028),
.B(n_2033),
.Y(n_2106)
);

INVx1_ASAP7_75t_SL g2107 ( 
.A(n_2069),
.Y(n_2107)
);

OR2x2_ASAP7_75t_L g2108 ( 
.A(n_2067),
.B(n_1879),
.Y(n_2108)
);

INVx1_ASAP7_75t_L g2109 ( 
.A(n_2074),
.Y(n_2109)
);

AOI21xp5_ASAP7_75t_L g2110 ( 
.A1(n_2066),
.A2(n_2006),
.B(n_2015),
.Y(n_2110)
);

INVx1_ASAP7_75t_L g2111 ( 
.A(n_2078),
.Y(n_2111)
);

INVx2_ASAP7_75t_L g2112 ( 
.A(n_2018),
.Y(n_2112)
);

NOR2xp33_ASAP7_75t_L g2113 ( 
.A(n_2051),
.B(n_1946),
.Y(n_2113)
);

O2A1O1Ixp33_ASAP7_75t_L g2114 ( 
.A1(n_2005),
.A2(n_1989),
.B(n_1922),
.C(n_1939),
.Y(n_2114)
);

AO21x2_ASAP7_75t_L g2115 ( 
.A1(n_2058),
.A2(n_1970),
.B(n_1953),
.Y(n_2115)
);

INVx1_ASAP7_75t_L g2116 ( 
.A(n_2081),
.Y(n_2116)
);

INVx1_ASAP7_75t_L g2117 ( 
.A(n_2082),
.Y(n_2117)
);

AND2x2_ASAP7_75t_L g2118 ( 
.A(n_2043),
.B(n_1944),
.Y(n_2118)
);

OAI21x1_ASAP7_75t_L g2119 ( 
.A1(n_2063),
.A2(n_1967),
.B(n_1931),
.Y(n_2119)
);

AND2x4_ASAP7_75t_L g2120 ( 
.A(n_2059),
.B(n_1944),
.Y(n_2120)
);

AO21x2_ASAP7_75t_L g2121 ( 
.A1(n_2076),
.A2(n_1930),
.B(n_1967),
.Y(n_2121)
);

INVx1_ASAP7_75t_L g2122 ( 
.A(n_2062),
.Y(n_2122)
);

AOI21xp5_ASAP7_75t_L g2123 ( 
.A1(n_2035),
.A2(n_1979),
.B(n_1950),
.Y(n_2123)
);

INVx1_ASAP7_75t_SL g2124 ( 
.A(n_2022),
.Y(n_2124)
);

INVx2_ASAP7_75t_L g2125 ( 
.A(n_2052),
.Y(n_2125)
);

INVx2_ASAP7_75t_L g2126 ( 
.A(n_2052),
.Y(n_2126)
);

OA21x2_ASAP7_75t_L g2127 ( 
.A1(n_2056),
.A2(n_1976),
.B(n_1968),
.Y(n_2127)
);

OAI21x1_ASAP7_75t_L g2128 ( 
.A1(n_2040),
.A2(n_1949),
.B(n_1924),
.Y(n_2128)
);

AND2x2_ASAP7_75t_L g2129 ( 
.A(n_2079),
.B(n_1948),
.Y(n_2129)
);

AND2x4_ASAP7_75t_L g2130 ( 
.A(n_2059),
.B(n_733),
.Y(n_2130)
);

AOI22xp33_ASAP7_75t_L g2131 ( 
.A1(n_2070),
.A2(n_64),
.B1(n_62),
.B2(n_63),
.Y(n_2131)
);

INVx2_ASAP7_75t_L g2132 ( 
.A(n_2001),
.Y(n_2132)
);

NAND2xp5_ASAP7_75t_L g2133 ( 
.A(n_2077),
.B(n_64),
.Y(n_2133)
);

NAND2xp5_ASAP7_75t_SL g2134 ( 
.A(n_2086),
.B(n_2034),
.Y(n_2134)
);

INVx2_ASAP7_75t_SL g2135 ( 
.A(n_2093),
.Y(n_2135)
);

BUFx2_ASAP7_75t_L g2136 ( 
.A(n_2097),
.Y(n_2136)
);

INVx5_ASAP7_75t_L g2137 ( 
.A(n_2093),
.Y(n_2137)
);

INVx3_ASAP7_75t_L g2138 ( 
.A(n_2084),
.Y(n_2138)
);

AND2x2_ASAP7_75t_L g2139 ( 
.A(n_2118),
.B(n_2065),
.Y(n_2139)
);

OA21x2_ASAP7_75t_L g2140 ( 
.A1(n_2123),
.A2(n_2024),
.B(n_2057),
.Y(n_2140)
);

AOI21xp5_ASAP7_75t_L g2141 ( 
.A1(n_2094),
.A2(n_2064),
.B(n_2003),
.Y(n_2141)
);

AOI21xp5_ASAP7_75t_L g2142 ( 
.A1(n_2110),
.A2(n_2017),
.B(n_2004),
.Y(n_2142)
);

AOI22xp5_ASAP7_75t_L g2143 ( 
.A1(n_2083),
.A2(n_2071),
.B1(n_2010),
.B2(n_2000),
.Y(n_2143)
);

INVx2_ASAP7_75t_L g2144 ( 
.A(n_2100),
.Y(n_2144)
);

AO21x2_ASAP7_75t_L g2145 ( 
.A1(n_2099),
.A2(n_2027),
.B(n_2073),
.Y(n_2145)
);

AOI22xp5_ASAP7_75t_L g2146 ( 
.A1(n_2083),
.A2(n_2031),
.B1(n_2061),
.B2(n_2054),
.Y(n_2146)
);

OR2x2_ASAP7_75t_L g2147 ( 
.A(n_2087),
.B(n_2042),
.Y(n_2147)
);

INVx3_ASAP7_75t_L g2148 ( 
.A(n_2125),
.Y(n_2148)
);

NAND2x1p5_ASAP7_75t_L g2149 ( 
.A(n_2107),
.B(n_2128),
.Y(n_2149)
);

INVx2_ASAP7_75t_L g2150 ( 
.A(n_2112),
.Y(n_2150)
);

NAND2x1_ASAP7_75t_L g2151 ( 
.A(n_2091),
.B(n_2021),
.Y(n_2151)
);

INVx1_ASAP7_75t_L g2152 ( 
.A(n_2092),
.Y(n_2152)
);

AOI21x1_ASAP7_75t_L g2153 ( 
.A1(n_2103),
.A2(n_2032),
.B(n_2016),
.Y(n_2153)
);

INVx3_ASAP7_75t_L g2154 ( 
.A(n_2126),
.Y(n_2154)
);

INVx1_ASAP7_75t_L g2155 ( 
.A(n_2098),
.Y(n_2155)
);

BUFx12f_ASAP7_75t_L g2156 ( 
.A(n_2120),
.Y(n_2156)
);

HB1xp67_ASAP7_75t_L g2157 ( 
.A(n_2109),
.Y(n_2157)
);

AO21x2_ASAP7_75t_L g2158 ( 
.A1(n_2105),
.A2(n_2032),
.B(n_2042),
.Y(n_2158)
);

INVx2_ASAP7_75t_L g2159 ( 
.A(n_2111),
.Y(n_2159)
);

NAND2xp5_ASAP7_75t_L g2160 ( 
.A(n_2106),
.B(n_2019),
.Y(n_2160)
);

AOI22xp5_ASAP7_75t_L g2161 ( 
.A1(n_2090),
.A2(n_2075),
.B1(n_2014),
.B2(n_2002),
.Y(n_2161)
);

AO31x2_ASAP7_75t_L g2162 ( 
.A1(n_2116),
.A2(n_2016),
.A3(n_2050),
.B(n_2008),
.Y(n_2162)
);

NAND2xp5_ASAP7_75t_L g2163 ( 
.A(n_2132),
.B(n_2014),
.Y(n_2163)
);

AO21x2_ASAP7_75t_L g2164 ( 
.A1(n_2089),
.A2(n_2050),
.B(n_2045),
.Y(n_2164)
);

AND2x4_ASAP7_75t_L g2165 ( 
.A(n_2088),
.B(n_2048),
.Y(n_2165)
);

BUFx2_ASAP7_75t_L g2166 ( 
.A(n_2117),
.Y(n_2166)
);

INVx2_ASAP7_75t_L g2167 ( 
.A(n_2102),
.Y(n_2167)
);

OA21x2_ASAP7_75t_L g2168 ( 
.A1(n_2119),
.A2(n_65),
.B(n_66),
.Y(n_2168)
);

INVx2_ASAP7_75t_L g2169 ( 
.A(n_2108),
.Y(n_2169)
);

AND2x4_ASAP7_75t_L g2170 ( 
.A(n_2130),
.B(n_2025),
.Y(n_2170)
);

AOI21xp5_ASAP7_75t_L g2171 ( 
.A1(n_2095),
.A2(n_735),
.B(n_734),
.Y(n_2171)
);

BUFx2_ASAP7_75t_L g2172 ( 
.A(n_2101),
.Y(n_2172)
);

AOI21xp5_ASAP7_75t_L g2173 ( 
.A1(n_2085),
.A2(n_737),
.B(n_736),
.Y(n_2173)
);

OA21x2_ASAP7_75t_L g2174 ( 
.A1(n_2108),
.A2(n_65),
.B(n_66),
.Y(n_2174)
);

AOI21xp5_ASAP7_75t_L g2175 ( 
.A1(n_2114),
.A2(n_741),
.B(n_738),
.Y(n_2175)
);

BUFx3_ASAP7_75t_L g2176 ( 
.A(n_2113),
.Y(n_2176)
);

O2A1O1Ixp33_ASAP7_75t_L g2177 ( 
.A1(n_2133),
.A2(n_70),
.B(n_68),
.C(n_69),
.Y(n_2177)
);

AND2x2_ASAP7_75t_L g2178 ( 
.A(n_2122),
.B(n_68),
.Y(n_2178)
);

OAI21x1_ASAP7_75t_L g2179 ( 
.A1(n_2127),
.A2(n_745),
.B(n_742),
.Y(n_2179)
);

OA21x2_ASAP7_75t_L g2180 ( 
.A1(n_2131),
.A2(n_70),
.B(n_71),
.Y(n_2180)
);

NAND2xp5_ASAP7_75t_L g2181 ( 
.A(n_2104),
.B(n_2096),
.Y(n_2181)
);

INVx1_ASAP7_75t_L g2182 ( 
.A(n_2121),
.Y(n_2182)
);

AND2x2_ASAP7_75t_L g2183 ( 
.A(n_2124),
.B(n_72),
.Y(n_2183)
);

AO31x2_ASAP7_75t_L g2184 ( 
.A1(n_2115),
.A2(n_74),
.A3(n_72),
.B(n_73),
.Y(n_2184)
);

BUFx6f_ASAP7_75t_L g2185 ( 
.A(n_2129),
.Y(n_2185)
);

INVx2_ASAP7_75t_L g2186 ( 
.A(n_2100),
.Y(n_2186)
);

BUFx2_ASAP7_75t_L g2187 ( 
.A(n_2169),
.Y(n_2187)
);

INVx1_ASAP7_75t_L g2188 ( 
.A(n_2157),
.Y(n_2188)
);

INVx1_ASAP7_75t_L g2189 ( 
.A(n_2152),
.Y(n_2189)
);

NAND2xp5_ASAP7_75t_L g2190 ( 
.A(n_2136),
.B(n_73),
.Y(n_2190)
);

AND2x4_ASAP7_75t_L g2191 ( 
.A(n_2150),
.B(n_2166),
.Y(n_2191)
);

INVx2_ASAP7_75t_L g2192 ( 
.A(n_2159),
.Y(n_2192)
);

AND2x2_ASAP7_75t_L g2193 ( 
.A(n_2139),
.B(n_74),
.Y(n_2193)
);

INVx1_ASAP7_75t_L g2194 ( 
.A(n_2155),
.Y(n_2194)
);

HB1xp67_ASAP7_75t_L g2195 ( 
.A(n_2147),
.Y(n_2195)
);

HB1xp67_ASAP7_75t_L g2196 ( 
.A(n_2186),
.Y(n_2196)
);

INVx1_ASAP7_75t_L g2197 ( 
.A(n_2144),
.Y(n_2197)
);

INVx3_ASAP7_75t_L g2198 ( 
.A(n_2156),
.Y(n_2198)
);

INVx2_ASAP7_75t_SL g2199 ( 
.A(n_2137),
.Y(n_2199)
);

INVx1_ASAP7_75t_L g2200 ( 
.A(n_2167),
.Y(n_2200)
);

AND2x2_ASAP7_75t_L g2201 ( 
.A(n_2138),
.B(n_75),
.Y(n_2201)
);

BUFx2_ASAP7_75t_L g2202 ( 
.A(n_2172),
.Y(n_2202)
);

AND2x4_ASAP7_75t_L g2203 ( 
.A(n_2148),
.B(n_746),
.Y(n_2203)
);

INVx2_ASAP7_75t_SL g2204 ( 
.A(n_2137),
.Y(n_2204)
);

INVx2_ASAP7_75t_L g2205 ( 
.A(n_2182),
.Y(n_2205)
);

INVx1_ASAP7_75t_L g2206 ( 
.A(n_2162),
.Y(n_2206)
);

INVx1_ASAP7_75t_L g2207 ( 
.A(n_2162),
.Y(n_2207)
);

INVx1_ASAP7_75t_L g2208 ( 
.A(n_2184),
.Y(n_2208)
);

HB1xp67_ASAP7_75t_L g2209 ( 
.A(n_2149),
.Y(n_2209)
);

INVx1_ASAP7_75t_L g2210 ( 
.A(n_2184),
.Y(n_2210)
);

NAND2xp5_ASAP7_75t_L g2211 ( 
.A(n_2181),
.B(n_76),
.Y(n_2211)
);

INVx2_ASAP7_75t_L g2212 ( 
.A(n_2154),
.Y(n_2212)
);

INVx1_ASAP7_75t_L g2213 ( 
.A(n_2158),
.Y(n_2213)
);

NAND2xp5_ASAP7_75t_L g2214 ( 
.A(n_2134),
.B(n_77),
.Y(n_2214)
);

AO21x2_ASAP7_75t_L g2215 ( 
.A1(n_2142),
.A2(n_77),
.B(n_78),
.Y(n_2215)
);

INVxp67_ASAP7_75t_L g2216 ( 
.A(n_2163),
.Y(n_2216)
);

INVx1_ASAP7_75t_L g2217 ( 
.A(n_2151),
.Y(n_2217)
);

INVx1_ASAP7_75t_L g2218 ( 
.A(n_2153),
.Y(n_2218)
);

BUFx3_ASAP7_75t_L g2219 ( 
.A(n_2135),
.Y(n_2219)
);

AO21x2_ASAP7_75t_L g2220 ( 
.A1(n_2173),
.A2(n_78),
.B(n_79),
.Y(n_2220)
);

INVx1_ASAP7_75t_L g2221 ( 
.A(n_2174),
.Y(n_2221)
);

BUFx2_ASAP7_75t_L g2222 ( 
.A(n_2165),
.Y(n_2222)
);

AO21x2_ASAP7_75t_L g2223 ( 
.A1(n_2145),
.A2(n_2171),
.B(n_2175),
.Y(n_2223)
);

HB1xp67_ASAP7_75t_L g2224 ( 
.A(n_2164),
.Y(n_2224)
);

AND2x2_ASAP7_75t_L g2225 ( 
.A(n_2176),
.B(n_80),
.Y(n_2225)
);

HB1xp67_ASAP7_75t_L g2226 ( 
.A(n_2168),
.Y(n_2226)
);

AND2x2_ASAP7_75t_L g2227 ( 
.A(n_2160),
.B(n_80),
.Y(n_2227)
);

INVx4_ASAP7_75t_SL g2228 ( 
.A(n_2185),
.Y(n_2228)
);

INVx3_ASAP7_75t_L g2229 ( 
.A(n_2185),
.Y(n_2229)
);

AND2x2_ASAP7_75t_L g2230 ( 
.A(n_2183),
.B(n_81),
.Y(n_2230)
);

AND2x2_ASAP7_75t_L g2231 ( 
.A(n_2178),
.B(n_81),
.Y(n_2231)
);

HB1xp67_ASAP7_75t_L g2232 ( 
.A(n_2140),
.Y(n_2232)
);

INVx1_ASAP7_75t_L g2233 ( 
.A(n_2179),
.Y(n_2233)
);

INVx2_ASAP7_75t_L g2234 ( 
.A(n_2180),
.Y(n_2234)
);

INVx2_ASAP7_75t_L g2235 ( 
.A(n_2170),
.Y(n_2235)
);

INVx1_ASAP7_75t_L g2236 ( 
.A(n_2177),
.Y(n_2236)
);

OAI21x1_ASAP7_75t_L g2237 ( 
.A1(n_2141),
.A2(n_748),
.B(n_747),
.Y(n_2237)
);

AND2x2_ASAP7_75t_L g2238 ( 
.A(n_2161),
.B(n_82),
.Y(n_2238)
);

INVx2_ASAP7_75t_L g2239 ( 
.A(n_2146),
.Y(n_2239)
);

INVx1_ASAP7_75t_L g2240 ( 
.A(n_2143),
.Y(n_2240)
);

INVx2_ASAP7_75t_SL g2241 ( 
.A(n_2137),
.Y(n_2241)
);

AND2x2_ASAP7_75t_L g2242 ( 
.A(n_2136),
.B(n_82),
.Y(n_2242)
);

HB1xp67_ASAP7_75t_L g2243 ( 
.A(n_2169),
.Y(n_2243)
);

INVx1_ASAP7_75t_L g2244 ( 
.A(n_2157),
.Y(n_2244)
);

AND2x4_ASAP7_75t_L g2245 ( 
.A(n_2136),
.B(n_749),
.Y(n_2245)
);

OAI21x1_ASAP7_75t_L g2246 ( 
.A1(n_2142),
.A2(n_751),
.B(n_750),
.Y(n_2246)
);

AND2x2_ASAP7_75t_L g2247 ( 
.A(n_2136),
.B(n_83),
.Y(n_2247)
);

INVx1_ASAP7_75t_L g2248 ( 
.A(n_2157),
.Y(n_2248)
);

HB1xp67_ASAP7_75t_L g2249 ( 
.A(n_2169),
.Y(n_2249)
);

BUFx6f_ASAP7_75t_L g2250 ( 
.A(n_2137),
.Y(n_2250)
);

NAND2xp5_ASAP7_75t_L g2251 ( 
.A(n_2169),
.B(n_83),
.Y(n_2251)
);

INVx2_ASAP7_75t_L g2252 ( 
.A(n_2159),
.Y(n_2252)
);

INVx3_ASAP7_75t_L g2253 ( 
.A(n_2156),
.Y(n_2253)
);

BUFx3_ASAP7_75t_L g2254 ( 
.A(n_2135),
.Y(n_2254)
);

INVx3_ASAP7_75t_L g2255 ( 
.A(n_2156),
.Y(n_2255)
);

BUFx2_ASAP7_75t_L g2256 ( 
.A(n_2169),
.Y(n_2256)
);

INVx1_ASAP7_75t_L g2257 ( 
.A(n_2157),
.Y(n_2257)
);

AO31x2_ASAP7_75t_L g2258 ( 
.A1(n_2142),
.A2(n_86),
.A3(n_84),
.B(n_85),
.Y(n_2258)
);

HB1xp67_ASAP7_75t_L g2259 ( 
.A(n_2169),
.Y(n_2259)
);

INVx2_ASAP7_75t_L g2260 ( 
.A(n_2159),
.Y(n_2260)
);

BUFx2_ASAP7_75t_L g2261 ( 
.A(n_2169),
.Y(n_2261)
);

INVx1_ASAP7_75t_L g2262 ( 
.A(n_2157),
.Y(n_2262)
);

INVx1_ASAP7_75t_L g2263 ( 
.A(n_2189),
.Y(n_2263)
);

INVx2_ASAP7_75t_L g2264 ( 
.A(n_2187),
.Y(n_2264)
);

OAI221xp5_ASAP7_75t_L g2265 ( 
.A1(n_2236),
.A2(n_87),
.B1(n_85),
.B2(n_86),
.C(n_88),
.Y(n_2265)
);

OAI21xp33_ASAP7_75t_L g2266 ( 
.A1(n_2239),
.A2(n_87),
.B(n_88),
.Y(n_2266)
);

HB1xp67_ASAP7_75t_L g2267 ( 
.A(n_2195),
.Y(n_2267)
);

AOI22xp33_ASAP7_75t_L g2268 ( 
.A1(n_2240),
.A2(n_91),
.B1(n_89),
.B2(n_90),
.Y(n_2268)
);

AOI22xp33_ASAP7_75t_L g2269 ( 
.A1(n_2215),
.A2(n_92),
.B1(n_90),
.B2(n_91),
.Y(n_2269)
);

INVx2_ASAP7_75t_L g2270 ( 
.A(n_2187),
.Y(n_2270)
);

AOI21xp5_ASAP7_75t_L g2271 ( 
.A1(n_2223),
.A2(n_754),
.B(n_753),
.Y(n_2271)
);

OAI22xp33_ASAP7_75t_L g2272 ( 
.A1(n_2214),
.A2(n_94),
.B1(n_92),
.B2(n_93),
.Y(n_2272)
);

AOI221xp5_ASAP7_75t_L g2273 ( 
.A1(n_2232),
.A2(n_2221),
.B1(n_2226),
.B2(n_2234),
.C(n_2211),
.Y(n_2273)
);

OA21x2_ASAP7_75t_L g2274 ( 
.A1(n_2217),
.A2(n_93),
.B(n_94),
.Y(n_2274)
);

INVx1_ASAP7_75t_L g2275 ( 
.A(n_2194),
.Y(n_2275)
);

AOI22xp33_ASAP7_75t_L g2276 ( 
.A1(n_2238),
.A2(n_97),
.B1(n_95),
.B2(n_96),
.Y(n_2276)
);

INVx1_ASAP7_75t_L g2277 ( 
.A(n_2196),
.Y(n_2277)
);

AOI22xp33_ASAP7_75t_SL g2278 ( 
.A1(n_2220),
.A2(n_97),
.B1(n_98),
.B2(n_96),
.Y(n_2278)
);

INVx1_ASAP7_75t_L g2279 ( 
.A(n_2188),
.Y(n_2279)
);

AOI221xp5_ASAP7_75t_L g2280 ( 
.A1(n_2190),
.A2(n_100),
.B1(n_95),
.B2(n_99),
.C(n_101),
.Y(n_2280)
);

AOI22xp33_ASAP7_75t_SL g2281 ( 
.A1(n_2246),
.A2(n_101),
.B1(n_102),
.B2(n_100),
.Y(n_2281)
);

INVxp67_ASAP7_75t_L g2282 ( 
.A(n_2202),
.Y(n_2282)
);

AND2x2_ASAP7_75t_L g2283 ( 
.A(n_2256),
.B(n_99),
.Y(n_2283)
);

NAND4xp25_ASAP7_75t_L g2284 ( 
.A(n_2251),
.B(n_104),
.C(n_102),
.D(n_103),
.Y(n_2284)
);

INVx2_ASAP7_75t_L g2285 ( 
.A(n_2256),
.Y(n_2285)
);

INVx2_ASAP7_75t_L g2286 ( 
.A(n_2261),
.Y(n_2286)
);

OAI21x1_ASAP7_75t_L g2287 ( 
.A1(n_2213),
.A2(n_103),
.B(n_105),
.Y(n_2287)
);

AOI22xp5_ASAP7_75t_L g2288 ( 
.A1(n_2216),
.A2(n_107),
.B1(n_105),
.B2(n_106),
.Y(n_2288)
);

AND2x2_ASAP7_75t_L g2289 ( 
.A(n_2261),
.B(n_106),
.Y(n_2289)
);

OAI211xp5_ASAP7_75t_L g2290 ( 
.A1(n_2218),
.A2(n_109),
.B(n_107),
.C(n_108),
.Y(n_2290)
);

NAND2xp5_ASAP7_75t_L g2291 ( 
.A(n_2243),
.B(n_109),
.Y(n_2291)
);

AND2x4_ASAP7_75t_L g2292 ( 
.A(n_2191),
.B(n_110),
.Y(n_2292)
);

AOI22xp33_ASAP7_75t_SL g2293 ( 
.A1(n_2237),
.A2(n_112),
.B1(n_113),
.B2(n_111),
.Y(n_2293)
);

INVx5_ASAP7_75t_L g2294 ( 
.A(n_2250),
.Y(n_2294)
);

AOI22xp5_ASAP7_75t_L g2295 ( 
.A1(n_2222),
.A2(n_112),
.B1(n_110),
.B2(n_111),
.Y(n_2295)
);

INVx1_ASAP7_75t_L g2296 ( 
.A(n_2244),
.Y(n_2296)
);

OAI22xp33_ASAP7_75t_SL g2297 ( 
.A1(n_2209),
.A2(n_115),
.B1(n_113),
.B2(n_114),
.Y(n_2297)
);

AOI221xp5_ASAP7_75t_L g2298 ( 
.A1(n_2248),
.A2(n_118),
.B1(n_115),
.B2(n_117),
.C(n_119),
.Y(n_2298)
);

INVx1_ASAP7_75t_L g2299 ( 
.A(n_2257),
.Y(n_2299)
);

OAI221xp5_ASAP7_75t_L g2300 ( 
.A1(n_2235),
.A2(n_2229),
.B1(n_2199),
.B2(n_2241),
.C(n_2204),
.Y(n_2300)
);

OAI21x1_ASAP7_75t_L g2301 ( 
.A1(n_2206),
.A2(n_120),
.B(n_121),
.Y(n_2301)
);

AND2x4_ASAP7_75t_L g2302 ( 
.A(n_2212),
.B(n_120),
.Y(n_2302)
);

OAI22xp5_ASAP7_75t_L g2303 ( 
.A1(n_2250),
.A2(n_123),
.B1(n_121),
.B2(n_122),
.Y(n_2303)
);

AOI22xp33_ASAP7_75t_L g2304 ( 
.A1(n_2227),
.A2(n_124),
.B1(n_122),
.B2(n_123),
.Y(n_2304)
);

BUFx4f_ASAP7_75t_SL g2305 ( 
.A(n_2198),
.Y(n_2305)
);

OAI21x1_ASAP7_75t_L g2306 ( 
.A1(n_2207),
.A2(n_124),
.B(n_125),
.Y(n_2306)
);

AND2x2_ASAP7_75t_L g2307 ( 
.A(n_2249),
.B(n_125),
.Y(n_2307)
);

OAI211xp5_ASAP7_75t_L g2308 ( 
.A1(n_2242),
.A2(n_128),
.B(n_126),
.C(n_127),
.Y(n_2308)
);

OAI221xp5_ASAP7_75t_L g2309 ( 
.A1(n_2262),
.A2(n_128),
.B1(n_126),
.B2(n_127),
.C(n_129),
.Y(n_2309)
);

AOI22xp5_ASAP7_75t_L g2310 ( 
.A1(n_2233),
.A2(n_131),
.B1(n_129),
.B2(n_130),
.Y(n_2310)
);

CKINVDCx11_ASAP7_75t_R g2311 ( 
.A(n_2228),
.Y(n_2311)
);

OR2x6_ASAP7_75t_L g2312 ( 
.A(n_2245),
.B(n_130),
.Y(n_2312)
);

AOI22xp33_ASAP7_75t_L g2313 ( 
.A1(n_2230),
.A2(n_133),
.B1(n_131),
.B2(n_132),
.Y(n_2313)
);

OA21x2_ASAP7_75t_L g2314 ( 
.A1(n_2208),
.A2(n_132),
.B(n_133),
.Y(n_2314)
);

AOI21xp5_ASAP7_75t_L g2315 ( 
.A1(n_2210),
.A2(n_758),
.B(n_755),
.Y(n_2315)
);

INVx1_ASAP7_75t_L g2316 ( 
.A(n_2192),
.Y(n_2316)
);

INVx2_ASAP7_75t_L g2317 ( 
.A(n_2252),
.Y(n_2317)
);

AND2x2_ASAP7_75t_L g2318 ( 
.A(n_2259),
.B(n_134),
.Y(n_2318)
);

INVx2_ASAP7_75t_L g2319 ( 
.A(n_2260),
.Y(n_2319)
);

OAI22xp5_ASAP7_75t_L g2320 ( 
.A1(n_2219),
.A2(n_136),
.B1(n_134),
.B2(n_135),
.Y(n_2320)
);

INVx1_ASAP7_75t_L g2321 ( 
.A(n_2197),
.Y(n_2321)
);

OAI221xp5_ASAP7_75t_L g2322 ( 
.A1(n_2253),
.A2(n_138),
.B1(n_136),
.B2(n_137),
.C(n_139),
.Y(n_2322)
);

AOI221xp5_ASAP7_75t_L g2323 ( 
.A1(n_2247),
.A2(n_139),
.B1(n_137),
.B2(n_138),
.C(n_140),
.Y(n_2323)
);

AOI221xp5_ASAP7_75t_L g2324 ( 
.A1(n_2193),
.A2(n_142),
.B1(n_140),
.B2(n_141),
.C(n_143),
.Y(n_2324)
);

AOI221xp5_ASAP7_75t_L g2325 ( 
.A1(n_2231),
.A2(n_143),
.B1(n_141),
.B2(n_142),
.C(n_144),
.Y(n_2325)
);

AOI22xp33_ASAP7_75t_L g2326 ( 
.A1(n_2255),
.A2(n_146),
.B1(n_144),
.B2(n_145),
.Y(n_2326)
);

BUFx2_ASAP7_75t_L g2327 ( 
.A(n_2228),
.Y(n_2327)
);

OAI22xp5_ASAP7_75t_L g2328 ( 
.A1(n_2254),
.A2(n_147),
.B1(n_145),
.B2(n_146),
.Y(n_2328)
);

AOI222xp33_ASAP7_75t_L g2329 ( 
.A1(n_2225),
.A2(n_2201),
.B1(n_2200),
.B2(n_2203),
.C1(n_2258),
.C2(n_2224),
.Y(n_2329)
);

INVxp67_ASAP7_75t_L g2330 ( 
.A(n_2205),
.Y(n_2330)
);

HB1xp67_ASAP7_75t_L g2331 ( 
.A(n_2258),
.Y(n_2331)
);

INVx2_ASAP7_75t_L g2332 ( 
.A(n_2187),
.Y(n_2332)
);

NOR2xp33_ASAP7_75t_L g2333 ( 
.A(n_2216),
.B(n_147),
.Y(n_2333)
);

INVx2_ASAP7_75t_L g2334 ( 
.A(n_2187),
.Y(n_2334)
);

AOI22xp33_ASAP7_75t_SL g2335 ( 
.A1(n_2236),
.A2(n_150),
.B1(n_151),
.B2(n_149),
.Y(n_2335)
);

INVx2_ASAP7_75t_L g2336 ( 
.A(n_2187),
.Y(n_2336)
);

AOI221xp5_ASAP7_75t_L g2337 ( 
.A1(n_2236),
.A2(n_150),
.B1(n_148),
.B2(n_149),
.C(n_151),
.Y(n_2337)
);

NAND2xp5_ASAP7_75t_L g2338 ( 
.A(n_2243),
.B(n_152),
.Y(n_2338)
);

BUFx6f_ASAP7_75t_L g2339 ( 
.A(n_2250),
.Y(n_2339)
);

AOI22xp33_ASAP7_75t_L g2340 ( 
.A1(n_2239),
.A2(n_155),
.B1(n_153),
.B2(n_154),
.Y(n_2340)
);

OAI22xp33_ASAP7_75t_L g2341 ( 
.A1(n_2239),
.A2(n_157),
.B1(n_155),
.B2(n_156),
.Y(n_2341)
);

OAI33xp33_ASAP7_75t_L g2342 ( 
.A1(n_2236),
.A2(n_159),
.A3(n_161),
.B1(n_156),
.B2(n_157),
.B3(n_160),
.Y(n_2342)
);

OAI22xp33_ASAP7_75t_L g2343 ( 
.A1(n_2239),
.A2(n_162),
.B1(n_159),
.B2(n_160),
.Y(n_2343)
);

NAND2xp5_ASAP7_75t_L g2344 ( 
.A(n_2243),
.B(n_162),
.Y(n_2344)
);

OAI211xp5_ASAP7_75t_L g2345 ( 
.A1(n_2236),
.A2(n_165),
.B(n_163),
.C(n_164),
.Y(n_2345)
);

AOI221xp5_ASAP7_75t_L g2346 ( 
.A1(n_2236),
.A2(n_166),
.B1(n_164),
.B2(n_165),
.C(n_167),
.Y(n_2346)
);

AND2x2_ASAP7_75t_L g2347 ( 
.A(n_2202),
.B(n_166),
.Y(n_2347)
);

AND2x2_ASAP7_75t_L g2348 ( 
.A(n_2202),
.B(n_167),
.Y(n_2348)
);

AOI22xp5_ASAP7_75t_L g2349 ( 
.A1(n_2236),
.A2(n_170),
.B1(n_168),
.B2(n_169),
.Y(n_2349)
);

AOI22xp33_ASAP7_75t_L g2350 ( 
.A1(n_2239),
.A2(n_170),
.B1(n_168),
.B2(n_169),
.Y(n_2350)
);

AOI22xp33_ASAP7_75t_L g2351 ( 
.A1(n_2239),
.A2(n_173),
.B1(n_171),
.B2(n_172),
.Y(n_2351)
);

CKINVDCx20_ASAP7_75t_R g2352 ( 
.A(n_2222),
.Y(n_2352)
);

AOI22xp33_ASAP7_75t_L g2353 ( 
.A1(n_2239),
.A2(n_174),
.B1(n_172),
.B2(n_173),
.Y(n_2353)
);

NAND3xp33_ASAP7_75t_L g2354 ( 
.A(n_2236),
.B(n_174),
.C(n_175),
.Y(n_2354)
);

AOI22xp33_ASAP7_75t_L g2355 ( 
.A1(n_2239),
.A2(n_177),
.B1(n_175),
.B2(n_176),
.Y(n_2355)
);

NAND2x1_ASAP7_75t_L g2356 ( 
.A(n_2217),
.B(n_178),
.Y(n_2356)
);

INVx1_ASAP7_75t_L g2357 ( 
.A(n_2189),
.Y(n_2357)
);

HB1xp67_ASAP7_75t_L g2358 ( 
.A(n_2195),
.Y(n_2358)
);

AND2x2_ASAP7_75t_L g2359 ( 
.A(n_2202),
.B(n_178),
.Y(n_2359)
);

AOI22xp33_ASAP7_75t_L g2360 ( 
.A1(n_2239),
.A2(n_181),
.B1(n_179),
.B2(n_180),
.Y(n_2360)
);

OR2x2_ASAP7_75t_L g2361 ( 
.A(n_2277),
.B(n_179),
.Y(n_2361)
);

AND2x2_ASAP7_75t_L g2362 ( 
.A(n_2282),
.B(n_180),
.Y(n_2362)
);

INVx2_ASAP7_75t_L g2363 ( 
.A(n_2264),
.Y(n_2363)
);

NAND2xp5_ASAP7_75t_L g2364 ( 
.A(n_2273),
.B(n_182),
.Y(n_2364)
);

INVx2_ASAP7_75t_L g2365 ( 
.A(n_2270),
.Y(n_2365)
);

NOR2xp67_ASAP7_75t_SL g2366 ( 
.A(n_2294),
.B(n_183),
.Y(n_2366)
);

AOI22xp5_ASAP7_75t_L g2367 ( 
.A1(n_2337),
.A2(n_185),
.B1(n_183),
.B2(n_184),
.Y(n_2367)
);

INVx1_ASAP7_75t_L g2368 ( 
.A(n_2263),
.Y(n_2368)
);

INVxp67_ASAP7_75t_SL g2369 ( 
.A(n_2267),
.Y(n_2369)
);

AND2x2_ASAP7_75t_L g2370 ( 
.A(n_2285),
.B(n_184),
.Y(n_2370)
);

INVxp67_ASAP7_75t_SL g2371 ( 
.A(n_2358),
.Y(n_2371)
);

AND2x2_ASAP7_75t_L g2372 ( 
.A(n_2286),
.B(n_185),
.Y(n_2372)
);

INVx2_ASAP7_75t_L g2373 ( 
.A(n_2332),
.Y(n_2373)
);

AND2x2_ASAP7_75t_L g2374 ( 
.A(n_2334),
.B(n_2336),
.Y(n_2374)
);

NAND2xp5_ASAP7_75t_L g2375 ( 
.A(n_2279),
.B(n_186),
.Y(n_2375)
);

AND2x2_ASAP7_75t_L g2376 ( 
.A(n_2330),
.B(n_187),
.Y(n_2376)
);

OR2x2_ASAP7_75t_L g2377 ( 
.A(n_2296),
.B(n_187),
.Y(n_2377)
);

INVx1_ASAP7_75t_L g2378 ( 
.A(n_2275),
.Y(n_2378)
);

INVx1_ASAP7_75t_L g2379 ( 
.A(n_2357),
.Y(n_2379)
);

INVx1_ASAP7_75t_SL g2380 ( 
.A(n_2311),
.Y(n_2380)
);

NAND2xp5_ASAP7_75t_L g2381 ( 
.A(n_2299),
.B(n_188),
.Y(n_2381)
);

NOR2xp33_ASAP7_75t_L g2382 ( 
.A(n_2305),
.B(n_189),
.Y(n_2382)
);

INVx1_ASAP7_75t_L g2383 ( 
.A(n_2321),
.Y(n_2383)
);

OR2x2_ASAP7_75t_L g2384 ( 
.A(n_2316),
.B(n_189),
.Y(n_2384)
);

BUFx2_ASAP7_75t_L g2385 ( 
.A(n_2352),
.Y(n_2385)
);

INVx1_ASAP7_75t_L g2386 ( 
.A(n_2317),
.Y(n_2386)
);

NAND2xp5_ASAP7_75t_L g2387 ( 
.A(n_2329),
.B(n_190),
.Y(n_2387)
);

AND2x2_ASAP7_75t_L g2388 ( 
.A(n_2327),
.B(n_190),
.Y(n_2388)
);

INVx2_ASAP7_75t_L g2389 ( 
.A(n_2319),
.Y(n_2389)
);

INVx1_ASAP7_75t_L g2390 ( 
.A(n_2331),
.Y(n_2390)
);

INVx2_ASAP7_75t_L g2391 ( 
.A(n_2274),
.Y(n_2391)
);

INVx1_ASAP7_75t_L g2392 ( 
.A(n_2291),
.Y(n_2392)
);

INVx1_ASAP7_75t_L g2393 ( 
.A(n_2338),
.Y(n_2393)
);

INVx1_ASAP7_75t_L g2394 ( 
.A(n_2344),
.Y(n_2394)
);

INVxp67_ASAP7_75t_SL g2395 ( 
.A(n_2274),
.Y(n_2395)
);

INVx2_ASAP7_75t_L g2396 ( 
.A(n_2283),
.Y(n_2396)
);

AND2x2_ASAP7_75t_L g2397 ( 
.A(n_2289),
.B(n_2307),
.Y(n_2397)
);

INVxp67_ASAP7_75t_SL g2398 ( 
.A(n_2314),
.Y(n_2398)
);

AND2x2_ASAP7_75t_L g2399 ( 
.A(n_2318),
.B(n_191),
.Y(n_2399)
);

AND2x2_ASAP7_75t_L g2400 ( 
.A(n_2294),
.B(n_191),
.Y(n_2400)
);

INVx1_ASAP7_75t_L g2401 ( 
.A(n_2314),
.Y(n_2401)
);

INVx2_ASAP7_75t_L g2402 ( 
.A(n_2292),
.Y(n_2402)
);

OR2x2_ASAP7_75t_L g2403 ( 
.A(n_2300),
.B(n_192),
.Y(n_2403)
);

AND2x2_ASAP7_75t_L g2404 ( 
.A(n_2294),
.B(n_192),
.Y(n_2404)
);

AND2x4_ASAP7_75t_SL g2405 ( 
.A(n_2339),
.B(n_193),
.Y(n_2405)
);

AND2x2_ASAP7_75t_L g2406 ( 
.A(n_2347),
.B(n_193),
.Y(n_2406)
);

INVx1_ASAP7_75t_L g2407 ( 
.A(n_2287),
.Y(n_2407)
);

NAND2xp5_ASAP7_75t_L g2408 ( 
.A(n_2333),
.B(n_194),
.Y(n_2408)
);

NAND2xp5_ASAP7_75t_L g2409 ( 
.A(n_2348),
.B(n_2359),
.Y(n_2409)
);

NAND2xp5_ASAP7_75t_L g2410 ( 
.A(n_2302),
.B(n_194),
.Y(n_2410)
);

INVx1_ASAP7_75t_L g2411 ( 
.A(n_2301),
.Y(n_2411)
);

AND2x2_ASAP7_75t_L g2412 ( 
.A(n_2339),
.B(n_195),
.Y(n_2412)
);

NOR2xp33_ASAP7_75t_L g2413 ( 
.A(n_2284),
.B(n_195),
.Y(n_2413)
);

NAND2xp5_ASAP7_75t_L g2414 ( 
.A(n_2297),
.B(n_196),
.Y(n_2414)
);

INVx1_ASAP7_75t_L g2415 ( 
.A(n_2306),
.Y(n_2415)
);

NAND2xp5_ASAP7_75t_L g2416 ( 
.A(n_2272),
.B(n_196),
.Y(n_2416)
);

AND2x2_ASAP7_75t_L g2417 ( 
.A(n_2312),
.B(n_197),
.Y(n_2417)
);

INVx2_ASAP7_75t_L g2418 ( 
.A(n_2356),
.Y(n_2418)
);

INVx1_ASAP7_75t_L g2419 ( 
.A(n_2354),
.Y(n_2419)
);

INVx2_ASAP7_75t_L g2420 ( 
.A(n_2312),
.Y(n_2420)
);

AND2x2_ASAP7_75t_L g2421 ( 
.A(n_2295),
.B(n_197),
.Y(n_2421)
);

NAND2xp5_ASAP7_75t_L g2422 ( 
.A(n_2271),
.B(n_198),
.Y(n_2422)
);

INVx1_ASAP7_75t_L g2423 ( 
.A(n_2310),
.Y(n_2423)
);

AND2x4_ASAP7_75t_L g2424 ( 
.A(n_2288),
.B(n_198),
.Y(n_2424)
);

AOI22xp33_ASAP7_75t_L g2425 ( 
.A1(n_2346),
.A2(n_2265),
.B1(n_2342),
.B2(n_2266),
.Y(n_2425)
);

INVx1_ASAP7_75t_L g2426 ( 
.A(n_2290),
.Y(n_2426)
);

INVx2_ASAP7_75t_L g2427 ( 
.A(n_2309),
.Y(n_2427)
);

AOI22xp33_ASAP7_75t_L g2428 ( 
.A1(n_2280),
.A2(n_201),
.B1(n_199),
.B2(n_200),
.Y(n_2428)
);

INVx1_ASAP7_75t_L g2429 ( 
.A(n_2349),
.Y(n_2429)
);

AND2x2_ASAP7_75t_L g2430 ( 
.A(n_2276),
.B(n_201),
.Y(n_2430)
);

INVx2_ASAP7_75t_L g2431 ( 
.A(n_2322),
.Y(n_2431)
);

AND2x4_ASAP7_75t_L g2432 ( 
.A(n_2315),
.B(n_202),
.Y(n_2432)
);

INVx2_ASAP7_75t_L g2433 ( 
.A(n_2320),
.Y(n_2433)
);

OAI22xp5_ASAP7_75t_L g2434 ( 
.A1(n_2269),
.A2(n_205),
.B1(n_202),
.B2(n_204),
.Y(n_2434)
);

INVx1_ASAP7_75t_L g2435 ( 
.A(n_2345),
.Y(n_2435)
);

AOI22xp33_ASAP7_75t_L g2436 ( 
.A1(n_2278),
.A2(n_207),
.B1(n_204),
.B2(n_206),
.Y(n_2436)
);

AND2x2_ASAP7_75t_L g2437 ( 
.A(n_2293),
.B(n_206),
.Y(n_2437)
);

INVx1_ASAP7_75t_L g2438 ( 
.A(n_2308),
.Y(n_2438)
);

AND2x2_ASAP7_75t_L g2439 ( 
.A(n_2281),
.B(n_207),
.Y(n_2439)
);

INVx1_ASAP7_75t_L g2440 ( 
.A(n_2328),
.Y(n_2440)
);

INVx2_ASAP7_75t_L g2441 ( 
.A(n_2303),
.Y(n_2441)
);

INVx1_ASAP7_75t_L g2442 ( 
.A(n_2341),
.Y(n_2442)
);

NAND2xp5_ASAP7_75t_L g2443 ( 
.A(n_2323),
.B(n_208),
.Y(n_2443)
);

INVx1_ASAP7_75t_L g2444 ( 
.A(n_2343),
.Y(n_2444)
);

AND2x2_ASAP7_75t_L g2445 ( 
.A(n_2304),
.B(n_208),
.Y(n_2445)
);

NAND2xp5_ASAP7_75t_L g2446 ( 
.A(n_2324),
.B(n_209),
.Y(n_2446)
);

AOI222xp33_ASAP7_75t_L g2447 ( 
.A1(n_2325),
.A2(n_211),
.B1(n_213),
.B2(n_209),
.C1(n_210),
.C2(n_212),
.Y(n_2447)
);

INVx2_ASAP7_75t_L g2448 ( 
.A(n_2335),
.Y(n_2448)
);

INVx2_ASAP7_75t_L g2449 ( 
.A(n_2298),
.Y(n_2449)
);

AOI221xp5_ASAP7_75t_L g2450 ( 
.A1(n_2268),
.A2(n_212),
.B1(n_210),
.B2(n_211),
.C(n_214),
.Y(n_2450)
);

INVx1_ASAP7_75t_L g2451 ( 
.A(n_2313),
.Y(n_2451)
);

INVxp67_ASAP7_75t_L g2452 ( 
.A(n_2326),
.Y(n_2452)
);

NOR2xp67_ASAP7_75t_L g2453 ( 
.A(n_2340),
.B(n_215),
.Y(n_2453)
);

NOR2xp67_ASAP7_75t_L g2454 ( 
.A(n_2350),
.B(n_215),
.Y(n_2454)
);

BUFx3_ASAP7_75t_L g2455 ( 
.A(n_2351),
.Y(n_2455)
);

AND2x2_ASAP7_75t_L g2456 ( 
.A(n_2360),
.B(n_216),
.Y(n_2456)
);

OR2x2_ASAP7_75t_L g2457 ( 
.A(n_2353),
.B(n_216),
.Y(n_2457)
);

INVx3_ASAP7_75t_L g2458 ( 
.A(n_2355),
.Y(n_2458)
);

INVx2_ASAP7_75t_SL g2459 ( 
.A(n_2294),
.Y(n_2459)
);

AND2x2_ASAP7_75t_L g2460 ( 
.A(n_2282),
.B(n_217),
.Y(n_2460)
);

BUFx2_ASAP7_75t_L g2461 ( 
.A(n_2327),
.Y(n_2461)
);

INVx1_ASAP7_75t_L g2462 ( 
.A(n_2263),
.Y(n_2462)
);

INVx1_ASAP7_75t_L g2463 ( 
.A(n_2263),
.Y(n_2463)
);

INVx1_ASAP7_75t_L g2464 ( 
.A(n_2263),
.Y(n_2464)
);

INVx2_ASAP7_75t_L g2465 ( 
.A(n_2264),
.Y(n_2465)
);

NAND2xp5_ASAP7_75t_L g2466 ( 
.A(n_2273),
.B(n_217),
.Y(n_2466)
);

INVx2_ASAP7_75t_L g2467 ( 
.A(n_2264),
.Y(n_2467)
);

AND2x2_ASAP7_75t_L g2468 ( 
.A(n_2282),
.B(n_218),
.Y(n_2468)
);

AND2x2_ASAP7_75t_L g2469 ( 
.A(n_2282),
.B(n_219),
.Y(n_2469)
);

OR2x2_ASAP7_75t_L g2470 ( 
.A(n_2277),
.B(n_219),
.Y(n_2470)
);

INVx2_ASAP7_75t_L g2471 ( 
.A(n_2264),
.Y(n_2471)
);

INVx1_ASAP7_75t_L g2472 ( 
.A(n_2263),
.Y(n_2472)
);

AND2x2_ASAP7_75t_L g2473 ( 
.A(n_2282),
.B(n_220),
.Y(n_2473)
);

NAND2xp5_ASAP7_75t_L g2474 ( 
.A(n_2273),
.B(n_221),
.Y(n_2474)
);

AND2x2_ASAP7_75t_L g2475 ( 
.A(n_2282),
.B(n_221),
.Y(n_2475)
);

INVx2_ASAP7_75t_L g2476 ( 
.A(n_2264),
.Y(n_2476)
);

INVx2_ASAP7_75t_L g2477 ( 
.A(n_2264),
.Y(n_2477)
);

AND2x2_ASAP7_75t_L g2478 ( 
.A(n_2282),
.B(n_222),
.Y(n_2478)
);

INVx1_ASAP7_75t_L g2479 ( 
.A(n_2263),
.Y(n_2479)
);

INVx1_ASAP7_75t_L g2480 ( 
.A(n_2263),
.Y(n_2480)
);

INVx1_ASAP7_75t_L g2481 ( 
.A(n_2263),
.Y(n_2481)
);

BUFx2_ASAP7_75t_L g2482 ( 
.A(n_2327),
.Y(n_2482)
);

INVx1_ASAP7_75t_L g2483 ( 
.A(n_2263),
.Y(n_2483)
);

INVx1_ASAP7_75t_SL g2484 ( 
.A(n_2311),
.Y(n_2484)
);

INVx2_ASAP7_75t_L g2485 ( 
.A(n_2264),
.Y(n_2485)
);

INVx1_ASAP7_75t_L g2486 ( 
.A(n_2383),
.Y(n_2486)
);

AND2x2_ASAP7_75t_L g2487 ( 
.A(n_2461),
.B(n_223),
.Y(n_2487)
);

OR2x2_ASAP7_75t_L g2488 ( 
.A(n_2369),
.B(n_223),
.Y(n_2488)
);

AND2x2_ASAP7_75t_L g2489 ( 
.A(n_2461),
.B(n_224),
.Y(n_2489)
);

INVx2_ASAP7_75t_L g2490 ( 
.A(n_2482),
.Y(n_2490)
);

INVx1_ASAP7_75t_L g2491 ( 
.A(n_2368),
.Y(n_2491)
);

AND2x2_ASAP7_75t_L g2492 ( 
.A(n_2482),
.B(n_224),
.Y(n_2492)
);

NAND2xp5_ASAP7_75t_L g2493 ( 
.A(n_2419),
.B(n_225),
.Y(n_2493)
);

INVx1_ASAP7_75t_L g2494 ( 
.A(n_2378),
.Y(n_2494)
);

AND2x2_ASAP7_75t_L g2495 ( 
.A(n_2374),
.B(n_225),
.Y(n_2495)
);

INVxp67_ASAP7_75t_SL g2496 ( 
.A(n_2418),
.Y(n_2496)
);

NAND2xp5_ASAP7_75t_L g2497 ( 
.A(n_2407),
.B(n_226),
.Y(n_2497)
);

INVx2_ASAP7_75t_L g2498 ( 
.A(n_2459),
.Y(n_2498)
);

OAI21xp5_ASAP7_75t_SL g2499 ( 
.A1(n_2425),
.A2(n_226),
.B(n_227),
.Y(n_2499)
);

INVx1_ASAP7_75t_L g2500 ( 
.A(n_2379),
.Y(n_2500)
);

AND2x2_ASAP7_75t_L g2501 ( 
.A(n_2371),
.B(n_227),
.Y(n_2501)
);

INVx1_ASAP7_75t_L g2502 ( 
.A(n_2462),
.Y(n_2502)
);

INVx2_ASAP7_75t_L g2503 ( 
.A(n_2389),
.Y(n_2503)
);

INVx2_ASAP7_75t_L g2504 ( 
.A(n_2363),
.Y(n_2504)
);

AND2x4_ASAP7_75t_L g2505 ( 
.A(n_2420),
.B(n_228),
.Y(n_2505)
);

AND2x2_ASAP7_75t_L g2506 ( 
.A(n_2396),
.B(n_228),
.Y(n_2506)
);

INVx2_ASAP7_75t_L g2507 ( 
.A(n_2365),
.Y(n_2507)
);

OR2x2_ASAP7_75t_L g2508 ( 
.A(n_2392),
.B(n_229),
.Y(n_2508)
);

INVx1_ASAP7_75t_L g2509 ( 
.A(n_2463),
.Y(n_2509)
);

AND2x2_ASAP7_75t_L g2510 ( 
.A(n_2385),
.B(n_229),
.Y(n_2510)
);

AND2x4_ASAP7_75t_SL g2511 ( 
.A(n_2400),
.B(n_230),
.Y(n_2511)
);

INVx2_ASAP7_75t_L g2512 ( 
.A(n_2373),
.Y(n_2512)
);

AND2x4_ASAP7_75t_SL g2513 ( 
.A(n_2404),
.B(n_230),
.Y(n_2513)
);

OR2x2_ASAP7_75t_L g2514 ( 
.A(n_2393),
.B(n_231),
.Y(n_2514)
);

INVx1_ASAP7_75t_L g2515 ( 
.A(n_2464),
.Y(n_2515)
);

AND2x2_ASAP7_75t_L g2516 ( 
.A(n_2397),
.B(n_231),
.Y(n_2516)
);

AND2x2_ASAP7_75t_L g2517 ( 
.A(n_2394),
.B(n_232),
.Y(n_2517)
);

NAND2xp5_ASAP7_75t_L g2518 ( 
.A(n_2411),
.B(n_232),
.Y(n_2518)
);

INVx1_ASAP7_75t_L g2519 ( 
.A(n_2472),
.Y(n_2519)
);

INVx1_ASAP7_75t_L g2520 ( 
.A(n_2479),
.Y(n_2520)
);

INVx1_ASAP7_75t_L g2521 ( 
.A(n_2480),
.Y(n_2521)
);

AND2x4_ASAP7_75t_L g2522 ( 
.A(n_2402),
.B(n_233),
.Y(n_2522)
);

INVx2_ASAP7_75t_L g2523 ( 
.A(n_2465),
.Y(n_2523)
);

NOR2xp33_ASAP7_75t_L g2524 ( 
.A(n_2380),
.B(n_2484),
.Y(n_2524)
);

AND2x2_ASAP7_75t_L g2525 ( 
.A(n_2467),
.B(n_233),
.Y(n_2525)
);

BUFx3_ASAP7_75t_L g2526 ( 
.A(n_2388),
.Y(n_2526)
);

INVx1_ASAP7_75t_L g2527 ( 
.A(n_2481),
.Y(n_2527)
);

NAND2xp5_ASAP7_75t_L g2528 ( 
.A(n_2415),
.B(n_234),
.Y(n_2528)
);

NAND2xp5_ASAP7_75t_L g2529 ( 
.A(n_2387),
.B(n_235),
.Y(n_2529)
);

OA211x2_ASAP7_75t_L g2530 ( 
.A1(n_2364),
.A2(n_237),
.B(n_235),
.C(n_236),
.Y(n_2530)
);

INVx2_ASAP7_75t_L g2531 ( 
.A(n_2471),
.Y(n_2531)
);

AOI221xp5_ASAP7_75t_L g2532 ( 
.A1(n_2466),
.A2(n_238),
.B1(n_236),
.B2(n_237),
.C(n_239),
.Y(n_2532)
);

INVx2_ASAP7_75t_L g2533 ( 
.A(n_2476),
.Y(n_2533)
);

NAND2xp5_ASAP7_75t_L g2534 ( 
.A(n_2395),
.B(n_238),
.Y(n_2534)
);

HB1xp67_ASAP7_75t_L g2535 ( 
.A(n_2391),
.Y(n_2535)
);

NAND2xp5_ASAP7_75t_L g2536 ( 
.A(n_2423),
.B(n_239),
.Y(n_2536)
);

AND2x2_ASAP7_75t_L g2537 ( 
.A(n_2477),
.B(n_240),
.Y(n_2537)
);

NAND3xp33_ASAP7_75t_L g2538 ( 
.A(n_2474),
.B(n_240),
.C(n_241),
.Y(n_2538)
);

AND2x2_ASAP7_75t_L g2539 ( 
.A(n_2485),
.B(n_241),
.Y(n_2539)
);

HB1xp67_ASAP7_75t_L g2540 ( 
.A(n_2401),
.Y(n_2540)
);

OR2x2_ASAP7_75t_L g2541 ( 
.A(n_2398),
.B(n_242),
.Y(n_2541)
);

INVx1_ASAP7_75t_L g2542 ( 
.A(n_2483),
.Y(n_2542)
);

AND2x2_ASAP7_75t_L g2543 ( 
.A(n_2370),
.B(n_242),
.Y(n_2543)
);

INVx1_ASAP7_75t_L g2544 ( 
.A(n_2390),
.Y(n_2544)
);

INVx1_ASAP7_75t_L g2545 ( 
.A(n_2386),
.Y(n_2545)
);

NAND2xp5_ASAP7_75t_L g2546 ( 
.A(n_2376),
.B(n_243),
.Y(n_2546)
);

INVx1_ASAP7_75t_L g2547 ( 
.A(n_2384),
.Y(n_2547)
);

AND2x2_ASAP7_75t_L g2548 ( 
.A(n_2372),
.B(n_243),
.Y(n_2548)
);

AND2x2_ASAP7_75t_L g2549 ( 
.A(n_2409),
.B(n_244),
.Y(n_2549)
);

NAND3xp33_ASAP7_75t_L g2550 ( 
.A(n_2447),
.B(n_245),
.C(n_246),
.Y(n_2550)
);

AND2x2_ASAP7_75t_L g2551 ( 
.A(n_2362),
.B(n_245),
.Y(n_2551)
);

NAND2xp5_ASAP7_75t_L g2552 ( 
.A(n_2429),
.B(n_247),
.Y(n_2552)
);

INVx2_ASAP7_75t_L g2553 ( 
.A(n_2403),
.Y(n_2553)
);

AND2x2_ASAP7_75t_L g2554 ( 
.A(n_2460),
.B(n_247),
.Y(n_2554)
);

AOI22xp33_ASAP7_75t_L g2555 ( 
.A1(n_2427),
.A2(n_250),
.B1(n_248),
.B2(n_249),
.Y(n_2555)
);

AND2x2_ASAP7_75t_L g2556 ( 
.A(n_2468),
.B(n_248),
.Y(n_2556)
);

NAND2xp5_ASAP7_75t_L g2557 ( 
.A(n_2375),
.B(n_249),
.Y(n_2557)
);

OR2x2_ASAP7_75t_L g2558 ( 
.A(n_2361),
.B(n_250),
.Y(n_2558)
);

INVx1_ASAP7_75t_L g2559 ( 
.A(n_2377),
.Y(n_2559)
);

AND2x2_ASAP7_75t_L g2560 ( 
.A(n_2469),
.B(n_251),
.Y(n_2560)
);

NAND2xp5_ASAP7_75t_L g2561 ( 
.A(n_2381),
.B(n_251),
.Y(n_2561)
);

OR2x2_ASAP7_75t_L g2562 ( 
.A(n_2470),
.B(n_252),
.Y(n_2562)
);

AND2x2_ASAP7_75t_L g2563 ( 
.A(n_2473),
.B(n_252),
.Y(n_2563)
);

NOR2x1_ASAP7_75t_L g2564 ( 
.A(n_2475),
.B(n_253),
.Y(n_2564)
);

NAND2xp5_ASAP7_75t_L g2565 ( 
.A(n_2442),
.B(n_253),
.Y(n_2565)
);

INVx1_ASAP7_75t_L g2566 ( 
.A(n_2478),
.Y(n_2566)
);

INVx2_ASAP7_75t_SL g2567 ( 
.A(n_2412),
.Y(n_2567)
);

AND2x2_ASAP7_75t_L g2568 ( 
.A(n_2444),
.B(n_254),
.Y(n_2568)
);

NAND2xp5_ASAP7_75t_L g2569 ( 
.A(n_2440),
.B(n_254),
.Y(n_2569)
);

NAND2xp67_ASAP7_75t_L g2570 ( 
.A(n_2431),
.B(n_255),
.Y(n_2570)
);

AND2x2_ASAP7_75t_L g2571 ( 
.A(n_2441),
.B(n_255),
.Y(n_2571)
);

AND2x2_ASAP7_75t_L g2572 ( 
.A(n_2433),
.B(n_256),
.Y(n_2572)
);

INVx1_ASAP7_75t_L g2573 ( 
.A(n_2426),
.Y(n_2573)
);

NAND2x1p5_ASAP7_75t_L g2574 ( 
.A(n_2366),
.B(n_256),
.Y(n_2574)
);

AND2x2_ASAP7_75t_L g2575 ( 
.A(n_2399),
.B(n_2406),
.Y(n_2575)
);

INVx2_ASAP7_75t_L g2576 ( 
.A(n_2417),
.Y(n_2576)
);

BUFx2_ASAP7_75t_L g2577 ( 
.A(n_2438),
.Y(n_2577)
);

INVx1_ASAP7_75t_L g2578 ( 
.A(n_2451),
.Y(n_2578)
);

HB1xp67_ASAP7_75t_L g2579 ( 
.A(n_2435),
.Y(n_2579)
);

AND2x2_ASAP7_75t_L g2580 ( 
.A(n_2448),
.B(n_257),
.Y(n_2580)
);

NAND2xp5_ASAP7_75t_L g2581 ( 
.A(n_2458),
.B(n_257),
.Y(n_2581)
);

AND2x2_ASAP7_75t_L g2582 ( 
.A(n_2455),
.B(n_258),
.Y(n_2582)
);

OR2x2_ASAP7_75t_L g2583 ( 
.A(n_2408),
.B(n_2414),
.Y(n_2583)
);

AND2x2_ASAP7_75t_L g2584 ( 
.A(n_2452),
.B(n_259),
.Y(n_2584)
);

AND2x2_ASAP7_75t_L g2585 ( 
.A(n_2382),
.B(n_260),
.Y(n_2585)
);

AND2x2_ASAP7_75t_L g2586 ( 
.A(n_2410),
.B(n_2449),
.Y(n_2586)
);

NAND2xp5_ASAP7_75t_L g2587 ( 
.A(n_2422),
.B(n_260),
.Y(n_2587)
);

AND2x2_ASAP7_75t_L g2588 ( 
.A(n_2432),
.B(n_261),
.Y(n_2588)
);

AND2x2_ASAP7_75t_L g2589 ( 
.A(n_2424),
.B(n_262),
.Y(n_2589)
);

INVx2_ASAP7_75t_L g2590 ( 
.A(n_2405),
.Y(n_2590)
);

INVx2_ASAP7_75t_L g2591 ( 
.A(n_2421),
.Y(n_2591)
);

AOI221xp5_ASAP7_75t_L g2592 ( 
.A1(n_2413),
.A2(n_264),
.B1(n_262),
.B2(n_263),
.C(n_265),
.Y(n_2592)
);

AND2x2_ASAP7_75t_L g2593 ( 
.A(n_2437),
.B(n_264),
.Y(n_2593)
);

OR2x2_ASAP7_75t_L g2594 ( 
.A(n_2416),
.B(n_265),
.Y(n_2594)
);

INVx1_ASAP7_75t_L g2595 ( 
.A(n_2439),
.Y(n_2595)
);

INVx2_ASAP7_75t_L g2596 ( 
.A(n_2457),
.Y(n_2596)
);

AND2x2_ASAP7_75t_L g2597 ( 
.A(n_2430),
.B(n_266),
.Y(n_2597)
);

INVx1_ASAP7_75t_L g2598 ( 
.A(n_2446),
.Y(n_2598)
);

OR2x2_ASAP7_75t_L g2599 ( 
.A(n_2443),
.B(n_266),
.Y(n_2599)
);

AND2x2_ASAP7_75t_L g2600 ( 
.A(n_2445),
.B(n_267),
.Y(n_2600)
);

OR2x6_ASAP7_75t_L g2601 ( 
.A(n_2453),
.B(n_268),
.Y(n_2601)
);

INVxp67_ASAP7_75t_L g2602 ( 
.A(n_2456),
.Y(n_2602)
);

AND2x2_ASAP7_75t_L g2603 ( 
.A(n_2454),
.B(n_268),
.Y(n_2603)
);

AND2x2_ASAP7_75t_L g2604 ( 
.A(n_2367),
.B(n_2436),
.Y(n_2604)
);

INVx2_ASAP7_75t_L g2605 ( 
.A(n_2434),
.Y(n_2605)
);

AND2x4_ASAP7_75t_L g2606 ( 
.A(n_2428),
.B(n_269),
.Y(n_2606)
);

INVx2_ASAP7_75t_L g2607 ( 
.A(n_2450),
.Y(n_2607)
);

AND2x2_ASAP7_75t_L g2608 ( 
.A(n_2461),
.B(n_269),
.Y(n_2608)
);

AND2x2_ASAP7_75t_L g2609 ( 
.A(n_2461),
.B(n_270),
.Y(n_2609)
);

INVx2_ASAP7_75t_L g2610 ( 
.A(n_2461),
.Y(n_2610)
);

AND2x4_ASAP7_75t_L g2611 ( 
.A(n_2459),
.B(n_270),
.Y(n_2611)
);

AND2x2_ASAP7_75t_L g2612 ( 
.A(n_2461),
.B(n_272),
.Y(n_2612)
);

INVx3_ASAP7_75t_L g2613 ( 
.A(n_2459),
.Y(n_2613)
);

HB1xp67_ASAP7_75t_L g2614 ( 
.A(n_2461),
.Y(n_2614)
);

INVx1_ASAP7_75t_L g2615 ( 
.A(n_2383),
.Y(n_2615)
);

INVx3_ASAP7_75t_L g2616 ( 
.A(n_2459),
.Y(n_2616)
);

OAI221xp5_ASAP7_75t_L g2617 ( 
.A1(n_2387),
.A2(n_274),
.B1(n_272),
.B2(n_273),
.C(n_275),
.Y(n_2617)
);

NAND2xp5_ASAP7_75t_L g2618 ( 
.A(n_2419),
.B(n_273),
.Y(n_2618)
);

INVx1_ASAP7_75t_L g2619 ( 
.A(n_2383),
.Y(n_2619)
);

CKINVDCx16_ASAP7_75t_R g2620 ( 
.A(n_2385),
.Y(n_2620)
);

AND2x2_ASAP7_75t_L g2621 ( 
.A(n_2461),
.B(n_275),
.Y(n_2621)
);

INVx2_ASAP7_75t_L g2622 ( 
.A(n_2461),
.Y(n_2622)
);

HB1xp67_ASAP7_75t_L g2623 ( 
.A(n_2461),
.Y(n_2623)
);

OR2x2_ASAP7_75t_L g2624 ( 
.A(n_2369),
.B(n_276),
.Y(n_2624)
);

AND2x2_ASAP7_75t_L g2625 ( 
.A(n_2461),
.B(n_277),
.Y(n_2625)
);

AND2x2_ASAP7_75t_L g2626 ( 
.A(n_2461),
.B(n_277),
.Y(n_2626)
);

AND2x2_ASAP7_75t_L g2627 ( 
.A(n_2461),
.B(n_278),
.Y(n_2627)
);

BUFx2_ASAP7_75t_L g2628 ( 
.A(n_2461),
.Y(n_2628)
);

AND2x4_ASAP7_75t_L g2629 ( 
.A(n_2459),
.B(n_278),
.Y(n_2629)
);

INVx2_ASAP7_75t_L g2630 ( 
.A(n_2461),
.Y(n_2630)
);

HB1xp67_ASAP7_75t_L g2631 ( 
.A(n_2461),
.Y(n_2631)
);

INVx1_ASAP7_75t_L g2632 ( 
.A(n_2383),
.Y(n_2632)
);

OA21x2_ASAP7_75t_L g2633 ( 
.A1(n_2398),
.A2(n_279),
.B(n_280),
.Y(n_2633)
);

INVx1_ASAP7_75t_L g2634 ( 
.A(n_2383),
.Y(n_2634)
);

INVx3_ASAP7_75t_L g2635 ( 
.A(n_2459),
.Y(n_2635)
);

OR2x2_ASAP7_75t_L g2636 ( 
.A(n_2369),
.B(n_279),
.Y(n_2636)
);

AND2x2_ASAP7_75t_L g2637 ( 
.A(n_2461),
.B(n_280),
.Y(n_2637)
);

AND2x2_ASAP7_75t_L g2638 ( 
.A(n_2461),
.B(n_281),
.Y(n_2638)
);

NOR3xp33_ASAP7_75t_L g2639 ( 
.A(n_2387),
.B(n_282),
.C(n_283),
.Y(n_2639)
);

INVx1_ASAP7_75t_L g2640 ( 
.A(n_2383),
.Y(n_2640)
);

AND2x2_ASAP7_75t_L g2641 ( 
.A(n_2461),
.B(n_283),
.Y(n_2641)
);

AND2x2_ASAP7_75t_L g2642 ( 
.A(n_2461),
.B(n_284),
.Y(n_2642)
);

AND2x2_ASAP7_75t_L g2643 ( 
.A(n_2461),
.B(n_284),
.Y(n_2643)
);

AND2x2_ASAP7_75t_L g2644 ( 
.A(n_2461),
.B(n_285),
.Y(n_2644)
);

NAND2xp5_ASAP7_75t_L g2645 ( 
.A(n_2419),
.B(n_285),
.Y(n_2645)
);

NAND2xp5_ASAP7_75t_L g2646 ( 
.A(n_2419),
.B(n_286),
.Y(n_2646)
);

NAND2x1p5_ASAP7_75t_L g2647 ( 
.A(n_2385),
.B(n_287),
.Y(n_2647)
);

AND2x2_ASAP7_75t_L g2648 ( 
.A(n_2461),
.B(n_287),
.Y(n_2648)
);

HB1xp67_ASAP7_75t_L g2649 ( 
.A(n_2461),
.Y(n_2649)
);

OR2x2_ASAP7_75t_L g2650 ( 
.A(n_2369),
.B(n_288),
.Y(n_2650)
);

NAND2xp5_ASAP7_75t_L g2651 ( 
.A(n_2419),
.B(n_288),
.Y(n_2651)
);

NAND3xp33_ASAP7_75t_L g2652 ( 
.A(n_2364),
.B(n_290),
.C(n_291),
.Y(n_2652)
);

INVx1_ASAP7_75t_L g2653 ( 
.A(n_2383),
.Y(n_2653)
);

INVx1_ASAP7_75t_L g2654 ( 
.A(n_2383),
.Y(n_2654)
);

INVx1_ASAP7_75t_L g2655 ( 
.A(n_2383),
.Y(n_2655)
);

OAI221xp5_ASAP7_75t_SL g2656 ( 
.A1(n_2387),
.A2(n_292),
.B1(n_290),
.B2(n_291),
.C(n_293),
.Y(n_2656)
);

AOI22xp33_ASAP7_75t_L g2657 ( 
.A1(n_2607),
.A2(n_296),
.B1(n_292),
.B2(n_294),
.Y(n_2657)
);

OAI31xp33_ASAP7_75t_L g2658 ( 
.A1(n_2617),
.A2(n_298),
.A3(n_296),
.B(n_297),
.Y(n_2658)
);

INVx3_ASAP7_75t_L g2659 ( 
.A(n_2620),
.Y(n_2659)
);

NAND3xp33_ASAP7_75t_L g2660 ( 
.A(n_2550),
.B(n_297),
.C(n_298),
.Y(n_2660)
);

OAI221xp5_ASAP7_75t_L g2661 ( 
.A1(n_2499),
.A2(n_301),
.B1(n_299),
.B2(n_300),
.C(n_302),
.Y(n_2661)
);

INVx2_ASAP7_75t_L g2662 ( 
.A(n_2628),
.Y(n_2662)
);

AOI221xp5_ASAP7_75t_L g2663 ( 
.A1(n_2639),
.A2(n_301),
.B1(n_299),
.B2(n_300),
.C(n_302),
.Y(n_2663)
);

INVxp67_ASAP7_75t_SL g2664 ( 
.A(n_2614),
.Y(n_2664)
);

AOI22xp5_ASAP7_75t_L g2665 ( 
.A1(n_2577),
.A2(n_306),
.B1(n_303),
.B2(n_305),
.Y(n_2665)
);

AND2x2_ASAP7_75t_L g2666 ( 
.A(n_2613),
.B(n_303),
.Y(n_2666)
);

OAI22xp5_ASAP7_75t_L g2667 ( 
.A1(n_2577),
.A2(n_308),
.B1(n_306),
.B2(n_307),
.Y(n_2667)
);

AOI22xp33_ASAP7_75t_L g2668 ( 
.A1(n_2604),
.A2(n_310),
.B1(n_308),
.B2(n_309),
.Y(n_2668)
);

INVx3_ASAP7_75t_L g2669 ( 
.A(n_2616),
.Y(n_2669)
);

AOI22xp33_ASAP7_75t_L g2670 ( 
.A1(n_2605),
.A2(n_311),
.B1(n_309),
.B2(n_310),
.Y(n_2670)
);

AOI22xp5_ASAP7_75t_L g2671 ( 
.A1(n_2579),
.A2(n_313),
.B1(n_311),
.B2(n_312),
.Y(n_2671)
);

AOI22xp5_ASAP7_75t_L g2672 ( 
.A1(n_2578),
.A2(n_2553),
.B1(n_2532),
.B2(n_2598),
.Y(n_2672)
);

AOI221xp5_ASAP7_75t_L g2673 ( 
.A1(n_2656),
.A2(n_315),
.B1(n_312),
.B2(n_314),
.C(n_316),
.Y(n_2673)
);

INVx3_ASAP7_75t_L g2674 ( 
.A(n_2635),
.Y(n_2674)
);

NAND2xp5_ASAP7_75t_L g2675 ( 
.A(n_2586),
.B(n_314),
.Y(n_2675)
);

INVx1_ASAP7_75t_L g2676 ( 
.A(n_2623),
.Y(n_2676)
);

INVx1_ASAP7_75t_L g2677 ( 
.A(n_2631),
.Y(n_2677)
);

INVx1_ASAP7_75t_L g2678 ( 
.A(n_2649),
.Y(n_2678)
);

INVx1_ASAP7_75t_L g2679 ( 
.A(n_2540),
.Y(n_2679)
);

AND2x2_ASAP7_75t_L g2680 ( 
.A(n_2573),
.B(n_315),
.Y(n_2680)
);

OR2x2_ASAP7_75t_L g2681 ( 
.A(n_2591),
.B(n_317),
.Y(n_2681)
);

OAI22xp5_ASAP7_75t_SL g2682 ( 
.A1(n_2601),
.A2(n_319),
.B1(n_317),
.B2(n_318),
.Y(n_2682)
);

OR2x2_ASAP7_75t_L g2683 ( 
.A(n_2559),
.B(n_318),
.Y(n_2683)
);

INVx4_ASAP7_75t_L g2684 ( 
.A(n_2611),
.Y(n_2684)
);

OAI221xp5_ASAP7_75t_SL g2685 ( 
.A1(n_2592),
.A2(n_322),
.B1(n_320),
.B2(n_321),
.C(n_323),
.Y(n_2685)
);

AND2x4_ASAP7_75t_L g2686 ( 
.A(n_2498),
.B(n_320),
.Y(n_2686)
);

AND2x2_ASAP7_75t_L g2687 ( 
.A(n_2596),
.B(n_321),
.Y(n_2687)
);

HB1xp67_ASAP7_75t_L g2688 ( 
.A(n_2490),
.Y(n_2688)
);

INVx1_ASAP7_75t_L g2689 ( 
.A(n_2486),
.Y(n_2689)
);

INVx1_ASAP7_75t_L g2690 ( 
.A(n_2491),
.Y(n_2690)
);

AND2x2_ASAP7_75t_L g2691 ( 
.A(n_2576),
.B(n_322),
.Y(n_2691)
);

AOI33xp33_ASAP7_75t_L g2692 ( 
.A1(n_2555),
.A2(n_325),
.A3(n_327),
.B1(n_323),
.B2(n_324),
.B3(n_326),
.Y(n_2692)
);

NAND2xp5_ASAP7_75t_L g2693 ( 
.A(n_2547),
.B(n_324),
.Y(n_2693)
);

OA21x2_ASAP7_75t_L g2694 ( 
.A1(n_2496),
.A2(n_327),
.B(n_328),
.Y(n_2694)
);

INVx1_ASAP7_75t_L g2695 ( 
.A(n_2494),
.Y(n_2695)
);

AND2x2_ASAP7_75t_L g2696 ( 
.A(n_2610),
.B(n_328),
.Y(n_2696)
);

AND2x2_ASAP7_75t_L g2697 ( 
.A(n_2622),
.B(n_329),
.Y(n_2697)
);

HB1xp67_ASAP7_75t_L g2698 ( 
.A(n_2630),
.Y(n_2698)
);

AND2x2_ASAP7_75t_L g2699 ( 
.A(n_2567),
.B(n_329),
.Y(n_2699)
);

INVx1_ASAP7_75t_L g2700 ( 
.A(n_2500),
.Y(n_2700)
);

NAND2xp5_ASAP7_75t_L g2701 ( 
.A(n_2566),
.B(n_330),
.Y(n_2701)
);

OR2x2_ASAP7_75t_L g2702 ( 
.A(n_2504),
.B(n_330),
.Y(n_2702)
);

INVx1_ASAP7_75t_L g2703 ( 
.A(n_2502),
.Y(n_2703)
);

AOI211xp5_ASAP7_75t_L g2704 ( 
.A1(n_2538),
.A2(n_333),
.B(n_331),
.C(n_332),
.Y(n_2704)
);

AOI221xp5_ASAP7_75t_SL g2705 ( 
.A1(n_2534),
.A2(n_333),
.B1(n_331),
.B2(n_332),
.C(n_334),
.Y(n_2705)
);

INVx1_ASAP7_75t_L g2706 ( 
.A(n_2509),
.Y(n_2706)
);

AND2x2_ASAP7_75t_L g2707 ( 
.A(n_2595),
.B(n_334),
.Y(n_2707)
);

AND2x2_ASAP7_75t_L g2708 ( 
.A(n_2526),
.B(n_335),
.Y(n_2708)
);

OR2x2_ASAP7_75t_L g2709 ( 
.A(n_2507),
.B(n_2512),
.Y(n_2709)
);

AND2x4_ASAP7_75t_L g2710 ( 
.A(n_2590),
.B(n_335),
.Y(n_2710)
);

NAND2xp5_ASAP7_75t_L g2711 ( 
.A(n_2602),
.B(n_336),
.Y(n_2711)
);

INVx1_ASAP7_75t_L g2712 ( 
.A(n_2515),
.Y(n_2712)
);

BUFx2_ASAP7_75t_L g2713 ( 
.A(n_2487),
.Y(n_2713)
);

INVx1_ASAP7_75t_L g2714 ( 
.A(n_2519),
.Y(n_2714)
);

AND2x4_ASAP7_75t_L g2715 ( 
.A(n_2524),
.B(n_336),
.Y(n_2715)
);

AO21x2_ASAP7_75t_L g2716 ( 
.A1(n_2535),
.A2(n_337),
.B(n_338),
.Y(n_2716)
);

OR2x2_ASAP7_75t_L g2717 ( 
.A(n_2523),
.B(n_337),
.Y(n_2717)
);

INVx2_ASAP7_75t_L g2718 ( 
.A(n_2531),
.Y(n_2718)
);

AND2x4_ASAP7_75t_L g2719 ( 
.A(n_2575),
.B(n_338),
.Y(n_2719)
);

INVx3_ASAP7_75t_L g2720 ( 
.A(n_2629),
.Y(n_2720)
);

INVx1_ASAP7_75t_L g2721 ( 
.A(n_2520),
.Y(n_2721)
);

INVx2_ASAP7_75t_L g2722 ( 
.A(n_2533),
.Y(n_2722)
);

INVx1_ASAP7_75t_L g2723 ( 
.A(n_2521),
.Y(n_2723)
);

INVx2_ASAP7_75t_L g2724 ( 
.A(n_2503),
.Y(n_2724)
);

INVxp67_ASAP7_75t_L g2725 ( 
.A(n_2541),
.Y(n_2725)
);

INVx1_ASAP7_75t_L g2726 ( 
.A(n_2527),
.Y(n_2726)
);

INVx2_ASAP7_75t_L g2727 ( 
.A(n_2542),
.Y(n_2727)
);

BUFx3_ASAP7_75t_L g2728 ( 
.A(n_2505),
.Y(n_2728)
);

AOI22xp33_ASAP7_75t_L g2729 ( 
.A1(n_2606),
.A2(n_341),
.B1(n_339),
.B2(n_340),
.Y(n_2729)
);

INVx1_ASAP7_75t_L g2730 ( 
.A(n_2615),
.Y(n_2730)
);

AND2x4_ASAP7_75t_L g2731 ( 
.A(n_2489),
.B(n_340),
.Y(n_2731)
);

INVx1_ASAP7_75t_L g2732 ( 
.A(n_2619),
.Y(n_2732)
);

OR2x2_ASAP7_75t_L g2733 ( 
.A(n_2544),
.B(n_341),
.Y(n_2733)
);

INVx2_ASAP7_75t_L g2734 ( 
.A(n_2632),
.Y(n_2734)
);

INVx2_ASAP7_75t_L g2735 ( 
.A(n_2634),
.Y(n_2735)
);

INVx2_ASAP7_75t_L g2736 ( 
.A(n_2640),
.Y(n_2736)
);

NAND4xp25_ASAP7_75t_L g2737 ( 
.A(n_2530),
.B(n_345),
.C(n_346),
.D(n_344),
.Y(n_2737)
);

CKINVDCx5p33_ASAP7_75t_R g2738 ( 
.A(n_2601),
.Y(n_2738)
);

AND2x2_ASAP7_75t_L g2739 ( 
.A(n_2495),
.B(n_342),
.Y(n_2739)
);

AOI22xp33_ASAP7_75t_L g2740 ( 
.A1(n_2652),
.A2(n_345),
.B1(n_342),
.B2(n_344),
.Y(n_2740)
);

INVx2_ASAP7_75t_SL g2741 ( 
.A(n_2492),
.Y(n_2741)
);

BUFx3_ASAP7_75t_L g2742 ( 
.A(n_2511),
.Y(n_2742)
);

AOI222xp33_ASAP7_75t_SL g2743 ( 
.A1(n_2653),
.A2(n_2654),
.B1(n_2655),
.B2(n_2545),
.C1(n_2529),
.C2(n_2599),
.Y(n_2743)
);

INVx1_ASAP7_75t_L g2744 ( 
.A(n_2633),
.Y(n_2744)
);

INVx3_ASAP7_75t_L g2745 ( 
.A(n_2522),
.Y(n_2745)
);

INVx3_ASAP7_75t_L g2746 ( 
.A(n_2608),
.Y(n_2746)
);

AND2x4_ASAP7_75t_L g2747 ( 
.A(n_2609),
.B(n_348),
.Y(n_2747)
);

INVx1_ASAP7_75t_L g2748 ( 
.A(n_2633),
.Y(n_2748)
);

INVx2_ASAP7_75t_L g2749 ( 
.A(n_2525),
.Y(n_2749)
);

OR2x2_ASAP7_75t_L g2750 ( 
.A(n_2583),
.B(n_348),
.Y(n_2750)
);

BUFx3_ASAP7_75t_L g2751 ( 
.A(n_2513),
.Y(n_2751)
);

AND2x4_ASAP7_75t_L g2752 ( 
.A(n_2612),
.B(n_349),
.Y(n_2752)
);

OR2x2_ASAP7_75t_L g2753 ( 
.A(n_2488),
.B(n_349),
.Y(n_2753)
);

AND2x2_ASAP7_75t_L g2754 ( 
.A(n_2517),
.B(n_350),
.Y(n_2754)
);

INVx1_ASAP7_75t_SL g2755 ( 
.A(n_2621),
.Y(n_2755)
);

OAI31xp33_ASAP7_75t_L g2756 ( 
.A1(n_2574),
.A2(n_353),
.A3(n_351),
.B(n_352),
.Y(n_2756)
);

INVx3_ASAP7_75t_L g2757 ( 
.A(n_2625),
.Y(n_2757)
);

AOI33xp33_ASAP7_75t_L g2758 ( 
.A1(n_2582),
.A2(n_353),
.A3(n_355),
.B1(n_351),
.B2(n_352),
.B3(n_354),
.Y(n_2758)
);

INVx1_ASAP7_75t_L g2759 ( 
.A(n_2508),
.Y(n_2759)
);

AO221x2_ASAP7_75t_L g2760 ( 
.A1(n_2581),
.A2(n_356),
.B1(n_354),
.B2(n_355),
.C(n_357),
.Y(n_2760)
);

INVx1_ASAP7_75t_L g2761 ( 
.A(n_2514),
.Y(n_2761)
);

INVx1_ASAP7_75t_SL g2762 ( 
.A(n_2626),
.Y(n_2762)
);

OR2x2_ASAP7_75t_L g2763 ( 
.A(n_2624),
.B(n_356),
.Y(n_2763)
);

INVx2_ASAP7_75t_L g2764 ( 
.A(n_2537),
.Y(n_2764)
);

HB1xp67_ASAP7_75t_L g2765 ( 
.A(n_2627),
.Y(n_2765)
);

AND4x1_ASAP7_75t_L g2766 ( 
.A(n_2564),
.B(n_359),
.C(n_357),
.D(n_358),
.Y(n_2766)
);

AND2x4_ASAP7_75t_L g2767 ( 
.A(n_2637),
.B(n_358),
.Y(n_2767)
);

OR2x2_ASAP7_75t_L g2768 ( 
.A(n_2636),
.B(n_359),
.Y(n_2768)
);

INVx1_ASAP7_75t_L g2769 ( 
.A(n_2539),
.Y(n_2769)
);

AND2x4_ASAP7_75t_L g2770 ( 
.A(n_2638),
.B(n_360),
.Y(n_2770)
);

NAND2xp5_ASAP7_75t_L g2771 ( 
.A(n_2641),
.B(n_361),
.Y(n_2771)
);

AND2x4_ASAP7_75t_L g2772 ( 
.A(n_2642),
.B(n_362),
.Y(n_2772)
);

AND2x2_ASAP7_75t_L g2773 ( 
.A(n_2516),
.B(n_362),
.Y(n_2773)
);

AND2x2_ASAP7_75t_L g2774 ( 
.A(n_2568),
.B(n_363),
.Y(n_2774)
);

INVx1_ASAP7_75t_L g2775 ( 
.A(n_2650),
.Y(n_2775)
);

AOI221xp5_ASAP7_75t_L g2776 ( 
.A1(n_2497),
.A2(n_365),
.B1(n_363),
.B2(n_364),
.C(n_366),
.Y(n_2776)
);

OAI22xp5_ASAP7_75t_L g2777 ( 
.A1(n_2518),
.A2(n_368),
.B1(n_366),
.B2(n_367),
.Y(n_2777)
);

AOI31xp67_ASAP7_75t_L g2778 ( 
.A1(n_2528),
.A2(n_370),
.A3(n_367),
.B(n_369),
.Y(n_2778)
);

AOI21xp5_ASAP7_75t_L g2779 ( 
.A1(n_2587),
.A2(n_369),
.B(n_370),
.Y(n_2779)
);

AND2x2_ASAP7_75t_L g2780 ( 
.A(n_2659),
.B(n_2571),
.Y(n_2780)
);

INVx1_ASAP7_75t_L g2781 ( 
.A(n_2733),
.Y(n_2781)
);

NAND2xp5_ASAP7_75t_L g2782 ( 
.A(n_2713),
.B(n_2746),
.Y(n_2782)
);

INVx3_ASAP7_75t_L g2783 ( 
.A(n_2684),
.Y(n_2783)
);

INVx1_ASAP7_75t_L g2784 ( 
.A(n_2664),
.Y(n_2784)
);

INVx1_ASAP7_75t_L g2785 ( 
.A(n_2679),
.Y(n_2785)
);

OR2x2_ASAP7_75t_L g2786 ( 
.A(n_2765),
.B(n_2569),
.Y(n_2786)
);

INVx1_ASAP7_75t_L g2787 ( 
.A(n_2727),
.Y(n_2787)
);

HB1xp67_ASAP7_75t_L g2788 ( 
.A(n_2757),
.Y(n_2788)
);

AND2x2_ASAP7_75t_L g2789 ( 
.A(n_2669),
.B(n_2584),
.Y(n_2789)
);

NAND2xp5_ASAP7_75t_L g2790 ( 
.A(n_2755),
.B(n_2643),
.Y(n_2790)
);

OR2x2_ASAP7_75t_L g2791 ( 
.A(n_2762),
.B(n_2493),
.Y(n_2791)
);

AND2x2_ASAP7_75t_L g2792 ( 
.A(n_2674),
.B(n_2572),
.Y(n_2792)
);

AND2x2_ASAP7_75t_L g2793 ( 
.A(n_2741),
.B(n_2549),
.Y(n_2793)
);

INVx3_ASAP7_75t_L g2794 ( 
.A(n_2742),
.Y(n_2794)
);

INVx2_ASAP7_75t_L g2795 ( 
.A(n_2720),
.Y(n_2795)
);

HB1xp67_ASAP7_75t_L g2796 ( 
.A(n_2662),
.Y(n_2796)
);

NOR2x1_ASAP7_75t_L g2797 ( 
.A(n_2716),
.B(n_2644),
.Y(n_2797)
);

AND2x2_ASAP7_75t_L g2798 ( 
.A(n_2749),
.B(n_2648),
.Y(n_2798)
);

NAND2xp5_ASAP7_75t_L g2799 ( 
.A(n_2764),
.B(n_2769),
.Y(n_2799)
);

NAND2xp5_ASAP7_75t_SL g2800 ( 
.A(n_2738),
.B(n_2647),
.Y(n_2800)
);

AND2x2_ASAP7_75t_L g2801 ( 
.A(n_2775),
.B(n_2580),
.Y(n_2801)
);

NAND2xp5_ASAP7_75t_L g2802 ( 
.A(n_2725),
.B(n_2618),
.Y(n_2802)
);

AND2x2_ASAP7_75t_L g2803 ( 
.A(n_2759),
.B(n_2510),
.Y(n_2803)
);

INVx1_ASAP7_75t_L g2804 ( 
.A(n_2734),
.Y(n_2804)
);

OR2x2_ASAP7_75t_L g2805 ( 
.A(n_2761),
.B(n_2645),
.Y(n_2805)
);

INVx2_ASAP7_75t_L g2806 ( 
.A(n_2751),
.Y(n_2806)
);

AND2x2_ASAP7_75t_L g2807 ( 
.A(n_2745),
.B(n_2588),
.Y(n_2807)
);

AND2x2_ASAP7_75t_L g2808 ( 
.A(n_2728),
.B(n_2688),
.Y(n_2808)
);

INVx3_ASAP7_75t_L g2809 ( 
.A(n_2686),
.Y(n_2809)
);

AND2x2_ASAP7_75t_L g2810 ( 
.A(n_2698),
.B(n_2589),
.Y(n_2810)
);

AND2x2_ASAP7_75t_L g2811 ( 
.A(n_2676),
.B(n_2551),
.Y(n_2811)
);

INVx1_ASAP7_75t_L g2812 ( 
.A(n_2735),
.Y(n_2812)
);

AND2x2_ASAP7_75t_L g2813 ( 
.A(n_2677),
.B(n_2678),
.Y(n_2813)
);

INVx2_ASAP7_75t_L g2814 ( 
.A(n_2702),
.Y(n_2814)
);

NOR2xp33_ASAP7_75t_L g2815 ( 
.A(n_2750),
.B(n_2646),
.Y(n_2815)
);

AND2x4_ASAP7_75t_SL g2816 ( 
.A(n_2715),
.B(n_2501),
.Y(n_2816)
);

AND2x2_ASAP7_75t_L g2817 ( 
.A(n_2707),
.B(n_2554),
.Y(n_2817)
);

NAND2xp5_ASAP7_75t_L g2818 ( 
.A(n_2672),
.B(n_2651),
.Y(n_2818)
);

INVx1_ASAP7_75t_L g2819 ( 
.A(n_2736),
.Y(n_2819)
);

AND2x2_ASAP7_75t_L g2820 ( 
.A(n_2774),
.B(n_2687),
.Y(n_2820)
);

INVxp67_ASAP7_75t_L g2821 ( 
.A(n_2694),
.Y(n_2821)
);

INVx1_ASAP7_75t_L g2822 ( 
.A(n_2689),
.Y(n_2822)
);

INVx1_ASAP7_75t_L g2823 ( 
.A(n_2690),
.Y(n_2823)
);

AND2x2_ASAP7_75t_L g2824 ( 
.A(n_2680),
.B(n_2556),
.Y(n_2824)
);

INVxp67_ASAP7_75t_L g2825 ( 
.A(n_2743),
.Y(n_2825)
);

AND2x2_ASAP7_75t_L g2826 ( 
.A(n_2718),
.B(n_2560),
.Y(n_2826)
);

AND2x2_ASAP7_75t_L g2827 ( 
.A(n_2722),
.B(n_2563),
.Y(n_2827)
);

OR2x2_ASAP7_75t_L g2828 ( 
.A(n_2709),
.B(n_2536),
.Y(n_2828)
);

INVx1_ASAP7_75t_SL g2829 ( 
.A(n_2731),
.Y(n_2829)
);

INVx1_ASAP7_75t_L g2830 ( 
.A(n_2695),
.Y(n_2830)
);

INVx1_ASAP7_75t_L g2831 ( 
.A(n_2700),
.Y(n_2831)
);

INVx1_ASAP7_75t_L g2832 ( 
.A(n_2703),
.Y(n_2832)
);

INVx1_ASAP7_75t_L g2833 ( 
.A(n_2706),
.Y(n_2833)
);

AND2x2_ASAP7_75t_L g2834 ( 
.A(n_2724),
.B(n_2593),
.Y(n_2834)
);

AND2x2_ASAP7_75t_L g2835 ( 
.A(n_2696),
.B(n_2585),
.Y(n_2835)
);

AND2x4_ASAP7_75t_L g2836 ( 
.A(n_2666),
.B(n_2506),
.Y(n_2836)
);

NOR2x1_ASAP7_75t_L g2837 ( 
.A(n_2744),
.B(n_2594),
.Y(n_2837)
);

AND2x2_ASAP7_75t_L g2838 ( 
.A(n_2697),
.B(n_2597),
.Y(n_2838)
);

AND2x2_ASAP7_75t_L g2839 ( 
.A(n_2719),
.B(n_2754),
.Y(n_2839)
);

NOR2xp33_ASAP7_75t_L g2840 ( 
.A(n_2794),
.B(n_2693),
.Y(n_2840)
);

AND2x2_ASAP7_75t_L g2841 ( 
.A(n_2806),
.B(n_2710),
.Y(n_2841)
);

AND2x2_ASAP7_75t_L g2842 ( 
.A(n_2780),
.B(n_2699),
.Y(n_2842)
);

NAND2xp5_ASAP7_75t_L g2843 ( 
.A(n_2829),
.B(n_2779),
.Y(n_2843)
);

INVx2_ASAP7_75t_L g2844 ( 
.A(n_2783),
.Y(n_2844)
);

OR2x2_ASAP7_75t_L g2845 ( 
.A(n_2790),
.B(n_2748),
.Y(n_2845)
);

INVx1_ASAP7_75t_L g2846 ( 
.A(n_2784),
.Y(n_2846)
);

O2A1O1Ixp33_ASAP7_75t_L g2847 ( 
.A1(n_2825),
.A2(n_2661),
.B(n_2685),
.C(n_2667),
.Y(n_2847)
);

INVx2_ASAP7_75t_L g2848 ( 
.A(n_2808),
.Y(n_2848)
);

AND2x2_ASAP7_75t_L g2849 ( 
.A(n_2820),
.B(n_2708),
.Y(n_2849)
);

NOR2xp67_ASAP7_75t_L g2850 ( 
.A(n_2809),
.B(n_2733),
.Y(n_2850)
);

AND2x2_ASAP7_75t_L g2851 ( 
.A(n_2789),
.B(n_2739),
.Y(n_2851)
);

INVx2_ASAP7_75t_L g2852 ( 
.A(n_2839),
.Y(n_2852)
);

INVx2_ASAP7_75t_L g2853 ( 
.A(n_2816),
.Y(n_2853)
);

INVx1_ASAP7_75t_L g2854 ( 
.A(n_2781),
.Y(n_2854)
);

AND2x2_ASAP7_75t_L g2855 ( 
.A(n_2792),
.B(n_2747),
.Y(n_2855)
);

INVx1_ASAP7_75t_L g2856 ( 
.A(n_2781),
.Y(n_2856)
);

INVx1_ASAP7_75t_L g2857 ( 
.A(n_2788),
.Y(n_2857)
);

INVx1_ASAP7_75t_L g2858 ( 
.A(n_2796),
.Y(n_2858)
);

INVx2_ASAP7_75t_L g2859 ( 
.A(n_2807),
.Y(n_2859)
);

HB1xp67_ASAP7_75t_L g2860 ( 
.A(n_2810),
.Y(n_2860)
);

INVx1_ASAP7_75t_L g2861 ( 
.A(n_2799),
.Y(n_2861)
);

INVx1_ASAP7_75t_L g2862 ( 
.A(n_2814),
.Y(n_2862)
);

OR2x2_ASAP7_75t_L g2863 ( 
.A(n_2782),
.B(n_2681),
.Y(n_2863)
);

OR2x2_ASAP7_75t_L g2864 ( 
.A(n_2786),
.B(n_2675),
.Y(n_2864)
);

NAND2x1p5_ASAP7_75t_L g2865 ( 
.A(n_2797),
.B(n_2766),
.Y(n_2865)
);

INVx1_ASAP7_75t_L g2866 ( 
.A(n_2813),
.Y(n_2866)
);

INVx1_ASAP7_75t_L g2867 ( 
.A(n_2787),
.Y(n_2867)
);

NAND2xp5_ASAP7_75t_L g2868 ( 
.A(n_2835),
.B(n_2760),
.Y(n_2868)
);

INVx1_ASAP7_75t_L g2869 ( 
.A(n_2804),
.Y(n_2869)
);

NOR2xp33_ASAP7_75t_L g2870 ( 
.A(n_2800),
.B(n_2701),
.Y(n_2870)
);

INVx1_ASAP7_75t_L g2871 ( 
.A(n_2812),
.Y(n_2871)
);

INVx1_ASAP7_75t_L g2872 ( 
.A(n_2856),
.Y(n_2872)
);

INVx1_ASAP7_75t_L g2873 ( 
.A(n_2856),
.Y(n_2873)
);

AOI21xp5_ASAP7_75t_L g2874 ( 
.A1(n_2865),
.A2(n_2818),
.B(n_2847),
.Y(n_2874)
);

INVx2_ASAP7_75t_L g2875 ( 
.A(n_2841),
.Y(n_2875)
);

NAND2xp5_ASAP7_75t_L g2876 ( 
.A(n_2850),
.B(n_2803),
.Y(n_2876)
);

INVx1_ASAP7_75t_L g2877 ( 
.A(n_2860),
.Y(n_2877)
);

INVx1_ASAP7_75t_SL g2878 ( 
.A(n_2849),
.Y(n_2878)
);

INVx1_ASAP7_75t_L g2879 ( 
.A(n_2854),
.Y(n_2879)
);

INVx1_ASAP7_75t_L g2880 ( 
.A(n_2858),
.Y(n_2880)
);

XNOR2xp5_ASAP7_75t_L g2881 ( 
.A(n_2842),
.B(n_2836),
.Y(n_2881)
);

O2A1O1Ixp5_ASAP7_75t_L g2882 ( 
.A1(n_2844),
.A2(n_2785),
.B(n_2795),
.C(n_2819),
.Y(n_2882)
);

AOI22xp5_ASAP7_75t_L g2883 ( 
.A1(n_2870),
.A2(n_2821),
.B1(n_2673),
.B2(n_2837),
.Y(n_2883)
);

NOR2xp33_ASAP7_75t_L g2884 ( 
.A(n_2868),
.B(n_2838),
.Y(n_2884)
);

AOI21xp33_ASAP7_75t_SL g2885 ( 
.A1(n_2843),
.A2(n_2660),
.B(n_2791),
.Y(n_2885)
);

AND2x2_ASAP7_75t_L g2886 ( 
.A(n_2853),
.B(n_2798),
.Y(n_2886)
);

INVx1_ASAP7_75t_L g2887 ( 
.A(n_2857),
.Y(n_2887)
);

NAND2x1p5_ASAP7_75t_L g2888 ( 
.A(n_2848),
.B(n_2603),
.Y(n_2888)
);

OR2x2_ASAP7_75t_L g2889 ( 
.A(n_2866),
.B(n_2828),
.Y(n_2889)
);

INVx1_ASAP7_75t_L g2890 ( 
.A(n_2846),
.Y(n_2890)
);

NAND2xp5_ASAP7_75t_SL g2891 ( 
.A(n_2855),
.B(n_2836),
.Y(n_2891)
);

INVx1_ASAP7_75t_L g2892 ( 
.A(n_2877),
.Y(n_2892)
);

OAI22xp5_ASAP7_75t_L g2893 ( 
.A1(n_2883),
.A2(n_2874),
.B1(n_2878),
.B2(n_2881),
.Y(n_2893)
);

NAND2xp5_ASAP7_75t_L g2894 ( 
.A(n_2886),
.B(n_2851),
.Y(n_2894)
);

AND2x2_ASAP7_75t_SL g2895 ( 
.A(n_2876),
.B(n_2840),
.Y(n_2895)
);

NOR2xp33_ASAP7_75t_SL g2896 ( 
.A(n_2888),
.B(n_2756),
.Y(n_2896)
);

INVx1_ASAP7_75t_L g2897 ( 
.A(n_2872),
.Y(n_2897)
);

INVx1_ASAP7_75t_L g2898 ( 
.A(n_2873),
.Y(n_2898)
);

OAI22xp5_ASAP7_75t_L g2899 ( 
.A1(n_2884),
.A2(n_2665),
.B1(n_2671),
.B2(n_2863),
.Y(n_2899)
);

HB1xp67_ASAP7_75t_L g2900 ( 
.A(n_2891),
.Y(n_2900)
);

NAND2xp5_ASAP7_75t_L g2901 ( 
.A(n_2875),
.B(n_2852),
.Y(n_2901)
);

INVx1_ASAP7_75t_L g2902 ( 
.A(n_2901),
.Y(n_2902)
);

INVx2_ASAP7_75t_SL g2903 ( 
.A(n_2900),
.Y(n_2903)
);

NAND2xp5_ASAP7_75t_L g2904 ( 
.A(n_2895),
.B(n_2811),
.Y(n_2904)
);

INVx2_ASAP7_75t_L g2905 ( 
.A(n_2894),
.Y(n_2905)
);

INVx1_ASAP7_75t_L g2906 ( 
.A(n_2892),
.Y(n_2906)
);

OAI22xp33_ASAP7_75t_L g2907 ( 
.A1(n_2896),
.A2(n_2737),
.B1(n_2885),
.B2(n_2845),
.Y(n_2907)
);

INVx2_ASAP7_75t_L g2908 ( 
.A(n_2897),
.Y(n_2908)
);

OAI21xp5_ASAP7_75t_L g2909 ( 
.A1(n_2893),
.A2(n_2882),
.B(n_2859),
.Y(n_2909)
);

AOI322xp5_ASAP7_75t_L g2910 ( 
.A1(n_2898),
.A2(n_2887),
.A3(n_2880),
.B1(n_2705),
.B2(n_2861),
.C1(n_2890),
.C2(n_2879),
.Y(n_2910)
);

AOI21xp5_ASAP7_75t_L g2911 ( 
.A1(n_2907),
.A2(n_2899),
.B(n_2802),
.Y(n_2911)
);

OAI21xp33_ASAP7_75t_L g2912 ( 
.A1(n_2903),
.A2(n_2862),
.B(n_2889),
.Y(n_2912)
);

NAND3xp33_ASAP7_75t_SL g2913 ( 
.A(n_2909),
.B(n_2910),
.C(n_2904),
.Y(n_2913)
);

AOI221xp5_ASAP7_75t_L g2914 ( 
.A1(n_2906),
.A2(n_2871),
.B1(n_2869),
.B2(n_2867),
.C(n_2830),
.Y(n_2914)
);

AOI221xp5_ASAP7_75t_L g2915 ( 
.A1(n_2902),
.A2(n_2831),
.B1(n_2833),
.B2(n_2832),
.C(n_2823),
.Y(n_2915)
);

OA21x2_ASAP7_75t_L g2916 ( 
.A1(n_2908),
.A2(n_2822),
.B(n_2711),
.Y(n_2916)
);

NOR3xp33_ASAP7_75t_L g2917 ( 
.A(n_2905),
.B(n_2864),
.C(n_2815),
.Y(n_2917)
);

OAI221xp5_ASAP7_75t_L g2918 ( 
.A1(n_2909),
.A2(n_2658),
.B1(n_2663),
.B2(n_2704),
.C(n_2776),
.Y(n_2918)
);

INVx1_ASAP7_75t_L g2919 ( 
.A(n_2903),
.Y(n_2919)
);

NOR2xp33_ASAP7_75t_L g2920 ( 
.A(n_2907),
.B(n_2801),
.Y(n_2920)
);

OA22x2_ASAP7_75t_SL g2921 ( 
.A1(n_2902),
.A2(n_2714),
.B1(n_2721),
.B2(n_2712),
.Y(n_2921)
);

NAND2xp5_ASAP7_75t_L g2922 ( 
.A(n_2907),
.B(n_2793),
.Y(n_2922)
);

NAND4xp75_ASAP7_75t_L g2923 ( 
.A(n_2903),
.B(n_2691),
.C(n_2771),
.D(n_2565),
.Y(n_2923)
);

NAND2xp33_ASAP7_75t_SL g2924 ( 
.A(n_2903),
.B(n_2805),
.Y(n_2924)
);

AOI21xp5_ASAP7_75t_L g2925 ( 
.A1(n_2907),
.A2(n_2682),
.B(n_2552),
.Y(n_2925)
);

NAND2xp5_ASAP7_75t_L g2926 ( 
.A(n_2907),
.B(n_2824),
.Y(n_2926)
);

AOI322xp5_ASAP7_75t_L g2927 ( 
.A1(n_2907),
.A2(n_2668),
.A3(n_2670),
.B1(n_2657),
.B2(n_2729),
.C1(n_2740),
.C2(n_2600),
.Y(n_2927)
);

AOI222xp33_ASAP7_75t_L g2928 ( 
.A1(n_2907),
.A2(n_2777),
.B1(n_2557),
.B2(n_2561),
.C1(n_2834),
.C2(n_2827),
.Y(n_2928)
);

AOI22xp5_ASAP7_75t_L g2929 ( 
.A1(n_2913),
.A2(n_2826),
.B1(n_2817),
.B2(n_2723),
.Y(n_2929)
);

AOI21xp5_ASAP7_75t_L g2930 ( 
.A1(n_2924),
.A2(n_2683),
.B(n_2717),
.Y(n_2930)
);

NAND2xp5_ASAP7_75t_L g2931 ( 
.A(n_2919),
.B(n_2925),
.Y(n_2931)
);

INVx1_ASAP7_75t_SL g2932 ( 
.A(n_2916),
.Y(n_2932)
);

OAI31xp33_ASAP7_75t_L g2933 ( 
.A1(n_2918),
.A2(n_2753),
.A3(n_2768),
.B(n_2763),
.Y(n_2933)
);

AOI22xp5_ASAP7_75t_L g2934 ( 
.A1(n_2920),
.A2(n_2917),
.B1(n_2912),
.B2(n_2923),
.Y(n_2934)
);

AOI22xp5_ASAP7_75t_L g2935 ( 
.A1(n_2922),
.A2(n_2730),
.B1(n_2732),
.B2(n_2726),
.Y(n_2935)
);

AOI21xp33_ASAP7_75t_L g2936 ( 
.A1(n_2926),
.A2(n_2562),
.B(n_2558),
.Y(n_2936)
);

AOI221xp5_ASAP7_75t_L g2937 ( 
.A1(n_2911),
.A2(n_2767),
.B1(n_2772),
.B2(n_2770),
.C(n_2752),
.Y(n_2937)
);

OAI21xp5_ASAP7_75t_L g2938 ( 
.A1(n_2914),
.A2(n_2773),
.B(n_2546),
.Y(n_2938)
);

INVxp67_ASAP7_75t_L g2939 ( 
.A(n_2916),
.Y(n_2939)
);

AOI211x1_ASAP7_75t_SL g2940 ( 
.A1(n_2921),
.A2(n_2758),
.B(n_2778),
.C(n_2692),
.Y(n_2940)
);

OAI21xp33_ASAP7_75t_SL g2941 ( 
.A1(n_2928),
.A2(n_2548),
.B(n_2543),
.Y(n_2941)
);

NOR2xp33_ASAP7_75t_L g2942 ( 
.A(n_2915),
.B(n_2570),
.Y(n_2942)
);

AOI21xp5_ASAP7_75t_L g2943 ( 
.A1(n_2927),
.A2(n_371),
.B(n_372),
.Y(n_2943)
);

INVx1_ASAP7_75t_L g2944 ( 
.A(n_2919),
.Y(n_2944)
);

OR2x2_ASAP7_75t_L g2945 ( 
.A(n_2924),
.B(n_371),
.Y(n_2945)
);

AOI221xp5_ASAP7_75t_L g2946 ( 
.A1(n_2913),
.A2(n_374),
.B1(n_376),
.B2(n_373),
.C(n_375),
.Y(n_2946)
);

AOI221xp5_ASAP7_75t_L g2947 ( 
.A1(n_2913),
.A2(n_374),
.B1(n_377),
.B2(n_373),
.C(n_376),
.Y(n_2947)
);

OAI22xp5_ASAP7_75t_L g2948 ( 
.A1(n_2918),
.A2(n_378),
.B1(n_372),
.B2(n_377),
.Y(n_2948)
);

A2O1A1Ixp33_ASAP7_75t_SL g2949 ( 
.A1(n_2944),
.A2(n_380),
.B(n_378),
.C(n_379),
.Y(n_2949)
);

INVx1_ASAP7_75t_L g2950 ( 
.A(n_2945),
.Y(n_2950)
);

INVx1_ASAP7_75t_L g2951 ( 
.A(n_2931),
.Y(n_2951)
);

INVx1_ASAP7_75t_SL g2952 ( 
.A(n_2932),
.Y(n_2952)
);

AOI22xp33_ASAP7_75t_L g2953 ( 
.A1(n_2946),
.A2(n_382),
.B1(n_380),
.B2(n_381),
.Y(n_2953)
);

XOR2xp5_ASAP7_75t_L g2954 ( 
.A(n_2934),
.B(n_381),
.Y(n_2954)
);

INVx1_ASAP7_75t_L g2955 ( 
.A(n_2939),
.Y(n_2955)
);

INVx1_ASAP7_75t_SL g2956 ( 
.A(n_2930),
.Y(n_2956)
);

OAI21xp5_ASAP7_75t_SL g2957 ( 
.A1(n_2929),
.A2(n_382),
.B(n_383),
.Y(n_2957)
);

INVx2_ASAP7_75t_SL g2958 ( 
.A(n_2935),
.Y(n_2958)
);

INVx3_ASAP7_75t_L g2959 ( 
.A(n_2937),
.Y(n_2959)
);

AOI22xp5_ASAP7_75t_L g2960 ( 
.A1(n_2941),
.A2(n_385),
.B1(n_383),
.B2(n_384),
.Y(n_2960)
);

AOI22xp5_ASAP7_75t_L g2961 ( 
.A1(n_2942),
.A2(n_2947),
.B1(n_2948),
.B2(n_2943),
.Y(n_2961)
);

AOI221xp5_ASAP7_75t_L g2962 ( 
.A1(n_2936),
.A2(n_386),
.B1(n_384),
.B2(n_385),
.C(n_387),
.Y(n_2962)
);

AOI22xp5_ASAP7_75t_L g2963 ( 
.A1(n_2938),
.A2(n_388),
.B1(n_386),
.B2(n_387),
.Y(n_2963)
);

A2O1A1Ixp33_ASAP7_75t_L g2964 ( 
.A1(n_2933),
.A2(n_390),
.B(n_388),
.C(n_389),
.Y(n_2964)
);

OAI211xp5_ASAP7_75t_L g2965 ( 
.A1(n_2940),
.A2(n_397),
.B(n_405),
.C(n_389),
.Y(n_2965)
);

AOI222xp33_ASAP7_75t_L g2966 ( 
.A1(n_2939),
.A2(n_392),
.B1(n_394),
.B2(n_390),
.C1(n_391),
.C2(n_393),
.Y(n_2966)
);

O2A1O1Ixp33_ASAP7_75t_L g2967 ( 
.A1(n_2939),
.A2(n_394),
.B(n_391),
.C(n_393),
.Y(n_2967)
);

INVx1_ASAP7_75t_L g2968 ( 
.A(n_2945),
.Y(n_2968)
);

AOI21xp5_ASAP7_75t_L g2969 ( 
.A1(n_2932),
.A2(n_395),
.B(n_396),
.Y(n_2969)
);

NOR2x1_ASAP7_75t_L g2970 ( 
.A(n_2950),
.B(n_396),
.Y(n_2970)
);

INVx2_ASAP7_75t_L g2971 ( 
.A(n_2968),
.Y(n_2971)
);

NAND3xp33_ASAP7_75t_L g2972 ( 
.A(n_2964),
.B(n_397),
.C(n_398),
.Y(n_2972)
);

OAI321xp33_ASAP7_75t_L g2973 ( 
.A1(n_2961),
.A2(n_400),
.A3(n_402),
.B1(n_398),
.B2(n_399),
.C(n_401),
.Y(n_2973)
);

AOI321xp33_ASAP7_75t_L g2974 ( 
.A1(n_2951),
.A2(n_402),
.A3(n_404),
.B1(n_399),
.B2(n_400),
.C(n_403),
.Y(n_2974)
);

INVx1_ASAP7_75t_L g2975 ( 
.A(n_2955),
.Y(n_2975)
);

AOI211xp5_ASAP7_75t_L g2976 ( 
.A1(n_2965),
.A2(n_405),
.B(n_403),
.C(n_404),
.Y(n_2976)
);

AOI22xp5_ASAP7_75t_L g2977 ( 
.A1(n_2956),
.A2(n_408),
.B1(n_406),
.B2(n_407),
.Y(n_2977)
);

AOI22xp33_ASAP7_75t_L g2978 ( 
.A1(n_2959),
.A2(n_410),
.B1(n_406),
.B2(n_409),
.Y(n_2978)
);

NAND4xp25_ASAP7_75t_L g2979 ( 
.A(n_2960),
.B(n_411),
.C(n_409),
.D(n_410),
.Y(n_2979)
);

AOI211xp5_ASAP7_75t_SL g2980 ( 
.A1(n_2959),
.A2(n_413),
.B(n_411),
.C(n_412),
.Y(n_2980)
);

NAND2xp5_ASAP7_75t_L g2981 ( 
.A(n_2952),
.B(n_412),
.Y(n_2981)
);

OAI211xp5_ASAP7_75t_L g2982 ( 
.A1(n_2957),
.A2(n_2954),
.B(n_2969),
.C(n_2953),
.Y(n_2982)
);

OAI21xp5_ASAP7_75t_SL g2983 ( 
.A1(n_2963),
.A2(n_413),
.B(n_414),
.Y(n_2983)
);

AOI221xp5_ASAP7_75t_L g2984 ( 
.A1(n_2958),
.A2(n_416),
.B1(n_414),
.B2(n_415),
.C(n_417),
.Y(n_2984)
);

NAND2xp5_ASAP7_75t_L g2985 ( 
.A(n_2966),
.B(n_416),
.Y(n_2985)
);

XNOR2xp5_ASAP7_75t_L g2986 ( 
.A(n_2962),
.B(n_417),
.Y(n_2986)
);

XNOR2x1_ASAP7_75t_L g2987 ( 
.A(n_2949),
.B(n_418),
.Y(n_2987)
);

XOR2x2_ASAP7_75t_L g2988 ( 
.A(n_2967),
.B(n_418),
.Y(n_2988)
);

NAND3xp33_ASAP7_75t_SL g2989 ( 
.A(n_2956),
.B(n_419),
.C(n_420),
.Y(n_2989)
);

NAND2xp5_ASAP7_75t_L g2990 ( 
.A(n_2956),
.B(n_420),
.Y(n_2990)
);

NAND3xp33_ASAP7_75t_SL g2991 ( 
.A(n_2956),
.B(n_421),
.C(n_422),
.Y(n_2991)
);

INVx1_ASAP7_75t_L g2992 ( 
.A(n_2950),
.Y(n_2992)
);

AOI211xp5_ASAP7_75t_L g2993 ( 
.A1(n_2965),
.A2(n_425),
.B(n_421),
.C(n_423),
.Y(n_2993)
);

HB1xp67_ASAP7_75t_L g2994 ( 
.A(n_2956),
.Y(n_2994)
);

INVxp67_ASAP7_75t_L g2995 ( 
.A(n_2950),
.Y(n_2995)
);

NOR2x1_ASAP7_75t_SL g2996 ( 
.A(n_2950),
.B(n_425),
.Y(n_2996)
);

AOI22xp5_ASAP7_75t_L g2997 ( 
.A1(n_2956),
.A2(n_428),
.B1(n_426),
.B2(n_427),
.Y(n_2997)
);

AOI211xp5_ASAP7_75t_L g2998 ( 
.A1(n_2965),
.A2(n_429),
.B(n_427),
.C(n_428),
.Y(n_2998)
);

OAI22xp5_ASAP7_75t_L g2999 ( 
.A1(n_2956),
.A2(n_431),
.B1(n_429),
.B2(n_430),
.Y(n_2999)
);

NAND2xp5_ASAP7_75t_L g3000 ( 
.A(n_2956),
.B(n_431),
.Y(n_3000)
);

HB1xp67_ASAP7_75t_L g3001 ( 
.A(n_2956),
.Y(n_3001)
);

AOI31xp33_ASAP7_75t_L g3002 ( 
.A1(n_2956),
.A2(n_440),
.A3(n_448),
.B(n_432),
.Y(n_3002)
);

NOR2x1_ASAP7_75t_L g3003 ( 
.A(n_2950),
.B(n_432),
.Y(n_3003)
);

INVx1_ASAP7_75t_SL g3004 ( 
.A(n_2956),
.Y(n_3004)
);

INVx1_ASAP7_75t_SL g3005 ( 
.A(n_2956),
.Y(n_3005)
);

INVx1_ASAP7_75t_L g3006 ( 
.A(n_2950),
.Y(n_3006)
);

AOI221xp5_ASAP7_75t_L g3007 ( 
.A1(n_2965),
.A2(n_435),
.B1(n_433),
.B2(n_434),
.C(n_436),
.Y(n_3007)
);

XNOR2x1_ASAP7_75t_L g3008 ( 
.A(n_2954),
.B(n_433),
.Y(n_3008)
);

NAND3xp33_ASAP7_75t_L g3009 ( 
.A(n_2964),
.B(n_434),
.C(n_435),
.Y(n_3009)
);

INVx1_ASAP7_75t_L g3010 ( 
.A(n_2996),
.Y(n_3010)
);

INVx2_ASAP7_75t_L g3011 ( 
.A(n_2970),
.Y(n_3011)
);

NOR2xp33_ASAP7_75t_L g3012 ( 
.A(n_2979),
.B(n_437),
.Y(n_3012)
);

INVx2_ASAP7_75t_L g3013 ( 
.A(n_3003),
.Y(n_3013)
);

AND3x4_ASAP7_75t_L g3014 ( 
.A(n_2971),
.B(n_437),
.C(n_438),
.Y(n_3014)
);

INVx1_ASAP7_75t_L g3015 ( 
.A(n_3002),
.Y(n_3015)
);

NOR2x1_ASAP7_75t_L g3016 ( 
.A(n_2989),
.B(n_438),
.Y(n_3016)
);

NOR2x1_ASAP7_75t_L g3017 ( 
.A(n_2991),
.B(n_439),
.Y(n_3017)
);

NOR2x1_ASAP7_75t_L g3018 ( 
.A(n_2987),
.B(n_439),
.Y(n_3018)
);

NOR2x1_ASAP7_75t_L g3019 ( 
.A(n_3008),
.B(n_440),
.Y(n_3019)
);

OR2x2_ASAP7_75t_L g3020 ( 
.A(n_2981),
.B(n_441),
.Y(n_3020)
);

OA22x2_ASAP7_75t_L g3021 ( 
.A1(n_2983),
.A2(n_444),
.B1(n_442),
.B2(n_443),
.Y(n_3021)
);

INVx1_ASAP7_75t_L g3022 ( 
.A(n_2990),
.Y(n_3022)
);

AOI31xp33_ASAP7_75t_L g3023 ( 
.A1(n_2980),
.A2(n_2976),
.A3(n_2998),
.B(n_2993),
.Y(n_3023)
);

NAND2xp5_ASAP7_75t_L g3024 ( 
.A(n_3007),
.B(n_442),
.Y(n_3024)
);

AND2x4_ASAP7_75t_L g3025 ( 
.A(n_2992),
.B(n_3006),
.Y(n_3025)
);

INVx1_ASAP7_75t_L g3026 ( 
.A(n_3000),
.Y(n_3026)
);

NOR2x1_ASAP7_75t_L g3027 ( 
.A(n_2999),
.B(n_443),
.Y(n_3027)
);

INVx1_ASAP7_75t_L g3028 ( 
.A(n_2988),
.Y(n_3028)
);

INVx2_ASAP7_75t_L g3029 ( 
.A(n_2975),
.Y(n_3029)
);

INVxp67_ASAP7_75t_SL g3030 ( 
.A(n_2994),
.Y(n_3030)
);

INVx1_ASAP7_75t_SL g3031 ( 
.A(n_3004),
.Y(n_3031)
);

AO22x1_ASAP7_75t_L g3032 ( 
.A1(n_3001),
.A2(n_446),
.B1(n_444),
.B2(n_445),
.Y(n_3032)
);

OAI211xp5_ASAP7_75t_SL g3033 ( 
.A1(n_2995),
.A2(n_447),
.B(n_445),
.C(n_446),
.Y(n_3033)
);

NOR2xp33_ASAP7_75t_L g3034 ( 
.A(n_2982),
.B(n_447),
.Y(n_3034)
);

INVx1_ASAP7_75t_L g3035 ( 
.A(n_2986),
.Y(n_3035)
);

INVx1_ASAP7_75t_L g3036 ( 
.A(n_2977),
.Y(n_3036)
);

INVx1_ASAP7_75t_L g3037 ( 
.A(n_2997),
.Y(n_3037)
);

NAND2xp5_ASAP7_75t_L g3038 ( 
.A(n_2978),
.B(n_448),
.Y(n_3038)
);

OR2x2_ASAP7_75t_L g3039 ( 
.A(n_2985),
.B(n_450),
.Y(n_3039)
);

OR2x2_ASAP7_75t_L g3040 ( 
.A(n_3005),
.B(n_450),
.Y(n_3040)
);

AOI22xp5_ASAP7_75t_L g3041 ( 
.A1(n_2972),
.A2(n_453),
.B1(n_451),
.B2(n_452),
.Y(n_3041)
);

NAND2xp5_ASAP7_75t_SL g3042 ( 
.A(n_2973),
.B(n_451),
.Y(n_3042)
);

OAI22xp5_ASAP7_75t_SL g3043 ( 
.A1(n_3009),
.A2(n_454),
.B1(n_452),
.B2(n_453),
.Y(n_3043)
);

NOR2x1_ASAP7_75t_L g3044 ( 
.A(n_2974),
.B(n_454),
.Y(n_3044)
);

INVx1_ASAP7_75t_L g3045 ( 
.A(n_2984),
.Y(n_3045)
);

NOR2x1_ASAP7_75t_L g3046 ( 
.A(n_2989),
.B(n_455),
.Y(n_3046)
);

INVx2_ASAP7_75t_L g3047 ( 
.A(n_2996),
.Y(n_3047)
);

INVx2_ASAP7_75t_L g3048 ( 
.A(n_2996),
.Y(n_3048)
);

AOI22xp33_ASAP7_75t_L g3049 ( 
.A1(n_2971),
.A2(n_457),
.B1(n_455),
.B2(n_456),
.Y(n_3049)
);

NAND2xp5_ASAP7_75t_L g3050 ( 
.A(n_2980),
.B(n_457),
.Y(n_3050)
);

AND2x2_ASAP7_75t_L g3051 ( 
.A(n_2971),
.B(n_458),
.Y(n_3051)
);

NOR3xp33_ASAP7_75t_L g3052 ( 
.A(n_2995),
.B(n_459),
.C(n_460),
.Y(n_3052)
);

INVx2_ASAP7_75t_SL g3053 ( 
.A(n_2970),
.Y(n_3053)
);

INVx2_ASAP7_75t_SL g3054 ( 
.A(n_2970),
.Y(n_3054)
);

NOR2xp33_ASAP7_75t_L g3055 ( 
.A(n_3010),
.B(n_461),
.Y(n_3055)
);

INVx1_ASAP7_75t_L g3056 ( 
.A(n_3047),
.Y(n_3056)
);

NAND2xp5_ASAP7_75t_L g3057 ( 
.A(n_3032),
.B(n_461),
.Y(n_3057)
);

NAND2xp5_ASAP7_75t_L g3058 ( 
.A(n_3053),
.B(n_462),
.Y(n_3058)
);

HB1xp67_ASAP7_75t_L g3059 ( 
.A(n_3048),
.Y(n_3059)
);

INVxp67_ASAP7_75t_L g3060 ( 
.A(n_3016),
.Y(n_3060)
);

INVx1_ASAP7_75t_L g3061 ( 
.A(n_3051),
.Y(n_3061)
);

HB1xp67_ASAP7_75t_L g3062 ( 
.A(n_3054),
.Y(n_3062)
);

XOR2x1_ASAP7_75t_L g3063 ( 
.A(n_3011),
.B(n_462),
.Y(n_3063)
);

XNOR2xp5_ASAP7_75t_L g3064 ( 
.A(n_3014),
.B(n_463),
.Y(n_3064)
);

XOR2xp5_ASAP7_75t_L g3065 ( 
.A(n_3044),
.B(n_463),
.Y(n_3065)
);

INVx1_ASAP7_75t_L g3066 ( 
.A(n_3021),
.Y(n_3066)
);

AND2x2_ASAP7_75t_L g3067 ( 
.A(n_3018),
.B(n_464),
.Y(n_3067)
);

INVx1_ASAP7_75t_L g3068 ( 
.A(n_3050),
.Y(n_3068)
);

NOR2x1_ASAP7_75t_L g3069 ( 
.A(n_3013),
.B(n_464),
.Y(n_3069)
);

NAND2x1p5_ASAP7_75t_L g3070 ( 
.A(n_3019),
.B(n_465),
.Y(n_3070)
);

NAND2x1p5_ASAP7_75t_L g3071 ( 
.A(n_3025),
.B(n_465),
.Y(n_3071)
);

OAI21x1_ASAP7_75t_SL g3072 ( 
.A1(n_3017),
.A2(n_466),
.B(n_467),
.Y(n_3072)
);

AOI22xp5_ASAP7_75t_L g3073 ( 
.A1(n_3031),
.A2(n_468),
.B1(n_466),
.B2(n_467),
.Y(n_3073)
);

NOR2x1_ASAP7_75t_L g3074 ( 
.A(n_3015),
.B(n_469),
.Y(n_3074)
);

NAND2x1p5_ASAP7_75t_L g3075 ( 
.A(n_3046),
.B(n_3027),
.Y(n_3075)
);

NOR3xp33_ASAP7_75t_L g3076 ( 
.A(n_3034),
.B(n_477),
.C(n_469),
.Y(n_3076)
);

NOR2x1p5_ASAP7_75t_L g3077 ( 
.A(n_3030),
.B(n_470),
.Y(n_3077)
);

INVx1_ASAP7_75t_L g3078 ( 
.A(n_3040),
.Y(n_3078)
);

NOR2x1_ASAP7_75t_L g3079 ( 
.A(n_3033),
.B(n_470),
.Y(n_3079)
);

NAND2xp5_ASAP7_75t_L g3080 ( 
.A(n_3052),
.B(n_471),
.Y(n_3080)
);

INVx1_ASAP7_75t_L g3081 ( 
.A(n_3043),
.Y(n_3081)
);

INVx1_ASAP7_75t_L g3082 ( 
.A(n_3020),
.Y(n_3082)
);

INVxp67_ASAP7_75t_SL g3083 ( 
.A(n_3042),
.Y(n_3083)
);

AOI22xp33_ASAP7_75t_SL g3084 ( 
.A1(n_3029),
.A2(n_474),
.B1(n_472),
.B2(n_473),
.Y(n_3084)
);

AND2x4_ASAP7_75t_L g3085 ( 
.A(n_3022),
.B(n_473),
.Y(n_3085)
);

NAND4xp75_ASAP7_75t_L g3086 ( 
.A(n_3028),
.B(n_476),
.C(n_474),
.D(n_475),
.Y(n_3086)
);

NOR2x1_ASAP7_75t_L g3087 ( 
.A(n_3039),
.B(n_476),
.Y(n_3087)
);

AND2x2_ASAP7_75t_SL g3088 ( 
.A(n_3012),
.B(n_477),
.Y(n_3088)
);

INVx1_ASAP7_75t_L g3089 ( 
.A(n_3024),
.Y(n_3089)
);

NOR2x1p5_ASAP7_75t_L g3090 ( 
.A(n_3038),
.B(n_478),
.Y(n_3090)
);

XNOR2x1_ASAP7_75t_L g3091 ( 
.A(n_3036),
.B(n_479),
.Y(n_3091)
);

INVx2_ASAP7_75t_L g3092 ( 
.A(n_3026),
.Y(n_3092)
);

OR2x2_ASAP7_75t_L g3093 ( 
.A(n_3037),
.B(n_480),
.Y(n_3093)
);

AOI211x1_ASAP7_75t_L g3094 ( 
.A1(n_3023),
.A2(n_482),
.B(n_480),
.C(n_481),
.Y(n_3094)
);

INVxp67_ASAP7_75t_SL g3095 ( 
.A(n_3041),
.Y(n_3095)
);

NOR2xp67_ASAP7_75t_L g3096 ( 
.A(n_3045),
.B(n_3035),
.Y(n_3096)
);

NOR2x1_ASAP7_75t_L g3097 ( 
.A(n_3049),
.B(n_481),
.Y(n_3097)
);

NAND2xp5_ASAP7_75t_SL g3098 ( 
.A(n_3047),
.B(n_482),
.Y(n_3098)
);

NAND4xp75_ASAP7_75t_L g3099 ( 
.A(n_3018),
.B(n_485),
.C(n_483),
.D(n_484),
.Y(n_3099)
);

AND2x4_ASAP7_75t_L g3100 ( 
.A(n_3047),
.B(n_484),
.Y(n_3100)
);

INVx1_ASAP7_75t_L g3101 ( 
.A(n_3010),
.Y(n_3101)
);

AND2x4_ASAP7_75t_L g3102 ( 
.A(n_3047),
.B(n_485),
.Y(n_3102)
);

INVx2_ASAP7_75t_SL g3103 ( 
.A(n_3047),
.Y(n_3103)
);

NAND4xp75_ASAP7_75t_L g3104 ( 
.A(n_3018),
.B(n_488),
.C(n_486),
.D(n_487),
.Y(n_3104)
);

OR2x2_ASAP7_75t_L g3105 ( 
.A(n_3047),
.B(n_486),
.Y(n_3105)
);

NOR2xp67_ASAP7_75t_L g3106 ( 
.A(n_3053),
.B(n_489),
.Y(n_3106)
);

INVx2_ASAP7_75t_L g3107 ( 
.A(n_3047),
.Y(n_3107)
);

AOI22xp5_ASAP7_75t_L g3108 ( 
.A1(n_3031),
.A2(n_491),
.B1(n_487),
.B2(n_489),
.Y(n_3108)
);

INVx1_ASAP7_75t_L g3109 ( 
.A(n_3010),
.Y(n_3109)
);

NAND2xp5_ASAP7_75t_L g3110 ( 
.A(n_3032),
.B(n_491),
.Y(n_3110)
);

INVx2_ASAP7_75t_L g3111 ( 
.A(n_3047),
.Y(n_3111)
);

AOI22xp5_ASAP7_75t_L g3112 ( 
.A1(n_3103),
.A2(n_3056),
.B1(n_3109),
.B2(n_3101),
.Y(n_3112)
);

NAND2xp5_ASAP7_75t_SL g3113 ( 
.A(n_3106),
.B(n_492),
.Y(n_3113)
);

NAND4xp25_ASAP7_75t_L g3114 ( 
.A(n_3096),
.B(n_495),
.C(n_493),
.D(n_494),
.Y(n_3114)
);

AOI211xp5_ASAP7_75t_L g3115 ( 
.A1(n_3059),
.A2(n_495),
.B(n_493),
.C(n_494),
.Y(n_3115)
);

OAI211xp5_ASAP7_75t_L g3116 ( 
.A1(n_3094),
.A2(n_498),
.B(n_496),
.C(n_497),
.Y(n_3116)
);

AOI22xp5_ASAP7_75t_L g3117 ( 
.A1(n_3107),
.A2(n_499),
.B1(n_496),
.B2(n_497),
.Y(n_3117)
);

OAI22xp5_ASAP7_75t_L g3118 ( 
.A1(n_3060),
.A2(n_501),
.B1(n_499),
.B2(n_500),
.Y(n_3118)
);

INVx1_ASAP7_75t_L g3119 ( 
.A(n_3063),
.Y(n_3119)
);

NOR2xp33_ASAP7_75t_SL g3120 ( 
.A(n_3099),
.B(n_500),
.Y(n_3120)
);

NAND4xp25_ASAP7_75t_L g3121 ( 
.A(n_3079),
.B(n_503),
.C(n_501),
.D(n_502),
.Y(n_3121)
);

AOI211x1_ASAP7_75t_L g3122 ( 
.A1(n_3066),
.A2(n_3067),
.B(n_3058),
.C(n_3081),
.Y(n_3122)
);

AOI22xp5_ASAP7_75t_L g3123 ( 
.A1(n_3111),
.A2(n_504),
.B1(n_502),
.B2(n_503),
.Y(n_3123)
);

OA22x2_ASAP7_75t_L g3124 ( 
.A1(n_3072),
.A2(n_507),
.B1(n_505),
.B2(n_506),
.Y(n_3124)
);

O2A1O1Ixp5_ASAP7_75t_L g3125 ( 
.A1(n_3083),
.A2(n_507),
.B(n_505),
.C(n_506),
.Y(n_3125)
);

XNOR2xp5_ASAP7_75t_L g3126 ( 
.A(n_3065),
.B(n_508),
.Y(n_3126)
);

OAI211xp5_ASAP7_75t_SL g3127 ( 
.A1(n_3068),
.A2(n_511),
.B(n_509),
.C(n_510),
.Y(n_3127)
);

O2A1O1Ixp33_ASAP7_75t_L g3128 ( 
.A1(n_3062),
.A2(n_511),
.B(n_509),
.C(n_510),
.Y(n_3128)
);

NOR3x2_ASAP7_75t_L g3129 ( 
.A(n_3104),
.B(n_3086),
.C(n_3105),
.Y(n_3129)
);

NAND2xp5_ASAP7_75t_L g3130 ( 
.A(n_3100),
.B(n_512),
.Y(n_3130)
);

INVx2_ASAP7_75t_L g3131 ( 
.A(n_3071),
.Y(n_3131)
);

AOI211xp5_ASAP7_75t_L g3132 ( 
.A1(n_3076),
.A2(n_3057),
.B(n_3110),
.C(n_3098),
.Y(n_3132)
);

AOI221xp5_ASAP7_75t_L g3133 ( 
.A1(n_3095),
.A2(n_514),
.B1(n_512),
.B2(n_513),
.C(n_515),
.Y(n_3133)
);

OAI22xp33_ASAP7_75t_L g3134 ( 
.A1(n_3093),
.A2(n_516),
.B1(n_513),
.B2(n_515),
.Y(n_3134)
);

AOI22xp5_ASAP7_75t_L g3135 ( 
.A1(n_3064),
.A2(n_519),
.B1(n_516),
.B2(n_517),
.Y(n_3135)
);

AOI22xp5_ASAP7_75t_L g3136 ( 
.A1(n_3091),
.A2(n_521),
.B1(n_519),
.B2(n_520),
.Y(n_3136)
);

OAI211xp5_ASAP7_75t_SL g3137 ( 
.A1(n_3078),
.A2(n_523),
.B(n_520),
.C(n_522),
.Y(n_3137)
);

OAI221xp5_ASAP7_75t_L g3138 ( 
.A1(n_3075),
.A2(n_524),
.B1(n_522),
.B2(n_523),
.C(n_525),
.Y(n_3138)
);

NAND3x1_ASAP7_75t_SL g3139 ( 
.A(n_3069),
.B(n_524),
.C(n_526),
.Y(n_3139)
);

OAI31xp33_ASAP7_75t_L g3140 ( 
.A1(n_3070),
.A2(n_3077),
.A3(n_3090),
.B(n_3061),
.Y(n_3140)
);

AND2x4_ASAP7_75t_L g3141 ( 
.A(n_3074),
.B(n_526),
.Y(n_3141)
);

AOI221xp5_ASAP7_75t_L g3142 ( 
.A1(n_3092),
.A2(n_529),
.B1(n_527),
.B2(n_528),
.C(n_530),
.Y(n_3142)
);

AOI21xp5_ASAP7_75t_L g3143 ( 
.A1(n_3080),
.A2(n_527),
.B(n_528),
.Y(n_3143)
);

AOI221xp5_ASAP7_75t_L g3144 ( 
.A1(n_3089),
.A2(n_531),
.B1(n_529),
.B2(n_530),
.C(n_532),
.Y(n_3144)
);

AOI211xp5_ASAP7_75t_SL g3145 ( 
.A1(n_3082),
.A2(n_3055),
.B(n_3108),
.C(n_3073),
.Y(n_3145)
);

INVx1_ASAP7_75t_L g3146 ( 
.A(n_3102),
.Y(n_3146)
);

NOR3xp33_ASAP7_75t_L g3147 ( 
.A(n_3087),
.B(n_531),
.C(n_532),
.Y(n_3147)
);

NAND3x1_ASAP7_75t_L g3148 ( 
.A(n_3097),
.B(n_533),
.C(n_534),
.Y(n_3148)
);

OA22x2_ASAP7_75t_L g3149 ( 
.A1(n_3085),
.A2(n_535),
.B1(n_533),
.B2(n_534),
.Y(n_3149)
);

AOI211xp5_ASAP7_75t_L g3150 ( 
.A1(n_3088),
.A2(n_537),
.B(n_535),
.C(n_536),
.Y(n_3150)
);

NAND4xp25_ASAP7_75t_L g3151 ( 
.A(n_3084),
.B(n_538),
.C(n_536),
.D(n_537),
.Y(n_3151)
);

INVx1_ASAP7_75t_L g3152 ( 
.A(n_3063),
.Y(n_3152)
);

NAND3xp33_ASAP7_75t_L g3153 ( 
.A(n_3094),
.B(n_538),
.C(n_539),
.Y(n_3153)
);

AND2x4_ASAP7_75t_L g3154 ( 
.A(n_3106),
.B(n_539),
.Y(n_3154)
);

INVx1_ASAP7_75t_L g3155 ( 
.A(n_3063),
.Y(n_3155)
);

OAI221xp5_ASAP7_75t_SL g3156 ( 
.A1(n_3060),
.A2(n_542),
.B1(n_540),
.B2(n_541),
.C(n_543),
.Y(n_3156)
);

NOR2xp67_ASAP7_75t_L g3157 ( 
.A(n_3060),
.B(n_540),
.Y(n_3157)
);

AOI22xp5_ASAP7_75t_L g3158 ( 
.A1(n_3103),
.A2(n_544),
.B1(n_542),
.B2(n_543),
.Y(n_3158)
);

XOR2xp5_ASAP7_75t_L g3159 ( 
.A(n_3064),
.B(n_544),
.Y(n_3159)
);

NAND2xp5_ASAP7_75t_L g3160 ( 
.A(n_3106),
.B(n_545),
.Y(n_3160)
);

OAI211xp5_ASAP7_75t_L g3161 ( 
.A1(n_3094),
.A2(n_547),
.B(n_545),
.C(n_546),
.Y(n_3161)
);

AOI221xp5_ASAP7_75t_L g3162 ( 
.A1(n_3101),
.A2(n_549),
.B1(n_547),
.B2(n_548),
.C(n_550),
.Y(n_3162)
);

AOI211xp5_ASAP7_75t_L g3163 ( 
.A1(n_3106),
.A2(n_551),
.B(n_549),
.C(n_550),
.Y(n_3163)
);

AND2x4_ASAP7_75t_L g3164 ( 
.A(n_3154),
.B(n_551),
.Y(n_3164)
);

NOR3xp33_ASAP7_75t_L g3165 ( 
.A(n_3139),
.B(n_552),
.C(n_553),
.Y(n_3165)
);

XNOR2xp5_ASAP7_75t_L g3166 ( 
.A(n_3159),
.B(n_552),
.Y(n_3166)
);

INVx1_ASAP7_75t_L g3167 ( 
.A(n_3149),
.Y(n_3167)
);

NOR3x1_ASAP7_75t_L g3168 ( 
.A(n_3153),
.B(n_553),
.C(n_554),
.Y(n_3168)
);

INVx3_ASAP7_75t_L g3169 ( 
.A(n_3154),
.Y(n_3169)
);

XNOR2xp5_ASAP7_75t_L g3170 ( 
.A(n_3126),
.B(n_3129),
.Y(n_3170)
);

AOI22xp33_ASAP7_75t_L g3171 ( 
.A1(n_3119),
.A2(n_556),
.B1(n_554),
.B2(n_555),
.Y(n_3171)
);

XOR2x1_ASAP7_75t_L g3172 ( 
.A(n_3141),
.B(n_555),
.Y(n_3172)
);

NAND2x1p5_ASAP7_75t_L g3173 ( 
.A(n_3152),
.B(n_557),
.Y(n_3173)
);

AND3x2_ASAP7_75t_L g3174 ( 
.A(n_3141),
.B(n_3147),
.C(n_3163),
.Y(n_3174)
);

XOR2x2_ASAP7_75t_L g3175 ( 
.A(n_3148),
.B(n_558),
.Y(n_3175)
);

AOI22xp33_ASAP7_75t_L g3176 ( 
.A1(n_3155),
.A2(n_560),
.B1(n_558),
.B2(n_559),
.Y(n_3176)
);

NOR3xp33_ASAP7_75t_L g3177 ( 
.A(n_3131),
.B(n_559),
.C(n_560),
.Y(n_3177)
);

XNOR2x2_ASAP7_75t_SL g3178 ( 
.A(n_3112),
.B(n_561),
.Y(n_3178)
);

AND4x1_ASAP7_75t_L g3179 ( 
.A(n_3140),
.B(n_563),
.C(n_561),
.D(n_562),
.Y(n_3179)
);

NAND5xp2_ASAP7_75t_L g3180 ( 
.A(n_3145),
.B(n_566),
.C(n_564),
.D(n_565),
.E(n_567),
.Y(n_3180)
);

AND3x2_ASAP7_75t_L g3181 ( 
.A(n_3150),
.B(n_565),
.C(n_566),
.Y(n_3181)
);

INVx1_ASAP7_75t_L g3182 ( 
.A(n_3124),
.Y(n_3182)
);

INVx1_ASAP7_75t_L g3183 ( 
.A(n_3160),
.Y(n_3183)
);

OAI21xp33_ASAP7_75t_L g3184 ( 
.A1(n_3120),
.A2(n_567),
.B(n_568),
.Y(n_3184)
);

INVx2_ASAP7_75t_L g3185 ( 
.A(n_3125),
.Y(n_3185)
);

XOR2x1_ASAP7_75t_L g3186 ( 
.A(n_3134),
.B(n_569),
.Y(n_3186)
);

NOR3xp33_ASAP7_75t_L g3187 ( 
.A(n_3146),
.B(n_569),
.C(n_570),
.Y(n_3187)
);

INVx3_ASAP7_75t_L g3188 ( 
.A(n_3130),
.Y(n_3188)
);

XNOR2x1_ASAP7_75t_L g3189 ( 
.A(n_3135),
.B(n_570),
.Y(n_3189)
);

INVx3_ASAP7_75t_L g3190 ( 
.A(n_3157),
.Y(n_3190)
);

INVx2_ASAP7_75t_L g3191 ( 
.A(n_3113),
.Y(n_3191)
);

XNOR2x1_ASAP7_75t_L g3192 ( 
.A(n_3136),
.B(n_571),
.Y(n_3192)
);

INVxp67_ASAP7_75t_SL g3193 ( 
.A(n_3128),
.Y(n_3193)
);

NAND3xp33_ASAP7_75t_L g3194 ( 
.A(n_3132),
.B(n_572),
.C(n_573),
.Y(n_3194)
);

INVx1_ASAP7_75t_L g3195 ( 
.A(n_3114),
.Y(n_3195)
);

XOR2x1_ASAP7_75t_L g3196 ( 
.A(n_3118),
.B(n_572),
.Y(n_3196)
);

OR3x2_ASAP7_75t_L g3197 ( 
.A(n_3121),
.B(n_573),
.C(n_574),
.Y(n_3197)
);

OR2x6_ASAP7_75t_L g3198 ( 
.A(n_3122),
.B(n_574),
.Y(n_3198)
);

INVx1_ASAP7_75t_L g3199 ( 
.A(n_3116),
.Y(n_3199)
);

INVx1_ASAP7_75t_L g3200 ( 
.A(n_3161),
.Y(n_3200)
);

NAND3xp33_ASAP7_75t_SL g3201 ( 
.A(n_3115),
.B(n_575),
.C(n_576),
.Y(n_3201)
);

INVx2_ASAP7_75t_L g3202 ( 
.A(n_3138),
.Y(n_3202)
);

OR3x1_ASAP7_75t_L g3203 ( 
.A(n_3151),
.B(n_575),
.C(n_576),
.Y(n_3203)
);

AOI22xp5_ASAP7_75t_L g3204 ( 
.A1(n_3137),
.A2(n_579),
.B1(n_577),
.B2(n_578),
.Y(n_3204)
);

BUFx3_ASAP7_75t_L g3205 ( 
.A(n_3169),
.Y(n_3205)
);

AOI21x1_ASAP7_75t_L g3206 ( 
.A1(n_3198),
.A2(n_3175),
.B(n_3164),
.Y(n_3206)
);

INVx2_ASAP7_75t_L g3207 ( 
.A(n_3172),
.Y(n_3207)
);

NOR2xp67_ASAP7_75t_L g3208 ( 
.A(n_3180),
.B(n_3158),
.Y(n_3208)
);

NOR2x1_ASAP7_75t_SL g3209 ( 
.A(n_3198),
.B(n_3127),
.Y(n_3209)
);

NOR2xp33_ASAP7_75t_SL g3210 ( 
.A(n_3184),
.B(n_3156),
.Y(n_3210)
);

INVx2_ASAP7_75t_L g3211 ( 
.A(n_3173),
.Y(n_3211)
);

NOR2xp33_ASAP7_75t_L g3212 ( 
.A(n_3179),
.B(n_3143),
.Y(n_3212)
);

NAND2x1p5_ASAP7_75t_L g3213 ( 
.A(n_3190),
.B(n_3117),
.Y(n_3213)
);

NOR3xp33_ASAP7_75t_L g3214 ( 
.A(n_3193),
.B(n_3133),
.C(n_3162),
.Y(n_3214)
);

XNOR2xp5_ASAP7_75t_L g3215 ( 
.A(n_3166),
.B(n_3123),
.Y(n_3215)
);

XNOR2xp5_ASAP7_75t_L g3216 ( 
.A(n_3170),
.B(n_3142),
.Y(n_3216)
);

NAND2xp5_ASAP7_75t_L g3217 ( 
.A(n_3181),
.B(n_3144),
.Y(n_3217)
);

NAND2xp5_ASAP7_75t_L g3218 ( 
.A(n_3165),
.B(n_577),
.Y(n_3218)
);

INVx1_ASAP7_75t_L g3219 ( 
.A(n_3203),
.Y(n_3219)
);

INVx1_ASAP7_75t_L g3220 ( 
.A(n_3197),
.Y(n_3220)
);

AOI21xp5_ASAP7_75t_L g3221 ( 
.A1(n_3178),
.A2(n_579),
.B(n_580),
.Y(n_3221)
);

XOR2x1_ASAP7_75t_L g3222 ( 
.A(n_3185),
.B(n_580),
.Y(n_3222)
);

XNOR2xp5_ASAP7_75t_L g3223 ( 
.A(n_3189),
.B(n_581),
.Y(n_3223)
);

HB1xp67_ASAP7_75t_L g3224 ( 
.A(n_3186),
.Y(n_3224)
);

NOR3xp33_ASAP7_75t_L g3225 ( 
.A(n_3199),
.B(n_582),
.C(n_584),
.Y(n_3225)
);

NAND2xp5_ASAP7_75t_L g3226 ( 
.A(n_3177),
.B(n_582),
.Y(n_3226)
);

XNOR2xp5_ASAP7_75t_L g3227 ( 
.A(n_3192),
.B(n_584),
.Y(n_3227)
);

INVx1_ASAP7_75t_L g3228 ( 
.A(n_3196),
.Y(n_3228)
);

INVx2_ASAP7_75t_L g3229 ( 
.A(n_3168),
.Y(n_3229)
);

INVx1_ASAP7_75t_L g3230 ( 
.A(n_3194),
.Y(n_3230)
);

AND2x4_ASAP7_75t_L g3231 ( 
.A(n_3182),
.B(n_585),
.Y(n_3231)
);

HB1xp67_ASAP7_75t_L g3232 ( 
.A(n_3167),
.Y(n_3232)
);

OAI22x1_ASAP7_75t_L g3233 ( 
.A1(n_3204),
.A2(n_587),
.B1(n_585),
.B2(n_586),
.Y(n_3233)
);

INVx1_ASAP7_75t_L g3234 ( 
.A(n_3200),
.Y(n_3234)
);

XOR2xp5_ASAP7_75t_L g3235 ( 
.A(n_3201),
.B(n_587),
.Y(n_3235)
);

XOR2xp5_ASAP7_75t_L g3236 ( 
.A(n_3195),
.B(n_588),
.Y(n_3236)
);

OAI22xp5_ASAP7_75t_SL g3237 ( 
.A1(n_3235),
.A2(n_3191),
.B1(n_3202),
.B2(n_3183),
.Y(n_3237)
);

OA21x2_ASAP7_75t_L g3238 ( 
.A1(n_3221),
.A2(n_3176),
.B(n_3171),
.Y(n_3238)
);

INVx1_ASAP7_75t_L g3239 ( 
.A(n_3236),
.Y(n_3239)
);

INVx3_ASAP7_75t_L g3240 ( 
.A(n_3205),
.Y(n_3240)
);

AOI21xp5_ASAP7_75t_L g3241 ( 
.A1(n_3209),
.A2(n_3188),
.B(n_3187),
.Y(n_3241)
);

NAND2xp5_ASAP7_75t_L g3242 ( 
.A(n_3231),
.B(n_3174),
.Y(n_3242)
);

INVx1_ASAP7_75t_L g3243 ( 
.A(n_3222),
.Y(n_3243)
);

INVx1_ASAP7_75t_L g3244 ( 
.A(n_3218),
.Y(n_3244)
);

OAI211xp5_ASAP7_75t_SL g3245 ( 
.A1(n_3234),
.A2(n_590),
.B(n_588),
.C(n_589),
.Y(n_3245)
);

INVx1_ASAP7_75t_L g3246 ( 
.A(n_3232),
.Y(n_3246)
);

OAI22xp5_ASAP7_75t_SL g3247 ( 
.A1(n_3228),
.A2(n_591),
.B1(n_589),
.B2(n_590),
.Y(n_3247)
);

OAI21x1_ASAP7_75t_L g3248 ( 
.A1(n_3206),
.A2(n_591),
.B(n_593),
.Y(n_3248)
);

INVx1_ASAP7_75t_L g3249 ( 
.A(n_3223),
.Y(n_3249)
);

NAND2xp5_ASAP7_75t_L g3250 ( 
.A(n_3225),
.B(n_594),
.Y(n_3250)
);

NOR2xp33_ASAP7_75t_SL g3251 ( 
.A(n_3224),
.B(n_594),
.Y(n_3251)
);

NAND2xp5_ASAP7_75t_SL g3252 ( 
.A(n_3246),
.B(n_3208),
.Y(n_3252)
);

INVx2_ASAP7_75t_L g3253 ( 
.A(n_3248),
.Y(n_3253)
);

INVx1_ASAP7_75t_L g3254 ( 
.A(n_3240),
.Y(n_3254)
);

BUFx2_ASAP7_75t_SL g3255 ( 
.A(n_3243),
.Y(n_3255)
);

OAI22xp5_ASAP7_75t_L g3256 ( 
.A1(n_3242),
.A2(n_3219),
.B1(n_3207),
.B2(n_3220),
.Y(n_3256)
);

OAI22xp5_ASAP7_75t_L g3257 ( 
.A1(n_3250),
.A2(n_3226),
.B1(n_3213),
.B2(n_3211),
.Y(n_3257)
);

NAND2xp5_ASAP7_75t_L g3258 ( 
.A(n_3251),
.B(n_3233),
.Y(n_3258)
);

INVx1_ASAP7_75t_L g3259 ( 
.A(n_3247),
.Y(n_3259)
);

INVxp67_ASAP7_75t_SL g3260 ( 
.A(n_3238),
.Y(n_3260)
);

NAND3xp33_ASAP7_75t_L g3261 ( 
.A(n_3241),
.B(n_3214),
.C(n_3227),
.Y(n_3261)
);

INVx1_ASAP7_75t_L g3262 ( 
.A(n_3237),
.Y(n_3262)
);

INVx1_ASAP7_75t_L g3263 ( 
.A(n_3245),
.Y(n_3263)
);

BUFx2_ASAP7_75t_L g3264 ( 
.A(n_3239),
.Y(n_3264)
);

OAI21xp5_ASAP7_75t_L g3265 ( 
.A1(n_3260),
.A2(n_3212),
.B(n_3216),
.Y(n_3265)
);

OA22x2_ASAP7_75t_L g3266 ( 
.A1(n_3262),
.A2(n_3215),
.B1(n_3230),
.B2(n_3229),
.Y(n_3266)
);

OAI22x1_ASAP7_75t_L g3267 ( 
.A1(n_3259),
.A2(n_3249),
.B1(n_3244),
.B2(n_3217),
.Y(n_3267)
);

INVx1_ASAP7_75t_L g3268 ( 
.A(n_3258),
.Y(n_3268)
);

AO22x1_ASAP7_75t_L g3269 ( 
.A1(n_3253),
.A2(n_3210),
.B1(n_597),
.B2(n_595),
.Y(n_3269)
);

OA22x2_ASAP7_75t_L g3270 ( 
.A1(n_3255),
.A2(n_597),
.B1(n_595),
.B2(n_596),
.Y(n_3270)
);

OAI22xp5_ASAP7_75t_L g3271 ( 
.A1(n_3254),
.A2(n_3261),
.B1(n_3263),
.B2(n_3264),
.Y(n_3271)
);

OAI22xp5_ASAP7_75t_L g3272 ( 
.A1(n_3252),
.A2(n_599),
.B1(n_596),
.B2(n_598),
.Y(n_3272)
);

OA21x2_ASAP7_75t_L g3273 ( 
.A1(n_3256),
.A2(n_3257),
.B(n_598),
.Y(n_3273)
);

BUFx2_ASAP7_75t_L g3274 ( 
.A(n_3253),
.Y(n_3274)
);

CKINVDCx20_ASAP7_75t_R g3275 ( 
.A(n_3264),
.Y(n_3275)
);

NAND2xp5_ASAP7_75t_L g3276 ( 
.A(n_3269),
.B(n_600),
.Y(n_3276)
);

INVx1_ASAP7_75t_L g3277 ( 
.A(n_3270),
.Y(n_3277)
);

INVx4_ASAP7_75t_L g3278 ( 
.A(n_3274),
.Y(n_3278)
);

INVxp67_ASAP7_75t_L g3279 ( 
.A(n_3273),
.Y(n_3279)
);

OAI21xp5_ASAP7_75t_L g3280 ( 
.A1(n_3265),
.A2(n_600),
.B(n_601),
.Y(n_3280)
);

OAI21x1_ASAP7_75t_SL g3281 ( 
.A1(n_3272),
.A2(n_601),
.B(n_602),
.Y(n_3281)
);

INVx1_ASAP7_75t_L g3282 ( 
.A(n_3275),
.Y(n_3282)
);

OAI22xp5_ASAP7_75t_L g3283 ( 
.A1(n_3268),
.A2(n_604),
.B1(n_602),
.B2(n_603),
.Y(n_3283)
);

AOI22xp5_ASAP7_75t_L g3284 ( 
.A1(n_3271),
.A2(n_605),
.B1(n_603),
.B2(n_604),
.Y(n_3284)
);

AOI21xp5_ASAP7_75t_L g3285 ( 
.A1(n_3267),
.A2(n_3266),
.B(n_605),
.Y(n_3285)
);

OAI21xp5_ASAP7_75t_L g3286 ( 
.A1(n_3265),
.A2(n_606),
.B(n_607),
.Y(n_3286)
);

AOI221xp5_ASAP7_75t_L g3287 ( 
.A1(n_3285),
.A2(n_608),
.B1(n_606),
.B2(n_607),
.C(n_609),
.Y(n_3287)
);

OAI22xp5_ASAP7_75t_L g3288 ( 
.A1(n_3282),
.A2(n_611),
.B1(n_609),
.B2(n_610),
.Y(n_3288)
);

OAI21xp33_ASAP7_75t_L g3289 ( 
.A1(n_3280),
.A2(n_610),
.B(n_611),
.Y(n_3289)
);

NAND2xp5_ASAP7_75t_SL g3290 ( 
.A(n_3278),
.B(n_612),
.Y(n_3290)
);

NOR2xp33_ASAP7_75t_L g3291 ( 
.A(n_3278),
.B(n_612),
.Y(n_3291)
);

INVxp33_ASAP7_75t_SL g3292 ( 
.A(n_3277),
.Y(n_3292)
);

OAI21xp5_ASAP7_75t_L g3293 ( 
.A1(n_3276),
.A2(n_613),
.B(n_614),
.Y(n_3293)
);

NAND2xp5_ASAP7_75t_L g3294 ( 
.A(n_3286),
.B(n_613),
.Y(n_3294)
);

NAND2xp5_ASAP7_75t_L g3295 ( 
.A(n_3284),
.B(n_614),
.Y(n_3295)
);

AOI21xp5_ASAP7_75t_L g3296 ( 
.A1(n_3292),
.A2(n_3279),
.B(n_3281),
.Y(n_3296)
);

AOI21xp5_ASAP7_75t_L g3297 ( 
.A1(n_3294),
.A2(n_3283),
.B(n_615),
.Y(n_3297)
);

AOI22xp33_ASAP7_75t_L g3298 ( 
.A1(n_3289),
.A2(n_617),
.B1(n_615),
.B2(n_616),
.Y(n_3298)
);

AOI22xp5_ASAP7_75t_L g3299 ( 
.A1(n_3287),
.A2(n_619),
.B1(n_616),
.B2(n_618),
.Y(n_3299)
);

INVx2_ASAP7_75t_L g3300 ( 
.A(n_3290),
.Y(n_3300)
);

AOI22xp5_ASAP7_75t_L g3301 ( 
.A1(n_3299),
.A2(n_3295),
.B1(n_3293),
.B2(n_3288),
.Y(n_3301)
);

AOI22xp33_ASAP7_75t_L g3302 ( 
.A1(n_3300),
.A2(n_3291),
.B1(n_621),
.B2(n_618),
.Y(n_3302)
);

AOI22xp33_ASAP7_75t_L g3303 ( 
.A1(n_3296),
.A2(n_622),
.B1(n_620),
.B2(n_621),
.Y(n_3303)
);

OAI21x1_ASAP7_75t_SL g3304 ( 
.A1(n_3301),
.A2(n_3297),
.B(n_3298),
.Y(n_3304)
);

OR2x6_ASAP7_75t_L g3305 ( 
.A(n_3302),
.B(n_620),
.Y(n_3305)
);

AOI21xp5_ASAP7_75t_L g3306 ( 
.A1(n_3304),
.A2(n_3303),
.B(n_622),
.Y(n_3306)
);

AOI211xp5_ASAP7_75t_L g3307 ( 
.A1(n_3306),
.A2(n_3305),
.B(n_625),
.C(n_623),
.Y(n_3307)
);


endmodule