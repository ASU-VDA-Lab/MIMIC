module real_aes_393_n_78 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_77, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_78);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_78;
wire n_480;
wire n_113;
wire n_476;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_522;
wire n_485;
wire n_222;
wire n_357;
wire n_287;
wire n_503;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_341;
wire n_232;
wire n_460;
wire n_401;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_320;
wire n_260;
wire n_97;
wire n_186;
wire n_138;
wire n_453;
wire n_379;
wire n_374;
wire n_235;
wire n_399;
wire n_378;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_145;
wire n_415;
wire n_227;
wire n_519;
wire n_92;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_292;
wire n_400;
wire n_116;
wire n_94;
wire n_289;
wire n_462;
wire n_280;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_408;
wire n_184;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_530;
wire n_104;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_506;
wire n_513;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_231;
wire n_102;
wire n_454;
wire n_122;
wire n_443;
wire n_534;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_204;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_331;
wire n_93;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_323;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_368;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_250;
wire n_85;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_402;
wire n_87;
wire n_171;
wire n_531;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_488;
wire n_501;
wire n_251;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_288;
wire n_147;
wire n_150;
wire n_404;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_158;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_109;
wire n_203;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_526;
wire n_155;
wire n_243;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_446;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_180;
wire n_212;
wire n_210;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_371;
wire n_103;
wire n_166;
wire n_224;
wire n_151;
wire n_130;
wire n_253;
wire n_459;
wire n_99;
wire n_440;
wire n_525;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_305;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_465;
wire n_473;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_340;
wire n_483;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_206;
wire n_307;
wire n_500;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_264;
wire n_237;
wire n_91;
AO22x2_ASAP7_75t_L g95 ( .A1(n_0), .A2(n_55), .B1(n_96), .B2(n_97), .Y(n_95) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_1), .B(n_224), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_2), .B(n_250), .Y(n_262) );
INVx1_ASAP7_75t_L g196 ( .A(n_3), .Y(n_196) );
AO22x2_ASAP7_75t_L g99 ( .A1(n_4), .A2(n_13), .B1(n_96), .B2(n_100), .Y(n_99) );
AND2x2_ASAP7_75t_L g253 ( .A(n_5), .B(n_254), .Y(n_253) );
AOI22xp5_ASAP7_75t_L g144 ( .A1(n_6), .A2(n_34), .B1(n_145), .B2(n_148), .Y(n_144) );
AND2x2_ASAP7_75t_L g264 ( .A(n_7), .B(n_265), .Y(n_264) );
INVx2_ASAP7_75t_L g213 ( .A(n_8), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_9), .B(n_250), .Y(n_319) );
AOI22xp5_ASAP7_75t_L g166 ( .A1(n_10), .A2(n_24), .B1(n_167), .B2(n_170), .Y(n_166) );
NAND2xp5_ASAP7_75t_SL g304 ( .A(n_11), .B(n_224), .Y(n_304) );
AOI22xp33_ASAP7_75t_L g216 ( .A1(n_12), .A2(n_71), .B1(n_217), .B2(n_224), .Y(n_216) );
OAI221xp5_ASAP7_75t_L g188 ( .A1(n_13), .A2(n_55), .B1(n_60), .B2(n_189), .C(n_191), .Y(n_188) );
OR2x2_ASAP7_75t_L g214 ( .A(n_14), .B(n_69), .Y(n_214) );
OA21x2_ASAP7_75t_L g243 ( .A1(n_14), .A2(n_69), .B(n_213), .Y(n_243) );
OAI22xp5_ASAP7_75t_SL g176 ( .A1(n_15), .A2(n_26), .B1(n_177), .B2(n_178), .Y(n_176) );
INVxp67_ASAP7_75t_L g178 ( .A(n_15), .Y(n_178) );
CKINVDCx20_ASAP7_75t_R g89 ( .A(n_16), .Y(n_89) );
INVx3_ASAP7_75t_L g96 ( .A(n_17), .Y(n_96) );
AO21x2_ASAP7_75t_L g314 ( .A1(n_18), .A2(n_254), .B(n_315), .Y(n_314) );
AOI21xp5_ASAP7_75t_L g259 ( .A1(n_19), .A2(n_232), .B(n_260), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_20), .B(n_250), .Y(n_299) );
INVx1_ASAP7_75t_L g534 ( .A(n_20), .Y(n_534) );
INVx1_ASAP7_75t_SL g104 ( .A(n_21), .Y(n_104) );
AOI22xp33_ASAP7_75t_L g152 ( .A1(n_22), .A2(n_48), .B1(n_153), .B2(n_158), .Y(n_152) );
INVx1_ASAP7_75t_L g198 ( .A(n_23), .Y(n_198) );
AND2x2_ASAP7_75t_L g222 ( .A(n_23), .B(n_223), .Y(n_222) );
AND2x2_ASAP7_75t_L g230 ( .A(n_23), .B(n_196), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_25), .B(n_224), .Y(n_263) );
INVx1_ASAP7_75t_L g177 ( .A(n_26), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_27), .B(n_250), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_28), .B(n_224), .Y(n_272) );
AOI22xp5_ASAP7_75t_L g128 ( .A1(n_29), .A2(n_33), .B1(n_129), .B2(n_134), .Y(n_128) );
AOI21xp5_ASAP7_75t_L g245 ( .A1(n_30), .A2(n_232), .B(n_246), .Y(n_245) );
AO22x2_ASAP7_75t_L g107 ( .A1(n_31), .A2(n_60), .B1(n_96), .B2(n_108), .Y(n_107) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_32), .B(n_248), .Y(n_276) );
NAND2xp5_ASAP7_75t_SL g316 ( .A(n_35), .B(n_224), .Y(n_316) );
INVx1_ASAP7_75t_L g220 ( .A(n_36), .Y(n_220) );
INVx1_ASAP7_75t_L g227 ( .A(n_36), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_37), .B(n_250), .Y(n_249) );
AOI22xp33_ASAP7_75t_L g160 ( .A1(n_38), .A2(n_70), .B1(n_161), .B2(n_163), .Y(n_160) );
AND2x2_ASAP7_75t_L g284 ( .A(n_39), .B(n_211), .Y(n_284) );
INVx1_ASAP7_75t_L g105 ( .A(n_40), .Y(n_105) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_41), .B(n_248), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_42), .B(n_248), .Y(n_298) );
NAND2xp5_ASAP7_75t_SL g252 ( .A(n_43), .B(n_224), .Y(n_252) );
AOI22xp5_ASAP7_75t_L g173 ( .A1(n_44), .A2(n_174), .B1(n_183), .B2(n_184), .Y(n_173) );
INVx1_ASAP7_75t_L g183 ( .A(n_44), .Y(n_183) );
NAND2xp5_ASAP7_75t_SL g286 ( .A(n_45), .B(n_224), .Y(n_286) );
AOI21xp5_ASAP7_75t_L g296 ( .A1(n_46), .A2(n_232), .B(n_297), .Y(n_296) );
AOI22xp5_ASAP7_75t_L g518 ( .A1(n_46), .A2(n_85), .B1(n_86), .B2(n_519), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_46), .Y(n_519) );
AND2x2_ASAP7_75t_L g310 ( .A(n_47), .B(n_212), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_49), .B(n_248), .Y(n_290) );
AOI22xp33_ASAP7_75t_L g117 ( .A1(n_50), .A2(n_76), .B1(n_118), .B2(n_124), .Y(n_117) );
AOI22xp5_ASAP7_75t_L g179 ( .A1(n_51), .A2(n_59), .B1(n_180), .B2(n_181), .Y(n_179) );
INVx1_ASAP7_75t_L g181 ( .A(n_51), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_52), .B(n_248), .Y(n_320) );
AOI22xp5_ASAP7_75t_L g525 ( .A1(n_53), .A2(n_85), .B1(n_86), .B2(n_526), .Y(n_525) );
CKINVDCx20_ASAP7_75t_R g526 ( .A(n_53), .Y(n_526) );
OAI22xp5_ASAP7_75t_SL g82 ( .A1(n_54), .A2(n_72), .B1(n_83), .B2(n_84), .Y(n_82) );
INVx1_ASAP7_75t_L g84 ( .A(n_54), .Y(n_84) );
AOI22xp5_ASAP7_75t_L g231 ( .A1(n_54), .A2(n_73), .B1(n_232), .B2(n_234), .Y(n_231) );
INVxp33_ASAP7_75t_L g193 ( .A(n_55), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_56), .B(n_250), .Y(n_307) );
INVx1_ASAP7_75t_L g223 ( .A(n_57), .Y(n_223) );
INVx1_ASAP7_75t_L g229 ( .A(n_57), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_58), .B(n_248), .Y(n_261) );
INVx1_ASAP7_75t_L g180 ( .A(n_59), .Y(n_180) );
INVxp67_ASAP7_75t_L g192 ( .A(n_60), .Y(n_192) );
AOI21xp5_ASAP7_75t_L g287 ( .A1(n_61), .A2(n_232), .B(n_288), .Y(n_287) );
AOI21xp5_ASAP7_75t_L g273 ( .A1(n_62), .A2(n_232), .B(n_274), .Y(n_273) );
AOI21xp5_ASAP7_75t_L g317 ( .A1(n_63), .A2(n_232), .B(n_318), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_64), .B(n_110), .Y(n_109) );
AND2x2_ASAP7_75t_L g301 ( .A(n_65), .B(n_212), .Y(n_301) );
NAND2xp5_ASAP7_75t_SL g210 ( .A(n_66), .B(n_211), .Y(n_210) );
AND2x2_ASAP7_75t_L g277 ( .A(n_67), .B(n_265), .Y(n_277) );
NAND2xp33_ASAP7_75t_SL g137 ( .A(n_68), .B(n_138), .Y(n_137) );
INVx1_ASAP7_75t_L g83 ( .A(n_72), .Y(n_83) );
AOI21xp5_ASAP7_75t_L g305 ( .A1(n_72), .A2(n_232), .B(n_306), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_74), .B(n_250), .Y(n_275) );
BUFx2_ASAP7_75t_L g309 ( .A(n_75), .Y(n_309) );
BUFx2_ASAP7_75t_SL g190 ( .A(n_77), .Y(n_190) );
AOI221xp5_ASAP7_75t_L g78 ( .A1(n_79), .A2(n_185), .B1(n_199), .B2(n_516), .C(n_517), .Y(n_78) );
XOR2xp5_ASAP7_75t_L g79 ( .A(n_80), .B(n_173), .Y(n_79) );
AOI22xp5_ASAP7_75t_L g80 ( .A1(n_81), .A2(n_82), .B1(n_85), .B2(n_86), .Y(n_80) );
CKINVDCx16_ASAP7_75t_R g81 ( .A(n_82), .Y(n_81) );
INVx1_ASAP7_75t_L g85 ( .A(n_86), .Y(n_85) );
OR2x2_ASAP7_75t_L g86 ( .A(n_87), .B(n_143), .Y(n_86) );
NAND4xp25_ASAP7_75t_L g87 ( .A(n_88), .B(n_117), .C(n_128), .D(n_137), .Y(n_87) );
OA21x2_ASAP7_75t_SL g88 ( .A1(n_89), .A2(n_90), .B(n_109), .Y(n_88) );
INVxp33_ASAP7_75t_L g90 ( .A(n_91), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_92), .Y(n_91) );
INVx3_ASAP7_75t_L g92 ( .A(n_93), .Y(n_92) );
AND2x2_ASAP7_75t_L g93 ( .A(n_94), .B(n_101), .Y(n_93) );
AND2x4_ASAP7_75t_L g150 ( .A(n_94), .B(n_151), .Y(n_150) );
AND2x2_ASAP7_75t_L g157 ( .A(n_94), .B(n_122), .Y(n_157) );
AND2x2_ASAP7_75t_L g94 ( .A(n_95), .B(n_98), .Y(n_94) );
INVx2_ASAP7_75t_L g116 ( .A(n_95), .Y(n_116) );
AND2x2_ASAP7_75t_L g132 ( .A(n_95), .B(n_99), .Y(n_132) );
INVx1_ASAP7_75t_L g97 ( .A(n_96), .Y(n_97) );
INVx2_ASAP7_75t_L g100 ( .A(n_96), .Y(n_100) );
OAI22x1_ASAP7_75t_L g102 ( .A1(n_96), .A2(n_103), .B1(n_104), .B2(n_105), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_96), .Y(n_103) );
INVx1_ASAP7_75t_L g108 ( .A(n_96), .Y(n_108) );
HB1xp67_ASAP7_75t_L g142 ( .A(n_98), .Y(n_142) );
INVx1_ASAP7_75t_L g98 ( .A(n_99), .Y(n_98) );
INVx1_ASAP7_75t_L g115 ( .A(n_99), .Y(n_115) );
AND2x4_ASAP7_75t_L g121 ( .A(n_99), .B(n_116), .Y(n_121) );
AND2x2_ASAP7_75t_L g136 ( .A(n_101), .B(n_121), .Y(n_136) );
AND2x4_ASAP7_75t_L g162 ( .A(n_101), .B(n_114), .Y(n_162) );
AND2x2_ASAP7_75t_L g101 ( .A(n_102), .B(n_106), .Y(n_101) );
AND2x2_ASAP7_75t_L g113 ( .A(n_102), .B(n_107), .Y(n_113) );
INVx2_ASAP7_75t_L g123 ( .A(n_102), .Y(n_123) );
HB1xp67_ASAP7_75t_L g133 ( .A(n_102), .Y(n_133) );
AND2x4_ASAP7_75t_L g151 ( .A(n_106), .B(n_123), .Y(n_151) );
INVx2_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
AND2x2_ASAP7_75t_L g122 ( .A(n_107), .B(n_123), .Y(n_122) );
BUFx2_ASAP7_75t_L g159 ( .A(n_107), .Y(n_159) );
INVx3_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
INVx6_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
AND2x2_ASAP7_75t_L g112 ( .A(n_113), .B(n_114), .Y(n_112) );
AND2x4_ASAP7_75t_L g126 ( .A(n_113), .B(n_127), .Y(n_126) );
AND2x4_ASAP7_75t_L g140 ( .A(n_113), .B(n_141), .Y(n_140) );
AND2x2_ASAP7_75t_L g147 ( .A(n_114), .B(n_122), .Y(n_147) );
AND2x4_ASAP7_75t_L g172 ( .A(n_114), .B(n_151), .Y(n_172) );
AND2x4_ASAP7_75t_L g114 ( .A(n_115), .B(n_116), .Y(n_114) );
INVxp67_ASAP7_75t_L g127 ( .A(n_116), .Y(n_127) );
BUFx2_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
BUFx6f_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
AND2x4_ASAP7_75t_L g120 ( .A(n_121), .B(n_122), .Y(n_120) );
AND2x4_ASAP7_75t_L g165 ( .A(n_121), .B(n_151), .Y(n_165) );
INVx2_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
INVx6_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
INVx3_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
INVx3_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
AND2x2_ASAP7_75t_L g131 ( .A(n_132), .B(n_133), .Y(n_131) );
AND2x4_ASAP7_75t_L g158 ( .A(n_132), .B(n_159), .Y(n_158) );
AND2x4_ASAP7_75t_L g169 ( .A(n_132), .B(n_151), .Y(n_169) );
BUFx6f_ASAP7_75t_SL g134 ( .A(n_135), .Y(n_134) );
BUFx3_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
BUFx6f_ASAP7_75t_SL g138 ( .A(n_139), .Y(n_138) );
BUFx3_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
INVx1_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
NAND4xp25_ASAP7_75t_L g143 ( .A(n_144), .B(n_152), .C(n_160), .D(n_166), .Y(n_143) );
BUFx3_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
BUFx2_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx2_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx8_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx1_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx2_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx2_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
BUFx3_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
BUFx6f_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
BUFx6f_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
BUFx6f_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
BUFx3_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
INVx2_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
INVx8_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
CKINVDCx20_ASAP7_75t_R g184 ( .A(n_174), .Y(n_184) );
AOI22xp5_ASAP7_75t_L g174 ( .A1(n_175), .A2(n_176), .B1(n_179), .B2(n_182), .Y(n_174) );
CKINVDCx20_ASAP7_75t_R g175 ( .A(n_176), .Y(n_175) );
CKINVDCx20_ASAP7_75t_R g182 ( .A(n_179), .Y(n_182) );
CKINVDCx20_ASAP7_75t_R g185 ( .A(n_186), .Y(n_185) );
CKINVDCx20_ASAP7_75t_R g186 ( .A(n_187), .Y(n_186) );
AND3x1_ASAP7_75t_SL g187 ( .A(n_188), .B(n_194), .C(n_197), .Y(n_187) );
INVxp67_ASAP7_75t_L g524 ( .A(n_188), .Y(n_524) );
CKINVDCx8_ASAP7_75t_R g189 ( .A(n_190), .Y(n_189) );
NOR2xp33_ASAP7_75t_L g191 ( .A(n_192), .B(n_193), .Y(n_191) );
CKINVDCx16_ASAP7_75t_R g522 ( .A(n_194), .Y(n_522) );
OAI21xp5_ASAP7_75t_L g531 ( .A1(n_194), .A2(n_532), .B(n_533), .Y(n_531) );
INVx1_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
AND2x2_ASAP7_75t_L g218 ( .A(n_195), .B(n_219), .Y(n_218) );
OR2x2_ASAP7_75t_SL g529 ( .A(n_195), .B(n_197), .Y(n_529) );
HB1xp67_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
AND2x2_ASAP7_75t_L g233 ( .A(n_196), .B(n_220), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_197), .B(n_524), .Y(n_523) );
INVx1_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
NOR2x1p5_ASAP7_75t_L g235 ( .A(n_198), .B(n_236), .Y(n_235) );
HB1xp67_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
OR2x6_ASAP7_75t_L g200 ( .A(n_201), .B(n_453), .Y(n_200) );
NAND3xp33_ASAP7_75t_L g201 ( .A(n_202), .B(n_369), .C(n_406), .Y(n_201) );
NOR3xp33_ASAP7_75t_L g202 ( .A(n_203), .B(n_337), .C(n_352), .Y(n_202) );
OAI221xp5_ASAP7_75t_L g203 ( .A1(n_204), .A2(n_281), .B1(n_311), .B2(n_323), .C(n_324), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
NAND2xp5_ASAP7_75t_SL g205 ( .A(n_206), .B(n_266), .Y(n_205) );
OAI22xp33_ASAP7_75t_SL g397 ( .A1(n_206), .A2(n_361), .B1(n_398), .B2(n_401), .Y(n_397) );
OR2x2_ASAP7_75t_L g206 ( .A(n_207), .B(n_238), .Y(n_206) );
OAI21xp33_ASAP7_75t_SL g407 ( .A1(n_207), .A2(n_408), .B(n_414), .Y(n_407) );
OR2x2_ASAP7_75t_L g436 ( .A(n_207), .B(n_268), .Y(n_436) );
AND2x2_ASAP7_75t_L g437 ( .A(n_207), .B(n_356), .Y(n_437) );
INVx2_ASAP7_75t_L g468 ( .A(n_207), .Y(n_468) );
INVx2_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_208), .B(n_328), .Y(n_449) );
INVx2_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
OR2x2_ASAP7_75t_L g323 ( .A(n_209), .B(n_241), .Y(n_323) );
BUFx3_ASAP7_75t_L g349 ( .A(n_209), .Y(n_349) );
AND2x2_ASAP7_75t_L g485 ( .A(n_209), .B(n_486), .Y(n_485) );
AND2x2_ASAP7_75t_L g508 ( .A(n_209), .B(n_269), .Y(n_508) );
AND2x4_ASAP7_75t_L g209 ( .A(n_210), .B(n_215), .Y(n_209) );
AND2x4_ASAP7_75t_L g280 ( .A(n_210), .B(n_215), .Y(n_280) );
AO21x2_ASAP7_75t_L g215 ( .A1(n_211), .A2(n_216), .B(n_231), .Y(n_215) );
CKINVDCx5p33_ASAP7_75t_R g257 ( .A(n_211), .Y(n_257) );
AOI21xp5_ASAP7_75t_L g271 ( .A1(n_211), .A2(n_272), .B(n_273), .Y(n_271) );
BUFx6f_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
AND2x2_ASAP7_75t_SL g212 ( .A(n_213), .B(n_214), .Y(n_212) );
AND2x4_ASAP7_75t_L g291 ( .A(n_213), .B(n_214), .Y(n_291) );
AND2x4_ASAP7_75t_L g217 ( .A(n_218), .B(n_221), .Y(n_217) );
INVx1_ASAP7_75t_L g533 ( .A(n_218), .Y(n_533) );
INVx2_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
AND2x4_ASAP7_75t_L g250 ( .A(n_220), .B(n_228), .Y(n_250) );
BUFx3_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
AND2x6_ASAP7_75t_L g232 ( .A(n_222), .B(n_233), .Y(n_232) );
INVx2_ASAP7_75t_L g237 ( .A(n_223), .Y(n_237) );
AND2x6_ASAP7_75t_L g248 ( .A(n_223), .B(n_226), .Y(n_248) );
AND2x4_ASAP7_75t_L g224 ( .A(n_225), .B(n_230), .Y(n_224) );
AND2x4_ASAP7_75t_L g225 ( .A(n_226), .B(n_228), .Y(n_225) );
INVx2_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
INVx2_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
INVx5_ASAP7_75t_L g251 ( .A(n_230), .Y(n_251) );
AND2x4_ASAP7_75t_L g234 ( .A(n_233), .B(n_235), .Y(n_234) );
HB1xp67_ASAP7_75t_L g516 ( .A(n_234), .Y(n_516) );
HB1xp67_ASAP7_75t_L g532 ( .A(n_235), .Y(n_532) );
INVx3_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
INVx1_ASAP7_75t_SL g238 ( .A(n_239), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_239), .B(n_269), .Y(n_428) );
INVx1_ASAP7_75t_L g465 ( .A(n_239), .Y(n_465) );
AND2x2_ASAP7_75t_L g239 ( .A(n_240), .B(n_255), .Y(n_239) );
AND2x2_ASAP7_75t_L g279 ( .A(n_240), .B(n_280), .Y(n_279) );
INVx1_ASAP7_75t_L g486 ( .A(n_240), .Y(n_486) );
INVx2_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
INVx2_ASAP7_75t_L g329 ( .A(n_241), .Y(n_329) );
AND2x2_ASAP7_75t_L g330 ( .A(n_241), .B(n_255), .Y(n_330) );
AND2x2_ASAP7_75t_L g351 ( .A(n_241), .B(n_270), .Y(n_351) );
AND2x2_ASAP7_75t_L g433 ( .A(n_241), .B(n_256), .Y(n_433) );
AO21x2_ASAP7_75t_L g241 ( .A1(n_242), .A2(n_244), .B(n_253), .Y(n_241) );
INVx4_ASAP7_75t_L g254 ( .A(n_242), .Y(n_254) );
INVx3_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
BUFx4f_ASAP7_75t_L g265 ( .A(n_243), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_245), .B(n_252), .Y(n_244) );
AOI21xp5_ASAP7_75t_L g246 ( .A1(n_247), .A2(n_249), .B(n_251), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_248), .B(n_309), .Y(n_308) );
AOI21xp5_ASAP7_75t_L g260 ( .A1(n_251), .A2(n_261), .B(n_262), .Y(n_260) );
AOI21xp5_ASAP7_75t_L g274 ( .A1(n_251), .A2(n_275), .B(n_276), .Y(n_274) );
AOI21xp5_ASAP7_75t_L g288 ( .A1(n_251), .A2(n_289), .B(n_290), .Y(n_288) );
AOI21xp5_ASAP7_75t_L g297 ( .A1(n_251), .A2(n_298), .B(n_299), .Y(n_297) );
AOI21xp5_ASAP7_75t_L g306 ( .A1(n_251), .A2(n_307), .B(n_308), .Y(n_306) );
AOI21xp5_ASAP7_75t_L g318 ( .A1(n_251), .A2(n_319), .B(n_320), .Y(n_318) );
INVx3_ASAP7_75t_L g294 ( .A(n_254), .Y(n_294) );
AND2x4_ASAP7_75t_SL g326 ( .A(n_255), .B(n_270), .Y(n_326) );
INVx1_ASAP7_75t_L g357 ( .A(n_255), .Y(n_357) );
INVx2_ASAP7_75t_L g365 ( .A(n_255), .Y(n_365) );
HB1xp67_ASAP7_75t_L g389 ( .A(n_255), .Y(n_389) );
INVx3_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
HB1xp67_ASAP7_75t_L g278 ( .A(n_256), .Y(n_278) );
AOI21x1_ASAP7_75t_L g256 ( .A1(n_257), .A2(n_258), .B(n_264), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_259), .B(n_263), .Y(n_258) );
AOI21xp5_ASAP7_75t_L g303 ( .A1(n_265), .A2(n_304), .B(n_305), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_267), .B(n_279), .Y(n_266) );
AND2x2_ASAP7_75t_L g504 ( .A(n_267), .B(n_367), .Y(n_504) );
INVx1_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_269), .B(n_278), .Y(n_268) );
NAND2x1p5_ASAP7_75t_L g363 ( .A(n_269), .B(n_364), .Y(n_363) );
AND2x2_ASAP7_75t_L g415 ( .A(n_269), .B(n_330), .Y(n_415) );
AND2x2_ASAP7_75t_L g432 ( .A(n_269), .B(n_433), .Y(n_432) );
INVx4_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
AND2x4_ASAP7_75t_L g356 ( .A(n_270), .B(n_357), .Y(n_356) );
INVx1_ASAP7_75t_L g372 ( .A(n_270), .Y(n_372) );
AND2x2_ASAP7_75t_L g416 ( .A(n_270), .B(n_417), .Y(n_416) );
OR2x2_ASAP7_75t_L g423 ( .A(n_270), .B(n_424), .Y(n_423) );
NOR2x1_ASAP7_75t_L g438 ( .A(n_270), .B(n_329), .Y(n_438) );
BUFx2_ASAP7_75t_L g448 ( .A(n_270), .Y(n_448) );
AND2x2_ASAP7_75t_L g473 ( .A(n_270), .B(n_433), .Y(n_473) );
AND2x2_ASAP7_75t_L g494 ( .A(n_270), .B(n_495), .Y(n_494) );
OR2x6_ASAP7_75t_L g270 ( .A(n_271), .B(n_277), .Y(n_270) );
INVx1_ASAP7_75t_L g425 ( .A(n_278), .Y(n_425) );
NAND2xp5_ASAP7_75t_SL g371 ( .A(n_279), .B(n_372), .Y(n_371) );
AND2x2_ASAP7_75t_L g455 ( .A(n_279), .B(n_326), .Y(n_455) );
INVx3_ASAP7_75t_L g362 ( .A(n_280), .Y(n_362) );
AND2x2_ASAP7_75t_L g495 ( .A(n_280), .B(n_417), .Y(n_495) );
INVx1_ASAP7_75t_SL g281 ( .A(n_282), .Y(n_281) );
AOI22xp5_ASAP7_75t_L g324 ( .A1(n_282), .A2(n_325), .B1(n_330), .B2(n_331), .Y(n_324) );
AND2x2_ASAP7_75t_L g282 ( .A(n_283), .B(n_292), .Y(n_282) );
INVx4_ASAP7_75t_L g322 ( .A(n_283), .Y(n_322) );
INVx2_ASAP7_75t_L g359 ( .A(n_283), .Y(n_359) );
NAND2x1_ASAP7_75t_L g385 ( .A(n_283), .B(n_302), .Y(n_385) );
OR2x2_ASAP7_75t_L g400 ( .A(n_283), .B(n_335), .Y(n_400) );
OR2x2_ASAP7_75t_SL g427 ( .A(n_283), .B(n_399), .Y(n_427) );
AND2x2_ASAP7_75t_L g440 ( .A(n_283), .B(n_314), .Y(n_440) );
HB1xp67_ASAP7_75t_L g461 ( .A(n_283), .Y(n_461) );
OR2x6_ASAP7_75t_L g283 ( .A(n_284), .B(n_285), .Y(n_283) );
AOI21xp5_ASAP7_75t_L g285 ( .A1(n_286), .A2(n_287), .B(n_291), .Y(n_285) );
AOI21xp5_ASAP7_75t_L g315 ( .A1(n_291), .A2(n_316), .B(n_317), .Y(n_315) );
INVx2_ASAP7_75t_L g340 ( .A(n_292), .Y(n_340) );
AND2x2_ASAP7_75t_L g472 ( .A(n_292), .B(n_446), .Y(n_472) );
NOR2x1_ASAP7_75t_SL g292 ( .A(n_293), .B(n_302), .Y(n_292) );
AND2x2_ASAP7_75t_L g313 ( .A(n_293), .B(n_314), .Y(n_313) );
AND2x2_ASAP7_75t_L g489 ( .A(n_293), .B(n_412), .Y(n_489) );
AO21x1_ASAP7_75t_SL g293 ( .A1(n_294), .A2(n_295), .B(n_301), .Y(n_293) );
AO21x2_ASAP7_75t_L g336 ( .A1(n_294), .A2(n_295), .B(n_301), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_296), .B(n_300), .Y(n_295) );
OR2x2_ASAP7_75t_L g321 ( .A(n_302), .B(n_322), .Y(n_321) );
AND2x2_ASAP7_75t_L g332 ( .A(n_302), .B(n_322), .Y(n_332) );
AND2x2_ASAP7_75t_L g378 ( .A(n_302), .B(n_335), .Y(n_378) );
OR2x2_ASAP7_75t_L g399 ( .A(n_302), .B(n_314), .Y(n_399) );
INVx2_ASAP7_75t_SL g405 ( .A(n_302), .Y(n_405) );
AND2x2_ASAP7_75t_L g411 ( .A(n_302), .B(n_412), .Y(n_411) );
AND2x2_ASAP7_75t_L g421 ( .A(n_302), .B(n_404), .Y(n_421) );
BUFx2_ASAP7_75t_L g443 ( .A(n_302), .Y(n_443) );
OR2x6_ASAP7_75t_L g302 ( .A(n_303), .B(n_310), .Y(n_302) );
INVx2_ASAP7_75t_L g490 ( .A(n_311), .Y(n_490) );
OR2x2_ASAP7_75t_L g311 ( .A(n_312), .B(n_321), .Y(n_311) );
OR2x2_ASAP7_75t_L g515 ( .A(n_312), .B(n_359), .Y(n_515) );
INVx2_ASAP7_75t_SL g312 ( .A(n_313), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_313), .B(n_322), .Y(n_381) );
AND2x2_ASAP7_75t_L g452 ( .A(n_313), .B(n_332), .Y(n_452) );
INVx1_ASAP7_75t_L g334 ( .A(n_314), .Y(n_334) );
HB1xp67_ASAP7_75t_L g343 ( .A(n_314), .Y(n_343) );
INVx1_ASAP7_75t_L g376 ( .A(n_314), .Y(n_376) );
INVx2_ASAP7_75t_L g412 ( .A(n_314), .Y(n_412) );
NOR2xp67_ASAP7_75t_L g342 ( .A(n_322), .B(n_343), .Y(n_342) );
BUFx2_ASAP7_75t_L g402 ( .A(n_322), .Y(n_402) );
INVx2_ASAP7_75t_SL g478 ( .A(n_323), .Y(n_478) );
AOI22xp33_ASAP7_75t_L g379 ( .A1(n_325), .A2(n_380), .B1(n_382), .B2(n_386), .Y(n_379) );
AND2x2_ASAP7_75t_SL g325 ( .A(n_326), .B(n_327), .Y(n_325) );
AND2x2_ASAP7_75t_L g506 ( .A(n_326), .B(n_362), .Y(n_506) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
NOR2xp33_ASAP7_75t_L g451 ( .A(n_328), .B(n_372), .Y(n_451) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
AND2x2_ASAP7_75t_L g417 ( .A(n_329), .B(n_365), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_330), .B(n_467), .Y(n_466) );
INVx1_ASAP7_75t_L g360 ( .A(n_331), .Y(n_360) );
AOI221xp5_ASAP7_75t_L g474 ( .A1(n_331), .A2(n_475), .B1(n_479), .B2(n_481), .C(n_483), .Y(n_474) );
AND2x2_ASAP7_75t_L g331 ( .A(n_332), .B(n_333), .Y(n_331) );
AND2x2_ASAP7_75t_L g344 ( .A(n_332), .B(n_345), .Y(n_344) );
INVxp67_ASAP7_75t_SL g368 ( .A(n_332), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_332), .B(n_375), .Y(n_430) );
INVx1_ASAP7_75t_SL g426 ( .A(n_333), .Y(n_426) );
AOI221xp5_ASAP7_75t_SL g454 ( .A1(n_333), .A2(n_344), .B1(n_455), .B2(n_456), .C(n_459), .Y(n_454) );
AOI322xp5_ASAP7_75t_L g487 ( .A1(n_333), .A2(n_405), .A3(n_432), .B1(n_488), .B2(n_490), .C1(n_491), .C2(n_494), .Y(n_487) );
AND2x2_ASAP7_75t_L g333 ( .A(n_334), .B(n_335), .Y(n_333) );
BUFx2_ASAP7_75t_L g354 ( .A(n_334), .Y(n_354) );
HB1xp67_ASAP7_75t_L g346 ( .A(n_335), .Y(n_346) );
INVx2_ASAP7_75t_L g404 ( .A(n_335), .Y(n_404) );
AND2x2_ASAP7_75t_L g445 ( .A(n_335), .B(n_446), .Y(n_445) );
INVx3_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
OA21x2_ASAP7_75t_SL g337 ( .A1(n_338), .A2(n_344), .B(n_347), .Y(n_337) );
AOI211xp5_ASAP7_75t_L g507 ( .A1(n_338), .A2(n_508), .B(n_509), .C(n_513), .Y(n_507) );
INVx1_ASAP7_75t_SL g338 ( .A(n_339), .Y(n_338) );
OR2x2_ASAP7_75t_L g339 ( .A(n_340), .B(n_341), .Y(n_339) );
OR2x2_ASAP7_75t_L g396 ( .A(n_340), .B(n_358), .Y(n_396) );
OR2x2_ASAP7_75t_L g480 ( .A(n_340), .B(n_375), .Y(n_480) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
AND2x2_ASAP7_75t_L g420 ( .A(n_342), .B(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g498 ( .A(n_345), .Y(n_498) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
INVx1_ASAP7_75t_L g384 ( .A(n_346), .Y(n_384) );
INVx1_ASAP7_75t_SL g347 ( .A(n_348), .Y(n_347) );
OR2x2_ASAP7_75t_L g348 ( .A(n_349), .B(n_350), .Y(n_348) );
OR2x2_ASAP7_75t_L g353 ( .A(n_349), .B(n_354), .Y(n_353) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
AND2x2_ASAP7_75t_L g388 ( .A(n_351), .B(n_389), .Y(n_388) );
OAI322xp33_ASAP7_75t_L g352 ( .A1(n_353), .A2(n_355), .A3(n_358), .B1(n_360), .B2(n_361), .C1(n_366), .C2(n_368), .Y(n_352) );
INVx1_ASAP7_75t_L g394 ( .A(n_353), .Y(n_394) );
OR2x2_ASAP7_75t_L g366 ( .A(n_355), .B(n_367), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_355), .B(n_493), .Y(n_492) );
INVx2_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
INVx2_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
AND2x2_ASAP7_75t_L g377 ( .A(n_359), .B(n_378), .Y(n_377) );
OAI32xp33_ASAP7_75t_L g422 ( .A1(n_359), .A2(n_423), .A3(n_426), .B1(n_427), .B2(n_428), .Y(n_422) );
OR2x2_ASAP7_75t_L g361 ( .A(n_362), .B(n_363), .Y(n_361) );
INVx2_ASAP7_75t_L g367 ( .A(n_362), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_362), .B(n_425), .Y(n_424) );
NOR2x1_ASAP7_75t_L g464 ( .A(n_362), .B(n_465), .Y(n_464) );
AND2x2_ASAP7_75t_L g488 ( .A(n_362), .B(n_489), .Y(n_488) );
INVx1_ASAP7_75t_L g409 ( .A(n_363), .Y(n_409) );
INVx1_ASAP7_75t_SL g364 ( .A(n_365), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_367), .B(n_433), .Y(n_501) );
NOR2xp33_ASAP7_75t_L g369 ( .A(n_370), .B(n_390), .Y(n_369) );
OAI21xp33_ASAP7_75t_L g370 ( .A1(n_371), .A2(n_373), .B(n_379), .Y(n_370) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
AND2x4_ASAP7_75t_SL g374 ( .A(n_375), .B(n_377), .Y(n_374) );
INVx3_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
AND2x2_ASAP7_75t_L g439 ( .A(n_378), .B(n_440), .Y(n_439) );
INVx1_ASAP7_75t_SL g380 ( .A(n_381), .Y(n_380) );
OAI22xp5_ASAP7_75t_L g502 ( .A1(n_381), .A2(n_401), .B1(n_503), .B2(n_505), .Y(n_502) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
A2O1A1Ixp33_ASAP7_75t_L g429 ( .A1(n_383), .A2(n_430), .B(n_431), .C(n_434), .Y(n_429) );
OR2x2_ASAP7_75t_L g383 ( .A(n_384), .B(n_385), .Y(n_383) );
INVx3_ASAP7_75t_L g511 ( .A(n_385), .Y(n_511) );
INVx2_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
INVx2_ASAP7_75t_L g392 ( .A(n_389), .Y(n_392) );
AO21x1_ASAP7_75t_L g390 ( .A1(n_391), .A2(n_393), .B(n_397), .Y(n_390) );
HB1xp67_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
INVx2_ASAP7_75t_L g457 ( .A(n_392), .Y(n_457) );
AND2x2_ASAP7_75t_L g393 ( .A(n_394), .B(n_395), .Y(n_393) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
NOR2xp33_ASAP7_75t_L g483 ( .A(n_398), .B(n_484), .Y(n_483) );
OR2x2_ASAP7_75t_L g398 ( .A(n_399), .B(n_400), .Y(n_398) );
INVx1_ASAP7_75t_L g413 ( .A(n_400), .Y(n_413) );
OR2x2_ASAP7_75t_L g401 ( .A(n_402), .B(n_403), .Y(n_401) );
INVx1_ASAP7_75t_L g470 ( .A(n_403), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_404), .B(n_405), .Y(n_403) );
NOR3xp33_ASAP7_75t_L g406 ( .A(n_407), .B(n_429), .C(n_441), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_409), .B(n_410), .Y(n_408) );
OAI21xp5_ASAP7_75t_SL g471 ( .A1(n_410), .A2(n_472), .B(n_473), .Y(n_471) );
AND2x4_ASAP7_75t_L g410 ( .A(n_411), .B(n_413), .Y(n_410) );
INVx1_ASAP7_75t_L g446 ( .A(n_412), .Y(n_446) );
O2A1O1Ixp5_ASAP7_75t_SL g414 ( .A1(n_415), .A2(n_416), .B(n_418), .C(n_422), .Y(n_414) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx2_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
HB1xp67_ASAP7_75t_L g514 ( .A(n_424), .Y(n_514) );
INVx2_ASAP7_75t_L g499 ( .A(n_427), .Y(n_499) );
AOI21xp33_ASAP7_75t_L g513 ( .A1(n_428), .A2(n_514), .B(n_515), .Y(n_513) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g493 ( .A(n_433), .Y(n_493) );
OAI31xp33_ASAP7_75t_L g434 ( .A1(n_435), .A2(n_437), .A3(n_438), .B(n_439), .Y(n_434) );
INVx1_ASAP7_75t_SL g435 ( .A(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g512 ( .A(n_440), .Y(n_512) );
OAI21xp5_ASAP7_75t_L g441 ( .A1(n_442), .A2(n_447), .B(n_450), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_443), .B(n_444), .Y(n_442) );
BUFx2_ASAP7_75t_SL g444 ( .A(n_445), .Y(n_444) );
INVx1_ASAP7_75t_L g462 ( .A(n_445), .Y(n_462) );
AOI21xp33_ASAP7_75t_SL g509 ( .A1(n_447), .A2(n_510), .B(n_512), .Y(n_509) );
OR2x2_ASAP7_75t_L g447 ( .A(n_448), .B(n_449), .Y(n_447) );
INVx2_ASAP7_75t_L g477 ( .A(n_448), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_448), .B(n_468), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_448), .B(n_485), .Y(n_484) );
INVx2_ASAP7_75t_L g458 ( .A(n_449), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_451), .B(n_452), .Y(n_450) );
NAND5xp2_ASAP7_75t_L g453 ( .A(n_454), .B(n_474), .C(n_487), .D(n_496), .E(n_507), .Y(n_453) );
AND2x2_ASAP7_75t_L g456 ( .A(n_457), .B(n_458), .Y(n_456) );
OAI221xp5_ASAP7_75t_L g459 ( .A1(n_460), .A2(n_463), .B1(n_466), .B2(n_469), .C(n_471), .Y(n_459) );
OR2x2_ASAP7_75t_L g460 ( .A(n_461), .B(n_462), .Y(n_460) );
INVx1_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVxp67_ASAP7_75t_SL g467 ( .A(n_468), .Y(n_467) );
INVx1_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
INVxp67_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_477), .B(n_478), .Y(n_476) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx1_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
AOI21xp5_ASAP7_75t_L g496 ( .A1(n_497), .A2(n_500), .B(n_502), .Y(n_496) );
AND2x4_ASAP7_75t_L g497 ( .A(n_498), .B(n_499), .Y(n_497) );
INVx1_ASAP7_75t_SL g500 ( .A(n_501), .Y(n_500) );
INVx1_ASAP7_75t_SL g503 ( .A(n_504), .Y(n_503) );
INVxp67_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
INVx1_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
OAI222xp33_ASAP7_75t_L g517 ( .A1(n_518), .A2(n_520), .B1(n_525), .B2(n_527), .C1(n_530), .C2(n_534), .Y(n_517) );
HB1xp67_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
OR2x2_ASAP7_75t_L g521 ( .A(n_522), .B(n_523), .Y(n_521) );
CKINVDCx20_ASAP7_75t_R g527 ( .A(n_528), .Y(n_527) );
INVx2_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
CKINVDCx16_ASAP7_75t_R g530 ( .A(n_531), .Y(n_530) );
endmodule