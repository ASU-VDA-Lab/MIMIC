module fake_netlist_1_8700_n_25 (n_11, n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_25);
input n_11;
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_25;
wire n_20;
wire n_23;
wire n_22;
wire n_16;
wire n_13;
wire n_18;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
AND2x6_ASAP7_75t_L g12 ( .A(n_11), .B(n_6), .Y(n_12) );
INVx1_ASAP7_75t_L g13 ( .A(n_5), .Y(n_13) );
NAND2xp5_ASAP7_75t_L g14 ( .A(n_0), .B(n_10), .Y(n_14) );
INVx8_ASAP7_75t_L g15 ( .A(n_1), .Y(n_15) );
NAND2xp5_ASAP7_75t_SL g16 ( .A(n_3), .B(n_8), .Y(n_16) );
NAND2xp5_ASAP7_75t_L g17 ( .A(n_7), .B(n_9), .Y(n_17) );
HB1xp67_ASAP7_75t_L g18 ( .A(n_13), .Y(n_18) );
NAND2xp5_ASAP7_75t_L g19 ( .A(n_15), .B(n_2), .Y(n_19) );
INVx3_ASAP7_75t_L g20 ( .A(n_19), .Y(n_20) );
NAND2xp5_ASAP7_75t_L g21 ( .A(n_20), .B(n_18), .Y(n_21) );
AOI221xp5_ASAP7_75t_L g22 ( .A1(n_21), .A2(n_16), .B1(n_14), .B2(n_17), .C(n_12), .Y(n_22) );
NAND2x1p5_ASAP7_75t_L g23 ( .A(n_22), .B(n_12), .Y(n_23) );
HB1xp67_ASAP7_75t_L g24 ( .A(n_23), .Y(n_24) );
NOR2xp33_ASAP7_75t_SL g25 ( .A(n_24), .B(n_4), .Y(n_25) );
endmodule