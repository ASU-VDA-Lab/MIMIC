module fake_jpeg_2133_n_595 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_595);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_595;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_543;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_442;
wire n_299;
wire n_300;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx16f_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_9),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_12),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_7),
.Y(n_35)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

INVx1_ASAP7_75t_SL g37 ( 
.A(n_3),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_16),
.B(n_7),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_11),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_12),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

BUFx16f_ASAP7_75t_L g46 ( 
.A(n_11),
.Y(n_46)
);

BUFx16f_ASAP7_75t_L g47 ( 
.A(n_2),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_4),
.Y(n_48)
);

BUFx4f_ASAP7_75t_L g49 ( 
.A(n_13),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_3),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_16),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_11),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_11),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_7),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_1),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_4),
.Y(n_56)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_23),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_57),
.Y(n_135)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

BUFx2_ASAP7_75t_L g188 ( 
.A(n_58),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_23),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_59),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_23),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_60),
.Y(n_161)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_32),
.Y(n_61)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_61),
.Y(n_142)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_21),
.Y(n_62)
);

INVx4_ASAP7_75t_SL g209 ( 
.A(n_62),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_42),
.B(n_30),
.Y(n_63)
);

A2O1A1Ixp33_ASAP7_75t_L g179 ( 
.A1(n_63),
.A2(n_72),
.B(n_90),
.C(n_101),
.Y(n_179)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

BUFx2_ASAP7_75t_L g214 ( 
.A(n_64),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

INVx6_ASAP7_75t_L g171 ( 
.A(n_65),
.Y(n_171)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_32),
.Y(n_66)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_66),
.Y(n_143)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_27),
.Y(n_67)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_67),
.Y(n_128)
);

BUFx4f_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

INVx2_ASAP7_75t_SL g129 ( 
.A(n_68),
.Y(n_129)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_21),
.Y(n_69)
);

BUFx4f_ASAP7_75t_SL g174 ( 
.A(n_69),
.Y(n_174)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_27),
.Y(n_70)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_70),
.Y(n_148)
);

INVx3_ASAP7_75t_SL g71 ( 
.A(n_46),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_71),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_42),
.B(n_17),
.Y(n_72)
);

INVx6_ASAP7_75t_SL g73 ( 
.A(n_21),
.Y(n_73)
);

CKINVDCx6p67_ASAP7_75t_R g178 ( 
.A(n_73),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_38),
.Y(n_74)
);

INVx6_ASAP7_75t_L g173 ( 
.A(n_74),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_21),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_75),
.B(n_77),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_38),
.Y(n_76)
);

INVx6_ASAP7_75t_L g187 ( 
.A(n_76),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_51),
.B(n_17),
.Y(n_77)
);

BUFx5_ASAP7_75t_L g78 ( 
.A(n_46),
.Y(n_78)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_78),
.Y(n_130)
);

BUFx5_ASAP7_75t_L g79 ( 
.A(n_46),
.Y(n_79)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_79),
.Y(n_167)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_56),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g191 ( 
.A(n_80),
.Y(n_191)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_39),
.Y(n_81)
);

INVx5_ASAP7_75t_L g132 ( 
.A(n_81),
.Y(n_132)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_47),
.Y(n_82)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_82),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_47),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_83),
.B(n_111),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_43),
.Y(n_84)
);

INVx6_ASAP7_75t_L g192 ( 
.A(n_84),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_43),
.Y(n_85)
);

INVx3_ASAP7_75t_SL g144 ( 
.A(n_85),
.Y(n_144)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_19),
.Y(n_86)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_86),
.Y(n_137)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_39),
.Y(n_87)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_87),
.Y(n_138)
);

INVx11_ASAP7_75t_L g88 ( 
.A(n_39),
.Y(n_88)
);

INVx11_ASAP7_75t_L g134 ( 
.A(n_88),
.Y(n_134)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_19),
.Y(n_89)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_89),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_37),
.B(n_0),
.Y(n_90)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_36),
.Y(n_91)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_91),
.Y(n_170)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_56),
.Y(n_92)
);

INVx5_ASAP7_75t_L g140 ( 
.A(n_92),
.Y(n_140)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_49),
.Y(n_93)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_93),
.Y(n_160)
);

HB1xp67_ASAP7_75t_L g94 ( 
.A(n_47),
.Y(n_94)
);

INVx1_ASAP7_75t_SL g172 ( 
.A(n_94),
.Y(n_172)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_43),
.Y(n_95)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_95),
.Y(n_162)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_49),
.Y(n_96)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_96),
.Y(n_177)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_36),
.Y(n_97)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_97),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_54),
.Y(n_98)
);

INVx5_ASAP7_75t_L g181 ( 
.A(n_98),
.Y(n_181)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_54),
.Y(n_99)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_99),
.Y(n_180)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_47),
.Y(n_100)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_100),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_37),
.B(n_0),
.Y(n_101)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_54),
.Y(n_102)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_102),
.Y(n_183)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_56),
.Y(n_103)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_103),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_51),
.B(n_15),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_104),
.B(n_2),
.Y(n_153)
);

INVx11_ASAP7_75t_L g105 ( 
.A(n_52),
.Y(n_105)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_105),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_24),
.Y(n_106)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_106),
.Y(n_194)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_25),
.Y(n_107)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_107),
.Y(n_152)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_25),
.Y(n_108)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_108),
.Y(n_168)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_26),
.Y(n_109)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_109),
.Y(n_195)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_52),
.Y(n_110)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_110),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_29),
.B(n_0),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_22),
.B(n_1),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_112),
.B(n_120),
.Y(n_182)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_41),
.Y(n_113)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_113),
.Y(n_199)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_26),
.Y(n_114)
);

INVx4_ASAP7_75t_L g200 ( 
.A(n_114),
.Y(n_200)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_52),
.Y(n_115)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_115),
.Y(n_215)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_49),
.Y(n_116)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_116),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_24),
.Y(n_117)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_117),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_24),
.Y(n_118)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_118),
.Y(n_205)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_52),
.Y(n_119)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_119),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_29),
.B(n_1),
.Y(n_120)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_49),
.Y(n_121)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_121),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_33),
.Y(n_122)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_122),
.Y(n_220)
);

BUFx5_ASAP7_75t_L g123 ( 
.A(n_28),
.Y(n_123)
);

INVx4_ASAP7_75t_L g217 ( 
.A(n_123),
.Y(n_217)
);

BUFx8_ASAP7_75t_L g124 ( 
.A(n_28),
.Y(n_124)
);

BUFx5_ASAP7_75t_L g166 ( 
.A(n_124),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_33),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_125),
.B(n_64),
.Y(n_189)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_33),
.Y(n_126)
);

INVx1_ASAP7_75t_SL g201 ( 
.A(n_126),
.Y(n_201)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_41),
.Y(n_127)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_127),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_124),
.A2(n_120),
.B1(n_68),
.B2(n_114),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_131),
.A2(n_146),
.B1(n_164),
.B2(n_9),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_63),
.B(n_72),
.Y(n_133)
);

OR2x2_ASAP7_75t_L g250 ( 
.A(n_133),
.B(n_13),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_57),
.A2(n_50),
.B1(n_35),
.B2(n_34),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_141),
.A2(n_156),
.B1(n_184),
.B2(n_144),
.Y(n_291)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_109),
.A2(n_20),
.B1(n_53),
.B2(n_48),
.Y(n_146)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_94),
.Y(n_150)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_150),
.Y(n_223)
);

OR2x2_ASAP7_75t_L g151 ( 
.A(n_90),
.B(n_20),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_151),
.B(n_182),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_153),
.B(n_155),
.Y(n_233)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_71),
.Y(n_154)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_154),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_101),
.B(n_44),
.Y(n_155)
);

OAI22xp33_ASAP7_75t_L g156 ( 
.A1(n_95),
.A2(n_44),
.B1(n_53),
.B2(n_40),
.Y(n_156)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_119),
.Y(n_158)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_158),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_69),
.B(n_40),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_163),
.B(n_197),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_69),
.A2(n_45),
.B1(n_48),
.B2(n_50),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_106),
.Y(n_165)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_165),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_99),
.A2(n_55),
.B1(n_35),
.B2(n_34),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_102),
.A2(n_55),
.B1(n_31),
.B2(n_22),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_186),
.A2(n_198),
.B1(n_219),
.B2(n_8),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g234 ( 
.A(n_189),
.B(n_203),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_92),
.B(n_45),
.C(n_31),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_190),
.B(n_15),
.C(n_13),
.Y(n_251)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_117),
.Y(n_193)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_193),
.Y(n_246)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_118),
.Y(n_196)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_196),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_81),
.B(n_3),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_59),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_198)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_122),
.Y(n_206)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_206),
.Y(n_271)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_60),
.Y(n_207)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_207),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_87),
.B(n_5),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_210),
.B(n_211),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_65),
.B(n_5),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_74),
.B(n_5),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_213),
.B(n_216),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_76),
.B(n_6),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_84),
.B(n_8),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_218),
.B(n_12),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_85),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_219)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_160),
.Y(n_221)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_221),
.Y(n_332)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_132),
.Y(n_222)
);

BUFx2_ASAP7_75t_L g354 ( 
.A(n_222),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_182),
.A2(n_98),
.B1(n_110),
.B2(n_10),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g314 ( 
.A(n_224),
.B(n_251),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_L g333 ( 
.A1(n_225),
.A2(n_252),
.B1(n_288),
.B2(n_291),
.Y(n_333)
);

INVx6_ASAP7_75t_L g226 ( 
.A(n_157),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g300 ( 
.A(n_226),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_227),
.B(n_228),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_159),
.B(n_9),
.Y(n_228)
);

INVx6_ASAP7_75t_L g229 ( 
.A(n_157),
.Y(n_229)
);

INVx5_ASAP7_75t_L g324 ( 
.A(n_229),
.Y(n_324)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_161),
.Y(n_232)
);

INVx5_ASAP7_75t_L g350 ( 
.A(n_232),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_234),
.B(n_255),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_178),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_237),
.Y(n_351)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_161),
.Y(n_238)
);

INVx3_ASAP7_75t_L g312 ( 
.A(n_238),
.Y(n_312)
);

INVx3_ASAP7_75t_L g239 ( 
.A(n_138),
.Y(n_239)
);

INVx3_ASAP7_75t_L g326 ( 
.A(n_239),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_241),
.Y(n_306)
);

INVx3_ASAP7_75t_L g243 ( 
.A(n_172),
.Y(n_243)
);

INVx3_ASAP7_75t_L g337 ( 
.A(n_243),
.Y(n_337)
);

INVx8_ASAP7_75t_L g244 ( 
.A(n_178),
.Y(n_244)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_244),
.Y(n_342)
);

NOR2x1_ASAP7_75t_R g245 ( 
.A(n_176),
.B(n_12),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g320 ( 
.A(n_245),
.Y(n_320)
);

INVx4_ASAP7_75t_L g247 ( 
.A(n_129),
.Y(n_247)
);

INVx2_ASAP7_75t_SL g330 ( 
.A(n_247),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_248),
.B(n_250),
.Y(n_307)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_177),
.Y(n_249)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_249),
.Y(n_334)
);

AOI22xp33_ASAP7_75t_L g252 ( 
.A1(n_128),
.A2(n_144),
.B1(n_156),
.B2(n_181),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_202),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g355 ( 
.A(n_253),
.Y(n_355)
);

OAI21xp5_ASAP7_75t_SL g254 ( 
.A1(n_176),
.A2(n_14),
.B(n_159),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_254),
.B(n_250),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_137),
.B(n_14),
.Y(n_255)
);

BUFx4f_ASAP7_75t_SL g256 ( 
.A(n_178),
.Y(n_256)
);

CKINVDCx16_ASAP7_75t_R g319 ( 
.A(n_256),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_151),
.B(n_14),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_258),
.B(n_259),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_179),
.B(n_14),
.Y(n_259)
);

AND2x2_ASAP7_75t_L g260 ( 
.A(n_203),
.B(n_129),
.Y(n_260)
);

CKINVDCx16_ASAP7_75t_R g335 ( 
.A(n_260),
.Y(n_335)
);

BUFx12f_ASAP7_75t_L g261 ( 
.A(n_169),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_261),
.B(n_263),
.Y(n_341)
);

AOI22xp33_ASAP7_75t_SL g262 ( 
.A1(n_217),
.A2(n_152),
.B1(n_199),
.B2(n_168),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_SL g352 ( 
.A1(n_262),
.A2(n_281),
.B1(n_285),
.B2(n_292),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_139),
.B(n_197),
.Y(n_263)
);

INVx3_ASAP7_75t_L g264 ( 
.A(n_140),
.Y(n_264)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_264),
.Y(n_301)
);

BUFx3_ASAP7_75t_L g265 ( 
.A(n_130),
.Y(n_265)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_265),
.Y(n_305)
);

INVx4_ASAP7_75t_L g266 ( 
.A(n_170),
.Y(n_266)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_266),
.Y(n_310)
);

AND2x2_ASAP7_75t_L g267 ( 
.A(n_148),
.B(n_143),
.Y(n_267)
);

CKINVDCx16_ASAP7_75t_R g347 ( 
.A(n_267),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_189),
.B(n_147),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_268),
.A2(n_284),
.B1(n_297),
.B2(n_298),
.Y(n_343)
);

INVx6_ASAP7_75t_L g269 ( 
.A(n_135),
.Y(n_269)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_269),
.Y(n_311)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_131),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_270),
.Y(n_302)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_212),
.Y(n_272)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_272),
.Y(n_325)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_171),
.Y(n_273)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_273),
.Y(n_327)
);

INVx3_ASAP7_75t_L g274 ( 
.A(n_175),
.Y(n_274)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_274),
.Y(n_338)
);

AND2x2_ASAP7_75t_L g275 ( 
.A(n_142),
.B(n_145),
.Y(n_275)
);

AND2x2_ASAP7_75t_L g356 ( 
.A(n_275),
.B(n_279),
.Y(n_356)
);

INVx2_ASAP7_75t_SL g276 ( 
.A(n_214),
.Y(n_276)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_276),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_214),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_278),
.Y(n_303)
);

INVx1_ASAP7_75t_SL g279 ( 
.A(n_209),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_208),
.Y(n_280)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_280),
.Y(n_349)
);

INVx1_ASAP7_75t_SL g281 ( 
.A(n_209),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_136),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_282),
.Y(n_309)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_162),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_283),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_215),
.B(n_149),
.Y(n_284)
);

INVx4_ASAP7_75t_L g285 ( 
.A(n_167),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_210),
.B(n_180),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_286),
.B(n_293),
.Y(n_322)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_183),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_287),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_146),
.A2(n_164),
.B1(n_194),
.B2(n_204),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_188),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_289),
.Y(n_336)
);

HB1xp67_ASAP7_75t_L g290 ( 
.A(n_201),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_290),
.Y(n_353)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_205),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_220),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_135),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_294),
.B(n_295),
.Y(n_340)
);

BUFx12f_ASAP7_75t_L g295 ( 
.A(n_174),
.Y(n_295)
);

INVx13_ASAP7_75t_L g296 ( 
.A(n_174),
.Y(n_296)
);

NAND2x1_ASAP7_75t_L g318 ( 
.A(n_296),
.B(n_260),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_200),
.B(n_195),
.Y(n_297)
);

INVx1_ASAP7_75t_SL g298 ( 
.A(n_191),
.Y(n_298)
);

BUFx6f_ASAP7_75t_L g299 ( 
.A(n_171),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_299),
.B(n_238),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_270),
.A2(n_188),
.B1(n_191),
.B2(n_173),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g372 ( 
.A1(n_308),
.A2(n_323),
.B1(n_331),
.B2(n_256),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_241),
.A2(n_173),
.B1(n_187),
.B2(n_192),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_313),
.A2(n_316),
.B1(n_232),
.B2(n_247),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_252),
.A2(n_187),
.B1(n_192),
.B2(n_185),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_SL g317 ( 
.A1(n_235),
.A2(n_166),
.B(n_134),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_SL g361 ( 
.A1(n_317),
.A2(n_302),
.B(n_320),
.Y(n_361)
);

OR2x2_ASAP7_75t_L g400 ( 
.A(n_318),
.B(n_342),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_236),
.A2(n_242),
.B1(n_234),
.B2(n_251),
.Y(n_323)
);

AOI22xp33_ASAP7_75t_L g331 ( 
.A1(n_277),
.A2(n_257),
.B1(n_271),
.B2(n_246),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_233),
.B(n_267),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_339),
.B(n_346),
.C(n_266),
.Y(n_388)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_344),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_345),
.B(n_244),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_224),
.B(n_223),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_322),
.B(n_245),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_357),
.B(n_359),
.Y(n_405)
);

INVxp67_ASAP7_75t_L g358 ( 
.A(n_356),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_358),
.B(n_365),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_322),
.B(n_240),
.Y(n_359)
);

AOI21xp5_ASAP7_75t_L g360 ( 
.A1(n_306),
.A2(n_262),
.B(n_281),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_L g422 ( 
.A1(n_360),
.A2(n_362),
.B(n_381),
.Y(n_422)
);

OAI21xp33_ASAP7_75t_L g426 ( 
.A1(n_361),
.A2(n_370),
.B(n_376),
.Y(n_426)
);

AOI21xp5_ASAP7_75t_L g362 ( 
.A1(n_306),
.A2(n_279),
.B(n_298),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_314),
.A2(n_269),
.B1(n_299),
.B2(n_273),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g413 ( 
.A1(n_363),
.A2(n_399),
.B1(n_330),
.B2(n_319),
.Y(n_413)
);

INVxp67_ASAP7_75t_L g365 ( 
.A(n_356),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g366 ( 
.A(n_339),
.B(n_231),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_366),
.B(n_369),
.Y(n_414)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_348),
.Y(n_367)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_367),
.Y(n_402)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_348),
.Y(n_368)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_368),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_346),
.B(n_275),
.Y(n_369)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_301),
.Y(n_371)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_371),
.Y(n_415)
);

INVxp67_ASAP7_75t_L g411 ( 
.A(n_372),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_323),
.B(n_230),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_373),
.B(n_377),
.Y(n_419)
);

AND2x2_ASAP7_75t_L g374 ( 
.A(n_356),
.B(n_318),
.Y(n_374)
);

XNOR2x1_ASAP7_75t_SL g406 ( 
.A(n_374),
.B(n_378),
.Y(n_406)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_326),
.Y(n_375)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_375),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_304),
.B(n_256),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_314),
.B(n_222),
.Y(n_377)
);

AND2x2_ASAP7_75t_L g378 ( 
.A(n_318),
.B(n_239),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_326),
.Y(n_379)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_379),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_336),
.B(n_243),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_380),
.B(n_389),
.Y(n_432)
);

AOI21xp5_ASAP7_75t_L g381 ( 
.A1(n_314),
.A2(n_317),
.B(n_352),
.Y(n_381)
);

AND2x2_ASAP7_75t_L g382 ( 
.A(n_347),
.B(n_308),
.Y(n_382)
);

NAND2x1_ASAP7_75t_L g416 ( 
.A(n_382),
.B(n_400),
.Y(n_416)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_301),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_383),
.B(n_390),
.Y(n_404)
);

BUFx3_ASAP7_75t_L g384 ( 
.A(n_342),
.Y(n_384)
);

AOI22xp33_ASAP7_75t_SL g436 ( 
.A1(n_384),
.A2(n_386),
.B1(n_350),
.B2(n_337),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_SL g385 ( 
.A(n_345),
.B(n_274),
.Y(n_385)
);

XOR2xp5_ASAP7_75t_L g407 ( 
.A(n_385),
.B(n_388),
.Y(n_407)
);

AOI22xp33_ASAP7_75t_SL g386 ( 
.A1(n_313),
.A2(n_264),
.B1(n_295),
.B2(n_276),
.Y(n_386)
);

OAI21xp5_ASAP7_75t_SL g387 ( 
.A1(n_343),
.A2(n_296),
.B(n_295),
.Y(n_387)
);

INVxp67_ASAP7_75t_L g421 ( 
.A(n_387),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_341),
.B(n_261),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_325),
.Y(n_390)
);

OAI22xp33_ASAP7_75t_L g420 ( 
.A1(n_391),
.A2(n_315),
.B1(n_328),
.B2(n_324),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_L g392 ( 
.A1(n_333),
.A2(n_316),
.B1(n_320),
.B2(n_335),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_L g433 ( 
.A1(n_392),
.A2(n_395),
.B1(n_396),
.B2(n_310),
.Y(n_433)
);

INVxp67_ASAP7_75t_L g393 ( 
.A(n_329),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_393),
.B(n_398),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_353),
.B(n_285),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_394),
.B(n_397),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_344),
.A2(n_265),
.B1(n_229),
.B2(n_226),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_321),
.A2(n_261),
.B1(n_303),
.B2(n_307),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_325),
.Y(n_397)
);

INVxp67_ASAP7_75t_L g398 ( 
.A(n_343),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_311),
.A2(n_340),
.B1(n_309),
.B2(n_327),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_392),
.A2(n_311),
.B1(n_340),
.B2(n_327),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_L g437 ( 
.A1(n_401),
.A2(n_420),
.B1(n_391),
.B2(n_368),
.Y(n_437)
);

CKINVDCx16_ASAP7_75t_R g403 ( 
.A(n_380),
.Y(n_403)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_403),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_385),
.B(n_334),
.C(n_349),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_408),
.B(n_409),
.C(n_428),
.Y(n_451)
);

XOR2xp5_ASAP7_75t_L g409 ( 
.A(n_388),
.B(n_349),
.Y(n_409)
);

CKINVDCx16_ASAP7_75t_R g410 ( 
.A(n_394),
.Y(n_410)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_410),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_L g461 ( 
.A1(n_413),
.A2(n_429),
.B1(n_433),
.B2(n_395),
.Y(n_461)
);

OAI32xp33_ASAP7_75t_L g417 ( 
.A1(n_359),
.A2(n_338),
.A3(n_310),
.B1(n_330),
.B2(n_332),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_417),
.B(n_425),
.Y(n_440)
);

OA21x2_ASAP7_75t_L g425 ( 
.A1(n_382),
.A2(n_351),
.B(n_330),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_385),
.B(n_338),
.C(n_355),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_364),
.A2(n_312),
.B1(n_324),
.B2(n_354),
.Y(n_429)
);

OAI22x1_ASAP7_75t_L g430 ( 
.A1(n_382),
.A2(n_351),
.B1(n_354),
.B2(n_312),
.Y(n_430)
);

AOI22x1_ASAP7_75t_L g456 ( 
.A1(n_430),
.A2(n_422),
.B1(n_425),
.B2(n_401),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_399),
.Y(n_434)
);

INVxp67_ASAP7_75t_SL g465 ( 
.A(n_434),
.Y(n_465)
);

OA21x2_ASAP7_75t_L g435 ( 
.A1(n_382),
.A2(n_381),
.B(n_372),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_435),
.B(n_362),
.Y(n_457)
);

AOI22xp33_ASAP7_75t_SL g469 ( 
.A1(n_436),
.A2(n_378),
.B1(n_384),
.B2(n_375),
.Y(n_469)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_437),
.Y(n_471)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_404),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_441),
.B(n_448),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_404),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_SL g472 ( 
.A(n_442),
.B(n_447),
.Y(n_472)
);

XOR2xp5_ASAP7_75t_L g443 ( 
.A(n_407),
.B(n_409),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g482 ( 
.A(n_443),
.B(n_445),
.Y(n_482)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_412),
.Y(n_444)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_444),
.Y(n_479)
);

XNOR2xp5_ASAP7_75t_SL g445 ( 
.A(n_407),
.B(n_366),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_SL g446 ( 
.A1(n_411),
.A2(n_364),
.B1(n_373),
.B2(n_370),
.Y(n_446)
);

AOI22xp5_ASAP7_75t_L g485 ( 
.A1(n_446),
.A2(n_430),
.B1(n_423),
.B2(n_424),
.Y(n_485)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_427),
.Y(n_447)
);

OAI32xp33_ASAP7_75t_L g448 ( 
.A1(n_419),
.A2(n_369),
.A3(n_377),
.B1(n_357),
.B2(n_361),
.Y(n_448)
);

XOR2xp5_ASAP7_75t_L g449 ( 
.A(n_428),
.B(n_374),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_SL g490 ( 
.A(n_449),
.B(n_450),
.Y(n_490)
);

XNOR2xp5_ASAP7_75t_L g450 ( 
.A(n_414),
.B(n_408),
.Y(n_450)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_412),
.Y(n_452)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_452),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_SL g453 ( 
.A(n_403),
.B(n_396),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_SL g470 ( 
.A(n_453),
.B(n_459),
.Y(n_470)
);

XNOR2x1_ASAP7_75t_L g454 ( 
.A(n_406),
.B(n_416),
.Y(n_454)
);

AOI21xp5_ASAP7_75t_L g492 ( 
.A1(n_454),
.A2(n_456),
.B(n_416),
.Y(n_492)
);

XNOR2xp5_ASAP7_75t_L g455 ( 
.A(n_414),
.B(n_374),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_SL g497 ( 
.A(n_455),
.B(n_466),
.Y(n_497)
);

AOI22x1_ASAP7_75t_L g488 ( 
.A1(n_457),
.A2(n_416),
.B1(n_417),
.B2(n_402),
.Y(n_488)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_415),
.Y(n_458)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_458),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_432),
.B(n_376),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_415),
.Y(n_460)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_460),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_461),
.B(n_462),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_427),
.B(n_367),
.Y(n_462)
);

OAI21xp5_ASAP7_75t_SL g463 ( 
.A1(n_422),
.A2(n_387),
.B(n_360),
.Y(n_463)
);

OAI21xp5_ASAP7_75t_L g486 ( 
.A1(n_463),
.A2(n_469),
.B(n_400),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_432),
.B(n_389),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_SL g491 ( 
.A(n_464),
.B(n_402),
.Y(n_491)
);

CKINVDCx16_ASAP7_75t_R g466 ( 
.A(n_425),
.Y(n_466)
);

XOR2xp5_ASAP7_75t_L g467 ( 
.A(n_426),
.B(n_406),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_467),
.B(n_410),
.Y(n_474)
);

OAI22xp5_ASAP7_75t_L g468 ( 
.A1(n_434),
.A2(n_400),
.B1(n_378),
.B2(n_363),
.Y(n_468)
);

CKINVDCx14_ASAP7_75t_R g494 ( 
.A(n_468),
.Y(n_494)
);

XOR2xp5_ASAP7_75t_L g506 ( 
.A(n_474),
.B(n_467),
.Y(n_506)
);

OAI22xp5_ASAP7_75t_L g475 ( 
.A1(n_465),
.A2(n_435),
.B1(n_433),
.B2(n_425),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_L g516 ( 
.A1(n_475),
.A2(n_476),
.B1(n_478),
.B2(n_481),
.Y(n_516)
);

AOI22xp5_ASAP7_75t_SL g476 ( 
.A1(n_457),
.A2(n_421),
.B1(n_430),
.B2(n_435),
.Y(n_476)
);

CKINVDCx20_ASAP7_75t_R g477 ( 
.A(n_462),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_477),
.B(n_480),
.Y(n_501)
);

OAI22xp5_ASAP7_75t_L g478 ( 
.A1(n_456),
.A2(n_435),
.B1(n_413),
.B2(n_405),
.Y(n_478)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_440),
.Y(n_480)
);

OAI22xp5_ASAP7_75t_L g481 ( 
.A1(n_456),
.A2(n_405),
.B1(n_419),
.B2(n_429),
.Y(n_481)
);

INVx3_ASAP7_75t_L g484 ( 
.A(n_438),
.Y(n_484)
);

INVxp67_ASAP7_75t_L g512 ( 
.A(n_484),
.Y(n_512)
);

OAI22xp5_ASAP7_75t_SL g505 ( 
.A1(n_485),
.A2(n_498),
.B1(n_438),
.B2(n_439),
.Y(n_505)
);

AOI22xp5_ASAP7_75t_L g523 ( 
.A1(n_486),
.A2(n_379),
.B1(n_384),
.B2(n_305),
.Y(n_523)
);

CKINVDCx20_ASAP7_75t_R g487 ( 
.A(n_440),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_487),
.B(n_488),
.Y(n_507)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_491),
.Y(n_517)
);

AOI21xp33_ASAP7_75t_L g515 ( 
.A1(n_492),
.A2(n_448),
.B(n_458),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_441),
.B(n_431),
.Y(n_493)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_493),
.Y(n_519)
);

CKINVDCx16_ASAP7_75t_R g495 ( 
.A(n_446),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_SL g514 ( 
.A(n_495),
.B(n_463),
.Y(n_514)
);

AOI22xp5_ASAP7_75t_L g498 ( 
.A1(n_437),
.A2(n_431),
.B1(n_418),
.B2(n_397),
.Y(n_498)
);

XNOR2xp5_ASAP7_75t_L g500 ( 
.A(n_490),
.B(n_451),
.Y(n_500)
);

XOR2xp5_ASAP7_75t_L g527 ( 
.A(n_500),
.B(n_504),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_482),
.B(n_443),
.C(n_451),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g528 ( 
.A(n_502),
.B(n_503),
.C(n_511),
.Y(n_528)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_482),
.B(n_449),
.C(n_445),
.Y(n_503)
);

XNOR2xp5_ASAP7_75t_L g504 ( 
.A(n_483),
.B(n_450),
.Y(n_504)
);

AOI22xp5_ASAP7_75t_L g524 ( 
.A1(n_505),
.A2(n_522),
.B1(n_473),
.B2(n_475),
.Y(n_524)
);

XOR2xp5_ASAP7_75t_L g535 ( 
.A(n_506),
.B(n_509),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_470),
.B(n_472),
.Y(n_508)
);

CKINVDCx16_ASAP7_75t_R g538 ( 
.A(n_508),
.Y(n_538)
);

XNOR2xp5_ASAP7_75t_L g509 ( 
.A(n_483),
.B(n_455),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_470),
.B(n_439),
.Y(n_510)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_510),
.Y(n_526)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_497),
.B(n_454),
.C(n_452),
.Y(n_511)
);

INVxp67_ASAP7_75t_L g513 ( 
.A(n_484),
.Y(n_513)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_513),
.Y(n_529)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_514),
.Y(n_537)
);

XOR2xp5_ASAP7_75t_L g541 ( 
.A(n_515),
.B(n_518),
.Y(n_541)
);

XNOR2xp5_ASAP7_75t_SL g518 ( 
.A(n_492),
.B(n_460),
.Y(n_518)
);

CKINVDCx20_ASAP7_75t_R g520 ( 
.A(n_493),
.Y(n_520)
);

NOR3xp33_ASAP7_75t_L g536 ( 
.A(n_520),
.B(n_491),
.C(n_477),
.Y(n_536)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_494),
.B(n_444),
.C(n_371),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g534 ( 
.A(n_521),
.B(n_499),
.C(n_496),
.Y(n_534)
);

OAI22xp5_ASAP7_75t_SL g522 ( 
.A1(n_471),
.A2(n_418),
.B1(n_390),
.B2(n_383),
.Y(n_522)
);

OAI22xp5_ASAP7_75t_SL g525 ( 
.A1(n_523),
.A2(n_498),
.B1(n_471),
.B2(n_473),
.Y(n_525)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_524),
.Y(n_544)
);

AOI22xp5_ASAP7_75t_L g549 ( 
.A1(n_525),
.A2(n_532),
.B1(n_533),
.B2(n_481),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_504),
.B(n_517),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_SL g548 ( 
.A(n_530),
.B(n_531),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_521),
.B(n_509),
.Y(n_531)
);

AOI22xp5_ASAP7_75t_L g532 ( 
.A1(n_516),
.A2(n_489),
.B1(n_480),
.B2(n_487),
.Y(n_532)
);

OAI22xp5_ASAP7_75t_SL g533 ( 
.A1(n_519),
.A2(n_489),
.B1(n_476),
.B2(n_485),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_SL g545 ( 
.A(n_534),
.B(n_540),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_536),
.Y(n_546)
);

AND2x2_ASAP7_75t_L g539 ( 
.A(n_523),
.B(n_478),
.Y(n_539)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_539),
.Y(n_551)
);

MAJIxp5_ASAP7_75t_L g540 ( 
.A(n_500),
.B(n_486),
.C(n_488),
.Y(n_540)
);

MAJIxp5_ASAP7_75t_L g542 ( 
.A(n_527),
.B(n_528),
.C(n_502),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_SL g562 ( 
.A(n_542),
.B(n_543),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_538),
.B(n_505),
.Y(n_543)
);

MAJIxp5_ASAP7_75t_L g547 ( 
.A(n_527),
.B(n_503),
.C(n_511),
.Y(n_547)
);

AOI21xp5_ASAP7_75t_L g568 ( 
.A1(n_547),
.A2(n_479),
.B(n_305),
.Y(n_568)
);

OAI22xp5_ASAP7_75t_SL g558 ( 
.A1(n_549),
.A2(n_552),
.B1(n_554),
.B2(n_524),
.Y(n_558)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_534),
.Y(n_550)
);

AOI22xp5_ASAP7_75t_L g557 ( 
.A1(n_550),
.A2(n_553),
.B1(n_541),
.B2(n_537),
.Y(n_557)
);

AOI22xp5_ASAP7_75t_L g552 ( 
.A1(n_533),
.A2(n_507),
.B1(n_501),
.B2(n_522),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_529),
.Y(n_553)
);

AOI22xp5_ASAP7_75t_L g554 ( 
.A1(n_539),
.A2(n_507),
.B1(n_513),
.B2(n_512),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_SL g555 ( 
.A(n_526),
.B(n_512),
.Y(n_555)
);

CKINVDCx16_ASAP7_75t_R g569 ( 
.A(n_555),
.Y(n_569)
);

XNOR2xp5_ASAP7_75t_L g556 ( 
.A(n_541),
.B(n_528),
.Y(n_556)
);

XNOR2xp5_ASAP7_75t_L g559 ( 
.A(n_556),
.B(n_535),
.Y(n_559)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_557),
.Y(n_572)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_558),
.Y(n_576)
);

XNOR2xp5_ASAP7_75t_L g574 ( 
.A(n_559),
.B(n_560),
.Y(n_574)
);

XOR2xp5_ASAP7_75t_L g560 ( 
.A(n_549),
.B(n_535),
.Y(n_560)
);

AOI22xp5_ASAP7_75t_L g561 ( 
.A1(n_546),
.A2(n_525),
.B1(n_539),
.B2(n_532),
.Y(n_561)
);

HB1xp67_ASAP7_75t_L g575 ( 
.A(n_561),
.Y(n_575)
);

XOR2xp5_ASAP7_75t_L g563 ( 
.A(n_547),
.B(n_545),
.Y(n_563)
);

XOR2xp5_ASAP7_75t_L g570 ( 
.A(n_563),
.B(n_564),
.Y(n_570)
);

XOR2xp5_ASAP7_75t_L g564 ( 
.A(n_556),
.B(n_540),
.Y(n_564)
);

AOI22xp5_ASAP7_75t_SL g565 ( 
.A1(n_544),
.A2(n_518),
.B1(n_488),
.B2(n_506),
.Y(n_565)
);

MAJIxp5_ASAP7_75t_L g571 ( 
.A(n_565),
.B(n_552),
.C(n_551),
.Y(n_571)
);

XNOR2x1_ASAP7_75t_L g566 ( 
.A(n_554),
.B(n_499),
.Y(n_566)
);

NOR2xp33_ASAP7_75t_L g577 ( 
.A(n_566),
.B(n_567),
.Y(n_577)
);

XOR2xp5_ASAP7_75t_L g567 ( 
.A(n_544),
.B(n_496),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_L g578 ( 
.A(n_568),
.B(n_548),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_571),
.B(n_573),
.Y(n_580)
);

MAJIxp5_ASAP7_75t_L g573 ( 
.A(n_563),
.B(n_542),
.C(n_551),
.Y(n_573)
);

NOR2xp33_ASAP7_75t_L g581 ( 
.A(n_578),
.B(n_559),
.Y(n_581)
);

OAI21xp5_ASAP7_75t_L g579 ( 
.A1(n_572),
.A2(n_562),
.B(n_569),
.Y(n_579)
);

AOI21xp5_ASAP7_75t_L g587 ( 
.A1(n_579),
.A2(n_584),
.B(n_571),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_581),
.B(n_582),
.Y(n_586)
);

MAJIxp5_ASAP7_75t_L g582 ( 
.A(n_573),
.B(n_564),
.C(n_560),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_L g583 ( 
.A(n_575),
.B(n_567),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_583),
.B(n_574),
.Y(n_588)
);

OAI21xp5_ASAP7_75t_L g584 ( 
.A1(n_570),
.A2(n_565),
.B(n_566),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_SL g585 ( 
.A(n_580),
.B(n_576),
.Y(n_585)
);

OAI21x1_ASAP7_75t_SL g590 ( 
.A1(n_585),
.A2(n_587),
.B(n_588),
.Y(n_590)
);

INVxp67_ASAP7_75t_L g589 ( 
.A(n_586),
.Y(n_589)
);

NAND3xp33_ASAP7_75t_L g591 ( 
.A(n_589),
.B(n_577),
.C(n_570),
.Y(n_591)
);

MAJx2_ASAP7_75t_L g592 ( 
.A(n_591),
.B(n_590),
.C(n_479),
.Y(n_592)
);

AOI21xp5_ASAP7_75t_L g593 ( 
.A1(n_592),
.A2(n_337),
.B(n_355),
.Y(n_593)
);

MAJIxp5_ASAP7_75t_L g594 ( 
.A(n_593),
.B(n_300),
.C(n_332),
.Y(n_594)
);

AOI21xp5_ASAP7_75t_L g595 ( 
.A1(n_594),
.A2(n_350),
.B(n_300),
.Y(n_595)
);


endmodule