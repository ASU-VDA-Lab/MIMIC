module fake_ibex_532_n_2657 (n_151, n_85, n_395, n_84, n_64, n_171, n_103, n_389, n_204, n_274, n_387, n_130, n_177, n_76, n_273, n_309, n_330, n_9, n_328, n_293, n_341, n_372, n_124, n_37, n_256, n_418, n_193, n_446, n_108, n_350, n_165, n_452, n_86, n_70, n_255, n_175, n_398, n_59, n_28, n_125, n_304, n_191, n_5, n_62, n_71, n_153, n_194, n_249, n_334, n_312, n_478, n_239, n_94, n_134, n_432, n_371, n_403, n_423, n_357, n_88, n_412, n_457, n_142, n_226, n_336, n_258, n_40, n_90, n_17, n_74, n_449, n_176, n_58, n_43, n_216, n_33, n_421, n_475, n_166, n_163, n_114, n_236, n_34, n_376, n_377, n_15, n_24, n_189, n_280, n_317, n_340, n_375, n_105, n_187, n_1, n_154, n_182, n_196, n_326, n_327, n_89, n_50, n_144, n_170, n_270, n_346, n_383, n_113, n_117, n_417, n_471, n_265, n_158, n_259, n_276, n_339, n_470, n_210, n_348, n_220, n_91, n_481, n_287, n_54, n_243, n_19, n_228, n_147, n_251, n_384, n_373, n_458, n_244, n_73, n_343, n_310, n_426, n_323, n_469, n_143, n_106, n_386, n_8, n_224, n_183, n_67, n_453, n_333, n_110, n_306, n_400, n_47, n_169, n_10, n_21, n_242, n_278, n_316, n_16, n_404, n_60, n_7, n_109, n_127, n_121, n_465, n_48, n_325, n_57, n_301, n_434, n_296, n_120, n_168, n_155, n_315, n_441, n_13, n_122, n_116, n_370, n_431, n_0, n_289, n_12, n_150, n_286, n_321, n_133, n_51, n_215, n_279, n_49, n_374, n_235, n_464, n_22, n_136, n_261, n_459, n_30, n_367, n_221, n_437, n_355, n_474, n_407, n_102, n_52, n_448, n_99, n_466, n_269, n_156, n_126, n_356, n_25, n_104, n_45, n_420, n_141, n_222, n_186, n_349, n_454, n_295, n_331, n_230, n_96, n_185, n_388, n_352, n_290, n_174, n_467, n_427, n_157, n_219, n_246, n_31, n_442, n_146, n_207, n_438, n_167, n_128, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_358, n_205, n_139, n_429, n_275, n_98, n_129, n_267, n_245, n_229, n_209, n_472, n_347, n_473, n_445, n_335, n_413, n_82, n_263, n_27, n_353, n_359, n_299, n_87, n_262, n_433, n_75, n_439, n_137, n_338, n_173, n_477, n_363, n_402, n_180, n_369, n_201, n_14, n_351, n_368, n_456, n_257, n_77, n_44, n_401, n_66, n_305, n_307, n_192, n_140, n_480, n_416, n_365, n_4, n_6, n_100, n_179, n_354, n_206, n_392, n_329, n_447, n_26, n_188, n_200, n_444, n_199, n_410, n_308, n_463, n_411, n_135, n_283, n_366, n_397, n_111, n_36, n_18, n_322, n_53, n_227, n_115, n_11, n_248, n_92, n_451, n_101, n_190, n_138, n_409, n_214, n_238, n_332, n_211, n_218, n_314, n_132, n_277, n_337, n_479, n_225, n_360, n_272, n_23, n_468, n_223, n_381, n_382, n_95, n_405, n_415, n_285, n_288, n_247, n_320, n_379, n_55, n_291, n_318, n_63, n_161, n_237, n_29, n_203, n_268, n_440, n_148, n_2, n_342, n_233, n_385, n_414, n_430, n_118, n_378, n_422, n_164, n_38, n_198, n_264, n_217, n_324, n_391, n_78, n_20, n_69, n_390, n_39, n_178, n_303, n_362, n_93, n_162, n_240, n_282, n_61, n_266, n_42, n_294, n_112, n_46, n_284, n_80, n_172, n_250, n_460, n_476, n_461, n_313, n_345, n_408, n_119, n_361, n_455, n_419, n_72, n_319, n_195, n_212, n_311, n_406, n_97, n_197, n_181, n_131, n_123, n_260, n_462, n_302, n_450, n_443, n_344, n_393, n_436, n_428, n_297, n_435, n_41, n_252, n_396, n_83, n_32, n_107, n_149, n_399, n_254, n_213, n_424, n_271, n_241, n_68, n_292, n_394, n_79, n_81, n_35, n_364, n_159, n_202, n_231, n_298, n_160, n_184, n_56, n_232, n_380, n_281, n_425, n_2657);

input n_151;
input n_85;
input n_395;
input n_84;
input n_64;
input n_171;
input n_103;
input n_389;
input n_204;
input n_274;
input n_387;
input n_130;
input n_177;
input n_76;
input n_273;
input n_309;
input n_330;
input n_9;
input n_328;
input n_293;
input n_341;
input n_372;
input n_124;
input n_37;
input n_256;
input n_418;
input n_193;
input n_446;
input n_108;
input n_350;
input n_165;
input n_452;
input n_86;
input n_70;
input n_255;
input n_175;
input n_398;
input n_59;
input n_28;
input n_125;
input n_304;
input n_191;
input n_5;
input n_62;
input n_71;
input n_153;
input n_194;
input n_249;
input n_334;
input n_312;
input n_478;
input n_239;
input n_94;
input n_134;
input n_432;
input n_371;
input n_403;
input n_423;
input n_357;
input n_88;
input n_412;
input n_457;
input n_142;
input n_226;
input n_336;
input n_258;
input n_40;
input n_90;
input n_17;
input n_74;
input n_449;
input n_176;
input n_58;
input n_43;
input n_216;
input n_33;
input n_421;
input n_475;
input n_166;
input n_163;
input n_114;
input n_236;
input n_34;
input n_376;
input n_377;
input n_15;
input n_24;
input n_189;
input n_280;
input n_317;
input n_340;
input n_375;
input n_105;
input n_187;
input n_1;
input n_154;
input n_182;
input n_196;
input n_326;
input n_327;
input n_89;
input n_50;
input n_144;
input n_170;
input n_270;
input n_346;
input n_383;
input n_113;
input n_117;
input n_417;
input n_471;
input n_265;
input n_158;
input n_259;
input n_276;
input n_339;
input n_470;
input n_210;
input n_348;
input n_220;
input n_91;
input n_481;
input n_287;
input n_54;
input n_243;
input n_19;
input n_228;
input n_147;
input n_251;
input n_384;
input n_373;
input n_458;
input n_244;
input n_73;
input n_343;
input n_310;
input n_426;
input n_323;
input n_469;
input n_143;
input n_106;
input n_386;
input n_8;
input n_224;
input n_183;
input n_67;
input n_453;
input n_333;
input n_110;
input n_306;
input n_400;
input n_47;
input n_169;
input n_10;
input n_21;
input n_242;
input n_278;
input n_316;
input n_16;
input n_404;
input n_60;
input n_7;
input n_109;
input n_127;
input n_121;
input n_465;
input n_48;
input n_325;
input n_57;
input n_301;
input n_434;
input n_296;
input n_120;
input n_168;
input n_155;
input n_315;
input n_441;
input n_13;
input n_122;
input n_116;
input n_370;
input n_431;
input n_0;
input n_289;
input n_12;
input n_150;
input n_286;
input n_321;
input n_133;
input n_51;
input n_215;
input n_279;
input n_49;
input n_374;
input n_235;
input n_464;
input n_22;
input n_136;
input n_261;
input n_459;
input n_30;
input n_367;
input n_221;
input n_437;
input n_355;
input n_474;
input n_407;
input n_102;
input n_52;
input n_448;
input n_99;
input n_466;
input n_269;
input n_156;
input n_126;
input n_356;
input n_25;
input n_104;
input n_45;
input n_420;
input n_141;
input n_222;
input n_186;
input n_349;
input n_454;
input n_295;
input n_331;
input n_230;
input n_96;
input n_185;
input n_388;
input n_352;
input n_290;
input n_174;
input n_467;
input n_427;
input n_157;
input n_219;
input n_246;
input n_31;
input n_442;
input n_146;
input n_207;
input n_438;
input n_167;
input n_128;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_358;
input n_205;
input n_139;
input n_429;
input n_275;
input n_98;
input n_129;
input n_267;
input n_245;
input n_229;
input n_209;
input n_472;
input n_347;
input n_473;
input n_445;
input n_335;
input n_413;
input n_82;
input n_263;
input n_27;
input n_353;
input n_359;
input n_299;
input n_87;
input n_262;
input n_433;
input n_75;
input n_439;
input n_137;
input n_338;
input n_173;
input n_477;
input n_363;
input n_402;
input n_180;
input n_369;
input n_201;
input n_14;
input n_351;
input n_368;
input n_456;
input n_257;
input n_77;
input n_44;
input n_401;
input n_66;
input n_305;
input n_307;
input n_192;
input n_140;
input n_480;
input n_416;
input n_365;
input n_4;
input n_6;
input n_100;
input n_179;
input n_354;
input n_206;
input n_392;
input n_329;
input n_447;
input n_26;
input n_188;
input n_200;
input n_444;
input n_199;
input n_410;
input n_308;
input n_463;
input n_411;
input n_135;
input n_283;
input n_366;
input n_397;
input n_111;
input n_36;
input n_18;
input n_322;
input n_53;
input n_227;
input n_115;
input n_11;
input n_248;
input n_92;
input n_451;
input n_101;
input n_190;
input n_138;
input n_409;
input n_214;
input n_238;
input n_332;
input n_211;
input n_218;
input n_314;
input n_132;
input n_277;
input n_337;
input n_479;
input n_225;
input n_360;
input n_272;
input n_23;
input n_468;
input n_223;
input n_381;
input n_382;
input n_95;
input n_405;
input n_415;
input n_285;
input n_288;
input n_247;
input n_320;
input n_379;
input n_55;
input n_291;
input n_318;
input n_63;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_440;
input n_148;
input n_2;
input n_342;
input n_233;
input n_385;
input n_414;
input n_430;
input n_118;
input n_378;
input n_422;
input n_164;
input n_38;
input n_198;
input n_264;
input n_217;
input n_324;
input n_391;
input n_78;
input n_20;
input n_69;
input n_390;
input n_39;
input n_178;
input n_303;
input n_362;
input n_93;
input n_162;
input n_240;
input n_282;
input n_61;
input n_266;
input n_42;
input n_294;
input n_112;
input n_46;
input n_284;
input n_80;
input n_172;
input n_250;
input n_460;
input n_476;
input n_461;
input n_313;
input n_345;
input n_408;
input n_119;
input n_361;
input n_455;
input n_419;
input n_72;
input n_319;
input n_195;
input n_212;
input n_311;
input n_406;
input n_97;
input n_197;
input n_181;
input n_131;
input n_123;
input n_260;
input n_462;
input n_302;
input n_450;
input n_443;
input n_344;
input n_393;
input n_436;
input n_428;
input n_297;
input n_435;
input n_41;
input n_252;
input n_396;
input n_83;
input n_32;
input n_107;
input n_149;
input n_399;
input n_254;
input n_213;
input n_424;
input n_271;
input n_241;
input n_68;
input n_292;
input n_394;
input n_79;
input n_81;
input n_35;
input n_364;
input n_159;
input n_202;
input n_231;
input n_298;
input n_160;
input n_184;
input n_56;
input n_232;
input n_380;
input n_281;
input n_425;

output n_2657;

wire n_1084;
wire n_2594;
wire n_1474;
wire n_1295;
wire n_507;
wire n_1983;
wire n_992;
wire n_1582;
wire n_2201;
wire n_2512;
wire n_766;
wire n_2175;
wire n_2071;
wire n_1110;
wire n_2607;
wire n_1382;
wire n_2569;
wire n_1998;
wire n_1596;
wire n_926;
wire n_1079;
wire n_1100;
wire n_845;
wire n_2177;
wire n_1930;
wire n_2123;
wire n_1234;
wire n_2047;
wire n_1594;
wire n_1944;
wire n_2235;
wire n_1802;
wire n_2498;
wire n_773;
wire n_2038;
wire n_2504;
wire n_1469;
wire n_821;
wire n_2017;
wire n_873;
wire n_1227;
wire n_962;
wire n_1080;
wire n_909;
wire n_862;
wire n_2290;
wire n_957;
wire n_1652;
wire n_678;
wire n_969;
wire n_1859;
wire n_1954;
wire n_2183;
wire n_2074;
wire n_1883;
wire n_1125;
wire n_733;
wire n_2037;
wire n_622;
wire n_1226;
wire n_1034;
wire n_2383;
wire n_1765;
wire n_872;
wire n_2392;
wire n_1873;
wire n_1619;
wire n_1666;
wire n_2640;
wire n_494;
wire n_930;
wire n_1044;
wire n_1492;
wire n_1134;
wire n_1478;
wire n_1684;
wire n_1796;
wire n_1614;
wire n_2374;
wire n_2598;
wire n_1722;
wire n_911;
wire n_2023;
wire n_652;
wire n_781;
wire n_802;
wire n_2322;
wire n_1233;
wire n_2335;
wire n_2276;
wire n_1045;
wire n_1856;
wire n_500;
wire n_963;
wire n_1782;
wire n_2230;
wire n_2139;
wire n_531;
wire n_1308;
wire n_556;
wire n_1138;
wire n_498;
wire n_708;
wire n_1096;
wire n_2151;
wire n_2391;
wire n_1391;
wire n_884;
wire n_667;
wire n_2396;
wire n_850;
wire n_1971;
wire n_2485;
wire n_2479;
wire n_879;
wire n_2179;
wire n_1957;
wire n_2188;
wire n_723;
wire n_1144;
wire n_2359;
wire n_2360;
wire n_2506;
wire n_1392;
wire n_2158;
wire n_1268;
wire n_2571;
wire n_739;
wire n_2475;
wire n_853;
wire n_504;
wire n_948;
wire n_1752;
wire n_1829;
wire n_1338;
wire n_1730;
wire n_875;
wire n_1307;
wire n_1327;
wire n_2644;
wire n_876;
wire n_497;
wire n_711;
wire n_1840;
wire n_671;
wire n_989;
wire n_1908;
wire n_1668;
wire n_2343;
wire n_2605;
wire n_1641;
wire n_829;
wire n_2565;
wire n_825;
wire n_1480;
wire n_1463;
wire n_1823;
wire n_1681;
wire n_939;
wire n_1636;
wire n_1687;
wire n_655;
wire n_2192;
wire n_1766;
wire n_550;
wire n_1922;
wire n_2032;
wire n_641;
wire n_557;
wire n_1937;
wire n_2311;
wire n_893;
wire n_527;
wire n_1654;
wire n_496;
wire n_1258;
wire n_1344;
wire n_2208;
wire n_2198;
wire n_1929;
wire n_1749;
wire n_1680;
wire n_835;
wire n_1981;
wire n_1195;
wire n_824;
wire n_1945;
wire n_2638;
wire n_694;
wire n_523;
wire n_787;
wire n_2448;
wire n_614;
wire n_2015;
wire n_2537;
wire n_1130;
wire n_2643;
wire n_1228;
wire n_2336;
wire n_2163;
wire n_1081;
wire n_538;
wire n_2354;
wire n_1155;
wire n_1292;
wire n_2432;
wire n_1576;
wire n_1664;
wire n_2273;
wire n_518;
wire n_852;
wire n_1427;
wire n_1133;
wire n_2421;
wire n_1926;
wire n_904;
wire n_2363;
wire n_2003;
wire n_1970;
wire n_2621;
wire n_1778;
wire n_646;
wire n_2558;
wire n_2347;
wire n_1030;
wire n_1698;
wire n_1094;
wire n_2462;
wire n_1496;
wire n_1910;
wire n_715;
wire n_2333;
wire n_530;
wire n_1663;
wire n_2436;
wire n_1214;
wire n_1274;
wire n_2527;
wire n_1606;
wire n_769;
wire n_1595;
wire n_2164;
wire n_1509;
wire n_1618;
wire n_1648;
wire n_1886;
wire n_2269;
wire n_857;
wire n_765;
wire n_1070;
wire n_1841;
wire n_2472;
wire n_777;
wire n_1955;
wire n_917;
wire n_2249;
wire n_2413;
wire n_2362;
wire n_968;
wire n_1253;
wire n_1306;
wire n_1484;
wire n_1493;
wire n_2597;
wire n_1313;
wire n_558;
wire n_2090;
wire n_666;
wire n_2260;
wire n_1638;
wire n_2215;
wire n_1071;
wire n_1449;
wire n_1723;
wire n_1960;
wire n_793;
wire n_937;
wire n_2595;
wire n_2116;
wire n_1645;
wire n_973;
wire n_1038;
wire n_2280;
wire n_618;
wire n_1943;
wire n_1863;
wire n_1269;
wire n_2393;
wire n_662;
wire n_979;
wire n_1309;
wire n_1999;
wire n_1316;
wire n_1562;
wire n_1215;
wire n_629;
wire n_2480;
wire n_1445;
wire n_573;
wire n_2283;
wire n_2147;
wire n_1716;
wire n_1466;
wire n_1412;
wire n_1672;
wire n_1007;
wire n_2253;
wire n_643;
wire n_1276;
wire n_1637;
wire n_841;
wire n_772;
wire n_810;
wire n_1401;
wire n_1817;
wire n_2145;
wire n_2122;
wire n_1588;
wire n_2216;
wire n_1301;
wire n_2579;
wire n_2242;
wire n_869;
wire n_1620;
wire n_1561;
wire n_718;
wire n_2370;
wire n_553;
wire n_554;
wire n_2025;
wire n_1078;
wire n_2247;
wire n_1219;
wire n_713;
wire n_1865;
wire n_1252;
wire n_2022;
wire n_1170;
wire n_1927;
wire n_605;
wire n_539;
wire n_2373;
wire n_630;
wire n_1869;
wire n_567;
wire n_1853;
wire n_2275;
wire n_2189;
wire n_2482;
wire n_745;
wire n_2112;
wire n_1753;
wire n_562;
wire n_564;
wire n_1322;
wire n_2008;
wire n_1305;
wire n_2088;
wire n_795;
wire n_592;
wire n_1248;
wire n_2171;
wire n_762;
wire n_1388;
wire n_800;
wire n_2564;
wire n_706;
wire n_784;
wire n_684;
wire n_1653;
wire n_1375;
wire n_1356;
wire n_894;
wire n_1118;
wire n_692;
wire n_2591;
wire n_1881;
wire n_1969;
wire n_709;
wire n_1296;
wire n_499;
wire n_971;
wire n_1326;
wire n_702;
wire n_1350;
wire n_906;
wire n_2586;
wire n_1093;
wire n_1764;
wire n_2412;
wire n_978;
wire n_899;
wire n_579;
wire n_1799;
wire n_1019;
wire n_902;
wire n_1689;
wire n_1250;
wire n_2550;
wire n_1190;
wire n_1304;
wire n_744;
wire n_563;
wire n_2541;
wire n_1506;
wire n_881;
wire n_1702;
wire n_734;
wire n_1558;
wire n_1650;
wire n_1520;
wire n_1073;
wire n_1453;
wire n_1108;
wire n_2509;
wire n_1794;
wire n_1423;
wire n_1239;
wire n_2399;
wire n_1370;
wire n_1209;
wire n_1708;
wire n_2213;
wire n_551;
wire n_1616;
wire n_729;
wire n_1569;
wire n_1434;
wire n_603;
wire n_1649;
wire n_2389;
wire n_1936;
wire n_2114;
wire n_1717;
wire n_2107;
wire n_1609;
wire n_2257;
wire n_1613;
wire n_820;
wire n_805;
wire n_1988;
wire n_670;
wire n_1132;
wire n_892;
wire n_1467;
wire n_1803;
wire n_544;
wire n_2401;
wire n_1787;
wire n_2511;
wire n_1281;
wire n_1447;
wire n_2166;
wire n_2451;
wire n_2150;
wire n_695;
wire n_1549;
wire n_639;
wire n_2631;
wire n_1867;
wire n_1531;
wire n_1332;
wire n_482;
wire n_2292;
wire n_2334;
wire n_1424;
wire n_2444;
wire n_2625;
wire n_1742;
wire n_2350;
wire n_1818;
wire n_870;
wire n_2199;
wire n_1709;
wire n_1610;
wire n_2219;
wire n_1298;
wire n_1844;
wire n_1387;
wire n_2649;
wire n_609;
wire n_1040;
wire n_2203;
wire n_1159;
wire n_1368;
wire n_2281;
wire n_1154;
wire n_2539;
wire n_2431;
wire n_1701;
wire n_2084;
wire n_1243;
wire n_2387;
wire n_2646;
wire n_2397;
wire n_1121;
wire n_693;
wire n_2256;
wire n_606;
wire n_737;
wire n_2445;
wire n_1571;
wire n_1980;
wire n_2529;
wire n_2019;
wire n_1407;
wire n_1235;
wire n_1821;
wire n_1003;
wire n_889;
wire n_816;
wire n_1058;
wire n_1835;
wire n_1862;
wire n_2224;
wire n_2470;
wire n_2355;
wire n_1543;
wire n_823;
wire n_2233;
wire n_2499;
wire n_1504;
wire n_1519;
wire n_1425;
wire n_1781;
wire n_2069;
wire n_2602;
wire n_1441;
wire n_2028;
wire n_1924;
wire n_1921;
wire n_657;
wire n_1156;
wire n_1293;
wire n_1360;
wire n_749;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_819;
wire n_2070;
wire n_822;
wire n_1042;
wire n_1888;
wire n_743;
wire n_754;
wire n_1786;
wire n_2033;
wire n_1319;
wire n_1553;
wire n_1041;
wire n_1964;
wire n_1090;
wire n_1196;
wire n_1182;
wire n_1271;
wire n_2416;
wire n_1731;
wire n_1905;
wire n_1031;
wire n_2052;
wire n_981;
wire n_2425;
wire n_2118;
wire n_2259;
wire n_2162;
wire n_2236;
wire n_2377;
wire n_2577;
wire n_1591;
wire n_583;
wire n_2289;
wire n_2288;
wire n_1671;
wire n_1795;
wire n_1409;
wire n_1015;
wire n_663;
wire n_2101;
wire n_1377;
wire n_2473;
wire n_1583;
wire n_1521;
wire n_2632;
wire n_1152;
wire n_2456;
wire n_2264;
wire n_2076;
wire n_974;
wire n_1036;
wire n_2599;
wire n_1831;
wire n_864;
wire n_608;
wire n_1987;
wire n_959;
wire n_1106;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_1733;
wire n_1634;
wire n_1932;
wire n_1552;
wire n_1452;
wire n_1318;
wire n_1508;
wire n_2217;
wire n_738;
wire n_1217;
wire n_2655;
wire n_2454;
wire n_1715;
wire n_1189;
wire n_761;
wire n_748;
wire n_1713;
wire n_901;
wire n_1577;
wire n_2036;
wire n_1255;
wire n_1700;
wire n_2623;
wire n_2622;
wire n_1218;
wire n_2178;
wire n_1181;
wire n_1140;
wire n_1985;
wire n_1772;
wire n_1056;
wire n_2626;
wire n_1283;
wire n_1446;
wire n_2404;
wire n_1487;
wire n_2603;
wire n_840;
wire n_1203;
wire n_1421;
wire n_561;
wire n_2573;
wire n_846;
wire n_1793;
wire n_1237;
wire n_2424;
wire n_2390;
wire n_2423;
wire n_859;
wire n_1109;
wire n_965;
wire n_1633;
wire n_2580;
wire n_1711;
wire n_1051;
wire n_1008;
wire n_2375;
wire n_1498;
wire n_2312;
wire n_2572;
wire n_1053;
wire n_1656;
wire n_1207;
wire n_1076;
wire n_1735;
wire n_2063;
wire n_1032;
wire n_936;
wire n_1884;
wire n_2176;
wire n_1825;
wire n_1589;
wire n_2204;
wire n_2575;
wire n_1210;
wire n_2319;
wire n_591;
wire n_1933;
wire n_2522;
wire n_1996;
wire n_1510;
wire n_1201;
wire n_1842;
wire n_2132;
wire n_1246;
wire n_1677;
wire n_732;
wire n_1236;
wire n_832;
wire n_2297;
wire n_1792;
wire n_1712;
wire n_1984;
wire n_590;
wire n_1568;
wire n_1877;
wire n_1184;
wire n_1477;
wire n_2080;
wire n_2220;
wire n_2585;
wire n_1724;
wire n_2554;
wire n_1364;
wire n_1540;
wire n_1676;
wire n_1013;
wire n_2468;
wire n_929;
wire n_637;
wire n_1136;
wire n_1890;
wire n_1075;
wire n_1249;
wire n_1918;
wire n_574;
wire n_2606;
wire n_2549;
wire n_2461;
wire n_2006;
wire n_2440;
wire n_515;
wire n_1229;
wire n_1440;
wire n_1490;
wire n_2152;
wire n_907;
wire n_1179;
wire n_1990;
wire n_1153;
wire n_1751;
wire n_669;
wire n_2467;
wire n_2146;
wire n_2341;
wire n_1737;
wire n_521;
wire n_1117;
wire n_1273;
wire n_2547;
wire n_2616;
wire n_1748;
wire n_1083;
wire n_1014;
wire n_724;
wire n_938;
wire n_1178;
wire n_878;
wire n_2441;
wire n_2358;
wire n_2490;
wire n_594;
wire n_2361;
wire n_1566;
wire n_1464;
wire n_944;
wire n_1848;
wire n_623;
wire n_2062;
wire n_2277;
wire n_585;
wire n_2650;
wire n_1982;
wire n_2252;
wire n_2339;
wire n_1334;
wire n_1963;
wire n_483;
wire n_1695;
wire n_1418;
wire n_2402;
wire n_1137;
wire n_2552;
wire n_660;
wire n_2590;
wire n_524;
wire n_1977;
wire n_2294;
wire n_1200;
wire n_2295;
wire n_2530;
wire n_2379;
wire n_1120;
wire n_2300;
wire n_576;
wire n_1602;
wire n_1776;
wire n_2372;
wire n_2382;
wire n_1852;
wire n_1522;
wire n_2523;
wire n_2557;
wire n_1279;
wire n_2505;
wire n_931;
wire n_827;
wire n_607;
wire n_2481;
wire n_1064;
wire n_1408;
wire n_1028;
wire n_1264;
wire n_2287;
wire n_2102;
wire n_1935;
wire n_2046;
wire n_1146;
wire n_488;
wire n_705;
wire n_2142;
wire n_1548;
wire n_1682;
wire n_1608;
wire n_1009;
wire n_1260;
wire n_589;
wire n_1896;
wire n_1704;
wire n_2160;
wire n_2234;
wire n_847;
wire n_1436;
wire n_2600;
wire n_1069;
wire n_1485;
wire n_2239;
wire n_1465;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_1232;
wire n_1979;
wire n_2328;
wire n_679;
wire n_1345;
wire n_2434;
wire n_696;
wire n_837;
wire n_1590;
wire n_2332;
wire n_640;
wire n_954;
wire n_1628;
wire n_725;
wire n_1773;
wire n_596;
wire n_2133;
wire n_1545;
wire n_2369;
wire n_1471;
wire n_1738;
wire n_1115;
wire n_998;
wire n_1395;
wire n_1729;
wire n_2551;
wire n_801;
wire n_2094;
wire n_2613;
wire n_1479;
wire n_2306;
wire n_1046;
wire n_2419;
wire n_882;
wire n_942;
wire n_1627;
wire n_1431;
wire n_651;
wire n_721;
wire n_2525;
wire n_814;
wire n_1864;
wire n_943;
wire n_2568;
wire n_2629;
wire n_1086;
wire n_1523;
wire n_2197;
wire n_1756;
wire n_2010;
wire n_2097;
wire n_2241;
wire n_1470;
wire n_2098;
wire n_2109;
wire n_1761;
wire n_2648;
wire n_2458;
wire n_1836;
wire n_2398;
wire n_1593;
wire n_986;
wire n_495;
wire n_1420;
wire n_2651;
wire n_1750;
wire n_1775;
wire n_1699;
wire n_927;
wire n_1563;
wire n_615;
wire n_803;
wire n_2570;
wire n_1875;
wire n_1615;
wire n_2184;
wire n_2418;
wire n_1087;
wire n_757;
wire n_1539;
wire n_712;
wire n_1400;
wire n_1599;
wire n_1806;
wire n_650;
wire n_2635;
wire n_2469;
wire n_1575;
wire n_2209;
wire n_1448;
wire n_2077;
wire n_517;
wire n_2520;
wire n_817;
wire n_2193;
wire n_2612;
wire n_2095;
wire n_555;
wire n_2486;
wire n_2628;
wire n_2395;
wire n_951;
wire n_2521;
wire n_2053;
wire n_1580;
wire n_2124;
wire n_1574;
wire n_780;
wire n_2200;
wire n_502;
wire n_1705;
wire n_633;
wire n_2304;
wire n_1746;
wire n_726;
wire n_532;
wire n_1439;
wire n_2263;
wire n_2212;
wire n_2352;
wire n_863;
wire n_597;
wire n_2185;
wire n_1832;
wire n_1128;
wire n_2476;
wire n_2376;
wire n_1266;
wire n_1300;
wire n_807;
wire n_741;
wire n_2460;
wire n_2170;
wire n_1785;
wire n_486;
wire n_1870;
wire n_2484;
wire n_1405;
wire n_997;
wire n_2308;
wire n_1428;
wire n_2243;
wire n_2400;
wire n_891;
wire n_2507;
wire n_1528;
wire n_1495;
wire n_2463;
wire n_2654;
wire n_717;
wire n_1357;
wire n_2503;
wire n_2478;
wire n_1512;
wire n_2496;
wire n_668;
wire n_871;
wire n_1339;
wire n_1544;
wire n_1426;
wire n_2365;
wire n_485;
wire n_2245;
wire n_1315;
wire n_1413;
wire n_2464;
wire n_811;
wire n_808;
wire n_945;
wire n_2270;
wire n_1706;
wire n_1560;
wire n_1592;
wire n_1461;
wire n_2630;
wire n_903;
wire n_1967;
wire n_2340;
wire n_2117;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_2488;
wire n_1378;
wire n_2042;
wire n_1048;
wire n_774;
wire n_2459;
wire n_1925;
wire n_2439;
wire n_2106;
wire n_588;
wire n_1430;
wire n_2414;
wire n_1251;
wire n_1247;
wire n_2450;
wire n_528;
wire n_836;
wire n_1475;
wire n_2465;
wire n_1263;
wire n_1185;
wire n_1683;
wire n_1122;
wire n_890;
wire n_628;
wire n_874;
wire n_1505;
wire n_1163;
wire n_677;
wire n_1514;
wire n_964;
wire n_916;
wire n_2298;
wire n_503;
wire n_895;
wire n_687;
wire n_1035;
wire n_2427;
wire n_2045;
wire n_1535;
wire n_751;
wire n_2190;
wire n_1127;
wire n_932;
wire n_1972;
wire n_947;
wire n_1004;
wire n_831;
wire n_778;
wire n_1898;
wire n_1254;
wire n_1148;
wire n_540;
wire n_1667;
wire n_1104;
wire n_1845;
wire n_1011;
wire n_2205;
wire n_2524;
wire n_1437;
wire n_529;
wire n_626;
wire n_1707;
wire n_1941;
wire n_2422;
wire n_2064;
wire n_1679;
wire n_2342;
wire n_2301;
wire n_1497;
wire n_2002;
wire n_2055;
wire n_2385;
wire n_2545;
wire n_1578;
wire n_2050;
wire n_1143;
wire n_1783;
wire n_510;
wire n_2584;
wire n_972;
wire n_1815;
wire n_2500;
wire n_601;
wire n_610;
wire n_1917;
wire n_1444;
wire n_920;
wire n_664;
wire n_2442;
wire n_1067;
wire n_994;
wire n_2000;
wire n_2089;
wire n_1857;
wire n_1920;
wire n_545;
wire n_887;
wire n_1162;
wire n_1997;
wire n_2578;
wire n_1894;
wire n_2110;
wire n_1349;
wire n_961;
wire n_634;
wire n_991;
wire n_1223;
wire n_1331;
wire n_2127;
wire n_1323;
wire n_578;
wire n_1739;
wire n_1777;
wire n_1353;
wire n_2386;
wire n_1429;
wire n_2029;
wire n_2026;
wire n_1546;
wire n_1432;
wire n_2103;
wire n_1950;
wire n_1320;
wire n_996;
wire n_915;
wire n_2238;
wire n_1174;
wire n_1834;
wire n_1874;
wire n_1727;
wire n_1286;
wire n_1657;
wire n_1741;
wire n_542;
wire n_1294;
wire n_1601;
wire n_900;
wire n_1351;
wire n_2138;
wire n_647;
wire n_1380;
wire n_1367;
wire n_1291;
wire n_1914;
wire n_1458;
wire n_1694;
wire n_1460;
wire n_2041;
wire n_2271;
wire n_2356;
wire n_1830;
wire n_2261;
wire n_1629;
wire n_2011;
wire n_2620;
wire n_1826;
wire n_1855;
wire n_1662;
wire n_2105;
wire n_2187;
wire n_1340;
wire n_2562;
wire n_2642;
wire n_2647;
wire n_1626;
wire n_674;
wire n_2223;
wire n_1660;
wire n_1850;
wire n_1643;
wire n_1670;
wire n_1789;
wire n_552;
wire n_2415;
wire n_2344;
wire n_2317;
wire n_2556;
wire n_1112;
wire n_1267;
wire n_2384;
wire n_1384;
wire n_1376;
wire n_1537;
wire n_1858;
wire n_1816;
wire n_2446;
wire n_1612;
wire n_703;
wire n_2318;
wire n_1172;
wire n_1099;
wire n_598;
wire n_2141;
wire n_1422;
wire n_508;
wire n_1527;
wire n_1055;
wire n_1524;
wire n_673;
wire n_798;
wire n_1754;
wire n_1177;
wire n_1025;
wire n_1991;
wire n_2566;
wire n_2210;
wire n_1517;
wire n_690;
wire n_2502;
wire n_1225;
wire n_1962;
wire n_2346;
wire n_982;
wire n_1624;
wire n_785;
wire n_1952;
wire n_2180;
wire n_2087;
wire n_604;
wire n_1598;
wire n_2617;
wire n_977;
wire n_1895;
wire n_2250;
wire n_719;
wire n_1491;
wire n_1860;
wire n_716;
wire n_1810;
wire n_1763;
wire n_923;
wire n_642;
wire n_1607;
wire n_2075;
wire n_1625;
wire n_2610;
wire n_2420;
wire n_2380;
wire n_2240;
wire n_933;
wire n_2221;
wire n_1774;
wire n_1797;
wire n_2516;
wire n_2120;
wire n_1037;
wire n_1899;
wire n_2031;
wire n_1289;
wire n_838;
wire n_1348;
wire n_1021;
wire n_746;
wire n_1557;
wire n_1188;
wire n_1567;
wire n_2007;
wire n_742;
wire n_1191;
wire n_2004;
wire n_2024;
wire n_2086;
wire n_1503;
wire n_1052;
wire n_789;
wire n_1942;
wire n_656;
wire n_602;
wire n_2309;
wire n_842;
wire n_2274;
wire n_767;
wire n_1617;
wire n_1839;
wire n_1587;
wire n_2330;
wire n_2555;
wire n_2639;
wire n_636;
wire n_1259;
wire n_490;
wire n_2108;
wire n_2535;
wire n_595;
wire n_1001;
wire n_570;
wire n_2143;
wire n_2410;
wire n_1396;
wire n_1224;
wire n_1923;
wire n_2196;
wire n_2611;
wire n_1538;
wire n_487;
wire n_2528;
wire n_2548;
wire n_2633;
wire n_1017;
wire n_2244;
wire n_730;
wire n_2604;
wire n_2437;
wire n_2351;
wire n_2049;
wire n_1456;
wire n_1889;
wire n_625;
wire n_2113;
wire n_619;
wire n_1124;
wire n_611;
wire n_1690;
wire n_1673;
wire n_2018;
wire n_922;
wire n_1790;
wire n_851;
wire n_993;
wire n_2085;
wire n_2581;
wire n_1725;
wire n_2149;
wire n_2237;
wire n_2268;
wire n_2320;
wire n_1135;
wire n_2255;
wire n_2001;
wire n_1820;
wire n_1800;
wire n_541;
wire n_613;
wire n_659;
wire n_1494;
wire n_1550;
wire n_2060;
wire n_1066;
wire n_2214;
wire n_648;
wire n_571;
wire n_1169;
wire n_1726;
wire n_1946;
wire n_1938;
wire n_830;
wire n_1241;
wire n_2589;
wire n_1072;
wire n_2194;
wire n_1231;
wire n_1173;
wire n_1208;
wire n_1604;
wire n_1639;
wire n_826;
wire n_1976;
wire n_2154;
wire n_2035;
wire n_1337;
wire n_1906;
wire n_1647;
wire n_1901;
wire n_839;
wire n_768;
wire n_1278;
wire n_2059;
wire n_796;
wire n_797;
wire n_1006;
wire n_1238;
wire n_1415;
wire n_976;
wire n_1710;
wire n_1063;
wire n_2153;
wire n_2452;
wire n_1270;
wire n_834;
wire n_2457;
wire n_2144;
wire n_1476;
wire n_935;
wire n_1603;
wire n_925;
wire n_2592;
wire n_1054;
wire n_2027;
wire n_2072;
wire n_2012;
wire n_722;
wire n_2251;
wire n_1644;
wire n_1406;
wire n_1489;
wire n_1880;
wire n_1993;
wire n_2137;
wire n_804;
wire n_1455;
wire n_484;
wire n_1642;
wire n_1871;
wire n_2182;
wire n_2447;
wire n_1057;
wire n_1473;
wire n_516;
wire n_2125;
wire n_2426;
wire n_1403;
wire n_2181;
wire n_2587;
wire n_1149;
wire n_1176;
wire n_1502;
wire n_1605;
wire n_506;
wire n_868;
wire n_2099;
wire n_1202;
wire n_1065;
wire n_1897;
wire n_2477;
wire n_1457;
wire n_905;
wire n_2159;
wire n_975;
wire n_675;
wire n_624;
wire n_934;
wire n_520;
wire n_775;
wire n_512;
wire n_950;
wire n_685;
wire n_1222;
wire n_1630;
wire n_2286;
wire n_1879;
wire n_1959;
wire n_2563;
wire n_1198;
wire n_2206;
wire n_1311;
wire n_1261;
wire n_2299;
wire n_2078;
wire n_2265;
wire n_776;
wire n_1114;
wire n_818;
wire n_1167;
wire n_2531;
wire n_2315;
wire n_2157;
wire n_1282;
wire n_2067;
wire n_2517;
wire n_1321;
wire n_700;
wire n_1779;
wire n_2489;
wire n_1770;
wire n_1107;
wire n_1846;
wire n_2211;
wire n_1573;
wire n_525;
wire n_815;
wire n_919;
wire n_2272;
wire n_535;
wire n_1956;
wire n_681;
wire n_2608;
wire n_1718;
wire n_2225;
wire n_2546;
wire n_1411;
wire n_1139;
wire n_858;
wire n_1018;
wire n_2345;
wire n_1324;
wire n_1669;
wire n_1501;
wire n_782;
wire n_616;
wire n_1885;
wire n_1740;
wire n_1989;
wire n_1838;
wire n_833;
wire n_1343;
wire n_1801;
wire n_1371;
wire n_1513;
wire n_728;
wire n_2161;
wire n_2191;
wire n_2329;
wire n_1788;
wire n_2093;
wire n_2348;
wire n_786;
wire n_2576;
wire n_2417;
wire n_505;
wire n_2043;
wire n_2366;
wire n_1621;
wire n_2338;
wire n_1919;
wire n_1342;
wire n_501;
wire n_752;
wire n_2009;
wire n_2248;
wire n_958;
wire n_1175;
wire n_1416;
wire n_1659;
wire n_1221;
wire n_1047;
wire n_1878;
wire n_1515;
wire n_1374;
wire n_2438;
wire n_1435;
wire n_1688;
wire n_792;
wire n_1314;
wire n_1433;
wire n_2567;
wire n_575;
wire n_1242;
wire n_1119;
wire n_2229;
wire n_1085;
wire n_2388;
wire n_2222;
wire n_1907;
wire n_885;
wire n_1530;
wire n_513;
wire n_877;
wire n_2135;
wire n_1088;
wire n_896;
wire n_2624;
wire n_1813;
wire n_1451;
wire n_1005;
wire n_1102;
wire n_631;
wire n_794;
wire n_2471;
wire n_1288;
wire n_1275;
wire n_985;
wire n_1165;
wire n_897;
wire n_1622;
wire n_697;
wire n_1105;
wire n_1459;
wire n_912;
wire n_2232;
wire n_2455;
wire n_2121;
wire n_1893;
wire n_2519;
wire n_1570;
wire n_2231;
wire n_701;
wire n_995;
wire n_2278;
wire n_1000;
wire n_2284;
wire n_1931;
wire n_2433;
wire n_1256;
wire n_587;
wire n_1303;
wire n_1994;
wire n_1771;
wire n_1526;
wire n_764;
wire n_1507;
wire n_1206;
wire n_1809;
wire n_855;
wire n_2367;
wire n_812;
wire n_1961;
wire n_2553;
wire n_1050;
wire n_2218;
wire n_599;
wire n_1769;
wire n_2130;
wire n_1060;
wire n_1372;
wire n_1847;
wire n_756;
wire n_1565;
wire n_1257;
wire n_2325;
wire n_2406;
wire n_1632;
wire n_688;
wire n_1542;
wire n_946;
wire n_1586;
wire n_707;
wire n_1362;
wire n_1547;
wire n_1097;
wire n_2518;
wire n_1909;
wire n_2543;
wire n_2381;
wire n_621;
wire n_2313;
wire n_956;
wire n_790;
wire n_2495;
wire n_1541;
wire n_1812;
wire n_1951;
wire n_586;
wire n_1330;
wire n_638;
wire n_1697;
wire n_2128;
wire n_2574;
wire n_1872;
wire n_1940;
wire n_593;
wire n_1747;
wire n_1212;
wire n_1887;
wire n_1199;
wire n_2020;
wire n_1978;
wire n_2508;
wire n_2540;
wire n_1767;
wire n_1939;
wire n_2428;
wire n_1768;
wire n_1443;
wire n_2068;
wire n_2636;
wire n_1585;
wire n_1861;
wire n_2316;
wire n_1564;
wire n_1995;
wire n_1631;
wire n_2593;
wire n_1623;
wire n_861;
wire n_1828;
wire n_2364;
wire n_1389;
wire n_1131;
wire n_2641;
wire n_547;
wire n_1798;
wire n_727;
wire n_1077;
wire n_1554;
wire n_1584;
wire n_1481;
wire n_2021;
wire n_1928;
wire n_828;
wire n_1438;
wire n_1973;
wire n_2314;
wire n_2156;
wire n_2494;
wire n_753;
wire n_2126;
wire n_645;
wire n_1147;
wire n_747;
wire n_1363;
wire n_2228;
wire n_1691;
wire n_1098;
wire n_584;
wire n_1366;
wire n_1518;
wire n_1361;
wire n_1187;
wire n_2034;
wire n_1693;
wire n_698;
wire n_2411;
wire n_2081;
wire n_1892;
wire n_1061;
wire n_2266;
wire n_682;
wire n_2061;
wire n_1373;
wire n_2449;
wire n_1686;
wire n_2131;
wire n_2526;
wire n_1302;
wire n_2083;
wire n_886;
wire n_2119;
wire n_1010;
wire n_883;
wire n_2207;
wire n_2044;
wire n_2542;
wire n_755;
wire n_2091;
wire n_1029;
wire n_2394;
wire n_770;
wire n_1572;
wire n_1635;
wire n_941;
wire n_1245;
wire n_1317;
wire n_2615;
wire n_2487;
wire n_632;
wire n_1329;
wire n_2409;
wire n_2637;
wire n_2337;
wire n_854;
wire n_2405;
wire n_2601;
wire n_2513;
wire n_1369;
wire n_714;
wire n_1297;
wire n_1912;
wire n_1734;
wire n_1876;
wire n_2323;
wire n_740;
wire n_549;
wire n_533;
wire n_1811;
wire n_898;
wire n_928;
wire n_1285;
wire n_967;
wire n_2561;
wire n_736;
wire n_2491;
wire n_1529;
wire n_1381;
wire n_1824;
wire n_2254;
wire n_1597;
wire n_1161;
wire n_1103;
wire n_1486;
wire n_1068;
wire n_617;
wire n_1833;
wire n_2371;
wire n_914;
wire n_1986;
wire n_526;
wire n_1024;
wire n_1141;
wire n_1949;
wire n_1197;
wire n_2493;
wire n_2408;
wire n_2429;
wire n_1168;
wire n_865;
wire n_2115;
wire n_2013;
wire n_2140;
wire n_2134;
wire n_569;
wire n_2483;
wire n_2305;
wire n_600;
wire n_1556;
wire n_1192;
wire n_1646;
wire n_1290;
wire n_2514;
wire n_2466;
wire n_1759;
wire n_2048;
wire n_987;
wire n_1299;
wire n_750;
wire n_2096;
wire n_2129;
wire n_665;
wire n_1101;
wire n_2532;
wire n_2079;
wire n_2296;
wire n_1720;
wire n_880;
wire n_654;
wire n_1911;
wire n_2293;
wire n_731;
wire n_1336;
wire n_758;
wire n_1166;
wire n_710;
wire n_720;
wire n_1390;
wire n_1023;
wire n_568;
wire n_1358;
wire n_813;
wire n_2310;
wire n_1397;
wire n_1211;
wire n_1284;
wire n_2005;
wire n_1359;
wire n_1116;
wire n_1758;
wire n_791;
wire n_1532;
wire n_1419;
wire n_543;
wire n_580;
wire n_1784;
wire n_1685;
wire n_1992;
wire n_1082;
wire n_1213;
wire n_2596;
wire n_980;
wire n_1193;
wire n_849;
wire n_1488;
wire n_2227;
wire n_2652;
wire n_1074;
wire n_1379;
wire n_759;
wire n_1721;
wire n_2627;
wire n_1827;
wire n_953;
wire n_1180;
wire n_1462;
wire n_536;
wire n_2326;
wire n_1866;
wire n_1220;
wire n_1398;
wire n_2111;
wire n_2169;
wire n_1262;
wire n_1904;
wire n_1692;
wire n_2501;
wire n_2051;
wire n_1012;
wire n_1805;
wire n_960;
wire n_689;
wire n_1022;
wire n_1760;
wire n_676;
wire n_1240;
wire n_2173;
wire n_1183;
wire n_1204;
wire n_1151;
wire n_1814;
wire n_771;
wire n_999;
wire n_514;
wire n_2634;
wire n_1092;
wire n_1808;
wire n_560;
wire n_1658;
wire n_1386;
wire n_2588;
wire n_2492;
wire n_910;
wire n_2291;
wire n_635;
wire n_844;
wire n_2172;
wire n_1728;
wire n_1020;
wire n_783;
wire n_1142;
wire n_1385;
wire n_1062;
wire n_1230;
wire n_1027;
wire n_1516;
wire n_2533;
wire n_1499;
wire n_1500;
wire n_2155;
wire n_1868;
wire n_966;
wire n_2148;
wire n_2104;
wire n_949;
wire n_704;
wire n_2303;
wire n_2357;
wire n_2618;
wire n_2653;
wire n_924;
wire n_2331;
wire n_1600;
wire n_1661;
wire n_1965;
wire n_1757;
wire n_699;
wire n_2136;
wire n_2403;
wire n_918;
wire n_2056;
wire n_1913;
wire n_672;
wire n_2054;
wire n_1039;
wire n_2226;
wire n_2407;
wire n_1043;
wire n_1402;
wire n_2267;
wire n_735;
wire n_1450;
wire n_2082;
wire n_2302;
wire n_2453;
wire n_2560;
wire n_2092;
wire n_566;
wire n_581;
wire n_1472;
wire n_1365;
wire n_2443;
wire n_2279;
wire n_1089;
wire n_1536;
wire n_1049;
wire n_1719;
wire n_2066;
wire n_548;
wire n_1158;
wire n_1974;
wire n_763;
wire n_1882;
wire n_1915;
wire n_940;
wire n_1762;
wire n_2534;
wire n_1404;
wire n_546;
wire n_788;
wire n_1736;
wire n_1160;
wire n_1442;
wire n_658;
wire n_1948;
wire n_2168;
wire n_1216;
wire n_1891;
wire n_1026;
wire n_1454;
wire n_1033;
wire n_627;
wire n_990;
wire n_1383;
wire n_1968;
wire n_2057;
wire n_2609;
wire n_2378;
wire n_888;
wire n_1325;
wire n_2014;
wire n_582;
wire n_1483;
wire n_1703;
wire n_653;
wire n_1205;
wire n_1822;
wire n_843;
wire n_1953;
wire n_1059;
wire n_799;
wire n_691;
wire n_1804;
wire n_1581;
wire n_522;
wire n_534;
wire n_1837;
wire n_511;
wire n_1744;
wire n_1975;
wire n_1414;
wire n_2324;
wire n_2246;
wire n_1002;
wire n_1851;
wire n_1755;
wire n_2195;
wire n_1111;
wire n_1819;
wire n_1341;
wire n_1807;
wire n_2645;
wire n_2202;
wire n_1310;
wire n_1745;
wire n_1714;
wire n_612;
wire n_1958;
wire n_1611;
wire n_2559;
wire n_2262;
wire n_955;
wire n_1333;
wire n_1916;
wire n_2619;
wire n_2073;
wire n_952;
wire n_1675;
wire n_1947;
wire n_2165;
wire n_1640;
wire n_2016;
wire n_1551;
wire n_1145;
wire n_1533;
wire n_2307;
wire n_2515;
wire n_1511;
wire n_1791;
wire n_537;
wire n_1113;
wire n_1651;
wire n_1966;
wire n_2058;
wire n_1468;
wire n_2327;
wire n_2656;
wire n_913;
wire n_2353;
wire n_509;
wire n_1164;
wire n_2258;
wire n_1732;
wire n_2167;
wire n_1354;
wire n_2039;
wire n_1277;
wire n_1696;
wire n_1016;
wire n_680;
wire n_1355;
wire n_809;
wire n_2544;
wire n_856;
wire n_779;
wire n_2538;
wire n_2582;
wire n_1559;
wire n_2321;
wire n_1579;
wire n_1280;
wire n_493;
wire n_1335;
wire n_2285;
wire n_1934;
wire n_1900;
wire n_2040;
wire n_2174;
wire n_519;
wire n_1843;
wire n_2186;
wire n_2510;
wire n_2030;
wire n_2614;
wire n_2435;
wire n_1665;
wire n_2583;
wire n_1091;
wire n_1678;
wire n_1780;
wire n_1287;
wire n_1482;
wire n_860;
wire n_1525;
wire n_661;
wire n_848;
wire n_2100;
wire n_2349;
wire n_1902;
wire n_2536;
wire n_2474;
wire n_683;
wire n_1194;
wire n_1150;
wire n_620;
wire n_1399;
wire n_1903;
wire n_1674;
wire n_1849;
wire n_686;
wire n_572;
wire n_867;
wire n_983;
wire n_1417;
wire n_644;
wire n_577;
wire n_2282;
wire n_970;
wire n_491;
wire n_2430;
wire n_921;
wire n_489;
wire n_1534;
wire n_908;
wire n_1346;
wire n_565;
wire n_1123;
wire n_1272;
wire n_2497;
wire n_1393;
wire n_984;
wire n_1655;
wire n_1410;
wire n_988;
wire n_2368;
wire n_760;
wire n_1157;
wire n_806;
wire n_1186;
wire n_2065;
wire n_1743;
wire n_492;
wire n_649;
wire n_1854;
wire n_866;
wire n_559;

BUFx3_ASAP7_75t_L g482 ( 
.A(n_321),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_446),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_39),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_131),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_354),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_226),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_455),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_452),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_293),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_260),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_257),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_283),
.Y(n_493)
);

INVx1_ASAP7_75t_SL g494 ( 
.A(n_419),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_382),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_236),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_96),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_433),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_259),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_351),
.Y(n_500)
);

INVxp67_ASAP7_75t_L g501 ( 
.A(n_470),
.Y(n_501)
);

CKINVDCx20_ASAP7_75t_R g502 ( 
.A(n_8),
.Y(n_502)
);

BUFx6f_ASAP7_75t_L g503 ( 
.A(n_39),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_178),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_95),
.Y(n_505)
);

CKINVDCx20_ASAP7_75t_R g506 ( 
.A(n_37),
.Y(n_506)
);

BUFx6f_ASAP7_75t_L g507 ( 
.A(n_228),
.Y(n_507)
);

BUFx3_ASAP7_75t_L g508 ( 
.A(n_224),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_27),
.Y(n_509)
);

BUFx6f_ASAP7_75t_L g510 ( 
.A(n_386),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_76),
.Y(n_511)
);

INVxp67_ASAP7_75t_L g512 ( 
.A(n_441),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_333),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_270),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_89),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_308),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_114),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_164),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_368),
.Y(n_519)
);

INVx1_ASAP7_75t_SL g520 ( 
.A(n_211),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_258),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_14),
.Y(n_522)
);

BUFx5_ASAP7_75t_L g523 ( 
.A(n_265),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_463),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_215),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_254),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_266),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_181),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_91),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_153),
.Y(n_530)
);

INVx2_ASAP7_75t_SL g531 ( 
.A(n_5),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_292),
.Y(n_532)
);

CKINVDCx16_ASAP7_75t_R g533 ( 
.A(n_476),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_90),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_132),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_353),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_123),
.Y(n_537)
);

BUFx3_ASAP7_75t_L g538 ( 
.A(n_374),
.Y(n_538)
);

BUFx6f_ASAP7_75t_L g539 ( 
.A(n_437),
.Y(n_539)
);

BUFx10_ASAP7_75t_L g540 ( 
.A(n_359),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_415),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_98),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_373),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_197),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_305),
.Y(n_545)
);

BUFx2_ASAP7_75t_SL g546 ( 
.A(n_296),
.Y(n_546)
);

BUFx10_ASAP7_75t_L g547 ( 
.A(n_436),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_58),
.Y(n_548)
);

INVx1_ASAP7_75t_SL g549 ( 
.A(n_98),
.Y(n_549)
);

INVx1_ASAP7_75t_SL g550 ( 
.A(n_206),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_267),
.Y(n_551)
);

BUFx10_ASAP7_75t_L g552 ( 
.A(n_420),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_52),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_428),
.Y(n_554)
);

BUFx5_ASAP7_75t_L g555 ( 
.A(n_156),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_300),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_116),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_150),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_52),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_408),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_377),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_210),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_453),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_474),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_17),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_304),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_389),
.Y(n_567)
);

BUFx3_ASAP7_75t_L g568 ( 
.A(n_1),
.Y(n_568)
);

INVx1_ASAP7_75t_SL g569 ( 
.A(n_218),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_394),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_141),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_235),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_403),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_378),
.Y(n_574)
);

BUFx2_ASAP7_75t_L g575 ( 
.A(n_25),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_322),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_302),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_167),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_319),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_1),
.Y(n_580)
);

CKINVDCx20_ASAP7_75t_R g581 ( 
.A(n_393),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_360),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_268),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_102),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_451),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_15),
.Y(n_586)
);

BUFx10_ASAP7_75t_L g587 ( 
.A(n_464),
.Y(n_587)
);

INVx3_ASAP7_75t_L g588 ( 
.A(n_406),
.Y(n_588)
);

BUFx10_ASAP7_75t_L g589 ( 
.A(n_100),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_383),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_188),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_42),
.Y(n_592)
);

BUFx6f_ASAP7_75t_L g593 ( 
.A(n_295),
.Y(n_593)
);

INVx1_ASAP7_75t_SL g594 ( 
.A(n_218),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_192),
.Y(n_595)
);

INVx1_ASAP7_75t_SL g596 ( 
.A(n_228),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_66),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_272),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_276),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_279),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_479),
.Y(n_601)
);

CKINVDCx20_ASAP7_75t_R g602 ( 
.A(n_234),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_328),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_278),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_332),
.Y(n_605)
);

BUFx3_ASAP7_75t_L g606 ( 
.A(n_64),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_401),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_443),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_461),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_37),
.Y(n_610)
);

BUFx3_ASAP7_75t_L g611 ( 
.A(n_105),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_345),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_400),
.Y(n_613)
);

CKINVDCx20_ASAP7_75t_R g614 ( 
.A(n_23),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_87),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_326),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_190),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_148),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_456),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_291),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_226),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_36),
.Y(n_622)
);

BUFx10_ASAP7_75t_L g623 ( 
.A(n_104),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_429),
.Y(n_624)
);

CKINVDCx20_ASAP7_75t_R g625 ( 
.A(n_60),
.Y(n_625)
);

CKINVDCx20_ASAP7_75t_R g626 ( 
.A(n_320),
.Y(n_626)
);

BUFx10_ASAP7_75t_L g627 ( 
.A(n_63),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_195),
.Y(n_628)
);

INVxp67_ASAP7_75t_L g629 ( 
.A(n_426),
.Y(n_629)
);

INVx2_ASAP7_75t_SL g630 ( 
.A(n_2),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_50),
.Y(n_631)
);

CKINVDCx16_ASAP7_75t_R g632 ( 
.A(n_208),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_161),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_412),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_285),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_171),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_244),
.Y(n_637)
);

CKINVDCx20_ASAP7_75t_R g638 ( 
.A(n_425),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_202),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_3),
.Y(n_640)
);

CKINVDCx20_ASAP7_75t_R g641 ( 
.A(n_50),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_286),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_42),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_367),
.Y(n_644)
);

CKINVDCx20_ASAP7_75t_R g645 ( 
.A(n_69),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_318),
.Y(n_646)
);

CKINVDCx20_ASAP7_75t_R g647 ( 
.A(n_303),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_247),
.Y(n_648)
);

INVx1_ASAP7_75t_SL g649 ( 
.A(n_480),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_3),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_224),
.Y(n_651)
);

CKINVDCx16_ASAP7_75t_R g652 ( 
.A(n_127),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_361),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_105),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_126),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_273),
.Y(n_656)
);

CKINVDCx20_ASAP7_75t_R g657 ( 
.A(n_257),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_371),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_88),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_232),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_71),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_366),
.Y(n_662)
);

BUFx6f_ASAP7_75t_L g663 ( 
.A(n_89),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_325),
.Y(n_664)
);

INVx1_ASAP7_75t_SL g665 ( 
.A(n_206),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_191),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_237),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_191),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_264),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_450),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_88),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_432),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_421),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_338),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_15),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_54),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_196),
.Y(n_677)
);

BUFx3_ASAP7_75t_L g678 ( 
.A(n_460),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_212),
.Y(n_679)
);

INVx1_ASAP7_75t_SL g680 ( 
.A(n_467),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_301),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_237),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_121),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_240),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_123),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_380),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_457),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_227),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_233),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_239),
.Y(n_690)
);

BUFx10_ASAP7_75t_L g691 ( 
.A(n_284),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_110),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_198),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_147),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_337),
.Y(n_695)
);

INVx2_ASAP7_75t_SL g696 ( 
.A(n_14),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_236),
.Y(n_697)
);

INVx1_ASAP7_75t_SL g698 ( 
.A(n_201),
.Y(n_698)
);

BUFx3_ASAP7_75t_L g699 ( 
.A(n_402),
.Y(n_699)
);

BUFx3_ASAP7_75t_L g700 ( 
.A(n_329),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_472),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_160),
.Y(n_702)
);

INVx1_ASAP7_75t_SL g703 ( 
.A(n_84),
.Y(n_703)
);

BUFx6f_ASAP7_75t_L g704 ( 
.A(n_313),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_458),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_277),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_481),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_217),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_122),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_75),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_306),
.Y(n_711)
);

INVx1_ASAP7_75t_SL g712 ( 
.A(n_137),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_82),
.Y(n_713)
);

CKINVDCx16_ASAP7_75t_R g714 ( 
.A(n_448),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_381),
.Y(n_715)
);

INVxp67_ASAP7_75t_L g716 ( 
.A(n_151),
.Y(n_716)
);

CKINVDCx20_ASAP7_75t_R g717 ( 
.A(n_376),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_163),
.Y(n_718)
);

INVx1_ASAP7_75t_SL g719 ( 
.A(n_362),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_201),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_68),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_110),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_442),
.Y(n_723)
);

BUFx6f_ASAP7_75t_L g724 ( 
.A(n_468),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_356),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_162),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_0),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_466),
.Y(n_728)
);

INVx1_ASAP7_75t_SL g729 ( 
.A(n_157),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_299),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_256),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_199),
.Y(n_732)
);

INVx3_ASAP7_75t_L g733 ( 
.A(n_28),
.Y(n_733)
);

BUFx6f_ASAP7_75t_L g734 ( 
.A(n_142),
.Y(n_734)
);

BUFx10_ASAP7_75t_L g735 ( 
.A(n_275),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_58),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_176),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_76),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_177),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_122),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_307),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_316),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_186),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_10),
.Y(n_744)
);

BUFx2_ASAP7_75t_L g745 ( 
.A(n_22),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_26),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_330),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_143),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_255),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_172),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_70),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_245),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_235),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_5),
.Y(n_754)
);

CKINVDCx5p33_ASAP7_75t_R g755 ( 
.A(n_375),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_290),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_397),
.Y(n_757)
);

INVxp67_ASAP7_75t_SL g758 ( 
.A(n_155),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_242),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_127),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_144),
.Y(n_761)
);

CKINVDCx20_ASAP7_75t_R g762 ( 
.A(n_335),
.Y(n_762)
);

INVx2_ASAP7_75t_SL g763 ( 
.A(n_144),
.Y(n_763)
);

CKINVDCx5p33_ASAP7_75t_R g764 ( 
.A(n_465),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_92),
.Y(n_765)
);

BUFx2_ASAP7_75t_L g766 ( 
.A(n_227),
.Y(n_766)
);

CKINVDCx5p33_ASAP7_75t_R g767 ( 
.A(n_84),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_390),
.Y(n_768)
);

CKINVDCx5p33_ASAP7_75t_R g769 ( 
.A(n_348),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_215),
.Y(n_770)
);

BUFx8_ASAP7_75t_SL g771 ( 
.A(n_143),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_477),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_192),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_216),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_179),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_99),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_36),
.Y(n_777)
);

BUFx6f_ASAP7_75t_L g778 ( 
.A(n_242),
.Y(n_778)
);

CKINVDCx5p33_ASAP7_75t_R g779 ( 
.A(n_274),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_106),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_317),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_186),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_138),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_141),
.Y(n_784)
);

CKINVDCx20_ASAP7_75t_R g785 ( 
.A(n_63),
.Y(n_785)
);

CKINVDCx20_ASAP7_75t_R g786 ( 
.A(n_27),
.Y(n_786)
);

BUFx5_ASAP7_75t_L g787 ( 
.A(n_312),
.Y(n_787)
);

INVx1_ASAP7_75t_SL g788 ( 
.A(n_20),
.Y(n_788)
);

CKINVDCx5p33_ASAP7_75t_R g789 ( 
.A(n_166),
.Y(n_789)
);

CKINVDCx20_ASAP7_75t_R g790 ( 
.A(n_387),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_263),
.Y(n_791)
);

INVxp33_ASAP7_75t_SL g792 ( 
.A(n_202),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_67),
.Y(n_793)
);

CKINVDCx5p33_ASAP7_75t_R g794 ( 
.A(n_103),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_102),
.Y(n_795)
);

CKINVDCx5p33_ASAP7_75t_R g796 ( 
.A(n_79),
.Y(n_796)
);

CKINVDCx5p33_ASAP7_75t_R g797 ( 
.A(n_294),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_178),
.Y(n_798)
);

HB1xp67_ASAP7_75t_L g799 ( 
.A(n_96),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_147),
.Y(n_800)
);

CKINVDCx5p33_ASAP7_75t_R g801 ( 
.A(n_372),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_182),
.Y(n_802)
);

INVxp67_ASAP7_75t_SL g803 ( 
.A(n_733),
.Y(n_803)
);

INVxp67_ASAP7_75t_SL g804 ( 
.A(n_733),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_733),
.Y(n_805)
);

BUFx2_ASAP7_75t_L g806 ( 
.A(n_575),
.Y(n_806)
);

CKINVDCx20_ASAP7_75t_R g807 ( 
.A(n_771),
.Y(n_807)
);

CKINVDCx5p33_ASAP7_75t_R g808 ( 
.A(n_771),
.Y(n_808)
);

INVx3_ASAP7_75t_L g809 ( 
.A(n_508),
.Y(n_809)
);

HB1xp67_ASAP7_75t_L g810 ( 
.A(n_799),
.Y(n_810)
);

INVxp67_ASAP7_75t_SL g811 ( 
.A(n_508),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_531),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_531),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_630),
.Y(n_814)
);

NOR2xp33_ASAP7_75t_L g815 ( 
.A(n_588),
.B(n_0),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_630),
.Y(n_816)
);

CKINVDCx5p33_ASAP7_75t_R g817 ( 
.A(n_533),
.Y(n_817)
);

CKINVDCx20_ASAP7_75t_R g818 ( 
.A(n_632),
.Y(n_818)
);

NOR2xp67_ASAP7_75t_L g819 ( 
.A(n_696),
.B(n_2),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_696),
.Y(n_820)
);

CKINVDCx16_ASAP7_75t_R g821 ( 
.A(n_652),
.Y(n_821)
);

CKINVDCx20_ASAP7_75t_R g822 ( 
.A(n_502),
.Y(n_822)
);

CKINVDCx5p33_ASAP7_75t_R g823 ( 
.A(n_714),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_581),
.Y(n_824)
);

CKINVDCx5p33_ASAP7_75t_R g825 ( 
.A(n_581),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_763),
.Y(n_826)
);

CKINVDCx5p33_ASAP7_75t_R g827 ( 
.A(n_626),
.Y(n_827)
);

CKINVDCx20_ASAP7_75t_R g828 ( 
.A(n_502),
.Y(n_828)
);

INVx3_ASAP7_75t_L g829 ( 
.A(n_568),
.Y(n_829)
);

BUFx3_ASAP7_75t_L g830 ( 
.A(n_588),
.Y(n_830)
);

CKINVDCx5p33_ASAP7_75t_R g831 ( 
.A(n_626),
.Y(n_831)
);

NOR2xp67_ASAP7_75t_L g832 ( 
.A(n_763),
.B(n_716),
.Y(n_832)
);

CKINVDCx5p33_ASAP7_75t_R g833 ( 
.A(n_638),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_568),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_606),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_606),
.Y(n_836)
);

INVxp67_ASAP7_75t_SL g837 ( 
.A(n_611),
.Y(n_837)
);

CKINVDCx5p33_ASAP7_75t_R g838 ( 
.A(n_638),
.Y(n_838)
);

INVxp67_ASAP7_75t_SL g839 ( 
.A(n_745),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_484),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_484),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_654),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_654),
.Y(n_843)
);

NOR2xp33_ASAP7_75t_L g844 ( 
.A(n_588),
.B(n_4),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_697),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_697),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_721),
.Y(n_847)
);

NOR2xp33_ASAP7_75t_L g848 ( 
.A(n_483),
.B(n_4),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_721),
.Y(n_849)
);

CKINVDCx5p33_ASAP7_75t_R g850 ( 
.A(n_647),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_722),
.Y(n_851)
);

CKINVDCx5p33_ASAP7_75t_R g852 ( 
.A(n_647),
.Y(n_852)
);

CKINVDCx5p33_ASAP7_75t_R g853 ( 
.A(n_717),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_722),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_726),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_726),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_737),
.Y(n_857)
);

CKINVDCx20_ASAP7_75t_R g858 ( 
.A(n_506),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_737),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_749),
.Y(n_860)
);

CKINVDCx20_ASAP7_75t_R g861 ( 
.A(n_506),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_749),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_751),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_751),
.Y(n_864)
);

CKINVDCx20_ASAP7_75t_R g865 ( 
.A(n_602),
.Y(n_865)
);

CKINVDCx5p33_ASAP7_75t_R g866 ( 
.A(n_717),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_754),
.Y(n_867)
);

CKINVDCx20_ASAP7_75t_R g868 ( 
.A(n_602),
.Y(n_868)
);

INVxp67_ASAP7_75t_SL g869 ( 
.A(n_766),
.Y(n_869)
);

CKINVDCx14_ASAP7_75t_R g870 ( 
.A(n_540),
.Y(n_870)
);

NOR2xp33_ASAP7_75t_L g871 ( 
.A(n_486),
.B(n_6),
.Y(n_871)
);

CKINVDCx5p33_ASAP7_75t_R g872 ( 
.A(n_762),
.Y(n_872)
);

CKINVDCx5p33_ASAP7_75t_R g873 ( 
.A(n_762),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_555),
.Y(n_874)
);

CKINVDCx20_ASAP7_75t_R g875 ( 
.A(n_614),
.Y(n_875)
);

CKINVDCx5p33_ASAP7_75t_R g876 ( 
.A(n_790),
.Y(n_876)
);

INVxp67_ASAP7_75t_L g877 ( 
.A(n_589),
.Y(n_877)
);

CKINVDCx20_ASAP7_75t_R g878 ( 
.A(n_614),
.Y(n_878)
);

CKINVDCx5p33_ASAP7_75t_R g879 ( 
.A(n_790),
.Y(n_879)
);

CKINVDCx20_ASAP7_75t_R g880 ( 
.A(n_625),
.Y(n_880)
);

CKINVDCx5p33_ASAP7_75t_R g881 ( 
.A(n_504),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_754),
.Y(n_882)
);

INVxp67_ASAP7_75t_L g883 ( 
.A(n_589),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_555),
.Y(n_884)
);

CKINVDCx20_ASAP7_75t_R g885 ( 
.A(n_625),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_773),
.Y(n_886)
);

CKINVDCx5p33_ASAP7_75t_R g887 ( 
.A(n_504),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_773),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_800),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_800),
.Y(n_890)
);

INVxp67_ASAP7_75t_SL g891 ( 
.A(n_555),
.Y(n_891)
);

HB1xp67_ASAP7_75t_L g892 ( 
.A(n_505),
.Y(n_892)
);

NOR2xp67_ASAP7_75t_L g893 ( 
.A(n_487),
.B(n_6),
.Y(n_893)
);

CKINVDCx20_ASAP7_75t_R g894 ( 
.A(n_641),
.Y(n_894)
);

CKINVDCx20_ASAP7_75t_R g895 ( 
.A(n_641),
.Y(n_895)
);

INVxp67_ASAP7_75t_L g896 ( 
.A(n_589),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_555),
.Y(n_897)
);

INVxp67_ASAP7_75t_SL g898 ( 
.A(n_555),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_505),
.B(n_7),
.Y(n_899)
);

INVx2_ASAP7_75t_L g900 ( 
.A(n_555),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_555),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_497),
.Y(n_902)
);

NOR2xp67_ASAP7_75t_L g903 ( 
.A(n_509),
.B(n_515),
.Y(n_903)
);

CKINVDCx5p33_ASAP7_75t_R g904 ( 
.A(n_511),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_517),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_518),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_526),
.Y(n_907)
);

CKINVDCx5p33_ASAP7_75t_R g908 ( 
.A(n_511),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_528),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_529),
.Y(n_910)
);

BUFx3_ASAP7_75t_L g911 ( 
.A(n_482),
.Y(n_911)
);

INVx2_ASAP7_75t_L g912 ( 
.A(n_523),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_530),
.Y(n_913)
);

INVxp67_ASAP7_75t_L g914 ( 
.A(n_623),
.Y(n_914)
);

CKINVDCx16_ASAP7_75t_R g915 ( 
.A(n_623),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_542),
.Y(n_916)
);

INVx1_ASAP7_75t_SL g917 ( 
.A(n_522),
.Y(n_917)
);

NOR2xp33_ASAP7_75t_L g918 ( 
.A(n_498),
.B(n_7),
.Y(n_918)
);

CKINVDCx5p33_ASAP7_75t_R g919 ( 
.A(n_522),
.Y(n_919)
);

CKINVDCx16_ASAP7_75t_R g920 ( 
.A(n_623),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_562),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_571),
.Y(n_922)
);

BUFx2_ASAP7_75t_L g923 ( 
.A(n_525),
.Y(n_923)
);

NOR2xp67_ASAP7_75t_L g924 ( 
.A(n_580),
.B(n_8),
.Y(n_924)
);

CKINVDCx5p33_ASAP7_75t_R g925 ( 
.A(n_525),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_586),
.Y(n_926)
);

NOR2xp33_ASAP7_75t_L g927 ( 
.A(n_500),
.B(n_9),
.Y(n_927)
);

CKINVDCx20_ASAP7_75t_R g928 ( 
.A(n_645),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_595),
.Y(n_929)
);

NOR2xp33_ASAP7_75t_L g930 ( 
.A(n_516),
.B(n_9),
.Y(n_930)
);

NOR2xp33_ASAP7_75t_L g931 ( 
.A(n_532),
.B(n_10),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_597),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_615),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_618),
.Y(n_934)
);

CKINVDCx5p33_ASAP7_75t_R g935 ( 
.A(n_513),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_622),
.Y(n_936)
);

CKINVDCx5p33_ASAP7_75t_R g937 ( 
.A(n_513),
.Y(n_937)
);

AND2x2_ASAP7_75t_SL g938 ( 
.A(n_915),
.B(n_503),
.Y(n_938)
);

NAND2x1p5_ASAP7_75t_L g939 ( 
.A(n_923),
.B(n_631),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_830),
.Y(n_940)
);

HB1xp67_ASAP7_75t_L g941 ( 
.A(n_881),
.Y(n_941)
);

INVx2_ASAP7_75t_L g942 ( 
.A(n_874),
.Y(n_942)
);

INVx2_ASAP7_75t_L g943 ( 
.A(n_874),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_812),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_803),
.B(n_727),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_813),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_814),
.Y(n_947)
);

BUFx8_ASAP7_75t_L g948 ( 
.A(n_806),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_816),
.Y(n_949)
);

AND2x6_ASAP7_75t_L g950 ( 
.A(n_815),
.B(n_482),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_804),
.B(n_727),
.Y(n_951)
);

INVx3_ASAP7_75t_L g952 ( 
.A(n_809),
.Y(n_952)
);

AND2x4_ASAP7_75t_L g953 ( 
.A(n_820),
.B(n_648),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_826),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_805),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_809),
.Y(n_956)
);

AND2x2_ASAP7_75t_L g957 ( 
.A(n_870),
.B(n_627),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_809),
.Y(n_958)
);

AND2x2_ASAP7_75t_L g959 ( 
.A(n_810),
.B(n_627),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_829),
.Y(n_960)
);

BUFx6f_ASAP7_75t_L g961 ( 
.A(n_884),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_811),
.B(n_731),
.Y(n_962)
);

HB1xp67_ASAP7_75t_L g963 ( 
.A(n_881),
.Y(n_963)
);

BUFx2_ASAP7_75t_L g964 ( 
.A(n_887),
.Y(n_964)
);

INVxp67_ASAP7_75t_L g965 ( 
.A(n_892),
.Y(n_965)
);

INVxp67_ASAP7_75t_L g966 ( 
.A(n_917),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_829),
.Y(n_967)
);

INVx2_ASAP7_75t_L g968 ( 
.A(n_884),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_837),
.B(n_731),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_911),
.B(n_736),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_829),
.Y(n_971)
);

HB1xp67_ASAP7_75t_L g972 ( 
.A(n_887),
.Y(n_972)
);

OA21x2_ASAP7_75t_L g973 ( 
.A1(n_912),
.A2(n_514),
.B(n_488),
.Y(n_973)
);

BUFx3_ASAP7_75t_L g974 ( 
.A(n_834),
.Y(n_974)
);

BUFx6f_ASAP7_75t_L g975 ( 
.A(n_900),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_835),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_836),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_891),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_898),
.Y(n_979)
);

OAI22xp5_ASAP7_75t_SL g980 ( 
.A1(n_822),
.A2(n_657),
.B1(n_785),
.B2(n_645),
.Y(n_980)
);

AND2x4_ASAP7_75t_L g981 ( 
.A(n_832),
.B(n_650),
.Y(n_981)
);

INVx3_ASAP7_75t_L g982 ( 
.A(n_912),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_897),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_901),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_844),
.Y(n_985)
);

INVx2_ASAP7_75t_L g986 ( 
.A(n_900),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_902),
.Y(n_987)
);

INVx2_ASAP7_75t_L g988 ( 
.A(n_840),
.Y(n_988)
);

BUFx6f_ASAP7_75t_L g989 ( 
.A(n_841),
.Y(n_989)
);

NOR3xp33_ASAP7_75t_L g990 ( 
.A(n_821),
.B(n_758),
.C(n_549),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_839),
.B(n_738),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_905),
.Y(n_992)
);

NOR2xp33_ASAP7_75t_L g993 ( 
.A(n_877),
.B(n_501),
.Y(n_993)
);

HB1xp67_ASAP7_75t_L g994 ( 
.A(n_904),
.Y(n_994)
);

HB1xp67_ASAP7_75t_L g995 ( 
.A(n_904),
.Y(n_995)
);

INVx2_ASAP7_75t_L g996 ( 
.A(n_842),
.Y(n_996)
);

INVx2_ASAP7_75t_L g997 ( 
.A(n_843),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_906),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_907),
.Y(n_999)
);

INVx2_ASAP7_75t_L g1000 ( 
.A(n_845),
.Y(n_1000)
);

BUFx3_ASAP7_75t_L g1001 ( 
.A(n_846),
.Y(n_1001)
);

INVx2_ASAP7_75t_L g1002 ( 
.A(n_847),
.Y(n_1002)
);

AND2x2_ASAP7_75t_L g1003 ( 
.A(n_869),
.B(n_627),
.Y(n_1003)
);

AND2x2_ASAP7_75t_SL g1004 ( 
.A(n_920),
.B(n_503),
.Y(n_1004)
);

INVx2_ASAP7_75t_L g1005 ( 
.A(n_849),
.Y(n_1005)
);

BUFx8_ASAP7_75t_L g1006 ( 
.A(n_909),
.Y(n_1006)
);

AND2x2_ASAP7_75t_L g1007 ( 
.A(n_883),
.B(n_540),
.Y(n_1007)
);

BUFx2_ASAP7_75t_L g1008 ( 
.A(n_908),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_935),
.B(n_738),
.Y(n_1009)
);

INVx2_ASAP7_75t_L g1010 ( 
.A(n_851),
.Y(n_1010)
);

INVxp67_ASAP7_75t_L g1011 ( 
.A(n_908),
.Y(n_1011)
);

AND2x4_ASAP7_75t_L g1012 ( 
.A(n_903),
.B(n_651),
.Y(n_1012)
);

NOR2x1_ASAP7_75t_L g1013 ( 
.A(n_910),
.B(n_541),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_913),
.Y(n_1014)
);

OAI22xp5_ASAP7_75t_SL g1015 ( 
.A1(n_822),
.A2(n_785),
.B1(n_786),
.B2(n_657),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_937),
.B(n_743),
.Y(n_1016)
);

AND2x2_ASAP7_75t_L g1017 ( 
.A(n_896),
.B(n_540),
.Y(n_1017)
);

BUFx6f_ASAP7_75t_L g1018 ( 
.A(n_854),
.Y(n_1018)
);

INVx2_ASAP7_75t_L g1019 ( 
.A(n_855),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_914),
.B(n_743),
.Y(n_1020)
);

NOR2xp33_ASAP7_75t_L g1021 ( 
.A(n_916),
.B(n_512),
.Y(n_1021)
);

NOR2xp33_ASAP7_75t_L g1022 ( 
.A(n_921),
.B(n_629),
.Y(n_1022)
);

INVx6_ASAP7_75t_L g1023 ( 
.A(n_819),
.Y(n_1023)
);

AND2x4_ASAP7_75t_L g1024 ( 
.A(n_922),
.B(n_655),
.Y(n_1024)
);

AND2x2_ASAP7_75t_L g1025 ( 
.A(n_926),
.B(n_547),
.Y(n_1025)
);

AND2x4_ASAP7_75t_L g1026 ( 
.A(n_929),
.B(n_661),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_932),
.B(n_744),
.Y(n_1027)
);

INVx2_ASAP7_75t_L g1028 ( 
.A(n_856),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_933),
.Y(n_1029)
);

BUFx2_ASAP7_75t_L g1030 ( 
.A(n_919),
.Y(n_1030)
);

INVx2_ASAP7_75t_L g1031 ( 
.A(n_857),
.Y(n_1031)
);

INVx3_ASAP7_75t_L g1032 ( 
.A(n_859),
.Y(n_1032)
);

INVxp67_ASAP7_75t_L g1033 ( 
.A(n_919),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_934),
.B(n_744),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_936),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_860),
.B(n_746),
.Y(n_1036)
);

OA21x2_ASAP7_75t_L g1037 ( 
.A1(n_848),
.A2(n_514),
.B(n_488),
.Y(n_1037)
);

INVx2_ASAP7_75t_L g1038 ( 
.A(n_862),
.Y(n_1038)
);

BUFx2_ASAP7_75t_L g1039 ( 
.A(n_925),
.Y(n_1039)
);

INVx2_ASAP7_75t_L g1040 ( 
.A(n_863),
.Y(n_1040)
);

BUFx6f_ASAP7_75t_L g1041 ( 
.A(n_864),
.Y(n_1041)
);

AND2x2_ASAP7_75t_L g1042 ( 
.A(n_925),
.B(n_547),
.Y(n_1042)
);

BUFx12f_ASAP7_75t_L g1043 ( 
.A(n_817),
.Y(n_1043)
);

INVx2_ASAP7_75t_L g1044 ( 
.A(n_867),
.Y(n_1044)
);

OAI21x1_ASAP7_75t_L g1045 ( 
.A1(n_882),
.A2(n_609),
.B(n_603),
.Y(n_1045)
);

INVx2_ASAP7_75t_L g1046 ( 
.A(n_886),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_888),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_889),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_890),
.Y(n_1049)
);

INVx2_ASAP7_75t_L g1050 ( 
.A(n_871),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_893),
.Y(n_1051)
);

BUFx8_ASAP7_75t_L g1052 ( 
.A(n_808),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_924),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_918),
.Y(n_1054)
);

OA21x2_ASAP7_75t_L g1055 ( 
.A1(n_927),
.A2(n_609),
.B(n_603),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_930),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_SL g1057 ( 
.A(n_931),
.B(n_695),
.Y(n_1057)
);

HB1xp67_ASAP7_75t_L g1058 ( 
.A(n_823),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_SL g1059 ( 
.A(n_899),
.B(n_695),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_823),
.Y(n_1060)
);

BUFx8_ASAP7_75t_L g1061 ( 
.A(n_807),
.Y(n_1061)
);

INVx2_ASAP7_75t_L g1062 ( 
.A(n_818),
.Y(n_1062)
);

INVx2_ASAP7_75t_L g1063 ( 
.A(n_818),
.Y(n_1063)
);

NOR2xp33_ASAP7_75t_L g1064 ( 
.A(n_824),
.B(n_556),
.Y(n_1064)
);

INVx2_ASAP7_75t_L g1065 ( 
.A(n_825),
.Y(n_1065)
);

INVx2_ASAP7_75t_L g1066 ( 
.A(n_825),
.Y(n_1066)
);

INVx3_ASAP7_75t_L g1067 ( 
.A(n_827),
.Y(n_1067)
);

BUFx3_ASAP7_75t_L g1068 ( 
.A(n_833),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_827),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_831),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_831),
.Y(n_1071)
);

INVx2_ASAP7_75t_L g1072 ( 
.A(n_866),
.Y(n_1072)
);

INVx6_ASAP7_75t_L g1073 ( 
.A(n_838),
.Y(n_1073)
);

INVx3_ASAP7_75t_L g1074 ( 
.A(n_866),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_850),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_852),
.Y(n_1076)
);

AND2x6_ASAP7_75t_L g1077 ( 
.A(n_853),
.B(n_538),
.Y(n_1077)
);

AND2x4_ASAP7_75t_L g1078 ( 
.A(n_872),
.B(n_666),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_873),
.Y(n_1079)
);

OAI22xp5_ASAP7_75t_L g1080 ( 
.A1(n_876),
.A2(n_792),
.B1(n_796),
.B2(n_492),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_879),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_807),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_828),
.Y(n_1083)
);

INVx2_ASAP7_75t_L g1084 ( 
.A(n_828),
.Y(n_1084)
);

AND2x2_ASAP7_75t_L g1085 ( 
.A(n_858),
.B(n_547),
.Y(n_1085)
);

AND2x4_ASAP7_75t_L g1086 ( 
.A(n_928),
.B(n_668),
.Y(n_1086)
);

HB1xp67_ASAP7_75t_L g1087 ( 
.A(n_858),
.Y(n_1087)
);

AND2x2_ASAP7_75t_L g1088 ( 
.A(n_861),
.B(n_552),
.Y(n_1088)
);

INVx3_ASAP7_75t_L g1089 ( 
.A(n_865),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_865),
.B(n_796),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_895),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_868),
.B(n_797),
.Y(n_1092)
);

OR2x6_ASAP7_75t_L g1093 ( 
.A(n_868),
.B(n_546),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_875),
.Y(n_1094)
);

AO21x2_ASAP7_75t_L g1095 ( 
.A1(n_875),
.A2(n_563),
.B(n_561),
.Y(n_1095)
);

BUFx3_ASAP7_75t_L g1096 ( 
.A(n_878),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_895),
.Y(n_1097)
);

INVx2_ASAP7_75t_L g1098 ( 
.A(n_878),
.Y(n_1098)
);

BUFx2_ASAP7_75t_L g1099 ( 
.A(n_880),
.Y(n_1099)
);

INVx4_ASAP7_75t_L g1100 ( 
.A(n_880),
.Y(n_1100)
);

INVx2_ASAP7_75t_L g1101 ( 
.A(n_885),
.Y(n_1101)
);

AND2x4_ASAP7_75t_L g1102 ( 
.A(n_885),
.B(n_676),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_894),
.B(n_801),
.Y(n_1103)
);

BUFx6f_ASAP7_75t_L g1104 ( 
.A(n_894),
.Y(n_1104)
);

AND2x2_ASAP7_75t_L g1105 ( 
.A(n_870),
.B(n_552),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_803),
.B(n_801),
.Y(n_1106)
);

INVx5_ASAP7_75t_L g1107 ( 
.A(n_809),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_830),
.Y(n_1108)
);

BUFx6f_ASAP7_75t_L g1109 ( 
.A(n_830),
.Y(n_1109)
);

AND2x4_ASAP7_75t_L g1110 ( 
.A(n_803),
.B(n_679),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_803),
.B(n_519),
.Y(n_1111)
);

BUFx6f_ASAP7_75t_L g1112 ( 
.A(n_830),
.Y(n_1112)
);

INVx3_ASAP7_75t_L g1113 ( 
.A(n_830),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_803),
.B(n_519),
.Y(n_1114)
);

AND2x2_ASAP7_75t_L g1115 ( 
.A(n_870),
.B(n_552),
.Y(n_1115)
);

INVx3_ASAP7_75t_L g1116 ( 
.A(n_830),
.Y(n_1116)
);

INVx2_ASAP7_75t_L g1117 ( 
.A(n_874),
.Y(n_1117)
);

INVx2_ASAP7_75t_L g1118 ( 
.A(n_874),
.Y(n_1118)
);

BUFx6f_ASAP7_75t_L g1119 ( 
.A(n_830),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_SL g1120 ( 
.A(n_897),
.B(n_523),
.Y(n_1120)
);

INVx3_ASAP7_75t_L g1121 ( 
.A(n_830),
.Y(n_1121)
);

INVx2_ASAP7_75t_L g1122 ( 
.A(n_874),
.Y(n_1122)
);

AND2x2_ASAP7_75t_L g1123 ( 
.A(n_870),
.B(n_587),
.Y(n_1123)
);

BUFx6f_ASAP7_75t_L g1124 ( 
.A(n_830),
.Y(n_1124)
);

INVx2_ASAP7_75t_L g1125 ( 
.A(n_874),
.Y(n_1125)
);

CKINVDCx20_ASAP7_75t_R g1126 ( 
.A(n_822),
.Y(n_1126)
);

INVx2_ASAP7_75t_L g1127 ( 
.A(n_874),
.Y(n_1127)
);

INVx2_ASAP7_75t_L g1128 ( 
.A(n_874),
.Y(n_1128)
);

INVx2_ASAP7_75t_L g1129 ( 
.A(n_874),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_830),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_830),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_803),
.B(n_797),
.Y(n_1132)
);

HB1xp67_ASAP7_75t_L g1133 ( 
.A(n_923),
.Y(n_1133)
);

HB1xp67_ASAP7_75t_L g1134 ( 
.A(n_923),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_830),
.Y(n_1135)
);

BUFx6f_ASAP7_75t_L g1136 ( 
.A(n_830),
.Y(n_1136)
);

INVx2_ASAP7_75t_L g1137 ( 
.A(n_874),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_830),
.Y(n_1138)
);

AND2x2_ASAP7_75t_L g1139 ( 
.A(n_870),
.B(n_587),
.Y(n_1139)
);

AND2x2_ASAP7_75t_L g1140 ( 
.A(n_870),
.B(n_587),
.Y(n_1140)
);

AND2x2_ASAP7_75t_L g1141 ( 
.A(n_870),
.B(n_691),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_SL g1142 ( 
.A(n_897),
.B(n_523),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_803),
.B(n_521),
.Y(n_1143)
);

AND2x6_ASAP7_75t_L g1144 ( 
.A(n_830),
.B(n_538),
.Y(n_1144)
);

AOI22xp33_ASAP7_75t_L g1145 ( 
.A1(n_985),
.A2(n_792),
.B1(n_684),
.B2(n_685),
.Y(n_1145)
);

XOR2xp5_ASAP7_75t_L g1146 ( 
.A(n_1126),
.B(n_786),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_SL g1147 ( 
.A(n_978),
.B(n_791),
.Y(n_1147)
);

OAI21xp33_ASAP7_75t_SL g1148 ( 
.A1(n_1059),
.A2(n_693),
.B(n_683),
.Y(n_1148)
);

INVx2_ASAP7_75t_L g1149 ( 
.A(n_1045),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_944),
.Y(n_1150)
);

INVx2_ASAP7_75t_L g1151 ( 
.A(n_1045),
.Y(n_1151)
);

INVx2_ASAP7_75t_L g1152 ( 
.A(n_982),
.Y(n_1152)
);

BUFx3_ASAP7_75t_L g1153 ( 
.A(n_1109),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_946),
.Y(n_1154)
);

AOI22xp33_ASAP7_75t_L g1155 ( 
.A1(n_979),
.A2(n_732),
.B1(n_739),
.B2(n_718),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_947),
.Y(n_1156)
);

NOR2xp33_ASAP7_75t_L g1157 ( 
.A(n_1106),
.B(n_691),
.Y(n_1157)
);

BUFx2_ASAP7_75t_L g1158 ( 
.A(n_966),
.Y(n_1158)
);

XNOR2xp5_ASAP7_75t_L g1159 ( 
.A(n_1126),
.B(n_485),
.Y(n_1159)
);

HB1xp67_ASAP7_75t_L g1160 ( 
.A(n_1006),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_1111),
.B(n_521),
.Y(n_1161)
);

AND3x2_ASAP7_75t_L g1162 ( 
.A(n_964),
.B(n_752),
.C(n_740),
.Y(n_1162)
);

INVx2_ASAP7_75t_L g1163 ( 
.A(n_1109),
.Y(n_1163)
);

NAND2xp33_ASAP7_75t_SL g1164 ( 
.A(n_957),
.B(n_524),
.Y(n_1164)
);

AOI22xp33_ASAP7_75t_L g1165 ( 
.A1(n_1110),
.A2(n_761),
.B1(n_774),
.B2(n_760),
.Y(n_1165)
);

INVx3_ASAP7_75t_L g1166 ( 
.A(n_952),
.Y(n_1166)
);

NOR2xp33_ASAP7_75t_L g1167 ( 
.A(n_1114),
.B(n_691),
.Y(n_1167)
);

NOR2xp33_ASAP7_75t_L g1168 ( 
.A(n_1132),
.B(n_735),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_949),
.Y(n_1169)
);

INVx2_ASAP7_75t_L g1170 ( 
.A(n_1112),
.Y(n_1170)
);

INVx2_ASAP7_75t_SL g1171 ( 
.A(n_957),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_954),
.Y(n_1172)
);

AND2x4_ASAP7_75t_L g1173 ( 
.A(n_1025),
.B(n_775),
.Y(n_1173)
);

AOI22xp33_ASAP7_75t_L g1174 ( 
.A1(n_1110),
.A2(n_782),
.B1(n_783),
.B2(n_777),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_1143),
.B(n_524),
.Y(n_1175)
);

INVxp33_ASAP7_75t_L g1176 ( 
.A(n_1133),
.Y(n_1176)
);

BUFx6f_ASAP7_75t_L g1177 ( 
.A(n_1112),
.Y(n_1177)
);

AND2x6_ASAP7_75t_L g1178 ( 
.A(n_1025),
.B(n_678),
.Y(n_1178)
);

INVx2_ASAP7_75t_L g1179 ( 
.A(n_1119),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_962),
.B(n_725),
.Y(n_1180)
);

INVx2_ASAP7_75t_L g1181 ( 
.A(n_1119),
.Y(n_1181)
);

AND2x2_ASAP7_75t_L g1182 ( 
.A(n_959),
.B(n_496),
.Y(n_1182)
);

INVx2_ASAP7_75t_SL g1183 ( 
.A(n_1105),
.Y(n_1183)
);

NOR2xp33_ASAP7_75t_L g1184 ( 
.A(n_1054),
.B(n_735),
.Y(n_1184)
);

INVx2_ASAP7_75t_L g1185 ( 
.A(n_982),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_SL g1186 ( 
.A(n_1119),
.B(n_570),
.Y(n_1186)
);

BUFx6f_ASAP7_75t_L g1187 ( 
.A(n_1119),
.Y(n_1187)
);

XOR2xp5_ASAP7_75t_L g1188 ( 
.A(n_980),
.B(n_534),
.Y(n_1188)
);

INVx2_ASAP7_75t_L g1189 ( 
.A(n_982),
.Y(n_1189)
);

BUFx3_ASAP7_75t_L g1190 ( 
.A(n_1124),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_SL g1191 ( 
.A(n_1124),
.B(n_576),
.Y(n_1191)
);

INVx2_ASAP7_75t_SL g1192 ( 
.A(n_1105),
.Y(n_1192)
);

INVx2_ASAP7_75t_L g1193 ( 
.A(n_973),
.Y(n_1193)
);

INVx1_ASAP7_75t_SL g1194 ( 
.A(n_964),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_969),
.B(n_1056),
.Y(n_1195)
);

NOR2xp33_ASAP7_75t_L g1196 ( 
.A(n_1050),
.B(n_735),
.Y(n_1196)
);

NAND2xp33_ASAP7_75t_SL g1197 ( 
.A(n_1030),
.B(n_725),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_952),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_952),
.Y(n_1199)
);

BUFx3_ASAP7_75t_L g1200 ( 
.A(n_1124),
.Y(n_1200)
);

NOR2xp33_ASAP7_75t_L g1201 ( 
.A(n_1050),
.B(n_728),
.Y(n_1201)
);

INVx2_ASAP7_75t_L g1202 ( 
.A(n_973),
.Y(n_1202)
);

INVx5_ASAP7_75t_L g1203 ( 
.A(n_1144),
.Y(n_1203)
);

INVx2_ASAP7_75t_L g1204 ( 
.A(n_961),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_956),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_945),
.B(n_728),
.Y(n_1206)
);

INVx2_ASAP7_75t_L g1207 ( 
.A(n_961),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_958),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_960),
.Y(n_1209)
);

AOI22xp33_ASAP7_75t_L g1210 ( 
.A1(n_1110),
.A2(n_798),
.B1(n_793),
.B2(n_503),
.Y(n_1210)
);

BUFx6f_ASAP7_75t_L g1211 ( 
.A(n_1124),
.Y(n_1211)
);

INVx3_ASAP7_75t_L g1212 ( 
.A(n_1001),
.Y(n_1212)
);

INVx2_ASAP7_75t_L g1213 ( 
.A(n_961),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_967),
.Y(n_1214)
);

BUFx10_ASAP7_75t_L g1215 ( 
.A(n_938),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_971),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_974),
.Y(n_1217)
);

NOR2xp33_ASAP7_75t_L g1218 ( 
.A(n_951),
.B(n_730),
.Y(n_1218)
);

HB1xp67_ASAP7_75t_L g1219 ( 
.A(n_1006),
.Y(n_1219)
);

AND2x6_ASAP7_75t_L g1220 ( 
.A(n_1007),
.B(n_678),
.Y(n_1220)
);

BUFx2_ASAP7_75t_L g1221 ( 
.A(n_1030),
.Y(n_1221)
);

INVx2_ASAP7_75t_L g1222 ( 
.A(n_961),
.Y(n_1222)
);

INVx3_ASAP7_75t_L g1223 ( 
.A(n_1001),
.Y(n_1223)
);

BUFx6f_ASAP7_75t_L g1224 ( 
.A(n_1136),
.Y(n_1224)
);

OR2x6_ASAP7_75t_L g1225 ( 
.A(n_1093),
.B(n_503),
.Y(n_1225)
);

AND3x1_ASAP7_75t_L g1226 ( 
.A(n_990),
.B(n_590),
.C(n_577),
.Y(n_1226)
);

AOI22xp33_ASAP7_75t_L g1227 ( 
.A1(n_1024),
.A2(n_507),
.B1(n_734),
.B2(n_663),
.Y(n_1227)
);

BUFx3_ASAP7_75t_L g1228 ( 
.A(n_1136),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_SL g1229 ( 
.A(n_1136),
.B(n_599),
.Y(n_1229)
);

BUFx6f_ASAP7_75t_L g1230 ( 
.A(n_1136),
.Y(n_1230)
);

INVx2_ASAP7_75t_L g1231 ( 
.A(n_989),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_974),
.Y(n_1232)
);

BUFx4f_ASAP7_75t_L g1233 ( 
.A(n_938),
.Y(n_1233)
);

INVx2_ASAP7_75t_L g1234 ( 
.A(n_989),
.Y(n_1234)
);

INVxp67_ASAP7_75t_SL g1235 ( 
.A(n_1006),
.Y(n_1235)
);

INVx5_ASAP7_75t_L g1236 ( 
.A(n_1144),
.Y(n_1236)
);

NOR2xp33_ASAP7_75t_L g1237 ( 
.A(n_953),
.B(n_730),
.Y(n_1237)
);

INVx2_ASAP7_75t_L g1238 ( 
.A(n_989),
.Y(n_1238)
);

AND2x2_ASAP7_75t_L g1239 ( 
.A(n_1134),
.B(n_535),
.Y(n_1239)
);

AOI22xp33_ASAP7_75t_SL g1240 ( 
.A1(n_948),
.A2(n_544),
.B1(n_548),
.B2(n_537),
.Y(n_1240)
);

INVx2_ASAP7_75t_L g1241 ( 
.A(n_989),
.Y(n_1241)
);

CKINVDCx16_ASAP7_75t_R g1242 ( 
.A(n_1043),
.Y(n_1242)
);

AND2x6_ASAP7_75t_L g1243 ( 
.A(n_1007),
.B(n_699),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_L g1244 ( 
.A(n_953),
.B(n_742),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1113),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_SL g1246 ( 
.A(n_942),
.B(n_943),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1113),
.Y(n_1247)
);

BUFx3_ASAP7_75t_L g1248 ( 
.A(n_1144),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1113),
.Y(n_1249)
);

BUFx6f_ASAP7_75t_L g1250 ( 
.A(n_1018),
.Y(n_1250)
);

AND2x6_ASAP7_75t_L g1251 ( 
.A(n_1017),
.B(n_699),
.Y(n_1251)
);

INVx2_ASAP7_75t_L g1252 ( 
.A(n_975),
.Y(n_1252)
);

INVx5_ASAP7_75t_L g1253 ( 
.A(n_1144),
.Y(n_1253)
);

INVx2_ASAP7_75t_L g1254 ( 
.A(n_1018),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_SL g1255 ( 
.A(n_942),
.B(n_601),
.Y(n_1255)
);

NOR2xp33_ASAP7_75t_L g1256 ( 
.A(n_1059),
.B(n_742),
.Y(n_1256)
);

NOR2xp33_ASAP7_75t_L g1257 ( 
.A(n_993),
.B(n_613),
.Y(n_1257)
);

HB1xp67_ASAP7_75t_L g1258 ( 
.A(n_939),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_970),
.B(n_489),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1116),
.Y(n_1260)
);

BUFx6f_ASAP7_75t_L g1261 ( 
.A(n_1018),
.Y(n_1261)
);

INVx2_ASAP7_75t_L g1262 ( 
.A(n_1041),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_SL g1263 ( 
.A(n_943),
.B(n_624),
.Y(n_1263)
);

AOI22xp33_ASAP7_75t_L g1264 ( 
.A1(n_1024),
.A2(n_507),
.B1(n_734),
.B2(n_663),
.Y(n_1264)
);

BUFx2_ASAP7_75t_L g1265 ( 
.A(n_948),
.Y(n_1265)
);

AO22x2_ASAP7_75t_L g1266 ( 
.A1(n_1086),
.A2(n_520),
.B1(n_569),
.B2(n_550),
.Y(n_1266)
);

AOI22xp33_ASAP7_75t_SL g1267 ( 
.A1(n_948),
.A2(n_553),
.B1(n_558),
.B2(n_557),
.Y(n_1267)
);

AND2x2_ASAP7_75t_SL g1268 ( 
.A(n_1004),
.B(n_507),
.Y(n_1268)
);

HB1xp67_ASAP7_75t_L g1269 ( 
.A(n_939),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_SL g1270 ( 
.A(n_968),
.B(n_634),
.Y(n_1270)
);

NAND2xp33_ASAP7_75t_SL g1271 ( 
.A(n_1115),
.B(n_559),
.Y(n_1271)
);

AOI22xp5_ASAP7_75t_L g1272 ( 
.A1(n_1003),
.A2(n_565),
.B1(n_578),
.B2(n_572),
.Y(n_1272)
);

BUFx3_ASAP7_75t_L g1273 ( 
.A(n_1144),
.Y(n_1273)
);

AND2x2_ASAP7_75t_SL g1274 ( 
.A(n_1004),
.B(n_507),
.Y(n_1274)
);

AO22x2_ASAP7_75t_L g1275 ( 
.A1(n_1086),
.A2(n_594),
.B1(n_665),
.B2(n_596),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1116),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1121),
.Y(n_1277)
);

INVx2_ASAP7_75t_SL g1278 ( 
.A(n_1115),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1121),
.Y(n_1279)
);

HB1xp67_ASAP7_75t_L g1280 ( 
.A(n_1008),
.Y(n_1280)
);

OAI22xp33_ASAP7_75t_L g1281 ( 
.A1(n_1093),
.A2(n_584),
.B1(n_592),
.B2(n_591),
.Y(n_1281)
);

AND2x2_ASAP7_75t_L g1282 ( 
.A(n_1123),
.B(n_610),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1121),
.Y(n_1283)
);

INVx3_ASAP7_75t_L g1284 ( 
.A(n_1032),
.Y(n_1284)
);

INVx2_ASAP7_75t_L g1285 ( 
.A(n_975),
.Y(n_1285)
);

NOR2xp33_ASAP7_75t_L g1286 ( 
.A(n_993),
.B(n_635),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_L g1287 ( 
.A(n_1027),
.B(n_490),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1032),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1032),
.Y(n_1289)
);

INVx2_ASAP7_75t_SL g1290 ( 
.A(n_1123),
.Y(n_1290)
);

AO22x2_ASAP7_75t_L g1291 ( 
.A1(n_1086),
.A2(n_703),
.B1(n_712),
.B2(n_698),
.Y(n_1291)
);

CKINVDCx5p33_ASAP7_75t_R g1292 ( 
.A(n_1061),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1047),
.Y(n_1293)
);

NOR2xp33_ASAP7_75t_L g1294 ( 
.A(n_1017),
.B(n_642),
.Y(n_1294)
);

INVx3_ASAP7_75t_L g1295 ( 
.A(n_988),
.Y(n_1295)
);

AND2x6_ASAP7_75t_L g1296 ( 
.A(n_1139),
.B(n_700),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_SL g1297 ( 
.A(n_968),
.B(n_644),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1048),
.Y(n_1298)
);

BUFx6f_ASAP7_75t_L g1299 ( 
.A(n_1037),
.Y(n_1299)
);

OAI22xp33_ASAP7_75t_L g1300 ( 
.A1(n_1093),
.A2(n_617),
.B1(n_628),
.B2(n_621),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1049),
.Y(n_1301)
);

CKINVDCx20_ASAP7_75t_R g1302 ( 
.A(n_1015),
.Y(n_1302)
);

INVx2_ASAP7_75t_SL g1303 ( 
.A(n_1139),
.Y(n_1303)
);

INVx2_ASAP7_75t_L g1304 ( 
.A(n_986),
.Y(n_1304)
);

INVx2_ASAP7_75t_L g1305 ( 
.A(n_986),
.Y(n_1305)
);

INVx2_ASAP7_75t_L g1306 ( 
.A(n_1117),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_955),
.Y(n_1307)
);

INVx2_ASAP7_75t_SL g1308 ( 
.A(n_1140),
.Y(n_1308)
);

NOR2xp33_ASAP7_75t_L g1309 ( 
.A(n_1034),
.B(n_1020),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_SL g1310 ( 
.A(n_1117),
.B(n_646),
.Y(n_1310)
);

OAI22xp33_ASAP7_75t_SL g1311 ( 
.A1(n_1093),
.A2(n_636),
.B1(n_637),
.B2(n_633),
.Y(n_1311)
);

INVx2_ASAP7_75t_L g1312 ( 
.A(n_1118),
.Y(n_1312)
);

INVx2_ASAP7_75t_L g1313 ( 
.A(n_1118),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_SL g1314 ( 
.A(n_1122),
.B(n_653),
.Y(n_1314)
);

NOR2xp33_ASAP7_75t_L g1315 ( 
.A(n_1023),
.B(n_664),
.Y(n_1315)
);

BUFx8_ASAP7_75t_SL g1316 ( 
.A(n_1099),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_L g1317 ( 
.A(n_1024),
.B(n_491),
.Y(n_1317)
);

INVx1_ASAP7_75t_SL g1318 ( 
.A(n_1039),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_L g1319 ( 
.A(n_1026),
.B(n_987),
.Y(n_1319)
);

NOR2xp33_ASAP7_75t_L g1320 ( 
.A(n_1023),
.B(n_1026),
.Y(n_1320)
);

AND2x6_ASAP7_75t_L g1321 ( 
.A(n_1140),
.B(n_700),
.Y(n_1321)
);

AOI22xp33_ASAP7_75t_L g1322 ( 
.A1(n_1026),
.A2(n_734),
.B1(n_778),
.B2(n_663),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_988),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_L g1324 ( 
.A(n_992),
.B(n_493),
.Y(n_1324)
);

INVx2_ASAP7_75t_SL g1325 ( 
.A(n_1141),
.Y(n_1325)
);

NAND2xp5_ASAP7_75t_SL g1326 ( 
.A(n_1122),
.B(n_672),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_996),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_996),
.Y(n_1328)
);

NAND2xp5_ASAP7_75t_SL g1329 ( 
.A(n_1125),
.B(n_681),
.Y(n_1329)
);

NAND2xp5_ASAP7_75t_L g1330 ( 
.A(n_998),
.B(n_495),
.Y(n_1330)
);

NAND2xp5_ASAP7_75t_SL g1331 ( 
.A(n_1125),
.B(n_705),
.Y(n_1331)
);

CKINVDCx20_ASAP7_75t_R g1332 ( 
.A(n_1061),
.Y(n_1332)
);

AND2x4_ASAP7_75t_L g1333 ( 
.A(n_1141),
.B(n_729),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_997),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_997),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_SL g1336 ( 
.A(n_1127),
.B(n_707),
.Y(n_1336)
);

INVx2_ASAP7_75t_L g1337 ( 
.A(n_1000),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1000),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_L g1339 ( 
.A(n_999),
.B(n_499),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_L g1340 ( 
.A(n_1014),
.B(n_1029),
.Y(n_1340)
);

NAND2xp5_ASAP7_75t_L g1341 ( 
.A(n_1035),
.B(n_527),
.Y(n_1341)
);

INVx2_ASAP7_75t_L g1342 ( 
.A(n_1002),
.Y(n_1342)
);

AOI22xp33_ASAP7_75t_L g1343 ( 
.A1(n_1037),
.A2(n_663),
.B1(n_778),
.B2(n_734),
.Y(n_1343)
);

INVx2_ASAP7_75t_SL g1344 ( 
.A(n_1023),
.Y(n_1344)
);

BUFx6f_ASAP7_75t_L g1345 ( 
.A(n_1037),
.Y(n_1345)
);

NAND2xp5_ASAP7_75t_L g1346 ( 
.A(n_1021),
.B(n_536),
.Y(n_1346)
);

NOR2xp33_ASAP7_75t_L g1347 ( 
.A(n_1009),
.B(n_711),
.Y(n_1347)
);

AND2x2_ASAP7_75t_L g1348 ( 
.A(n_965),
.B(n_639),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1002),
.Y(n_1349)
);

NAND2xp5_ASAP7_75t_SL g1350 ( 
.A(n_1128),
.B(n_1129),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1005),
.Y(n_1351)
);

AO22x2_ASAP7_75t_L g1352 ( 
.A1(n_1102),
.A2(n_1100),
.B1(n_1012),
.B2(n_1053),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1005),
.Y(n_1353)
);

AOI22xp33_ASAP7_75t_L g1354 ( 
.A1(n_1055),
.A2(n_950),
.B1(n_1019),
.B2(n_1010),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_SL g1355 ( 
.A(n_1128),
.B(n_723),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1010),
.Y(n_1356)
);

NOR2xp33_ASAP7_75t_L g1357 ( 
.A(n_1016),
.B(n_756),
.Y(n_1357)
);

AND2x2_ASAP7_75t_L g1358 ( 
.A(n_1003),
.B(n_1042),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1019),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_L g1360 ( 
.A(n_1021),
.B(n_543),
.Y(n_1360)
);

INVx2_ASAP7_75t_L g1361 ( 
.A(n_1028),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1028),
.Y(n_1362)
);

NAND2xp5_ASAP7_75t_L g1363 ( 
.A(n_1022),
.B(n_545),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_SL g1364 ( 
.A(n_1129),
.B(n_523),
.Y(n_1364)
);

INVx11_ASAP7_75t_L g1365 ( 
.A(n_1052),
.Y(n_1365)
);

INVx3_ASAP7_75t_L g1366 ( 
.A(n_1031),
.Y(n_1366)
);

INVx2_ASAP7_75t_L g1367 ( 
.A(n_1031),
.Y(n_1367)
);

INVx3_ASAP7_75t_L g1368 ( 
.A(n_1038),
.Y(n_1368)
);

OR2x6_ASAP7_75t_L g1369 ( 
.A(n_1043),
.B(n_778),
.Y(n_1369)
);

CKINVDCx20_ASAP7_75t_R g1370 ( 
.A(n_1068),
.Y(n_1370)
);

INVx3_ASAP7_75t_L g1371 ( 
.A(n_1038),
.Y(n_1371)
);

BUFx6f_ASAP7_75t_L g1372 ( 
.A(n_1055),
.Y(n_1372)
);

INVxp67_ASAP7_75t_SL g1373 ( 
.A(n_941),
.Y(n_1373)
);

INVx3_ASAP7_75t_L g1374 ( 
.A(n_1040),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_SL g1375 ( 
.A(n_1137),
.B(n_983),
.Y(n_1375)
);

NAND2xp33_ASAP7_75t_R g1376 ( 
.A(n_1067),
.B(n_640),
.Y(n_1376)
);

INVx2_ASAP7_75t_SL g1377 ( 
.A(n_1042),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1040),
.Y(n_1378)
);

NOR2xp33_ASAP7_75t_L g1379 ( 
.A(n_1036),
.B(n_494),
.Y(n_1379)
);

OAI22xp5_ASAP7_75t_L g1380 ( 
.A1(n_991),
.A2(n_659),
.B1(n_660),
.B2(n_643),
.Y(n_1380)
);

AND2x2_ASAP7_75t_L g1381 ( 
.A(n_963),
.B(n_972),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1044),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1044),
.Y(n_1383)
);

INVx2_ASAP7_75t_L g1384 ( 
.A(n_1046),
.Y(n_1384)
);

INVx2_ASAP7_75t_L g1385 ( 
.A(n_1046),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_976),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_977),
.Y(n_1387)
);

BUFx3_ASAP7_75t_L g1388 ( 
.A(n_1077),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_SL g1389 ( 
.A(n_1137),
.B(n_523),
.Y(n_1389)
);

NAND2xp5_ASAP7_75t_L g1390 ( 
.A(n_940),
.B(n_551),
.Y(n_1390)
);

BUFx10_ASAP7_75t_L g1391 ( 
.A(n_1064),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1108),
.Y(n_1392)
);

INVx2_ASAP7_75t_L g1393 ( 
.A(n_1107),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_SL g1394 ( 
.A(n_984),
.B(n_1107),
.Y(n_1394)
);

INVx3_ASAP7_75t_L g1395 ( 
.A(n_1107),
.Y(n_1395)
);

OR2x2_ASAP7_75t_L g1396 ( 
.A(n_1090),
.B(n_788),
.Y(n_1396)
);

BUFx2_ASAP7_75t_L g1397 ( 
.A(n_994),
.Y(n_1397)
);

AOI22xp33_ASAP7_75t_L g1398 ( 
.A1(n_1358),
.A2(n_1095),
.B1(n_1077),
.B2(n_1102),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_SL g1399 ( 
.A(n_1158),
.B(n_1011),
.Y(n_1399)
);

INVx2_ASAP7_75t_L g1400 ( 
.A(n_1284),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_L g1401 ( 
.A(n_1309),
.B(n_1055),
.Y(n_1401)
);

AND2x2_ASAP7_75t_L g1402 ( 
.A(n_1194),
.B(n_995),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1150),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1154),
.Y(n_1404)
);

OAI221xp5_ASAP7_75t_L g1405 ( 
.A1(n_1145),
.A2(n_1080),
.B1(n_1092),
.B2(n_1103),
.C(n_1033),
.Y(n_1405)
);

INVx2_ASAP7_75t_SL g1406 ( 
.A(n_1318),
.Y(n_1406)
);

INVx2_ASAP7_75t_L g1407 ( 
.A(n_1284),
.Y(n_1407)
);

INVxp67_ASAP7_75t_SL g1408 ( 
.A(n_1280),
.Y(n_1408)
);

O2A1O1Ixp33_ASAP7_75t_L g1409 ( 
.A1(n_1195),
.A2(n_1065),
.B(n_1072),
.C(n_1066),
.Y(n_1409)
);

BUFx6f_ASAP7_75t_SL g1410 ( 
.A(n_1369),
.Y(n_1410)
);

INVx2_ASAP7_75t_L g1411 ( 
.A(n_1212),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_L g1412 ( 
.A(n_1309),
.B(n_1013),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_L g1413 ( 
.A(n_1319),
.B(n_1095),
.Y(n_1413)
);

INVxp67_ASAP7_75t_L g1414 ( 
.A(n_1280),
.Y(n_1414)
);

NOR2xp67_ASAP7_75t_L g1415 ( 
.A(n_1292),
.B(n_1058),
.Y(n_1415)
);

INVx2_ASAP7_75t_L g1416 ( 
.A(n_1212),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1156),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_L g1418 ( 
.A(n_1169),
.B(n_1172),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1340),
.Y(n_1419)
);

INVx2_ASAP7_75t_L g1420 ( 
.A(n_1223),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_SL g1421 ( 
.A(n_1388),
.B(n_1065),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_SL g1422 ( 
.A(n_1388),
.B(n_1203),
.Y(n_1422)
);

NAND2xp5_ASAP7_75t_L g1423 ( 
.A(n_1307),
.B(n_1095),
.Y(n_1423)
);

NAND2xp5_ASAP7_75t_L g1424 ( 
.A(n_1386),
.B(n_950),
.Y(n_1424)
);

INVx2_ASAP7_75t_L g1425 ( 
.A(n_1223),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1387),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1293),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1298),
.Y(n_1428)
);

NAND2xp5_ASAP7_75t_SL g1429 ( 
.A(n_1203),
.B(n_1066),
.Y(n_1429)
);

NAND2xp5_ASAP7_75t_L g1430 ( 
.A(n_1178),
.B(n_1173),
.Y(n_1430)
);

NAND2xp5_ASAP7_75t_L g1431 ( 
.A(n_1178),
.B(n_950),
.Y(n_1431)
);

AND2x2_ASAP7_75t_L g1432 ( 
.A(n_1221),
.B(n_1085),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_L g1433 ( 
.A(n_1178),
.B(n_950),
.Y(n_1433)
);

CKINVDCx5p33_ASAP7_75t_R g1434 ( 
.A(n_1365),
.Y(n_1434)
);

NOR2xp33_ASAP7_75t_L g1435 ( 
.A(n_1176),
.B(n_1060),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_L g1436 ( 
.A(n_1178),
.B(n_950),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1301),
.Y(n_1437)
);

AND2x4_ASAP7_75t_L g1438 ( 
.A(n_1235),
.B(n_1072),
.Y(n_1438)
);

NAND2xp5_ASAP7_75t_L g1439 ( 
.A(n_1173),
.B(n_1064),
.Y(n_1439)
);

INVx2_ASAP7_75t_L g1440 ( 
.A(n_1295),
.Y(n_1440)
);

BUFx3_ASAP7_75t_L g1441 ( 
.A(n_1332),
.Y(n_1441)
);

INVx2_ASAP7_75t_L g1442 ( 
.A(n_1295),
.Y(n_1442)
);

INVxp33_ASAP7_75t_L g1443 ( 
.A(n_1176),
.Y(n_1443)
);

NOR2xp33_ASAP7_75t_L g1444 ( 
.A(n_1377),
.B(n_1069),
.Y(n_1444)
);

NAND2x1p5_ASAP7_75t_L g1445 ( 
.A(n_1233),
.B(n_1067),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_SL g1446 ( 
.A(n_1203),
.B(n_1067),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1205),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1208),
.Y(n_1448)
);

INVx2_ASAP7_75t_L g1449 ( 
.A(n_1366),
.Y(n_1449)
);

NAND2xp5_ASAP7_75t_L g1450 ( 
.A(n_1201),
.B(n_981),
.Y(n_1450)
);

NAND2xp5_ASAP7_75t_L g1451 ( 
.A(n_1201),
.B(n_981),
.Y(n_1451)
);

INVx2_ASAP7_75t_L g1452 ( 
.A(n_1366),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1209),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1214),
.Y(n_1454)
);

AOI22xp5_ASAP7_75t_L g1455 ( 
.A1(n_1182),
.A2(n_1070),
.B1(n_1071),
.B2(n_1078),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1216),
.Y(n_1456)
);

BUFx3_ASAP7_75t_L g1457 ( 
.A(n_1265),
.Y(n_1457)
);

INVxp67_ASAP7_75t_SL g1458 ( 
.A(n_1248),
.Y(n_1458)
);

BUFx5_ASAP7_75t_L g1459 ( 
.A(n_1248),
.Y(n_1459)
);

NOR2xp33_ASAP7_75t_L g1460 ( 
.A(n_1183),
.B(n_1075),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_L g1461 ( 
.A(n_1210),
.B(n_1057),
.Y(n_1461)
);

NAND2xp5_ASAP7_75t_L g1462 ( 
.A(n_1210),
.B(n_1057),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1392),
.Y(n_1463)
);

NAND2xp5_ASAP7_75t_SL g1464 ( 
.A(n_1236),
.B(n_1074),
.Y(n_1464)
);

NAND2xp5_ASAP7_75t_L g1465 ( 
.A(n_1165),
.B(n_1130),
.Y(n_1465)
);

INVx2_ASAP7_75t_SL g1466 ( 
.A(n_1258),
.Y(n_1466)
);

NAND2xp5_ASAP7_75t_L g1467 ( 
.A(n_1165),
.B(n_1131),
.Y(n_1467)
);

AND2x4_ASAP7_75t_L g1468 ( 
.A(n_1160),
.B(n_1219),
.Y(n_1468)
);

NOR2xp33_ASAP7_75t_L g1469 ( 
.A(n_1192),
.B(n_1076),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_L g1470 ( 
.A(n_1174),
.B(n_1135),
.Y(n_1470)
);

NOR2xp33_ASAP7_75t_L g1471 ( 
.A(n_1278),
.B(n_1079),
.Y(n_1471)
);

NOR2xp33_ASAP7_75t_L g1472 ( 
.A(n_1290),
.B(n_1303),
.Y(n_1472)
);

INVx2_ASAP7_75t_SL g1473 ( 
.A(n_1258),
.Y(n_1473)
);

INVx2_ASAP7_75t_L g1474 ( 
.A(n_1368),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_L g1475 ( 
.A(n_1174),
.B(n_1138),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1288),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_L g1477 ( 
.A(n_1294),
.B(n_981),
.Y(n_1477)
);

NAND3xp33_ASAP7_75t_L g1478 ( 
.A(n_1218),
.B(n_1088),
.C(n_1085),
.Y(n_1478)
);

BUFx6f_ASAP7_75t_L g1479 ( 
.A(n_1273),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_L g1480 ( 
.A(n_1294),
.B(n_1012),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_SL g1481 ( 
.A(n_1236),
.B(n_1078),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1289),
.Y(n_1482)
);

NAND3xp33_ASAP7_75t_L g1483 ( 
.A(n_1145),
.B(n_1088),
.C(n_1081),
.Y(n_1483)
);

AND2x4_ASAP7_75t_L g1484 ( 
.A(n_1160),
.B(n_1012),
.Y(n_1484)
);

INVx1_ASAP7_75t_SL g1485 ( 
.A(n_1397),
.Y(n_1485)
);

A2O1A1Ixp33_ASAP7_75t_L g1486 ( 
.A1(n_1257),
.A2(n_1120),
.B(n_1142),
.C(n_1051),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1368),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1371),
.Y(n_1488)
);

INVx4_ASAP7_75t_L g1489 ( 
.A(n_1225),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1371),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1374),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_L g1492 ( 
.A(n_1220),
.B(n_1077),
.Y(n_1492)
);

INVx3_ASAP7_75t_L g1493 ( 
.A(n_1166),
.Y(n_1493)
);

OAI22xp33_ASAP7_75t_L g1494 ( 
.A1(n_1225),
.A2(n_1219),
.B1(n_1100),
.B2(n_1233),
.Y(n_1494)
);

INVx2_ASAP7_75t_L g1495 ( 
.A(n_1374),
.Y(n_1495)
);

AND2x2_ASAP7_75t_L g1496 ( 
.A(n_1381),
.B(n_1102),
.Y(n_1496)
);

AND2x4_ASAP7_75t_L g1497 ( 
.A(n_1225),
.B(n_1077),
.Y(n_1497)
);

INVx2_ASAP7_75t_L g1498 ( 
.A(n_1153),
.Y(n_1498)
);

AOI22xp5_ASAP7_75t_L g1499 ( 
.A1(n_1268),
.A2(n_1077),
.B1(n_1073),
.B2(n_1063),
.Y(n_1499)
);

NOR2xp33_ASAP7_75t_L g1500 ( 
.A(n_1308),
.B(n_1062),
.Y(n_1500)
);

INVx2_ASAP7_75t_L g1501 ( 
.A(n_1153),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1323),
.Y(n_1502)
);

NOR2xp33_ASAP7_75t_L g1503 ( 
.A(n_1325),
.B(n_1062),
.Y(n_1503)
);

INVx2_ASAP7_75t_L g1504 ( 
.A(n_1190),
.Y(n_1504)
);

INVx2_ASAP7_75t_L g1505 ( 
.A(n_1190),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1327),
.Y(n_1506)
);

NAND2xp5_ASAP7_75t_SL g1507 ( 
.A(n_1253),
.B(n_1273),
.Y(n_1507)
);

NOR2xp33_ASAP7_75t_L g1508 ( 
.A(n_1171),
.B(n_1282),
.Y(n_1508)
);

NOR2xp33_ASAP7_75t_L g1509 ( 
.A(n_1391),
.B(n_1063),
.Y(n_1509)
);

AOI22xp33_ASAP7_75t_L g1510 ( 
.A1(n_1268),
.A2(n_1142),
.B1(n_1120),
.B2(n_1098),
.Y(n_1510)
);

BUFx6f_ASAP7_75t_L g1511 ( 
.A(n_1253),
.Y(n_1511)
);

INVx2_ASAP7_75t_L g1512 ( 
.A(n_1200),
.Y(n_1512)
);

OAI21xp33_ASAP7_75t_L g1513 ( 
.A1(n_1196),
.A2(n_1286),
.B(n_1257),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_L g1514 ( 
.A(n_1220),
.B(n_1107),
.Y(n_1514)
);

INVx2_ASAP7_75t_L g1515 ( 
.A(n_1200),
.Y(n_1515)
);

NAND2xp5_ASAP7_75t_L g1516 ( 
.A(n_1220),
.B(n_667),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1328),
.Y(n_1517)
);

NAND2xp5_ASAP7_75t_L g1518 ( 
.A(n_1243),
.B(n_671),
.Y(n_1518)
);

AO221x1_ASAP7_75t_L g1519 ( 
.A1(n_1281),
.A2(n_1300),
.B1(n_1266),
.B2(n_1291),
.C(n_1275),
.Y(n_1519)
);

INVxp67_ASAP7_75t_L g1520 ( 
.A(n_1269),
.Y(n_1520)
);

NAND2xp5_ASAP7_75t_L g1521 ( 
.A(n_1243),
.B(n_675),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_L g1522 ( 
.A(n_1243),
.B(n_677),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_SL g1523 ( 
.A(n_1253),
.B(n_554),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1334),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_L g1525 ( 
.A(n_1243),
.B(n_1251),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_SL g1526 ( 
.A(n_1197),
.B(n_560),
.Y(n_1526)
);

INVx2_ASAP7_75t_L g1527 ( 
.A(n_1228),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1251),
.B(n_682),
.Y(n_1528)
);

INVx2_ASAP7_75t_L g1529 ( 
.A(n_1228),
.Y(n_1529)
);

NOR3xp33_ASAP7_75t_L g1530 ( 
.A(n_1300),
.B(n_1089),
.C(n_1083),
.Y(n_1530)
);

OAI22xp5_ASAP7_75t_L g1531 ( 
.A1(n_1354),
.A2(n_1098),
.B1(n_1101),
.B2(n_1084),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1335),
.Y(n_1532)
);

AOI22xp5_ASAP7_75t_L g1533 ( 
.A1(n_1274),
.A2(n_1373),
.B1(n_1348),
.B2(n_1320),
.Y(n_1533)
);

INVx2_ASAP7_75t_L g1534 ( 
.A(n_1304),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_SL g1535 ( 
.A(n_1333),
.B(n_564),
.Y(n_1535)
);

AOI22xp33_ASAP7_75t_L g1536 ( 
.A1(n_1274),
.A2(n_1091),
.B1(n_1097),
.B2(n_1094),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1338),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_SL g1538 ( 
.A(n_1244),
.B(n_566),
.Y(n_1538)
);

BUFx6f_ASAP7_75t_L g1539 ( 
.A(n_1299),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1349),
.Y(n_1540)
);

AND2x2_ASAP7_75t_L g1541 ( 
.A(n_1269),
.B(n_1096),
.Y(n_1541)
);

NOR2xp33_ASAP7_75t_L g1542 ( 
.A(n_1396),
.B(n_1089),
.Y(n_1542)
);

AOI22xp5_ASAP7_75t_L g1543 ( 
.A1(n_1320),
.A2(n_689),
.B1(n_690),
.B2(n_688),
.Y(n_1543)
);

NOR2xp33_ASAP7_75t_L g1544 ( 
.A(n_1239),
.B(n_1087),
.Y(n_1544)
);

OAI22xp33_ASAP7_75t_SL g1545 ( 
.A1(n_1369),
.A2(n_1096),
.B1(n_694),
.B2(n_702),
.Y(n_1545)
);

NOR2xp67_ASAP7_75t_SL g1546 ( 
.A(n_1242),
.B(n_692),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1351),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_L g1548 ( 
.A(n_1251),
.B(n_708),
.Y(n_1548)
);

INVx2_ASAP7_75t_L g1549 ( 
.A(n_1305),
.Y(n_1549)
);

NOR2xp33_ASAP7_75t_L g1550 ( 
.A(n_1272),
.B(n_1104),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_L g1551 ( 
.A(n_1251),
.B(n_1286),
.Y(n_1551)
);

NOR2xp33_ASAP7_75t_L g1552 ( 
.A(n_1271),
.B(n_1104),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1353),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1251),
.B(n_709),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1356),
.Y(n_1555)
);

BUFx6f_ASAP7_75t_L g1556 ( 
.A(n_1299),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_L g1557 ( 
.A(n_1347),
.B(n_710),
.Y(n_1557)
);

NOR2xp33_ASAP7_75t_L g1558 ( 
.A(n_1164),
.B(n_1104),
.Y(n_1558)
);

INVx3_ASAP7_75t_L g1559 ( 
.A(n_1166),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1359),
.Y(n_1560)
);

NAND2xp5_ASAP7_75t_SL g1561 ( 
.A(n_1311),
.B(n_1237),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1362),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_L g1563 ( 
.A(n_1357),
.B(n_1378),
.Y(n_1563)
);

NAND2xp33_ASAP7_75t_L g1564 ( 
.A(n_1296),
.B(n_1321),
.Y(n_1564)
);

BUFx6f_ASAP7_75t_L g1565 ( 
.A(n_1299),
.Y(n_1565)
);

INVx2_ASAP7_75t_L g1566 ( 
.A(n_1306),
.Y(n_1566)
);

INVx2_ASAP7_75t_L g1567 ( 
.A(n_1306),
.Y(n_1567)
);

OAI221xp5_ASAP7_75t_L g1568 ( 
.A1(n_1155),
.A2(n_713),
.B1(n_750),
.B2(n_748),
.C(n_720),
.Y(n_1568)
);

CKINVDCx5p33_ASAP7_75t_R g1569 ( 
.A(n_1316),
.Y(n_1569)
);

INVx1_ASAP7_75t_SL g1570 ( 
.A(n_1370),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1382),
.Y(n_1571)
);

NAND2xp5_ASAP7_75t_L g1572 ( 
.A(n_1196),
.B(n_753),
.Y(n_1572)
);

INVx3_ASAP7_75t_L g1573 ( 
.A(n_1395),
.Y(n_1573)
);

AND2x2_ASAP7_75t_L g1574 ( 
.A(n_1266),
.B(n_1082),
.Y(n_1574)
);

NOR2xp67_ASAP7_75t_L g1575 ( 
.A(n_1148),
.B(n_1052),
.Y(n_1575)
);

AOI22xp33_ASAP7_75t_L g1576 ( 
.A1(n_1275),
.A2(n_1291),
.B1(n_1321),
.B2(n_1296),
.Y(n_1576)
);

NAND2xp5_ASAP7_75t_L g1577 ( 
.A(n_1379),
.B(n_1357),
.Y(n_1577)
);

NOR2xp33_ASAP7_75t_L g1578 ( 
.A(n_1184),
.B(n_1052),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_L g1579 ( 
.A(n_1379),
.B(n_802),
.Y(n_1579)
);

AOI22xp33_ASAP7_75t_L g1580 ( 
.A1(n_1275),
.A2(n_778),
.B1(n_765),
.B2(n_767),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_L g1581 ( 
.A(n_1206),
.B(n_795),
.Y(n_1581)
);

AOI221xp5_ASAP7_75t_L g1582 ( 
.A1(n_1291),
.A2(n_776),
.B1(n_780),
.B2(n_770),
.C(n_759),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_L g1583 ( 
.A(n_1383),
.B(n_784),
.Y(n_1583)
);

BUFx6f_ASAP7_75t_SL g1584 ( 
.A(n_1369),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1198),
.Y(n_1585)
);

INVx4_ASAP7_75t_L g1586 ( 
.A(n_1296),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1199),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_SL g1588 ( 
.A(n_1215),
.B(n_567),
.Y(n_1588)
);

BUFx6f_ASAP7_75t_SL g1589 ( 
.A(n_1296),
.Y(n_1589)
);

OR2x2_ASAP7_75t_L g1590 ( 
.A(n_1146),
.B(n_789),
.Y(n_1590)
);

NOR2xp33_ASAP7_75t_L g1591 ( 
.A(n_1184),
.B(n_1344),
.Y(n_1591)
);

INVx2_ASAP7_75t_SL g1592 ( 
.A(n_1162),
.Y(n_1592)
);

BUFx3_ASAP7_75t_L g1593 ( 
.A(n_1393),
.Y(n_1593)
);

BUFx5_ASAP7_75t_L g1594 ( 
.A(n_1245),
.Y(n_1594)
);

INVx2_ASAP7_75t_L g1595 ( 
.A(n_1312),
.Y(n_1595)
);

INVx2_ASAP7_75t_SL g1596 ( 
.A(n_1162),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_SL g1597 ( 
.A(n_1215),
.B(n_573),
.Y(n_1597)
);

NOR2xp33_ASAP7_75t_L g1598 ( 
.A(n_1380),
.B(n_794),
.Y(n_1598)
);

BUFx6f_ASAP7_75t_L g1599 ( 
.A(n_1345),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1217),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1232),
.Y(n_1601)
);

OAI22xp5_ASAP7_75t_L g1602 ( 
.A1(n_1193),
.A2(n_579),
.B1(n_582),
.B2(n_574),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1202),
.B(n_787),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1345),
.B(n_1372),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1337),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_SL g1606 ( 
.A(n_1161),
.B(n_583),
.Y(n_1606)
);

INVx3_ASAP7_75t_L g1607 ( 
.A(n_1395),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_SL g1608 ( 
.A(n_1175),
.B(n_585),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1180),
.B(n_598),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_L g1610 ( 
.A(n_1157),
.B(n_600),
.Y(n_1610)
);

AND2x2_ASAP7_75t_L g1611 ( 
.A(n_1240),
.B(n_11),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1157),
.B(n_604),
.Y(n_1612)
);

INVx8_ASAP7_75t_L g1613 ( 
.A(n_1321),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_SL g1614 ( 
.A(n_1317),
.B(n_605),
.Y(n_1614)
);

O2A1O1Ixp33_ASAP7_75t_L g1615 ( 
.A1(n_1147),
.A2(n_680),
.B(n_719),
.C(n_649),
.Y(n_1615)
);

AOI22xp33_ASAP7_75t_L g1616 ( 
.A1(n_1321),
.A2(n_787),
.B1(n_608),
.B2(n_612),
.Y(n_1616)
);

INVx3_ASAP7_75t_L g1617 ( 
.A(n_1342),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1361),
.Y(n_1618)
);

BUFx3_ASAP7_75t_L g1619 ( 
.A(n_1352),
.Y(n_1619)
);

OR2x2_ASAP7_75t_L g1620 ( 
.A(n_1159),
.B(n_1188),
.Y(n_1620)
);

BUFx3_ASAP7_75t_L g1621 ( 
.A(n_1352),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_SL g1622 ( 
.A(n_1287),
.B(n_607),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1367),
.Y(n_1623)
);

NOR2xp67_ASAP7_75t_L g1624 ( 
.A(n_1315),
.B(n_11),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1384),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_L g1626 ( 
.A(n_1345),
.B(n_787),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1267),
.B(n_12),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_SL g1628 ( 
.A(n_1259),
.B(n_616),
.Y(n_1628)
);

AND2x4_ASAP7_75t_SL g1629 ( 
.A(n_1302),
.B(n_510),
.Y(n_1629)
);

NAND3xp33_ASAP7_75t_L g1630 ( 
.A(n_1376),
.B(n_620),
.C(n_619),
.Y(n_1630)
);

INVx8_ASAP7_75t_L g1631 ( 
.A(n_1345),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1385),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_L g1633 ( 
.A(n_1372),
.B(n_787),
.Y(n_1633)
);

INVx2_ASAP7_75t_SL g1634 ( 
.A(n_1147),
.Y(n_1634)
);

INVx2_ASAP7_75t_SL g1635 ( 
.A(n_1255),
.Y(n_1635)
);

INVx2_ASAP7_75t_SL g1636 ( 
.A(n_1255),
.Y(n_1636)
);

HB1xp67_ASAP7_75t_L g1637 ( 
.A(n_1256),
.Y(n_1637)
);

INVx2_ASAP7_75t_L g1638 ( 
.A(n_1312),
.Y(n_1638)
);

INVx2_ASAP7_75t_SL g1639 ( 
.A(n_1263),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_L g1640 ( 
.A(n_1313),
.B(n_656),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_L g1641 ( 
.A(n_1313),
.B(n_658),
.Y(n_1641)
);

NAND2xp5_ASAP7_75t_SL g1642 ( 
.A(n_1324),
.B(n_662),
.Y(n_1642)
);

INVxp67_ASAP7_75t_L g1643 ( 
.A(n_1256),
.Y(n_1643)
);

NOR2xp33_ASAP7_75t_L g1644 ( 
.A(n_1167),
.B(n_669),
.Y(n_1644)
);

NOR2xp33_ASAP7_75t_L g1645 ( 
.A(n_1167),
.B(n_670),
.Y(n_1645)
);

BUFx6f_ASAP7_75t_L g1646 ( 
.A(n_1177),
.Y(n_1646)
);

AOI22xp33_ASAP7_75t_L g1647 ( 
.A1(n_1168),
.A2(n_1315),
.B1(n_1375),
.B2(n_1270),
.Y(n_1647)
);

AOI22xp5_ASAP7_75t_L g1648 ( 
.A1(n_1226),
.A2(n_674),
.B1(n_686),
.B2(n_673),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_SL g1649 ( 
.A(n_1330),
.B(n_687),
.Y(n_1649)
);

AND2x2_ASAP7_75t_L g1650 ( 
.A(n_1168),
.B(n_13),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1247),
.Y(n_1651)
);

INVx4_ASAP7_75t_L g1652 ( 
.A(n_1250),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_L g1653 ( 
.A(n_1149),
.B(n_701),
.Y(n_1653)
);

AND2x6_ASAP7_75t_SL g1654 ( 
.A(n_1346),
.B(n_13),
.Y(n_1654)
);

NAND2xp5_ASAP7_75t_L g1655 ( 
.A(n_1149),
.B(n_706),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1249),
.Y(n_1656)
);

INVx1_ASAP7_75t_SL g1657 ( 
.A(n_1339),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_L g1658 ( 
.A(n_1151),
.B(n_715),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_L g1659 ( 
.A(n_1151),
.B(n_741),
.Y(n_1659)
);

INVx2_ASAP7_75t_L g1660 ( 
.A(n_1152),
.Y(n_1660)
);

INVx3_ASAP7_75t_L g1661 ( 
.A(n_1489),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1419),
.Y(n_1662)
);

OAI21xp5_ASAP7_75t_L g1663 ( 
.A1(n_1401),
.A2(n_1604),
.B(n_1577),
.Y(n_1663)
);

NOR2xp33_ASAP7_75t_L g1664 ( 
.A(n_1478),
.B(n_1360),
.Y(n_1664)
);

NOR2xp33_ASAP7_75t_L g1665 ( 
.A(n_1485),
.B(n_1363),
.Y(n_1665)
);

AOI21xp5_ASAP7_75t_L g1666 ( 
.A1(n_1424),
.A2(n_1350),
.B(n_1246),
.Y(n_1666)
);

INVx3_ASAP7_75t_L g1667 ( 
.A(n_1489),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_SL g1668 ( 
.A(n_1406),
.B(n_1341),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1403),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_SL g1670 ( 
.A(n_1414),
.B(n_1494),
.Y(n_1670)
);

INVx2_ASAP7_75t_L g1671 ( 
.A(n_1404),
.Y(n_1671)
);

OAI21xp5_ASAP7_75t_L g1672 ( 
.A1(n_1604),
.A2(n_1343),
.B(n_1246),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_L g1673 ( 
.A(n_1418),
.B(n_1390),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_SL g1674 ( 
.A(n_1468),
.B(n_1227),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1417),
.Y(n_1675)
);

NOR2xp33_ASAP7_75t_L g1676 ( 
.A(n_1443),
.B(n_1394),
.Y(n_1676)
);

BUFx6f_ASAP7_75t_L g1677 ( 
.A(n_1631),
.Y(n_1677)
);

NOR2xp33_ASAP7_75t_L g1678 ( 
.A(n_1405),
.B(n_1394),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1426),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_L g1680 ( 
.A(n_1418),
.B(n_1513),
.Y(n_1680)
);

OAI22xp33_ASAP7_75t_L g1681 ( 
.A1(n_1408),
.A2(n_1276),
.B1(n_1277),
.B2(n_1260),
.Y(n_1681)
);

OAI22xp5_ASAP7_75t_L g1682 ( 
.A1(n_1576),
.A2(n_1343),
.B1(n_1264),
.B2(n_1322),
.Y(n_1682)
);

NAND2xp5_ASAP7_75t_L g1683 ( 
.A(n_1480),
.B(n_1263),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1480),
.B(n_1270),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_L g1685 ( 
.A(n_1477),
.B(n_1297),
.Y(n_1685)
);

O2A1O1Ixp33_ASAP7_75t_L g1686 ( 
.A1(n_1561),
.A2(n_1310),
.B(n_1314),
.C(n_1297),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_SL g1687 ( 
.A(n_1468),
.B(n_1227),
.Y(n_1687)
);

INVxp67_ASAP7_75t_L g1688 ( 
.A(n_1402),
.Y(n_1688)
);

O2A1O1Ixp33_ASAP7_75t_L g1689 ( 
.A1(n_1531),
.A2(n_1314),
.B(n_1326),
.C(n_1310),
.Y(n_1689)
);

AOI21xp5_ASAP7_75t_L g1690 ( 
.A1(n_1563),
.A2(n_1283),
.B(n_1279),
.Y(n_1690)
);

INVx2_ASAP7_75t_L g1691 ( 
.A(n_1427),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_L g1692 ( 
.A(n_1477),
.B(n_1326),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_L g1693 ( 
.A(n_1637),
.B(n_1329),
.Y(n_1693)
);

AOI21xp5_ASAP7_75t_L g1694 ( 
.A1(n_1653),
.A2(n_1389),
.B(n_1364),
.Y(n_1694)
);

INVx2_ASAP7_75t_L g1695 ( 
.A(n_1428),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1437),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_L g1697 ( 
.A(n_1439),
.B(n_1329),
.Y(n_1697)
);

NOR2x1p5_ASAP7_75t_SL g1698 ( 
.A(n_1594),
.B(n_1204),
.Y(n_1698)
);

INVx2_ASAP7_75t_SL g1699 ( 
.A(n_1457),
.Y(n_1699)
);

HB1xp67_ASAP7_75t_L g1700 ( 
.A(n_1466),
.Y(n_1700)
);

NOR2xp33_ASAP7_75t_L g1701 ( 
.A(n_1483),
.B(n_1331),
.Y(n_1701)
);

AOI21xp5_ASAP7_75t_L g1702 ( 
.A1(n_1655),
.A2(n_1389),
.B(n_1364),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_L g1703 ( 
.A(n_1439),
.B(n_1331),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1463),
.Y(n_1704)
);

INVx2_ASAP7_75t_L g1705 ( 
.A(n_1534),
.Y(n_1705)
);

AOI21xp5_ASAP7_75t_L g1706 ( 
.A1(n_1655),
.A2(n_1207),
.B(n_1204),
.Y(n_1706)
);

AOI21xp5_ASAP7_75t_L g1707 ( 
.A1(n_1658),
.A2(n_1213),
.B(n_1207),
.Y(n_1707)
);

OAI21xp5_ASAP7_75t_L g1708 ( 
.A1(n_1626),
.A2(n_1355),
.B(n_1336),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_L g1709 ( 
.A(n_1657),
.B(n_1355),
.Y(n_1709)
);

AOI21x1_ASAP7_75t_L g1710 ( 
.A1(n_1633),
.A2(n_1191),
.B(n_1186),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1447),
.Y(n_1711)
);

NAND2xp5_ASAP7_75t_L g1712 ( 
.A(n_1412),
.B(n_1336),
.Y(n_1712)
);

O2A1O1Ixp33_ASAP7_75t_L g1713 ( 
.A1(n_1413),
.A2(n_1191),
.B(n_1229),
.C(n_1186),
.Y(n_1713)
);

NOR2xp33_ASAP7_75t_L g1714 ( 
.A(n_1544),
.B(n_1152),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_1412),
.B(n_1185),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_SL g1716 ( 
.A(n_1497),
.B(n_1264),
.Y(n_1716)
);

AOI21xp5_ASAP7_75t_L g1717 ( 
.A1(n_1658),
.A2(n_1222),
.B(n_1213),
.Y(n_1717)
);

AND2x2_ASAP7_75t_L g1718 ( 
.A(n_1432),
.B(n_1322),
.Y(n_1718)
);

OAI21xp33_ASAP7_75t_L g1719 ( 
.A1(n_1542),
.A2(n_1557),
.B(n_1435),
.Y(n_1719)
);

AOI21xp5_ASAP7_75t_L g1720 ( 
.A1(n_1659),
.A2(n_1633),
.B(n_1551),
.Y(n_1720)
);

AOI21xp5_ASAP7_75t_L g1721 ( 
.A1(n_1659),
.A2(n_1252),
.B(n_1222),
.Y(n_1721)
);

AOI22xp5_ASAP7_75t_L g1722 ( 
.A1(n_1496),
.A2(n_1229),
.B1(n_1189),
.B2(n_1185),
.Y(n_1722)
);

AOI21xp5_ASAP7_75t_L g1723 ( 
.A1(n_1551),
.A2(n_1285),
.B(n_1252),
.Y(n_1723)
);

NAND2xp5_ASAP7_75t_L g1724 ( 
.A(n_1643),
.B(n_1189),
.Y(n_1724)
);

AO21x1_ASAP7_75t_L g1725 ( 
.A1(n_1423),
.A2(n_1170),
.B(n_1163),
.Y(n_1725)
);

AOI21x1_ASAP7_75t_L g1726 ( 
.A1(n_1603),
.A2(n_1181),
.B(n_1179),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1448),
.Y(n_1727)
);

AOI22xp33_ASAP7_75t_L g1728 ( 
.A1(n_1519),
.A2(n_1234),
.B1(n_1238),
.B2(n_1231),
.Y(n_1728)
);

OAI22xp5_ASAP7_75t_L g1729 ( 
.A1(n_1413),
.A2(n_1187),
.B1(n_1211),
.B2(n_1177),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_SL g1730 ( 
.A(n_1497),
.B(n_747),
.Y(n_1730)
);

AOI21xp5_ASAP7_75t_L g1731 ( 
.A1(n_1409),
.A2(n_1254),
.B(n_1241),
.Y(n_1731)
);

NAND2xp5_ASAP7_75t_SL g1732 ( 
.A(n_1473),
.B(n_755),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_L g1733 ( 
.A(n_1450),
.B(n_1262),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1453),
.Y(n_1734)
);

O2A1O1Ixp33_ASAP7_75t_SL g1735 ( 
.A1(n_1486),
.A2(n_1261),
.B(n_1250),
.C(n_1187),
.Y(n_1735)
);

NAND2xp5_ASAP7_75t_L g1736 ( 
.A(n_1451),
.B(n_1177),
.Y(n_1736)
);

BUFx2_ASAP7_75t_L g1737 ( 
.A(n_1520),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1454),
.Y(n_1738)
);

INVx2_ASAP7_75t_L g1739 ( 
.A(n_1549),
.Y(n_1739)
);

BUFx2_ASAP7_75t_L g1740 ( 
.A(n_1570),
.Y(n_1740)
);

AOI21xp5_ASAP7_75t_L g1741 ( 
.A1(n_1431),
.A2(n_1436),
.B(n_1433),
.Y(n_1741)
);

AOI22xp33_ASAP7_75t_L g1742 ( 
.A1(n_1530),
.A2(n_1261),
.B1(n_1224),
.B2(n_1230),
.Y(n_1742)
);

NAND2xp5_ASAP7_75t_L g1743 ( 
.A(n_1456),
.B(n_1211),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_L g1744 ( 
.A(n_1455),
.B(n_1224),
.Y(n_1744)
);

OAI21xp5_ASAP7_75t_L g1745 ( 
.A1(n_1461),
.A2(n_764),
.B(n_757),
.Y(n_1745)
);

BUFx2_ASAP7_75t_L g1746 ( 
.A(n_1541),
.Y(n_1746)
);

NOR2xp33_ASAP7_75t_L g1747 ( 
.A(n_1484),
.B(n_781),
.Y(n_1747)
);

NAND2xp5_ASAP7_75t_L g1748 ( 
.A(n_1583),
.B(n_768),
.Y(n_1748)
);

NOR2xp33_ASAP7_75t_L g1749 ( 
.A(n_1484),
.B(n_779),
.Y(n_1749)
);

BUFx6f_ASAP7_75t_L g1750 ( 
.A(n_1631),
.Y(n_1750)
);

OAI22xp5_ASAP7_75t_L g1751 ( 
.A1(n_1398),
.A2(n_539),
.B1(n_593),
.B2(n_510),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1600),
.Y(n_1752)
);

NOR2xp33_ASAP7_75t_L g1753 ( 
.A(n_1509),
.B(n_769),
.Y(n_1753)
);

O2A1O1Ixp33_ASAP7_75t_L g1754 ( 
.A1(n_1574),
.A2(n_18),
.B(n_16),
.C(n_17),
.Y(n_1754)
);

NAND2xp5_ASAP7_75t_L g1755 ( 
.A(n_1583),
.B(n_772),
.Y(n_1755)
);

OAI321xp33_ASAP7_75t_L g1756 ( 
.A1(n_1580),
.A2(n_724),
.A3(n_704),
.B1(n_593),
.B2(n_539),
.C(n_510),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1601),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_L g1758 ( 
.A(n_1550),
.B(n_18),
.Y(n_1758)
);

AOI21xp5_ASAP7_75t_L g1759 ( 
.A1(n_1461),
.A2(n_724),
.B(n_704),
.Y(n_1759)
);

NAND2xp5_ASAP7_75t_L g1760 ( 
.A(n_1508),
.B(n_19),
.Y(n_1760)
);

NAND2xp5_ASAP7_75t_L g1761 ( 
.A(n_1438),
.B(n_20),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1502),
.Y(n_1762)
);

AO21x1_ASAP7_75t_L g1763 ( 
.A1(n_1564),
.A2(n_704),
.B(n_593),
.Y(n_1763)
);

NOR2xp33_ASAP7_75t_L g1764 ( 
.A(n_1399),
.B(n_21),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1506),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_L g1766 ( 
.A(n_1438),
.B(n_21),
.Y(n_1766)
);

INVx5_ASAP7_75t_L g1767 ( 
.A(n_1613),
.Y(n_1767)
);

AOI21xp5_ASAP7_75t_L g1768 ( 
.A1(n_1462),
.A2(n_724),
.B(n_261),
.Y(n_1768)
);

HB1xp67_ASAP7_75t_L g1769 ( 
.A(n_1410),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_L g1770 ( 
.A(n_1533),
.B(n_22),
.Y(n_1770)
);

AOI21x1_ASAP7_75t_L g1771 ( 
.A1(n_1624),
.A2(n_724),
.B(n_262),
.Y(n_1771)
);

HB1xp67_ASAP7_75t_L g1772 ( 
.A(n_1410),
.Y(n_1772)
);

A2O1A1Ixp33_ASAP7_75t_L g1773 ( 
.A1(n_1444),
.A2(n_25),
.B(n_23),
.C(n_24),
.Y(n_1773)
);

BUFx4f_ASAP7_75t_L g1774 ( 
.A(n_1613),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1517),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_L g1776 ( 
.A(n_1634),
.B(n_26),
.Y(n_1776)
);

NAND2xp5_ASAP7_75t_L g1777 ( 
.A(n_1465),
.B(n_1467),
.Y(n_1777)
);

OAI21xp5_ASAP7_75t_L g1778 ( 
.A1(n_1465),
.A2(n_28),
.B(n_29),
.Y(n_1778)
);

NOR2xp33_ASAP7_75t_L g1779 ( 
.A(n_1535),
.B(n_29),
.Y(n_1779)
);

INVx2_ASAP7_75t_L g1780 ( 
.A(n_1566),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1524),
.Y(n_1781)
);

NAND2xp5_ASAP7_75t_L g1782 ( 
.A(n_1467),
.B(n_30),
.Y(n_1782)
);

OR2x2_ASAP7_75t_L g1783 ( 
.A(n_1590),
.B(n_30),
.Y(n_1783)
);

BUFx4f_ASAP7_75t_L g1784 ( 
.A(n_1613),
.Y(n_1784)
);

OAI21xp5_ASAP7_75t_L g1785 ( 
.A1(n_1470),
.A2(n_31),
.B(n_32),
.Y(n_1785)
);

AOI21xp5_ASAP7_75t_L g1786 ( 
.A1(n_1640),
.A2(n_271),
.B(n_269),
.Y(n_1786)
);

CKINVDCx5p33_ASAP7_75t_R g1787 ( 
.A(n_1569),
.Y(n_1787)
);

AOI22xp5_ASAP7_75t_L g1788 ( 
.A1(n_1578),
.A2(n_33),
.B1(n_31),
.B2(n_32),
.Y(n_1788)
);

A2O1A1Ixp33_ASAP7_75t_L g1789 ( 
.A1(n_1615),
.A2(n_35),
.B(n_33),
.C(n_34),
.Y(n_1789)
);

NAND2xp5_ASAP7_75t_L g1790 ( 
.A(n_1470),
.B(n_34),
.Y(n_1790)
);

BUFx6f_ASAP7_75t_L g1791 ( 
.A(n_1631),
.Y(n_1791)
);

AOI22xp5_ASAP7_75t_L g1792 ( 
.A1(n_1460),
.A2(n_40),
.B1(n_35),
.B2(n_38),
.Y(n_1792)
);

NOR2xp33_ASAP7_75t_L g1793 ( 
.A(n_1598),
.B(n_38),
.Y(n_1793)
);

AOI22xp5_ASAP7_75t_L g1794 ( 
.A1(n_1469),
.A2(n_43),
.B1(n_40),
.B2(n_41),
.Y(n_1794)
);

AOI21xp5_ASAP7_75t_L g1795 ( 
.A1(n_1641),
.A2(n_281),
.B(n_280),
.Y(n_1795)
);

BUFx2_ASAP7_75t_L g1796 ( 
.A(n_1441),
.Y(n_1796)
);

NOR2xp33_ASAP7_75t_L g1797 ( 
.A(n_1471),
.B(n_41),
.Y(n_1797)
);

NAND2xp5_ASAP7_75t_L g1798 ( 
.A(n_1475),
.B(n_43),
.Y(n_1798)
);

OAI21xp5_ASAP7_75t_L g1799 ( 
.A1(n_1475),
.A2(n_44),
.B(n_45),
.Y(n_1799)
);

AOI21xp5_ASAP7_75t_L g1800 ( 
.A1(n_1641),
.A2(n_287),
.B(n_282),
.Y(n_1800)
);

BUFx2_ASAP7_75t_L g1801 ( 
.A(n_1619),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1532),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1537),
.Y(n_1803)
);

NAND2xp5_ASAP7_75t_L g1804 ( 
.A(n_1430),
.B(n_1579),
.Y(n_1804)
);

AND2x2_ASAP7_75t_L g1805 ( 
.A(n_1582),
.B(n_44),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1540),
.Y(n_1806)
);

O2A1O1Ixp33_ASAP7_75t_L g1807 ( 
.A1(n_1545),
.A2(n_47),
.B(n_45),
.C(n_46),
.Y(n_1807)
);

INVxp67_ASAP7_75t_L g1808 ( 
.A(n_1584),
.Y(n_1808)
);

NAND2xp5_ASAP7_75t_L g1809 ( 
.A(n_1430),
.B(n_46),
.Y(n_1809)
);

AOI22xp5_ASAP7_75t_L g1810 ( 
.A1(n_1584),
.A2(n_49),
.B1(n_47),
.B2(n_48),
.Y(n_1810)
);

BUFx6f_ASAP7_75t_L g1811 ( 
.A(n_1539),
.Y(n_1811)
);

OR2x6_ASAP7_75t_L g1812 ( 
.A(n_1586),
.B(n_48),
.Y(n_1812)
);

NOR2xp33_ASAP7_75t_L g1813 ( 
.A(n_1472),
.B(n_49),
.Y(n_1813)
);

INVx2_ASAP7_75t_L g1814 ( 
.A(n_1567),
.Y(n_1814)
);

AOI22xp5_ASAP7_75t_L g1815 ( 
.A1(n_1500),
.A2(n_54),
.B1(n_51),
.B2(n_53),
.Y(n_1815)
);

INVx4_ASAP7_75t_L g1816 ( 
.A(n_1434),
.Y(n_1816)
);

OR2x2_ASAP7_75t_L g1817 ( 
.A(n_1620),
.B(n_51),
.Y(n_1817)
);

OAI22xp5_ASAP7_75t_L g1818 ( 
.A1(n_1621),
.A2(n_1586),
.B1(n_1553),
.B2(n_1555),
.Y(n_1818)
);

OAI21xp5_ASAP7_75t_L g1819 ( 
.A1(n_1595),
.A2(n_53),
.B(n_55),
.Y(n_1819)
);

INVx2_ASAP7_75t_L g1820 ( 
.A(n_1638),
.Y(n_1820)
);

NAND2x1_ASAP7_75t_L g1821 ( 
.A(n_1652),
.B(n_288),
.Y(n_1821)
);

INVx4_ASAP7_75t_L g1822 ( 
.A(n_1589),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1547),
.Y(n_1823)
);

NAND2xp5_ASAP7_75t_L g1824 ( 
.A(n_1650),
.B(n_55),
.Y(n_1824)
);

OR2x2_ASAP7_75t_L g1825 ( 
.A(n_1568),
.B(n_56),
.Y(n_1825)
);

OAI21xp5_ASAP7_75t_L g1826 ( 
.A1(n_1476),
.A2(n_56),
.B(n_57),
.Y(n_1826)
);

NAND2xp5_ASAP7_75t_L g1827 ( 
.A(n_1482),
.B(n_57),
.Y(n_1827)
);

A2O1A1Ixp33_ASAP7_75t_L g1828 ( 
.A1(n_1591),
.A2(n_61),
.B(n_59),
.C(n_60),
.Y(n_1828)
);

NOR2xp33_ASAP7_75t_L g1829 ( 
.A(n_1503),
.B(n_59),
.Y(n_1829)
);

AND2x6_ASAP7_75t_L g1830 ( 
.A(n_1479),
.B(n_1525),
.Y(n_1830)
);

NAND2xp33_ASAP7_75t_L g1831 ( 
.A(n_1459),
.B(n_289),
.Y(n_1831)
);

NAND2xp5_ASAP7_75t_L g1832 ( 
.A(n_1581),
.B(n_62),
.Y(n_1832)
);

NOR2x2_ASAP7_75t_L g1833 ( 
.A(n_1546),
.B(n_62),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1560),
.Y(n_1834)
);

INVx2_ASAP7_75t_SL g1835 ( 
.A(n_1629),
.Y(n_1835)
);

AND2x2_ASAP7_75t_L g1836 ( 
.A(n_1611),
.B(n_64),
.Y(n_1836)
);

O2A1O1Ixp33_ASAP7_75t_L g1837 ( 
.A1(n_1572),
.A2(n_67),
.B(n_65),
.C(n_66),
.Y(n_1837)
);

OAI21xp5_ASAP7_75t_L g1838 ( 
.A1(n_1562),
.A2(n_65),
.B(n_68),
.Y(n_1838)
);

NOR2xp33_ASAP7_75t_L g1839 ( 
.A(n_1543),
.B(n_69),
.Y(n_1839)
);

NAND2xp5_ASAP7_75t_L g1840 ( 
.A(n_1575),
.B(n_70),
.Y(n_1840)
);

OAI21xp5_ASAP7_75t_L g1841 ( 
.A1(n_1571),
.A2(n_71),
.B(n_72),
.Y(n_1841)
);

HB1xp67_ASAP7_75t_L g1842 ( 
.A(n_1415),
.Y(n_1842)
);

NAND2xp5_ASAP7_75t_L g1843 ( 
.A(n_1651),
.B(n_73),
.Y(n_1843)
);

CKINVDCx5p33_ASAP7_75t_R g1844 ( 
.A(n_1654),
.Y(n_1844)
);

NOR2xp33_ASAP7_75t_L g1845 ( 
.A(n_1592),
.B(n_74),
.Y(n_1845)
);

AOI21xp5_ASAP7_75t_L g1846 ( 
.A1(n_1492),
.A2(n_298),
.B(n_297),
.Y(n_1846)
);

AOI21xp5_ASAP7_75t_L g1847 ( 
.A1(n_1421),
.A2(n_1609),
.B(n_1514),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_1656),
.Y(n_1848)
);

AOI21xp5_ASAP7_75t_L g1849 ( 
.A1(n_1514),
.A2(n_310),
.B(n_309),
.Y(n_1849)
);

INVx2_ASAP7_75t_L g1850 ( 
.A(n_1660),
.Y(n_1850)
);

BUFx2_ASAP7_75t_L g1851 ( 
.A(n_1596),
.Y(n_1851)
);

INVx3_ASAP7_75t_L g1852 ( 
.A(n_1479),
.Y(n_1852)
);

OAI21xp5_ASAP7_75t_L g1853 ( 
.A1(n_1605),
.A2(n_77),
.B(n_78),
.Y(n_1853)
);

INVx2_ASAP7_75t_L g1854 ( 
.A(n_1617),
.Y(n_1854)
);

BUFx3_ASAP7_75t_L g1855 ( 
.A(n_1593),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1618),
.Y(n_1856)
);

AOI21xp5_ASAP7_75t_L g1857 ( 
.A1(n_1525),
.A2(n_314),
.B(n_311),
.Y(n_1857)
);

NOR2x1_ASAP7_75t_L g1858 ( 
.A(n_1630),
.B(n_79),
.Y(n_1858)
);

AOI21xp5_ASAP7_75t_L g1859 ( 
.A1(n_1429),
.A2(n_1625),
.B(n_1623),
.Y(n_1859)
);

OAI21xp33_ASAP7_75t_L g1860 ( 
.A1(n_1644),
.A2(n_80),
.B(n_81),
.Y(n_1860)
);

NAND2xp5_ASAP7_75t_SL g1861 ( 
.A(n_1602),
.B(n_1499),
.Y(n_1861)
);

INVx1_ASAP7_75t_L g1862 ( 
.A(n_1632),
.Y(n_1862)
);

A2O1A1Ixp33_ASAP7_75t_L g1863 ( 
.A1(n_1647),
.A2(n_82),
.B(n_80),
.C(n_81),
.Y(n_1863)
);

INVxp67_ASAP7_75t_L g1864 ( 
.A(n_1627),
.Y(n_1864)
);

BUFx6f_ASAP7_75t_L g1865 ( 
.A(n_1539),
.Y(n_1865)
);

O2A1O1Ixp5_ASAP7_75t_L g1866 ( 
.A1(n_1446),
.A2(n_323),
.B(n_324),
.C(n_315),
.Y(n_1866)
);

BUFx4f_ASAP7_75t_L g1867 ( 
.A(n_1445),
.Y(n_1867)
);

NOR3xp33_ASAP7_75t_L g1868 ( 
.A(n_1645),
.B(n_83),
.C(n_85),
.Y(n_1868)
);

AOI21xp5_ASAP7_75t_L g1869 ( 
.A1(n_1538),
.A2(n_331),
.B(n_327),
.Y(n_1869)
);

OAI21xp5_ASAP7_75t_L g1870 ( 
.A1(n_1585),
.A2(n_1587),
.B(n_1488),
.Y(n_1870)
);

NAND2xp5_ASAP7_75t_L g1871 ( 
.A(n_1635),
.B(n_83),
.Y(n_1871)
);

AOI21xp5_ASAP7_75t_L g1872 ( 
.A1(n_1606),
.A2(n_336),
.B(n_334),
.Y(n_1872)
);

INVx4_ASAP7_75t_L g1873 ( 
.A(n_1589),
.Y(n_1873)
);

INVx2_ASAP7_75t_L g1874 ( 
.A(n_1617),
.Y(n_1874)
);

AOI21xp5_ASAP7_75t_L g1875 ( 
.A1(n_1608),
.A2(n_340),
.B(n_339),
.Y(n_1875)
);

INVx3_ASAP7_75t_L g1876 ( 
.A(n_1479),
.Y(n_1876)
);

NAND2xp5_ASAP7_75t_L g1877 ( 
.A(n_1536),
.B(n_85),
.Y(n_1877)
);

AOI21xp5_ASAP7_75t_L g1878 ( 
.A1(n_1614),
.A2(n_342),
.B(n_341),
.Y(n_1878)
);

AOI21xp5_ASAP7_75t_L g1879 ( 
.A1(n_1487),
.A2(n_1491),
.B(n_1490),
.Y(n_1879)
);

INVx3_ASAP7_75t_L g1880 ( 
.A(n_1511),
.Y(n_1880)
);

AND2x4_ASAP7_75t_L g1881 ( 
.A(n_1481),
.B(n_86),
.Y(n_1881)
);

NAND2xp5_ASAP7_75t_L g1882 ( 
.A(n_1552),
.B(n_86),
.Y(n_1882)
);

NAND2xp5_ASAP7_75t_SL g1883 ( 
.A(n_1516),
.B(n_87),
.Y(n_1883)
);

INVx4_ASAP7_75t_L g1884 ( 
.A(n_1511),
.Y(n_1884)
);

INVx2_ASAP7_75t_L g1885 ( 
.A(n_1440),
.Y(n_1885)
);

AOI21xp5_ASAP7_75t_L g1886 ( 
.A1(n_1622),
.A2(n_344),
.B(n_343),
.Y(n_1886)
);

NAND2xp5_ASAP7_75t_SL g1887 ( 
.A(n_1516),
.B(n_90),
.Y(n_1887)
);

INVx3_ASAP7_75t_L g1888 ( 
.A(n_1511),
.Y(n_1888)
);

CKINVDCx5p33_ASAP7_75t_R g1889 ( 
.A(n_1558),
.Y(n_1889)
);

A2O1A1Ixp33_ASAP7_75t_L g1890 ( 
.A1(n_1636),
.A2(n_93),
.B(n_91),
.C(n_92),
.Y(n_1890)
);

INVx2_ASAP7_75t_L g1891 ( 
.A(n_1442),
.Y(n_1891)
);

A2O1A1Ixp33_ASAP7_75t_L g1892 ( 
.A1(n_1639),
.A2(n_95),
.B(n_93),
.C(n_94),
.Y(n_1892)
);

NAND2xp5_ASAP7_75t_L g1893 ( 
.A(n_1445),
.B(n_94),
.Y(n_1893)
);

AOI33xp33_ASAP7_75t_L g1894 ( 
.A1(n_1648),
.A2(n_97),
.A3(n_99),
.B1(n_100),
.B2(n_101),
.B3(n_103),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1449),
.Y(n_1895)
);

INVx4_ASAP7_75t_L g1896 ( 
.A(n_1646),
.Y(n_1896)
);

O2A1O1Ixp33_ASAP7_75t_L g1897 ( 
.A1(n_1518),
.A2(n_104),
.B(n_97),
.C(n_101),
.Y(n_1897)
);

NAND2xp5_ASAP7_75t_SL g1898 ( 
.A(n_1518),
.B(n_106),
.Y(n_1898)
);

AND2x2_ASAP7_75t_L g1899 ( 
.A(n_1521),
.B(n_107),
.Y(n_1899)
);

AOI21xp5_ASAP7_75t_L g1900 ( 
.A1(n_1628),
.A2(n_347),
.B(n_346),
.Y(n_1900)
);

BUFx4f_ASAP7_75t_L g1901 ( 
.A(n_1573),
.Y(n_1901)
);

NOR2xp33_ASAP7_75t_L g1902 ( 
.A(n_1610),
.B(n_107),
.Y(n_1902)
);

NAND2xp5_ASAP7_75t_L g1903 ( 
.A(n_1612),
.B(n_108),
.Y(n_1903)
);

AOI21xp5_ASAP7_75t_L g1904 ( 
.A1(n_1464),
.A2(n_350),
.B(n_349),
.Y(n_1904)
);

BUFx4f_ASAP7_75t_L g1905 ( 
.A(n_1573),
.Y(n_1905)
);

NAND2xp5_ASAP7_75t_L g1906 ( 
.A(n_1522),
.B(n_108),
.Y(n_1906)
);

AOI21xp5_ASAP7_75t_L g1907 ( 
.A1(n_1642),
.A2(n_1649),
.B(n_1474),
.Y(n_1907)
);

INVx3_ASAP7_75t_L g1908 ( 
.A(n_1493),
.Y(n_1908)
);

AOI21xp5_ASAP7_75t_L g1909 ( 
.A1(n_1452),
.A2(n_355),
.B(n_352),
.Y(n_1909)
);

NAND2xp5_ASAP7_75t_SL g1910 ( 
.A(n_1528),
.B(n_109),
.Y(n_1910)
);

NAND2xp5_ASAP7_75t_L g1911 ( 
.A(n_1528),
.B(n_111),
.Y(n_1911)
);

OAI21xp5_ASAP7_75t_L g1912 ( 
.A1(n_1510),
.A2(n_112),
.B(n_113),
.Y(n_1912)
);

AOI21xp5_ASAP7_75t_L g1913 ( 
.A1(n_1495),
.A2(n_358),
.B(n_357),
.Y(n_1913)
);

OAI21xp5_ASAP7_75t_L g1914 ( 
.A1(n_1548),
.A2(n_112),
.B(n_113),
.Y(n_1914)
);

AOI21xp5_ASAP7_75t_L g1915 ( 
.A1(n_1548),
.A2(n_364),
.B(n_363),
.Y(n_1915)
);

NAND2xp5_ASAP7_75t_L g1916 ( 
.A(n_1554),
.B(n_114),
.Y(n_1916)
);

NOR2xp33_ASAP7_75t_SL g1917 ( 
.A(n_1539),
.B(n_365),
.Y(n_1917)
);

O2A1O1Ixp5_ASAP7_75t_L g1918 ( 
.A1(n_1422),
.A2(n_478),
.B(n_475),
.C(n_473),
.Y(n_1918)
);

AND2x2_ASAP7_75t_L g1919 ( 
.A(n_1554),
.B(n_115),
.Y(n_1919)
);

OAI21xp5_ASAP7_75t_L g1920 ( 
.A1(n_1400),
.A2(n_115),
.B(n_116),
.Y(n_1920)
);

NOR2xp33_ASAP7_75t_L g1921 ( 
.A(n_1526),
.B(n_117),
.Y(n_1921)
);

AOI21xp5_ASAP7_75t_L g1922 ( 
.A1(n_1507),
.A2(n_370),
.B(n_369),
.Y(n_1922)
);

INVx2_ASAP7_75t_SL g1923 ( 
.A(n_1588),
.Y(n_1923)
);

NAND2xp5_ASAP7_75t_L g1924 ( 
.A(n_1597),
.B(n_117),
.Y(n_1924)
);

NAND2xp33_ASAP7_75t_L g1925 ( 
.A(n_1459),
.B(n_1556),
.Y(n_1925)
);

NAND2xp5_ASAP7_75t_L g1926 ( 
.A(n_1407),
.B(n_118),
.Y(n_1926)
);

INVx2_ASAP7_75t_L g1927 ( 
.A(n_1498),
.Y(n_1927)
);

HB1xp67_ASAP7_75t_L g1928 ( 
.A(n_1411),
.Y(n_1928)
);

NOR2xp33_ASAP7_75t_L g1929 ( 
.A(n_1493),
.B(n_118),
.Y(n_1929)
);

INVx2_ASAP7_75t_L g1930 ( 
.A(n_1662),
.Y(n_1930)
);

BUFx4_ASAP7_75t_SL g1931 ( 
.A(n_1787),
.Y(n_1931)
);

BUFx2_ASAP7_75t_L g1932 ( 
.A(n_1812),
.Y(n_1932)
);

INVx2_ASAP7_75t_L g1933 ( 
.A(n_1671),
.Y(n_1933)
);

AND2x2_ASAP7_75t_L g1934 ( 
.A(n_1688),
.B(n_1559),
.Y(n_1934)
);

NOR2xp67_ASAP7_75t_L g1935 ( 
.A(n_1767),
.B(n_1652),
.Y(n_1935)
);

NAND2xp5_ASAP7_75t_L g1936 ( 
.A(n_1719),
.B(n_1559),
.Y(n_1936)
);

A2O1A1Ixp33_ASAP7_75t_L g1937 ( 
.A1(n_1664),
.A2(n_1416),
.B(n_1420),
.C(n_1425),
.Y(n_1937)
);

AOI21xp5_ASAP7_75t_L g1938 ( 
.A1(n_1735),
.A2(n_1565),
.B(n_1556),
.Y(n_1938)
);

AO32x1_ASAP7_75t_L g1939 ( 
.A1(n_1751),
.A2(n_1529),
.A3(n_1504),
.B1(n_1505),
.B2(n_1512),
.Y(n_1939)
);

NAND2xp5_ASAP7_75t_L g1940 ( 
.A(n_1864),
.B(n_1607),
.Y(n_1940)
);

A2O1A1Ixp33_ASAP7_75t_L g1941 ( 
.A1(n_1678),
.A2(n_1616),
.B(n_1527),
.C(n_1501),
.Y(n_1941)
);

O2A1O1Ixp33_ASAP7_75t_L g1942 ( 
.A1(n_1670),
.A2(n_1523),
.B(n_1515),
.C(n_1458),
.Y(n_1942)
);

INVx1_ASAP7_75t_L g1943 ( 
.A(n_1691),
.Y(n_1943)
);

INVx4_ASAP7_75t_L g1944 ( 
.A(n_1677),
.Y(n_1944)
);

NAND2xp5_ASAP7_75t_SL g1945 ( 
.A(n_1677),
.B(n_1599),
.Y(n_1945)
);

NOR2xp33_ASAP7_75t_L g1946 ( 
.A(n_1740),
.B(n_1594),
.Y(n_1946)
);

NAND2xp5_ASAP7_75t_L g1947 ( 
.A(n_1673),
.B(n_1594),
.Y(n_1947)
);

NAND2xp5_ASAP7_75t_L g1948 ( 
.A(n_1669),
.B(n_1594),
.Y(n_1948)
);

BUFx2_ASAP7_75t_L g1949 ( 
.A(n_1812),
.Y(n_1949)
);

NAND2xp5_ASAP7_75t_L g1950 ( 
.A(n_1675),
.B(n_1679),
.Y(n_1950)
);

INVx1_ASAP7_75t_L g1951 ( 
.A(n_1695),
.Y(n_1951)
);

NAND2xp5_ASAP7_75t_L g1952 ( 
.A(n_1696),
.B(n_1594),
.Y(n_1952)
);

HB1xp67_ASAP7_75t_L g1953 ( 
.A(n_1737),
.Y(n_1953)
);

NAND2xp5_ASAP7_75t_SL g1954 ( 
.A(n_1677),
.B(n_1599),
.Y(n_1954)
);

INVx1_ASAP7_75t_L g1955 ( 
.A(n_1704),
.Y(n_1955)
);

NAND2xp5_ASAP7_75t_L g1956 ( 
.A(n_1711),
.B(n_1594),
.Y(n_1956)
);

NAND2xp5_ASAP7_75t_L g1957 ( 
.A(n_1727),
.B(n_1734),
.Y(n_1957)
);

AND2x2_ASAP7_75t_L g1958 ( 
.A(n_1746),
.B(n_119),
.Y(n_1958)
);

NAND2xp5_ASAP7_75t_L g1959 ( 
.A(n_1738),
.B(n_1714),
.Y(n_1959)
);

INVx3_ASAP7_75t_L g1960 ( 
.A(n_1750),
.Y(n_1960)
);

O2A1O1Ixp33_ASAP7_75t_L g1961 ( 
.A1(n_1789),
.A2(n_1459),
.B(n_120),
.C(n_121),
.Y(n_1961)
);

INVx2_ASAP7_75t_L g1962 ( 
.A(n_1762),
.Y(n_1962)
);

A2O1A1Ixp33_ASAP7_75t_L g1963 ( 
.A1(n_1902),
.A2(n_1646),
.B(n_1459),
.C(n_125),
.Y(n_1963)
);

AOI22xp5_ASAP7_75t_L g1964 ( 
.A1(n_1805),
.A2(n_1459),
.B1(n_124),
.B2(n_125),
.Y(n_1964)
);

NOR2xp33_ASAP7_75t_L g1965 ( 
.A(n_1665),
.B(n_1459),
.Y(n_1965)
);

NOR2xp33_ASAP7_75t_SL g1966 ( 
.A(n_1816),
.B(n_119),
.Y(n_1966)
);

INVx1_ASAP7_75t_L g1967 ( 
.A(n_1752),
.Y(n_1967)
);

AND2x2_ASAP7_75t_L g1968 ( 
.A(n_1700),
.B(n_126),
.Y(n_1968)
);

AOI22xp5_ASAP7_75t_L g1969 ( 
.A1(n_1718),
.A2(n_128),
.B1(n_129),
.B2(n_130),
.Y(n_1969)
);

NAND2xp5_ASAP7_75t_L g1970 ( 
.A(n_1765),
.B(n_128),
.Y(n_1970)
);

OAI22xp5_ASAP7_75t_L g1971 ( 
.A1(n_1812),
.A2(n_129),
.B1(n_130),
.B2(n_131),
.Y(n_1971)
);

AOI21xp5_ASAP7_75t_L g1972 ( 
.A1(n_1720),
.A2(n_384),
.B(n_379),
.Y(n_1972)
);

INVx2_ASAP7_75t_L g1973 ( 
.A(n_1775),
.Y(n_1973)
);

INVx1_ASAP7_75t_L g1974 ( 
.A(n_1757),
.Y(n_1974)
);

NAND2xp5_ASAP7_75t_L g1975 ( 
.A(n_1781),
.B(n_132),
.Y(n_1975)
);

INVx2_ASAP7_75t_L g1976 ( 
.A(n_1802),
.Y(n_1976)
);

HB1xp67_ASAP7_75t_L g1977 ( 
.A(n_1699),
.Y(n_1977)
);

AOI221xp5_ASAP7_75t_L g1978 ( 
.A1(n_1839),
.A2(n_133),
.B1(n_134),
.B2(n_135),
.C(n_136),
.Y(n_1978)
);

INVxp33_ASAP7_75t_L g1979 ( 
.A(n_1796),
.Y(n_1979)
);

NAND2xp33_ASAP7_75t_SL g1980 ( 
.A(n_1750),
.B(n_133),
.Y(n_1980)
);

O2A1O1Ixp33_ASAP7_75t_L g1981 ( 
.A1(n_1807),
.A2(n_135),
.B(n_136),
.C(n_137),
.Y(n_1981)
);

O2A1O1Ixp33_ASAP7_75t_L g1982 ( 
.A1(n_1793),
.A2(n_138),
.B(n_139),
.C(n_140),
.Y(n_1982)
);

CKINVDCx14_ASAP7_75t_R g1983 ( 
.A(n_1816),
.Y(n_1983)
);

NAND3xp33_ASAP7_75t_SL g1984 ( 
.A(n_1844),
.B(n_139),
.C(n_140),
.Y(n_1984)
);

A2O1A1Ixp33_ASAP7_75t_SL g1985 ( 
.A1(n_1756),
.A2(n_142),
.B(n_145),
.C(n_146),
.Y(n_1985)
);

BUFx2_ASAP7_75t_L g1986 ( 
.A(n_1750),
.Y(n_1986)
);

O2A1O1Ixp33_ASAP7_75t_L g1987 ( 
.A1(n_1760),
.A2(n_145),
.B(n_146),
.C(n_148),
.Y(n_1987)
);

NAND2xp5_ASAP7_75t_L g1988 ( 
.A(n_1803),
.B(n_149),
.Y(n_1988)
);

NOR2xp33_ASAP7_75t_L g1989 ( 
.A(n_1817),
.B(n_149),
.Y(n_1989)
);

BUFx6f_ASAP7_75t_L g1990 ( 
.A(n_1791),
.Y(n_1990)
);

A2O1A1Ixp33_ASAP7_75t_SL g1991 ( 
.A1(n_1756),
.A2(n_1797),
.B(n_1829),
.C(n_1813),
.Y(n_1991)
);

INVx8_ASAP7_75t_L g1992 ( 
.A(n_1791),
.Y(n_1992)
);

CKINVDCx5p33_ASAP7_75t_R g1993 ( 
.A(n_1769),
.Y(n_1993)
);

BUFx6f_ASAP7_75t_L g1994 ( 
.A(n_1791),
.Y(n_1994)
);

NAND2xp5_ASAP7_75t_L g1995 ( 
.A(n_1806),
.B(n_150),
.Y(n_1995)
);

BUFx6f_ASAP7_75t_L g1996 ( 
.A(n_1811),
.Y(n_1996)
);

BUFx6f_ASAP7_75t_L g1997 ( 
.A(n_1811),
.Y(n_1997)
);

NOR2xp33_ASAP7_75t_L g1998 ( 
.A(n_1668),
.B(n_151),
.Y(n_1998)
);

AOI21xp5_ASAP7_75t_L g1999 ( 
.A1(n_1680),
.A2(n_388),
.B(n_385),
.Y(n_1999)
);

AOI21xp5_ASAP7_75t_L g2000 ( 
.A1(n_1680),
.A2(n_392),
.B(n_391),
.Y(n_2000)
);

BUFx3_ASAP7_75t_L g2001 ( 
.A(n_1855),
.Y(n_2001)
);

BUFx2_ASAP7_75t_L g2002 ( 
.A(n_1801),
.Y(n_2002)
);

NAND2xp5_ASAP7_75t_SL g2003 ( 
.A(n_1867),
.B(n_152),
.Y(n_2003)
);

INVx1_ASAP7_75t_L g2004 ( 
.A(n_1848),
.Y(n_2004)
);

BUFx6f_ASAP7_75t_L g2005 ( 
.A(n_1811),
.Y(n_2005)
);

NAND2xp5_ASAP7_75t_L g2006 ( 
.A(n_1823),
.B(n_1834),
.Y(n_2006)
);

INVx2_ASAP7_75t_L g2007 ( 
.A(n_1705),
.Y(n_2007)
);

BUFx6f_ASAP7_75t_L g2008 ( 
.A(n_1865),
.Y(n_2008)
);

BUFx6f_ASAP7_75t_L g2009 ( 
.A(n_1865),
.Y(n_2009)
);

INVx1_ASAP7_75t_L g2010 ( 
.A(n_1827),
.Y(n_2010)
);

INVx6_ASAP7_75t_L g2011 ( 
.A(n_1822),
.Y(n_2011)
);

BUFx12f_ASAP7_75t_L g2012 ( 
.A(n_1835),
.Y(n_2012)
);

CKINVDCx14_ASAP7_75t_R g2013 ( 
.A(n_1772),
.Y(n_2013)
);

OAI22xp5_ASAP7_75t_L g2014 ( 
.A1(n_1818),
.A2(n_152),
.B1(n_153),
.B2(n_154),
.Y(n_2014)
);

OAI21xp5_ASAP7_75t_L g2015 ( 
.A1(n_1682),
.A2(n_154),
.B(n_155),
.Y(n_2015)
);

INVx3_ASAP7_75t_L g2016 ( 
.A(n_1767),
.Y(n_2016)
);

AND2x4_ASAP7_75t_L g2017 ( 
.A(n_1767),
.B(n_157),
.Y(n_2017)
);

NOR2xp33_ASAP7_75t_L g2018 ( 
.A(n_1783),
.B(n_158),
.Y(n_2018)
);

BUFx3_ASAP7_75t_L g2019 ( 
.A(n_1851),
.Y(n_2019)
);

BUFx2_ASAP7_75t_L g2020 ( 
.A(n_1867),
.Y(n_2020)
);

NAND2xp5_ASAP7_75t_L g2021 ( 
.A(n_1836),
.B(n_159),
.Y(n_2021)
);

OAI21x1_ASAP7_75t_L g2022 ( 
.A1(n_1726),
.A2(n_471),
.B(n_469),
.Y(n_2022)
);

INVx3_ASAP7_75t_L g2023 ( 
.A(n_1767),
.Y(n_2023)
);

NAND2xp5_ASAP7_75t_L g2024 ( 
.A(n_1709),
.B(n_162),
.Y(n_2024)
);

NOR2xp33_ASAP7_75t_L g2025 ( 
.A(n_1747),
.B(n_163),
.Y(n_2025)
);

BUFx6f_ASAP7_75t_L g2026 ( 
.A(n_1865),
.Y(n_2026)
);

NAND2xp5_ASAP7_75t_SL g2027 ( 
.A(n_1901),
.B(n_164),
.Y(n_2027)
);

INVx3_ASAP7_75t_L g2028 ( 
.A(n_1774),
.Y(n_2028)
);

NAND2xp5_ASAP7_75t_L g2029 ( 
.A(n_1697),
.B(n_165),
.Y(n_2029)
);

OR2x6_ASAP7_75t_L g2030 ( 
.A(n_1822),
.B(n_165),
.Y(n_2030)
);

NAND2xp5_ASAP7_75t_L g2031 ( 
.A(n_1703),
.B(n_166),
.Y(n_2031)
);

INVx4_ASAP7_75t_L g2032 ( 
.A(n_1774),
.Y(n_2032)
);

BUFx10_ASAP7_75t_L g2033 ( 
.A(n_1881),
.Y(n_2033)
);

O2A1O1Ixp33_ASAP7_75t_L g2034 ( 
.A1(n_1868),
.A2(n_167),
.B(n_168),
.C(n_169),
.Y(n_2034)
);

A2O1A1Ixp33_ASAP7_75t_L g2035 ( 
.A1(n_1701),
.A2(n_168),
.B(n_169),
.C(n_170),
.Y(n_2035)
);

NAND2xp5_ASAP7_75t_SL g2036 ( 
.A(n_1901),
.B(n_170),
.Y(n_2036)
);

AOI22xp33_ASAP7_75t_L g2037 ( 
.A1(n_1825),
.A2(n_171),
.B1(n_172),
.B2(n_173),
.Y(n_2037)
);

NAND2xp5_ASAP7_75t_L g2038 ( 
.A(n_1856),
.B(n_173),
.Y(n_2038)
);

O2A1O1Ixp33_ASAP7_75t_L g2039 ( 
.A1(n_1832),
.A2(n_174),
.B(n_175),
.C(n_176),
.Y(n_2039)
);

NAND2xp5_ASAP7_75t_SL g2040 ( 
.A(n_1905),
.B(n_174),
.Y(n_2040)
);

AND2x4_ASAP7_75t_L g2041 ( 
.A(n_1873),
.B(n_175),
.Y(n_2041)
);

INVx1_ASAP7_75t_L g2042 ( 
.A(n_1827),
.Y(n_2042)
);

A2O1A1Ixp33_ASAP7_75t_L g2043 ( 
.A1(n_1686),
.A2(n_177),
.B(n_179),
.C(n_180),
.Y(n_2043)
);

NAND2xp5_ASAP7_75t_SL g2044 ( 
.A(n_1905),
.B(n_180),
.Y(n_2044)
);

NAND2xp5_ASAP7_75t_L g2045 ( 
.A(n_1862),
.B(n_181),
.Y(n_2045)
);

OAI22xp5_ASAP7_75t_L g2046 ( 
.A1(n_1663),
.A2(n_182),
.B1(n_183),
.B2(n_184),
.Y(n_2046)
);

NOR3xp33_ASAP7_75t_L g2047 ( 
.A(n_1840),
.B(n_183),
.C(n_184),
.Y(n_2047)
);

INVxp67_ASAP7_75t_SL g2048 ( 
.A(n_1674),
.Y(n_2048)
);

INVx1_ASAP7_75t_L g2049 ( 
.A(n_1843),
.Y(n_2049)
);

AOI22xp33_ASAP7_75t_L g2050 ( 
.A1(n_1764),
.A2(n_185),
.B1(n_187),
.B2(n_188),
.Y(n_2050)
);

NAND2xp5_ASAP7_75t_L g2051 ( 
.A(n_1804),
.B(n_185),
.Y(n_2051)
);

NAND2xp5_ASAP7_75t_L g2052 ( 
.A(n_1693),
.B(n_187),
.Y(n_2052)
);

NOR2xp33_ASAP7_75t_L g2053 ( 
.A(n_1749),
.B(n_189),
.Y(n_2053)
);

AO21x1_ASAP7_75t_L g2054 ( 
.A1(n_1751),
.A2(n_189),
.B(n_190),
.Y(n_2054)
);

AOI21xp5_ASAP7_75t_L g2055 ( 
.A1(n_1729),
.A2(n_462),
.B(n_459),
.Y(n_2055)
);

NOR2xp33_ASAP7_75t_R g2056 ( 
.A(n_1784),
.B(n_193),
.Y(n_2056)
);

NOR2xp33_ASAP7_75t_L g2057 ( 
.A(n_1808),
.B(n_193),
.Y(n_2057)
);

OAI22xp5_ASAP7_75t_SL g2058 ( 
.A1(n_1842),
.A2(n_194),
.B1(n_195),
.B2(n_196),
.Y(n_2058)
);

A2O1A1Ixp33_ASAP7_75t_L g2059 ( 
.A1(n_1912),
.A2(n_198),
.B(n_199),
.C(n_200),
.Y(n_2059)
);

O2A1O1Ixp33_ASAP7_75t_L g2060 ( 
.A1(n_1828),
.A2(n_200),
.B(n_203),
.C(n_204),
.Y(n_2060)
);

INVx1_ASAP7_75t_L g2061 ( 
.A(n_1843),
.Y(n_2061)
);

NOR3xp33_ASAP7_75t_SL g2062 ( 
.A(n_1889),
.B(n_203),
.C(n_204),
.Y(n_2062)
);

BUFx2_ASAP7_75t_L g2063 ( 
.A(n_1884),
.Y(n_2063)
);

NOR2x1_ASAP7_75t_SL g2064 ( 
.A(n_1873),
.B(n_205),
.Y(n_2064)
);

HB1xp67_ASAP7_75t_L g2065 ( 
.A(n_1739),
.Y(n_2065)
);

NAND2xp5_ASAP7_75t_SL g2066 ( 
.A(n_1745),
.B(n_205),
.Y(n_2066)
);

AOI21xp5_ASAP7_75t_L g2067 ( 
.A1(n_1706),
.A2(n_454),
.B(n_449),
.Y(n_2067)
);

NAND2xp5_ASAP7_75t_SL g2068 ( 
.A(n_1745),
.B(n_207),
.Y(n_2068)
);

O2A1O1Ixp33_ASAP7_75t_SL g2069 ( 
.A1(n_1821),
.A2(n_447),
.B(n_445),
.C(n_444),
.Y(n_2069)
);

NOR2xp33_ASAP7_75t_R g2070 ( 
.A(n_1661),
.B(n_1667),
.Y(n_2070)
);

BUFx8_ASAP7_75t_L g2071 ( 
.A(n_1923),
.Y(n_2071)
);

INVx1_ASAP7_75t_SL g2072 ( 
.A(n_1833),
.Y(n_2072)
);

AOI21xp5_ASAP7_75t_L g2073 ( 
.A1(n_1707),
.A2(n_1721),
.B(n_1717),
.Y(n_2073)
);

OAI22xp5_ASAP7_75t_L g2074 ( 
.A1(n_1777),
.A2(n_209),
.B1(n_210),
.B2(n_211),
.Y(n_2074)
);

NOR2xp33_ASAP7_75t_SL g2075 ( 
.A(n_1896),
.B(n_209),
.Y(n_2075)
);

O2A1O1Ixp33_ASAP7_75t_L g2076 ( 
.A1(n_1773),
.A2(n_212),
.B(n_213),
.C(n_214),
.Y(n_2076)
);

NAND2xp5_ASAP7_75t_SL g2077 ( 
.A(n_1681),
.B(n_213),
.Y(n_2077)
);

BUFx6f_ASAP7_75t_L g2078 ( 
.A(n_1896),
.Y(n_2078)
);

OR2x6_ASAP7_75t_L g2079 ( 
.A(n_1838),
.B(n_219),
.Y(n_2079)
);

O2A1O1Ixp33_ASAP7_75t_L g2080 ( 
.A1(n_1754),
.A2(n_1863),
.B(n_1903),
.C(n_1687),
.Y(n_2080)
);

NAND2xp5_ASAP7_75t_L g2081 ( 
.A(n_1712),
.B(n_219),
.Y(n_2081)
);

NOR2x1p5_ASAP7_75t_L g2082 ( 
.A(n_1661),
.B(n_220),
.Y(n_2082)
);

HB1xp67_ASAP7_75t_L g2083 ( 
.A(n_1780),
.Y(n_2083)
);

BUFx4f_ASAP7_75t_L g2084 ( 
.A(n_1667),
.Y(n_2084)
);

OAI22xp5_ASAP7_75t_L g2085 ( 
.A1(n_1777),
.A2(n_220),
.B1(n_221),
.B2(n_222),
.Y(n_2085)
);

INVx3_ASAP7_75t_L g2086 ( 
.A(n_1884),
.Y(n_2086)
);

O2A1O1Ixp33_ASAP7_75t_L g2087 ( 
.A1(n_1837),
.A2(n_222),
.B(n_223),
.C(n_225),
.Y(n_2087)
);

NOR2xp33_ASAP7_75t_R g2088 ( 
.A(n_1880),
.B(n_223),
.Y(n_2088)
);

NAND2xp5_ASAP7_75t_L g2089 ( 
.A(n_1779),
.B(n_225),
.Y(n_2089)
);

NAND2xp5_ASAP7_75t_L g2090 ( 
.A(n_1770),
.B(n_229),
.Y(n_2090)
);

O2A1O1Ixp33_ASAP7_75t_L g2091 ( 
.A1(n_1924),
.A2(n_229),
.B(n_230),
.C(n_231),
.Y(n_2091)
);

NAND2xp5_ASAP7_75t_L g2092 ( 
.A(n_1683),
.B(n_230),
.Y(n_2092)
);

NAND2xp5_ASAP7_75t_L g2093 ( 
.A(n_1684),
.B(n_231),
.Y(n_2093)
);

NOR2xp33_ASAP7_75t_L g2094 ( 
.A(n_1676),
.B(n_232),
.Y(n_2094)
);

AND2x6_ASAP7_75t_SL g2095 ( 
.A(n_1845),
.B(n_1921),
.Y(n_2095)
);

AOI21xp5_ASAP7_75t_L g2096 ( 
.A1(n_1861),
.A2(n_404),
.B(n_440),
.Y(n_2096)
);

AOI21xp5_ASAP7_75t_L g2097 ( 
.A1(n_1759),
.A2(n_399),
.B(n_439),
.Y(n_2097)
);

NAND2xp5_ASAP7_75t_L g2098 ( 
.A(n_1685),
.B(n_233),
.Y(n_2098)
);

INVx1_ASAP7_75t_L g2099 ( 
.A(n_1871),
.Y(n_2099)
);

O2A1O1Ixp33_ASAP7_75t_L g2100 ( 
.A1(n_1824),
.A2(n_234),
.B(n_238),
.C(n_239),
.Y(n_2100)
);

OR2x2_ASAP7_75t_L g2101 ( 
.A(n_1928),
.B(n_238),
.Y(n_2101)
);

BUFx12f_ASAP7_75t_L g2102 ( 
.A(n_1830),
.Y(n_2102)
);

NAND2xp5_ASAP7_75t_L g2103 ( 
.A(n_1692),
.B(n_1870),
.Y(n_2103)
);

INVx2_ASAP7_75t_L g2104 ( 
.A(n_1814),
.Y(n_2104)
);

A2O1A1Ixp33_ASAP7_75t_L g2105 ( 
.A1(n_1912),
.A2(n_240),
.B(n_241),
.C(n_243),
.Y(n_2105)
);

AOI21xp5_ASAP7_75t_L g2106 ( 
.A1(n_1847),
.A2(n_409),
.B(n_438),
.Y(n_2106)
);

INVx1_ASAP7_75t_L g2107 ( 
.A(n_1871),
.Y(n_2107)
);

NAND2xp5_ASAP7_75t_L g2108 ( 
.A(n_1870),
.B(n_241),
.Y(n_2108)
);

INVx2_ASAP7_75t_L g2109 ( 
.A(n_1820),
.Y(n_2109)
);

INVx2_ASAP7_75t_L g2110 ( 
.A(n_1850),
.Y(n_2110)
);

AOI21xp5_ASAP7_75t_L g2111 ( 
.A1(n_1694),
.A2(n_410),
.B(n_435),
.Y(n_2111)
);

AOI21xp5_ASAP7_75t_L g2112 ( 
.A1(n_1702),
.A2(n_407),
.B(n_434),
.Y(n_2112)
);

INVx2_ASAP7_75t_L g2113 ( 
.A(n_1885),
.Y(n_2113)
);

INVx2_ASAP7_75t_SL g2114 ( 
.A(n_1730),
.Y(n_2114)
);

NOR2xp33_ASAP7_75t_L g2115 ( 
.A(n_1732),
.B(n_246),
.Y(n_2115)
);

AND2x2_ASAP7_75t_SL g2116 ( 
.A(n_1894),
.B(n_246),
.Y(n_2116)
);

O2A1O1Ixp33_ASAP7_75t_L g2117 ( 
.A1(n_1890),
.A2(n_247),
.B(n_248),
.C(n_249),
.Y(n_2117)
);

BUFx6f_ASAP7_75t_L g2118 ( 
.A(n_1852),
.Y(n_2118)
);

INVx2_ASAP7_75t_L g2119 ( 
.A(n_1891),
.Y(n_2119)
);

NAND2xp5_ASAP7_75t_L g2120 ( 
.A(n_1715),
.B(n_248),
.Y(n_2120)
);

BUFx2_ASAP7_75t_L g2121 ( 
.A(n_1888),
.Y(n_2121)
);

INVx1_ASAP7_75t_L g2122 ( 
.A(n_1761),
.Y(n_2122)
);

NAND3xp33_ASAP7_75t_SL g2123 ( 
.A(n_1788),
.B(n_249),
.C(n_250),
.Y(n_2123)
);

A2O1A1Ixp33_ASAP7_75t_L g2124 ( 
.A1(n_1860),
.A2(n_250),
.B(n_251),
.C(n_252),
.Y(n_2124)
);

INVx3_ASAP7_75t_L g2125 ( 
.A(n_1888),
.Y(n_2125)
);

NAND2xp5_ASAP7_75t_L g2126 ( 
.A(n_1877),
.B(n_251),
.Y(n_2126)
);

NAND2xp5_ASAP7_75t_L g2127 ( 
.A(n_1748),
.B(n_252),
.Y(n_2127)
);

INVxp67_ASAP7_75t_L g2128 ( 
.A(n_1953),
.Y(n_2128)
);

AO21x2_ASAP7_75t_L g2129 ( 
.A1(n_2073),
.A2(n_1725),
.B(n_1771),
.Y(n_2129)
);

BUFx4f_ASAP7_75t_SL g2130 ( 
.A(n_2012),
.Y(n_2130)
);

OAI22xp5_ASAP7_75t_L g2131 ( 
.A1(n_2079),
.A2(n_1794),
.B1(n_1792),
.B2(n_1815),
.Y(n_2131)
);

O2A1O1Ixp33_ASAP7_75t_SL g2132 ( 
.A1(n_2059),
.A2(n_1892),
.B(n_1838),
.C(n_1841),
.Y(n_2132)
);

O2A1O1Ixp33_ASAP7_75t_SL g2133 ( 
.A1(n_2105),
.A2(n_1841),
.B(n_1853),
.C(n_1819),
.Y(n_2133)
);

INVx2_ASAP7_75t_SL g2134 ( 
.A(n_1992),
.Y(n_2134)
);

BUFx12f_ASAP7_75t_L g2135 ( 
.A(n_2030),
.Y(n_2135)
);

AOI21xp5_ASAP7_75t_L g2136 ( 
.A1(n_1991),
.A2(n_1831),
.B(n_1925),
.Y(n_2136)
);

INVx1_ASAP7_75t_SL g2137 ( 
.A(n_2020),
.Y(n_2137)
);

AOI21x1_ASAP7_75t_L g2138 ( 
.A1(n_1938),
.A2(n_1763),
.B(n_1768),
.Y(n_2138)
);

NAND2xp5_ASAP7_75t_L g2139 ( 
.A(n_1959),
.B(n_1766),
.Y(n_2139)
);

INVx3_ASAP7_75t_SL g2140 ( 
.A(n_1992),
.Y(n_2140)
);

A2O1A1Ixp33_ASAP7_75t_L g2141 ( 
.A1(n_1964),
.A2(n_1981),
.B(n_2080),
.C(n_2087),
.Y(n_2141)
);

AOI21xp33_ASAP7_75t_L g2142 ( 
.A1(n_1961),
.A2(n_1758),
.B(n_1882),
.Y(n_2142)
);

O2A1O1Ixp5_ASAP7_75t_SL g2143 ( 
.A1(n_2014),
.A2(n_1799),
.B(n_1778),
.C(n_1785),
.Y(n_2143)
);

AOI21xp5_ASAP7_75t_SL g2144 ( 
.A1(n_2079),
.A2(n_1853),
.B(n_1819),
.Y(n_2144)
);

INVx1_ASAP7_75t_L g2145 ( 
.A(n_1930),
.Y(n_2145)
);

NOR2xp67_ASAP7_75t_L g2146 ( 
.A(n_2032),
.B(n_1810),
.Y(n_2146)
);

OAI21xp5_ASAP7_75t_L g2147 ( 
.A1(n_2015),
.A2(n_1914),
.B(n_1689),
.Y(n_2147)
);

AO31x2_ASAP7_75t_L g2148 ( 
.A1(n_2054),
.A2(n_1782),
.A3(n_1790),
.B(n_1798),
.Y(n_2148)
);

NOR2xp67_ASAP7_75t_SL g2149 ( 
.A(n_2032),
.B(n_1826),
.Y(n_2149)
);

O2A1O1Ixp5_ASAP7_75t_SL g2150 ( 
.A1(n_2066),
.A2(n_2068),
.B(n_1971),
.C(n_2036),
.Y(n_2150)
);

AOI21xp5_ASAP7_75t_L g2151 ( 
.A1(n_1947),
.A2(n_1917),
.B(n_1672),
.Y(n_2151)
);

AOI21xp5_ASAP7_75t_SL g2152 ( 
.A1(n_2017),
.A2(n_2082),
.B(n_2124),
.Y(n_2152)
);

OAI22x1_ASAP7_75t_L g2153 ( 
.A1(n_2072),
.A2(n_1949),
.B1(n_1932),
.B2(n_1969),
.Y(n_2153)
);

NOR2xp33_ASAP7_75t_L g2154 ( 
.A(n_1979),
.B(n_1753),
.Y(n_2154)
);

INVx4_ASAP7_75t_L g2155 ( 
.A(n_1992),
.Y(n_2155)
);

HB1xp67_ASAP7_75t_L g2156 ( 
.A(n_2065),
.Y(n_2156)
);

OAI21xp5_ASAP7_75t_L g2157 ( 
.A1(n_2077),
.A2(n_1910),
.B(n_1898),
.Y(n_2157)
);

NAND3x1_ASAP7_75t_L g2158 ( 
.A(n_1969),
.B(n_1920),
.C(n_1858),
.Y(n_2158)
);

OA21x2_ASAP7_75t_L g2159 ( 
.A1(n_2022),
.A2(n_1742),
.B(n_1731),
.Y(n_2159)
);

OAI21x1_ASAP7_75t_SL g2160 ( 
.A1(n_2064),
.A2(n_1964),
.B(n_2046),
.Y(n_2160)
);

INVx1_ASAP7_75t_L g2161 ( 
.A(n_1955),
.Y(n_2161)
);

INVx5_ASAP7_75t_L g2162 ( 
.A(n_1990),
.Y(n_2162)
);

NOR2xp33_ASAP7_75t_L g2163 ( 
.A(n_2095),
.B(n_1755),
.Y(n_2163)
);

AOI22xp5_ASAP7_75t_L g2164 ( 
.A1(n_2094),
.A2(n_1716),
.B1(n_1929),
.B2(n_1919),
.Y(n_2164)
);

NOR2xp67_ASAP7_75t_L g2165 ( 
.A(n_1944),
.B(n_1893),
.Y(n_2165)
);

A2O1A1Ixp33_ASAP7_75t_L g2166 ( 
.A1(n_2060),
.A2(n_2076),
.B(n_1982),
.C(n_2034),
.Y(n_2166)
);

NAND2xp5_ASAP7_75t_L g2167 ( 
.A(n_1967),
.B(n_1895),
.Y(n_2167)
);

NAND3xp33_ASAP7_75t_L g2168 ( 
.A(n_2062),
.B(n_1897),
.C(n_1887),
.Y(n_2168)
);

NAND2x1_ASAP7_75t_L g2169 ( 
.A(n_2016),
.B(n_1852),
.Y(n_2169)
);

NAND2x1p5_ASAP7_75t_L g2170 ( 
.A(n_1944),
.B(n_1876),
.Y(n_2170)
);

OAI22xp33_ASAP7_75t_L g2171 ( 
.A1(n_1966),
.A2(n_1724),
.B1(n_1776),
.B2(n_1744),
.Y(n_2171)
);

INVx3_ASAP7_75t_L g2172 ( 
.A(n_2084),
.Y(n_2172)
);

BUFx3_ASAP7_75t_L g2173 ( 
.A(n_2001),
.Y(n_2173)
);

A2O1A1Ixp33_ASAP7_75t_L g2174 ( 
.A1(n_2117),
.A2(n_1907),
.B(n_1713),
.C(n_1899),
.Y(n_2174)
);

A2O1A1Ixp33_ASAP7_75t_L g2175 ( 
.A1(n_1965),
.A2(n_1698),
.B(n_1800),
.C(n_1795),
.Y(n_2175)
);

AND2x2_ASAP7_75t_L g2176 ( 
.A(n_1958),
.B(n_253),
.Y(n_2176)
);

AOI21xp5_ASAP7_75t_L g2177 ( 
.A1(n_1939),
.A2(n_1741),
.B(n_1786),
.Y(n_2177)
);

BUFx6f_ASAP7_75t_L g2178 ( 
.A(n_1990),
.Y(n_2178)
);

INVx3_ASAP7_75t_L g2179 ( 
.A(n_2084),
.Y(n_2179)
);

O2A1O1Ixp33_ASAP7_75t_L g2180 ( 
.A1(n_2025),
.A2(n_1883),
.B(n_1906),
.C(n_1911),
.Y(n_2180)
);

INVx1_ASAP7_75t_L g2181 ( 
.A(n_1974),
.Y(n_2181)
);

INVx2_ASAP7_75t_L g2182 ( 
.A(n_1933),
.Y(n_2182)
);

INVx2_ASAP7_75t_SL g2183 ( 
.A(n_1931),
.Y(n_2183)
);

AND2x4_ASAP7_75t_L g2184 ( 
.A(n_1935),
.B(n_1908),
.Y(n_2184)
);

INVx2_ASAP7_75t_L g2185 ( 
.A(n_1962),
.Y(n_2185)
);

BUFx3_ASAP7_75t_L g2186 ( 
.A(n_2019),
.Y(n_2186)
);

AO31x2_ASAP7_75t_L g2187 ( 
.A1(n_2103),
.A2(n_1666),
.A3(n_1915),
.B(n_1849),
.Y(n_2187)
);

BUFx3_ASAP7_75t_L g2188 ( 
.A(n_2071),
.Y(n_2188)
);

AOI21x1_ASAP7_75t_L g2189 ( 
.A1(n_2055),
.A2(n_1846),
.B(n_1916),
.Y(n_2189)
);

NOR2xp33_ASAP7_75t_SL g2190 ( 
.A(n_2075),
.B(n_1876),
.Y(n_2190)
);

INVxp67_ASAP7_75t_L g2191 ( 
.A(n_1977),
.Y(n_2191)
);

AOI21xp5_ASAP7_75t_L g2192 ( 
.A1(n_1939),
.A2(n_1723),
.B(n_1736),
.Y(n_2192)
);

AOI21xp5_ASAP7_75t_L g2193 ( 
.A1(n_1939),
.A2(n_1859),
.B(n_1690),
.Y(n_2193)
);

AOI21xp5_ASAP7_75t_L g2194 ( 
.A1(n_2106),
.A2(n_1857),
.B(n_1743),
.Y(n_2194)
);

O2A1O1Ixp33_ASAP7_75t_SL g2195 ( 
.A1(n_1985),
.A2(n_1809),
.B(n_1926),
.C(n_1886),
.Y(n_2195)
);

BUFx2_ASAP7_75t_L g2196 ( 
.A(n_2070),
.Y(n_2196)
);

BUFx6f_ASAP7_75t_L g2197 ( 
.A(n_1990),
.Y(n_2197)
);

NAND2xp5_ASAP7_75t_L g2198 ( 
.A(n_2004),
.B(n_1950),
.Y(n_2198)
);

BUFx3_ASAP7_75t_L g2199 ( 
.A(n_2071),
.Y(n_2199)
);

INVx1_ASAP7_75t_L g2200 ( 
.A(n_1957),
.Y(n_2200)
);

BUFx10_ASAP7_75t_L g2201 ( 
.A(n_2041),
.Y(n_2201)
);

AOI21xp5_ASAP7_75t_L g2202 ( 
.A1(n_1945),
.A2(n_1879),
.B(n_1708),
.Y(n_2202)
);

INVx4_ASAP7_75t_L g2203 ( 
.A(n_1994),
.Y(n_2203)
);

INVx2_ASAP7_75t_L g2204 ( 
.A(n_1973),
.Y(n_2204)
);

A2O1A1Ixp33_ASAP7_75t_L g2205 ( 
.A1(n_2039),
.A2(n_1878),
.B(n_1900),
.C(n_1875),
.Y(n_2205)
);

NAND2xp5_ASAP7_75t_L g2206 ( 
.A(n_2006),
.B(n_1874),
.Y(n_2206)
);

AOI21xp5_ASAP7_75t_L g2207 ( 
.A1(n_1954),
.A2(n_1708),
.B(n_1913),
.Y(n_2207)
);

CKINVDCx16_ASAP7_75t_R g2208 ( 
.A(n_2056),
.Y(n_2208)
);

AOI21xp5_ASAP7_75t_L g2209 ( 
.A1(n_1936),
.A2(n_1909),
.B(n_1866),
.Y(n_2209)
);

NOR4xp25_ASAP7_75t_L g2210 ( 
.A(n_1984),
.B(n_1854),
.C(n_1927),
.D(n_1908),
.Y(n_2210)
);

OAI21xp5_ASAP7_75t_L g2211 ( 
.A1(n_1941),
.A2(n_1722),
.B(n_1869),
.Y(n_2211)
);

NAND2x1p5_ASAP7_75t_L g2212 ( 
.A(n_2028),
.B(n_1922),
.Y(n_2212)
);

A2O1A1Ixp33_ASAP7_75t_L g2213 ( 
.A1(n_1987),
.A2(n_1872),
.B(n_1918),
.C(n_1904),
.Y(n_2213)
);

BUFx10_ASAP7_75t_L g2214 ( 
.A(n_2041),
.Y(n_2214)
);

AOI21xp5_ASAP7_75t_L g2215 ( 
.A1(n_1972),
.A2(n_1728),
.B(n_1733),
.Y(n_2215)
);

NOR2xp33_ASAP7_75t_L g2216 ( 
.A(n_2114),
.B(n_1993),
.Y(n_2216)
);

O2A1O1Ixp33_ASAP7_75t_L g2217 ( 
.A1(n_2053),
.A2(n_1710),
.B(n_1830),
.C(n_255),
.Y(n_2217)
);

AND2x4_ASAP7_75t_L g2218 ( 
.A(n_1935),
.B(n_1830),
.Y(n_2218)
);

OAI21x1_ASAP7_75t_L g2219 ( 
.A1(n_2097),
.A2(n_1830),
.B(n_416),
.Y(n_2219)
);

O2A1O1Ixp33_ASAP7_75t_SL g2220 ( 
.A1(n_2035),
.A2(n_253),
.B(n_254),
.C(n_256),
.Y(n_2220)
);

INVx2_ASAP7_75t_L g2221 ( 
.A(n_1976),
.Y(n_2221)
);

NAND2xp5_ASAP7_75t_L g2222 ( 
.A(n_2010),
.B(n_395),
.Y(n_2222)
);

BUFx6f_ASAP7_75t_L g2223 ( 
.A(n_1994),
.Y(n_2223)
);

OAI21x1_ASAP7_75t_L g2224 ( 
.A1(n_2067),
.A2(n_396),
.B(n_398),
.Y(n_2224)
);

AOI21xp5_ASAP7_75t_L g2225 ( 
.A1(n_2042),
.A2(n_405),
.B(n_411),
.Y(n_2225)
);

AND2x4_ASAP7_75t_L g2226 ( 
.A(n_2016),
.B(n_413),
.Y(n_2226)
);

NAND3x1_ASAP7_75t_L g2227 ( 
.A(n_1989),
.B(n_414),
.C(n_417),
.Y(n_2227)
);

O2A1O1Ixp33_ASAP7_75t_SL g2228 ( 
.A1(n_1963),
.A2(n_418),
.B(n_422),
.C(n_423),
.Y(n_2228)
);

AO32x2_ASAP7_75t_L g2229 ( 
.A1(n_2058),
.A2(n_424),
.A3(n_427),
.B1(n_430),
.B2(n_431),
.Y(n_2229)
);

NAND3xp33_ASAP7_75t_L g2230 ( 
.A(n_2047),
.B(n_1978),
.C(n_2050),
.Y(n_2230)
);

INVx1_ASAP7_75t_L g2231 ( 
.A(n_1943),
.Y(n_2231)
);

OAI21xp5_ASAP7_75t_L g2232 ( 
.A1(n_2127),
.A2(n_2043),
.B(n_2090),
.Y(n_2232)
);

AOI21xp5_ASAP7_75t_L g2233 ( 
.A1(n_2049),
.A2(n_2061),
.B(n_1952),
.Y(n_2233)
);

AOI21xp5_ASAP7_75t_L g2234 ( 
.A1(n_1948),
.A2(n_1956),
.B(n_2096),
.Y(n_2234)
);

BUFx8_ASAP7_75t_L g2235 ( 
.A(n_1986),
.Y(n_2235)
);

NAND2xp5_ASAP7_75t_L g2236 ( 
.A(n_1951),
.B(n_2122),
.Y(n_2236)
);

BUFx2_ASAP7_75t_L g2237 ( 
.A(n_1994),
.Y(n_2237)
);

AOI221x1_ASAP7_75t_L g2238 ( 
.A1(n_1980),
.A2(n_2123),
.B1(n_2074),
.B2(n_2085),
.C(n_2108),
.Y(n_2238)
);

O2A1O1Ixp33_ASAP7_75t_SL g2239 ( 
.A1(n_2003),
.A2(n_2044),
.B(n_2027),
.C(n_2040),
.Y(n_2239)
);

OAI22xp5_ASAP7_75t_L g2240 ( 
.A1(n_2037),
.A2(n_2116),
.B1(n_2018),
.B2(n_2021),
.Y(n_2240)
);

AOI21xp5_ASAP7_75t_L g2241 ( 
.A1(n_2099),
.A2(n_2107),
.B(n_2069),
.Y(n_2241)
);

AOI21xp5_ASAP7_75t_L g2242 ( 
.A1(n_2081),
.A2(n_2092),
.B(n_2098),
.Y(n_2242)
);

OAI21x1_ASAP7_75t_L g2243 ( 
.A1(n_2111),
.A2(n_2112),
.B(n_2000),
.Y(n_2243)
);

A2O1A1Ixp33_ASAP7_75t_L g2244 ( 
.A1(n_2100),
.A2(n_2091),
.B(n_2115),
.C(n_1998),
.Y(n_2244)
);

INVx2_ASAP7_75t_L g2245 ( 
.A(n_2007),
.Y(n_2245)
);

AO31x2_ASAP7_75t_L g2246 ( 
.A1(n_1937),
.A2(n_1999),
.A3(n_2093),
.B(n_2029),
.Y(n_2246)
);

CKINVDCx20_ASAP7_75t_R g2247 ( 
.A(n_2130),
.Y(n_2247)
);

INVx2_ASAP7_75t_L g2248 ( 
.A(n_2182),
.Y(n_2248)
);

INVx1_ASAP7_75t_L g2249 ( 
.A(n_2161),
.Y(n_2249)
);

INVx1_ASAP7_75t_L g2250 ( 
.A(n_2181),
.Y(n_2250)
);

INVx1_ASAP7_75t_L g2251 ( 
.A(n_2231),
.Y(n_2251)
);

INVx1_ASAP7_75t_L g2252 ( 
.A(n_2145),
.Y(n_2252)
);

OAI22xp33_ASAP7_75t_L g2253 ( 
.A1(n_2208),
.A2(n_2002),
.B1(n_2101),
.B2(n_2102),
.Y(n_2253)
);

CKINVDCx5p33_ASAP7_75t_R g2254 ( 
.A(n_2188),
.Y(n_2254)
);

AND2x2_ASAP7_75t_L g2255 ( 
.A(n_2156),
.B(n_2083),
.Y(n_2255)
);

AOI22xp33_ASAP7_75t_L g2256 ( 
.A1(n_2131),
.A2(n_2088),
.B1(n_2017),
.B2(n_2033),
.Y(n_2256)
);

AOI22xp33_ASAP7_75t_SL g2257 ( 
.A1(n_2160),
.A2(n_2033),
.B1(n_2013),
.B2(n_1983),
.Y(n_2257)
);

AOI22xp33_ASAP7_75t_SL g2258 ( 
.A1(n_2135),
.A2(n_1946),
.B1(n_2063),
.B2(n_2023),
.Y(n_2258)
);

INVx2_ASAP7_75t_L g2259 ( 
.A(n_2245),
.Y(n_2259)
);

INVx6_ASAP7_75t_L g2260 ( 
.A(n_2235),
.Y(n_2260)
);

INVx1_ASAP7_75t_L g2261 ( 
.A(n_2185),
.Y(n_2261)
);

CKINVDCx5p33_ASAP7_75t_R g2262 ( 
.A(n_2199),
.Y(n_2262)
);

INVx1_ASAP7_75t_L g2263 ( 
.A(n_2204),
.Y(n_2263)
);

INVx2_ASAP7_75t_L g2264 ( 
.A(n_2221),
.Y(n_2264)
);

AOI22xp33_ASAP7_75t_L g2265 ( 
.A1(n_2230),
.A2(n_2089),
.B1(n_2057),
.B2(n_1968),
.Y(n_2265)
);

OAI22xp5_ASAP7_75t_L g2266 ( 
.A1(n_2144),
.A2(n_2051),
.B1(n_2048),
.B2(n_2120),
.Y(n_2266)
);

OAI22xp5_ASAP7_75t_L g2267 ( 
.A1(n_2158),
.A2(n_2052),
.B1(n_2024),
.B2(n_2031),
.Y(n_2267)
);

BUFx4f_ASAP7_75t_L g2268 ( 
.A(n_2140),
.Y(n_2268)
);

NAND2x1p5_ASAP7_75t_L g2269 ( 
.A(n_2196),
.B(n_2028),
.Y(n_2269)
);

AOI22xp33_ASAP7_75t_L g2270 ( 
.A1(n_2163),
.A2(n_2126),
.B1(n_1934),
.B2(n_1995),
.Y(n_2270)
);

AOI22xp33_ASAP7_75t_L g2271 ( 
.A1(n_2153),
.A2(n_1975),
.B1(n_1988),
.B2(n_1970),
.Y(n_2271)
);

INVx1_ASAP7_75t_L g2272 ( 
.A(n_2236),
.Y(n_2272)
);

BUFx8_ASAP7_75t_SL g2273 ( 
.A(n_2173),
.Y(n_2273)
);

BUFx10_ASAP7_75t_L g2274 ( 
.A(n_2183),
.Y(n_2274)
);

INVx1_ASAP7_75t_L g2275 ( 
.A(n_2200),
.Y(n_2275)
);

INVx1_ASAP7_75t_L g2276 ( 
.A(n_2198),
.Y(n_2276)
);

OAI22xp5_ASAP7_75t_L g2277 ( 
.A1(n_2164),
.A2(n_2045),
.B1(n_2038),
.B2(n_2086),
.Y(n_2277)
);

INVx2_ASAP7_75t_L g2278 ( 
.A(n_2167),
.Y(n_2278)
);

INVx1_ASAP7_75t_L g2279 ( 
.A(n_2206),
.Y(n_2279)
);

INVx1_ASAP7_75t_L g2280 ( 
.A(n_2128),
.Y(n_2280)
);

BUFx12f_ASAP7_75t_L g2281 ( 
.A(n_2201),
.Y(n_2281)
);

INVx1_ASAP7_75t_L g2282 ( 
.A(n_2191),
.Y(n_2282)
);

INVx4_ASAP7_75t_L g2283 ( 
.A(n_2162),
.Y(n_2283)
);

BUFx6f_ASAP7_75t_L g2284 ( 
.A(n_2155),
.Y(n_2284)
);

CKINVDCx11_ASAP7_75t_R g2285 ( 
.A(n_2214),
.Y(n_2285)
);

INVx6_ASAP7_75t_L g2286 ( 
.A(n_2235),
.Y(n_2286)
);

INVx4_ASAP7_75t_L g2287 ( 
.A(n_2162),
.Y(n_2287)
);

INVx6_ASAP7_75t_L g2288 ( 
.A(n_2162),
.Y(n_2288)
);

CKINVDCx11_ASAP7_75t_R g2289 ( 
.A(n_2186),
.Y(n_2289)
);

INVx1_ASAP7_75t_L g2290 ( 
.A(n_2233),
.Y(n_2290)
);

CKINVDCx11_ASAP7_75t_R g2291 ( 
.A(n_2137),
.Y(n_2291)
);

CKINVDCx11_ASAP7_75t_R g2292 ( 
.A(n_2178),
.Y(n_2292)
);

INVx1_ASAP7_75t_L g2293 ( 
.A(n_2226),
.Y(n_2293)
);

OAI22xp33_ASAP7_75t_L g2294 ( 
.A1(n_2190),
.A2(n_1940),
.B1(n_2011),
.B2(n_1960),
.Y(n_2294)
);

CKINVDCx20_ASAP7_75t_R g2295 ( 
.A(n_2134),
.Y(n_2295)
);

INVx1_ASAP7_75t_L g2296 ( 
.A(n_2226),
.Y(n_2296)
);

NAND2xp5_ASAP7_75t_L g2297 ( 
.A(n_2139),
.B(n_2110),
.Y(n_2297)
);

AOI22xp33_ASAP7_75t_L g2298 ( 
.A1(n_2240),
.A2(n_2121),
.B1(n_2119),
.B2(n_2113),
.Y(n_2298)
);

INVx1_ASAP7_75t_L g2299 ( 
.A(n_2149),
.Y(n_2299)
);

BUFx2_ASAP7_75t_SL g2300 ( 
.A(n_2172),
.Y(n_2300)
);

BUFx3_ASAP7_75t_L g2301 ( 
.A(n_2237),
.Y(n_2301)
);

INVx2_ASAP7_75t_L g2302 ( 
.A(n_2178),
.Y(n_2302)
);

AOI22xp33_ASAP7_75t_L g2303 ( 
.A1(n_2168),
.A2(n_2125),
.B1(n_1960),
.B2(n_2104),
.Y(n_2303)
);

INVx1_ASAP7_75t_SL g2304 ( 
.A(n_2178),
.Y(n_2304)
);

BUFx12f_ASAP7_75t_L g2305 ( 
.A(n_2203),
.Y(n_2305)
);

INVx2_ASAP7_75t_SL g2306 ( 
.A(n_2179),
.Y(n_2306)
);

CKINVDCx6p67_ASAP7_75t_R g2307 ( 
.A(n_2218),
.Y(n_2307)
);

INVx1_ASAP7_75t_L g2308 ( 
.A(n_2184),
.Y(n_2308)
);

NAND2xp5_ASAP7_75t_L g2309 ( 
.A(n_2141),
.B(n_2109),
.Y(n_2309)
);

BUFx6f_ASAP7_75t_SL g2310 ( 
.A(n_2218),
.Y(n_2310)
);

OAI22xp33_ASAP7_75t_L g2311 ( 
.A1(n_2146),
.A2(n_2078),
.B1(n_2118),
.B2(n_1997),
.Y(n_2311)
);

BUFx12f_ASAP7_75t_L g2312 ( 
.A(n_2197),
.Y(n_2312)
);

INVx1_ASAP7_75t_L g2313 ( 
.A(n_2184),
.Y(n_2313)
);

INVx1_ASAP7_75t_L g2314 ( 
.A(n_2176),
.Y(n_2314)
);

AOI22xp33_ASAP7_75t_L g2315 ( 
.A1(n_2232),
.A2(n_2078),
.B1(n_2118),
.B2(n_1997),
.Y(n_2315)
);

AOI22xp33_ASAP7_75t_L g2316 ( 
.A1(n_2154),
.A2(n_2078),
.B1(n_2118),
.B2(n_1997),
.Y(n_2316)
);

OAI22xp33_ASAP7_75t_L g2317 ( 
.A1(n_2238),
.A2(n_2165),
.B1(n_2147),
.B2(n_2171),
.Y(n_2317)
);

BUFx8_ASAP7_75t_SL g2318 ( 
.A(n_2197),
.Y(n_2318)
);

AOI22xp33_ASAP7_75t_SL g2319 ( 
.A1(n_2152),
.A2(n_2009),
.B1(n_1996),
.B2(n_2005),
.Y(n_2319)
);

OAI22xp5_ASAP7_75t_L g2320 ( 
.A1(n_2166),
.A2(n_2227),
.B1(n_2244),
.B2(n_2242),
.Y(n_2320)
);

INVx1_ASAP7_75t_L g2321 ( 
.A(n_2222),
.Y(n_2321)
);

INVx1_ASAP7_75t_L g2322 ( 
.A(n_2169),
.Y(n_2322)
);

INVx1_ASAP7_75t_L g2323 ( 
.A(n_2220),
.Y(n_2323)
);

INVx6_ASAP7_75t_L g2324 ( 
.A(n_2223),
.Y(n_2324)
);

CKINVDCx11_ASAP7_75t_R g2325 ( 
.A(n_2223),
.Y(n_2325)
);

BUFx6f_ASAP7_75t_L g2326 ( 
.A(n_2223),
.Y(n_2326)
);

INVx1_ASAP7_75t_L g2327 ( 
.A(n_2170),
.Y(n_2327)
);

OAI22xp5_ASAP7_75t_L g2328 ( 
.A1(n_2217),
.A2(n_2241),
.B1(n_2174),
.B2(n_2157),
.Y(n_2328)
);

INVx1_ASAP7_75t_L g2329 ( 
.A(n_2239),
.Y(n_2329)
);

INVx5_ASAP7_75t_L g2330 ( 
.A(n_2229),
.Y(n_2330)
);

NAND2xp5_ASAP7_75t_L g2331 ( 
.A(n_2148),
.B(n_2009),
.Y(n_2331)
);

OAI21xp5_ASAP7_75t_L g2332 ( 
.A1(n_2143),
.A2(n_1942),
.B(n_1996),
.Y(n_2332)
);

AND2x2_ASAP7_75t_SL g2333 ( 
.A(n_2268),
.B(n_2210),
.Y(n_2333)
);

BUFx6f_ASAP7_75t_L g2334 ( 
.A(n_2326),
.Y(n_2334)
);

AOI21x1_ASAP7_75t_L g2335 ( 
.A1(n_2320),
.A2(n_2177),
.B(n_2138),
.Y(n_2335)
);

AO21x2_ASAP7_75t_L g2336 ( 
.A1(n_2332),
.A2(n_2192),
.B(n_2193),
.Y(n_2336)
);

INVx1_ASAP7_75t_L g2337 ( 
.A(n_2290),
.Y(n_2337)
);

INVx3_ASAP7_75t_L g2338 ( 
.A(n_2330),
.Y(n_2338)
);

INVx4_ASAP7_75t_L g2339 ( 
.A(n_2326),
.Y(n_2339)
);

AND2x2_ASAP7_75t_L g2340 ( 
.A(n_2331),
.B(n_2129),
.Y(n_2340)
);

INVx1_ASAP7_75t_L g2341 ( 
.A(n_2249),
.Y(n_2341)
);

INVx1_ASAP7_75t_L g2342 ( 
.A(n_2250),
.Y(n_2342)
);

INVx1_ASAP7_75t_L g2343 ( 
.A(n_2251),
.Y(n_2343)
);

AND2x2_ASAP7_75t_L g2344 ( 
.A(n_2331),
.B(n_2148),
.Y(n_2344)
);

BUFx2_ASAP7_75t_L g2345 ( 
.A(n_2330),
.Y(n_2345)
);

INVx1_ASAP7_75t_L g2346 ( 
.A(n_2252),
.Y(n_2346)
);

AND2x2_ASAP7_75t_L g2347 ( 
.A(n_2330),
.B(n_2148),
.Y(n_2347)
);

INVx3_ASAP7_75t_L g2348 ( 
.A(n_2330),
.Y(n_2348)
);

INVx1_ASAP7_75t_L g2349 ( 
.A(n_2248),
.Y(n_2349)
);

INVx1_ASAP7_75t_L g2350 ( 
.A(n_2259),
.Y(n_2350)
);

INVx1_ASAP7_75t_L g2351 ( 
.A(n_2264),
.Y(n_2351)
);

NAND2xp5_ASAP7_75t_L g2352 ( 
.A(n_2276),
.B(n_2133),
.Y(n_2352)
);

NAND2x1p5_ASAP7_75t_L g2353 ( 
.A(n_2304),
.B(n_1996),
.Y(n_2353)
);

INVx3_ASAP7_75t_L g2354 ( 
.A(n_2326),
.Y(n_2354)
);

INVx1_ASAP7_75t_L g2355 ( 
.A(n_2261),
.Y(n_2355)
);

INVx1_ASAP7_75t_L g2356 ( 
.A(n_2263),
.Y(n_2356)
);

INVx1_ASAP7_75t_L g2357 ( 
.A(n_2275),
.Y(n_2357)
);

BUFx2_ASAP7_75t_L g2358 ( 
.A(n_2312),
.Y(n_2358)
);

INVx2_ASAP7_75t_L g2359 ( 
.A(n_2299),
.Y(n_2359)
);

AOI21x1_ASAP7_75t_L g2360 ( 
.A1(n_2320),
.A2(n_2209),
.B(n_2136),
.Y(n_2360)
);

INVx1_ASAP7_75t_L g2361 ( 
.A(n_2297),
.Y(n_2361)
);

INVx1_ASAP7_75t_L g2362 ( 
.A(n_2297),
.Y(n_2362)
);

INVx1_ASAP7_75t_L g2363 ( 
.A(n_2309),
.Y(n_2363)
);

INVx1_ASAP7_75t_L g2364 ( 
.A(n_2309),
.Y(n_2364)
);

NOR2xp33_ASAP7_75t_L g2365 ( 
.A(n_2253),
.B(n_2216),
.Y(n_2365)
);

INVx2_ASAP7_75t_L g2366 ( 
.A(n_2302),
.Y(n_2366)
);

AOI22xp33_ASAP7_75t_L g2367 ( 
.A1(n_2256),
.A2(n_2142),
.B1(n_2211),
.B2(n_2215),
.Y(n_2367)
);

AOI22xp33_ASAP7_75t_L g2368 ( 
.A1(n_2277),
.A2(n_2265),
.B1(n_2257),
.B2(n_2314),
.Y(n_2368)
);

AND2x2_ASAP7_75t_L g2369 ( 
.A(n_2279),
.B(n_2187),
.Y(n_2369)
);

BUFx12f_ASAP7_75t_L g2370 ( 
.A(n_2289),
.Y(n_2370)
);

OR2x2_ASAP7_75t_L g2371 ( 
.A(n_2278),
.B(n_2187),
.Y(n_2371)
);

OAI21x1_ASAP7_75t_L g2372 ( 
.A1(n_2328),
.A2(n_2151),
.B(n_2243),
.Y(n_2372)
);

INVx1_ASAP7_75t_L g2373 ( 
.A(n_2272),
.Y(n_2373)
);

AND2x2_ASAP7_75t_L g2374 ( 
.A(n_2308),
.B(n_2187),
.Y(n_2374)
);

AND2x2_ASAP7_75t_L g2375 ( 
.A(n_2313),
.B(n_2255),
.Y(n_2375)
);

INVx1_ASAP7_75t_L g2376 ( 
.A(n_2293),
.Y(n_2376)
);

HB1xp67_ASAP7_75t_L g2377 ( 
.A(n_2304),
.Y(n_2377)
);

INVx1_ASAP7_75t_L g2378 ( 
.A(n_2296),
.Y(n_2378)
);

INVx3_ASAP7_75t_L g2379 ( 
.A(n_2324),
.Y(n_2379)
);

AOI21x1_ASAP7_75t_L g2380 ( 
.A1(n_2267),
.A2(n_2189),
.B(n_2202),
.Y(n_2380)
);

INVx2_ASAP7_75t_L g2381 ( 
.A(n_2322),
.Y(n_2381)
);

OAI21x1_ASAP7_75t_L g2382 ( 
.A1(n_2266),
.A2(n_2234),
.B(n_2194),
.Y(n_2382)
);

INVx1_ASAP7_75t_L g2383 ( 
.A(n_2323),
.Y(n_2383)
);

INVx2_ASAP7_75t_L g2384 ( 
.A(n_2324),
.Y(n_2384)
);

OAI22xp33_ASAP7_75t_L g2385 ( 
.A1(n_2307),
.A2(n_2229),
.B1(n_2225),
.B2(n_2212),
.Y(n_2385)
);

INVx1_ASAP7_75t_L g2386 ( 
.A(n_2329),
.Y(n_2386)
);

INVx1_ASAP7_75t_L g2387 ( 
.A(n_2341),
.Y(n_2387)
);

INVx2_ASAP7_75t_L g2388 ( 
.A(n_2371),
.Y(n_2388)
);

AND2x2_ASAP7_75t_L g2389 ( 
.A(n_2375),
.B(n_2280),
.Y(n_2389)
);

AO32x2_ASAP7_75t_L g2390 ( 
.A1(n_2339),
.A2(n_2266),
.A3(n_2267),
.B1(n_2277),
.B2(n_2306),
.Y(n_2390)
);

AOI21xp5_ASAP7_75t_L g2391 ( 
.A1(n_2385),
.A2(n_2294),
.B(n_2311),
.Y(n_2391)
);

AO32x2_ASAP7_75t_L g2392 ( 
.A1(n_2339),
.A2(n_2287),
.A3(n_2283),
.B1(n_2282),
.B2(n_2317),
.Y(n_2392)
);

INVx1_ASAP7_75t_L g2393 ( 
.A(n_2341),
.Y(n_2393)
);

AO32x2_ASAP7_75t_L g2394 ( 
.A1(n_2339),
.A2(n_2283),
.A3(n_2287),
.B1(n_2271),
.B2(n_2298),
.Y(n_2394)
);

INVx2_ASAP7_75t_L g2395 ( 
.A(n_2371),
.Y(n_2395)
);

NAND4xp25_ASAP7_75t_L g2396 ( 
.A(n_2368),
.B(n_2270),
.C(n_2303),
.D(n_2258),
.Y(n_2396)
);

NOR2xp33_ASAP7_75t_SL g2397 ( 
.A(n_2370),
.B(n_2268),
.Y(n_2397)
);

AOI21xp5_ASAP7_75t_L g2398 ( 
.A1(n_2385),
.A2(n_2319),
.B(n_2228),
.Y(n_2398)
);

AND2x2_ASAP7_75t_L g2399 ( 
.A(n_2375),
.B(n_2301),
.Y(n_2399)
);

AND2x4_ASAP7_75t_L g2400 ( 
.A(n_2338),
.B(n_2315),
.Y(n_2400)
);

AND2x2_ASAP7_75t_L g2401 ( 
.A(n_2369),
.B(n_2321),
.Y(n_2401)
);

INVx2_ASAP7_75t_L g2402 ( 
.A(n_2371),
.Y(n_2402)
);

AND2x2_ASAP7_75t_L g2403 ( 
.A(n_2369),
.B(n_2246),
.Y(n_2403)
);

OAI21x1_ASAP7_75t_SL g2404 ( 
.A1(n_2368),
.A2(n_2286),
.B(n_2260),
.Y(n_2404)
);

A2O1A1Ixp33_ASAP7_75t_L g2405 ( 
.A1(n_2365),
.A2(n_2327),
.B(n_2300),
.C(n_2284),
.Y(n_2405)
);

OR2x6_ASAP7_75t_L g2406 ( 
.A(n_2345),
.B(n_2286),
.Y(n_2406)
);

AOI221xp5_ASAP7_75t_L g2407 ( 
.A1(n_2373),
.A2(n_2132),
.B1(n_2180),
.B2(n_2254),
.C(n_2262),
.Y(n_2407)
);

AOI22x1_ASAP7_75t_SL g2408 ( 
.A1(n_2370),
.A2(n_2247),
.B1(n_2295),
.B2(n_2260),
.Y(n_2408)
);

OAI21xp5_ASAP7_75t_L g2409 ( 
.A1(n_2333),
.A2(n_2150),
.B(n_2269),
.Y(n_2409)
);

AND2x2_ASAP7_75t_L g2410 ( 
.A(n_2369),
.B(n_2246),
.Y(n_2410)
);

A2O1A1Ixp33_ASAP7_75t_L g2411 ( 
.A1(n_2365),
.A2(n_2284),
.B(n_2316),
.C(n_2219),
.Y(n_2411)
);

AND2x2_ASAP7_75t_L g2412 ( 
.A(n_2374),
.B(n_2246),
.Y(n_2412)
);

AND2x2_ASAP7_75t_L g2413 ( 
.A(n_2374),
.B(n_2159),
.Y(n_2413)
);

AOI211xp5_ASAP7_75t_L g2414 ( 
.A1(n_2358),
.A2(n_2284),
.B(n_2205),
.C(n_2195),
.Y(n_2414)
);

AND2x2_ASAP7_75t_L g2415 ( 
.A(n_2374),
.B(n_2159),
.Y(n_2415)
);

AND2x2_ASAP7_75t_SL g2416 ( 
.A(n_2345),
.B(n_2310),
.Y(n_2416)
);

OAI22xp5_ASAP7_75t_L g2417 ( 
.A1(n_2333),
.A2(n_2260),
.B1(n_2286),
.B2(n_2269),
.Y(n_2417)
);

OAI22xp5_ASAP7_75t_SL g2418 ( 
.A1(n_2370),
.A2(n_2281),
.B1(n_2305),
.B2(n_2273),
.Y(n_2418)
);

INVx1_ASAP7_75t_L g2419 ( 
.A(n_2342),
.Y(n_2419)
);

AND2x2_ASAP7_75t_L g2420 ( 
.A(n_2412),
.B(n_2347),
.Y(n_2420)
);

BUFx2_ASAP7_75t_L g2421 ( 
.A(n_2406),
.Y(n_2421)
);

OAI22xp5_ASAP7_75t_L g2422 ( 
.A1(n_2405),
.A2(n_2333),
.B1(n_2358),
.B2(n_2310),
.Y(n_2422)
);

OR2x2_ASAP7_75t_L g2423 ( 
.A(n_2388),
.B(n_2361),
.Y(n_2423)
);

INVx1_ASAP7_75t_L g2424 ( 
.A(n_2387),
.Y(n_2424)
);

INVx1_ASAP7_75t_L g2425 ( 
.A(n_2393),
.Y(n_2425)
);

INVx1_ASAP7_75t_SL g2426 ( 
.A(n_2399),
.Y(n_2426)
);

INVx2_ASAP7_75t_L g2427 ( 
.A(n_2388),
.Y(n_2427)
);

INVx1_ASAP7_75t_L g2428 ( 
.A(n_2419),
.Y(n_2428)
);

INVx1_ASAP7_75t_L g2429 ( 
.A(n_2395),
.Y(n_2429)
);

NOR2xp33_ASAP7_75t_L g2430 ( 
.A(n_2397),
.B(n_2291),
.Y(n_2430)
);

INVx3_ASAP7_75t_L g2431 ( 
.A(n_2406),
.Y(n_2431)
);

NOR2xp33_ASAP7_75t_L g2432 ( 
.A(n_2408),
.B(n_2274),
.Y(n_2432)
);

NOR2xp33_ASAP7_75t_L g2433 ( 
.A(n_2418),
.B(n_2274),
.Y(n_2433)
);

AND2x2_ASAP7_75t_L g2434 ( 
.A(n_2412),
.B(n_2347),
.Y(n_2434)
);

INVx1_ASAP7_75t_L g2435 ( 
.A(n_2395),
.Y(n_2435)
);

INVx1_ASAP7_75t_SL g2436 ( 
.A(n_2406),
.Y(n_2436)
);

INVx1_ASAP7_75t_L g2437 ( 
.A(n_2402),
.Y(n_2437)
);

INVx1_ASAP7_75t_SL g2438 ( 
.A(n_2389),
.Y(n_2438)
);

INVx2_ASAP7_75t_SL g2439 ( 
.A(n_2416),
.Y(n_2439)
);

AND2x2_ASAP7_75t_L g2440 ( 
.A(n_2401),
.B(n_2347),
.Y(n_2440)
);

AND2x4_ASAP7_75t_L g2441 ( 
.A(n_2402),
.B(n_2338),
.Y(n_2441)
);

AND2x2_ASAP7_75t_L g2442 ( 
.A(n_2401),
.B(n_2344),
.Y(n_2442)
);

AND2x4_ASAP7_75t_L g2443 ( 
.A(n_2403),
.B(n_2338),
.Y(n_2443)
);

INVx2_ASAP7_75t_L g2444 ( 
.A(n_2403),
.Y(n_2444)
);

INVx1_ASAP7_75t_L g2445 ( 
.A(n_2410),
.Y(n_2445)
);

INVx1_ASAP7_75t_L g2446 ( 
.A(n_2410),
.Y(n_2446)
);

AND2x2_ASAP7_75t_L g2447 ( 
.A(n_2413),
.B(n_2344),
.Y(n_2447)
);

INVx1_ASAP7_75t_L g2448 ( 
.A(n_2413),
.Y(n_2448)
);

AND2x2_ASAP7_75t_L g2449 ( 
.A(n_2444),
.B(n_2415),
.Y(n_2449)
);

INVx2_ASAP7_75t_SL g2450 ( 
.A(n_2421),
.Y(n_2450)
);

INVx1_ASAP7_75t_L g2451 ( 
.A(n_2444),
.Y(n_2451)
);

AND2x4_ASAP7_75t_SL g2452 ( 
.A(n_2431),
.B(n_2400),
.Y(n_2452)
);

INVx1_ASAP7_75t_L g2453 ( 
.A(n_2444),
.Y(n_2453)
);

AND2x2_ASAP7_75t_L g2454 ( 
.A(n_2447),
.B(n_2415),
.Y(n_2454)
);

BUFx2_ASAP7_75t_L g2455 ( 
.A(n_2421),
.Y(n_2455)
);

HB1xp67_ASAP7_75t_L g2456 ( 
.A(n_2427),
.Y(n_2456)
);

INVx2_ASAP7_75t_L g2457 ( 
.A(n_2427),
.Y(n_2457)
);

INVxp67_ASAP7_75t_SL g2458 ( 
.A(n_2427),
.Y(n_2458)
);

AOI22xp5_ASAP7_75t_L g2459 ( 
.A1(n_2432),
.A2(n_2396),
.B1(n_2407),
.B2(n_2333),
.Y(n_2459)
);

HB1xp67_ASAP7_75t_L g2460 ( 
.A(n_2429),
.Y(n_2460)
);

INVx1_ASAP7_75t_L g2461 ( 
.A(n_2448),
.Y(n_2461)
);

NAND2xp5_ASAP7_75t_L g2462 ( 
.A(n_2445),
.B(n_2344),
.Y(n_2462)
);

NAND4xp25_ASAP7_75t_L g2463 ( 
.A(n_2433),
.B(n_2417),
.C(n_2405),
.D(n_2409),
.Y(n_2463)
);

CKINVDCx5p33_ASAP7_75t_R g2464 ( 
.A(n_2430),
.Y(n_2464)
);

INVx1_ASAP7_75t_SL g2465 ( 
.A(n_2426),
.Y(n_2465)
);

AND2x2_ASAP7_75t_L g2466 ( 
.A(n_2447),
.B(n_2445),
.Y(n_2466)
);

AND2x2_ASAP7_75t_L g2467 ( 
.A(n_2446),
.B(n_2345),
.Y(n_2467)
);

INVx2_ASAP7_75t_SL g2468 ( 
.A(n_2431),
.Y(n_2468)
);

AOI21xp33_ASAP7_75t_L g2469 ( 
.A1(n_2422),
.A2(n_2404),
.B(n_2386),
.Y(n_2469)
);

AOI22xp33_ASAP7_75t_L g2470 ( 
.A1(n_2443),
.A2(n_2391),
.B1(n_2398),
.B2(n_2348),
.Y(n_2470)
);

NAND2xp33_ASAP7_75t_L g2471 ( 
.A(n_2439),
.B(n_2411),
.Y(n_2471)
);

AND2x2_ASAP7_75t_L g2472 ( 
.A(n_2446),
.B(n_2338),
.Y(n_2472)
);

AOI211xp5_ASAP7_75t_L g2473 ( 
.A1(n_2439),
.A2(n_2411),
.B(n_2414),
.C(n_2373),
.Y(n_2473)
);

AND2x2_ASAP7_75t_L g2474 ( 
.A(n_2448),
.B(n_2338),
.Y(n_2474)
);

INVx1_ASAP7_75t_SL g2475 ( 
.A(n_2426),
.Y(n_2475)
);

HB1xp67_ASAP7_75t_L g2476 ( 
.A(n_2429),
.Y(n_2476)
);

INVx1_ASAP7_75t_L g2477 ( 
.A(n_2435),
.Y(n_2477)
);

HB1xp67_ASAP7_75t_L g2478 ( 
.A(n_2435),
.Y(n_2478)
);

INVx2_ASAP7_75t_L g2479 ( 
.A(n_2437),
.Y(n_2479)
);

AND2x2_ASAP7_75t_L g2480 ( 
.A(n_2455),
.B(n_2420),
.Y(n_2480)
);

AND2x2_ASAP7_75t_L g2481 ( 
.A(n_2455),
.B(n_2420),
.Y(n_2481)
);

AND2x2_ASAP7_75t_L g2482 ( 
.A(n_2450),
.B(n_2434),
.Y(n_2482)
);

NAND2xp5_ASAP7_75t_L g2483 ( 
.A(n_2461),
.B(n_2460),
.Y(n_2483)
);

AND2x4_ASAP7_75t_L g2484 ( 
.A(n_2450),
.B(n_2431),
.Y(n_2484)
);

AND2x2_ASAP7_75t_L g2485 ( 
.A(n_2450),
.B(n_2434),
.Y(n_2485)
);

HB1xp67_ASAP7_75t_L g2486 ( 
.A(n_2460),
.Y(n_2486)
);

INVx2_ASAP7_75t_L g2487 ( 
.A(n_2457),
.Y(n_2487)
);

INVx1_ASAP7_75t_L g2488 ( 
.A(n_2476),
.Y(n_2488)
);

AND2x2_ASAP7_75t_L g2489 ( 
.A(n_2454),
.B(n_2442),
.Y(n_2489)
);

INVx2_ASAP7_75t_L g2490 ( 
.A(n_2457),
.Y(n_2490)
);

INVx3_ASAP7_75t_L g2491 ( 
.A(n_2452),
.Y(n_2491)
);

NOR2x1_ASAP7_75t_L g2492 ( 
.A(n_2463),
.B(n_2431),
.Y(n_2492)
);

NOR2xp33_ASAP7_75t_L g2493 ( 
.A(n_2459),
.B(n_2438),
.Y(n_2493)
);

INVx3_ASAP7_75t_L g2494 ( 
.A(n_2452),
.Y(n_2494)
);

NAND2x1p5_ASAP7_75t_SL g2495 ( 
.A(n_2468),
.B(n_2463),
.Y(n_2495)
);

NAND2xp5_ASAP7_75t_L g2496 ( 
.A(n_2493),
.B(n_2470),
.Y(n_2496)
);

AND2x2_ASAP7_75t_L g2497 ( 
.A(n_2492),
.B(n_2466),
.Y(n_2497)
);

INVx2_ASAP7_75t_L g2498 ( 
.A(n_2487),
.Y(n_2498)
);

AND2x2_ASAP7_75t_L g2499 ( 
.A(n_2492),
.B(n_2466),
.Y(n_2499)
);

INVx2_ASAP7_75t_L g2500 ( 
.A(n_2487),
.Y(n_2500)
);

INVx2_ASAP7_75t_L g2501 ( 
.A(n_2487),
.Y(n_2501)
);

AND2x2_ASAP7_75t_L g2502 ( 
.A(n_2491),
.B(n_2494),
.Y(n_2502)
);

AND2x2_ASAP7_75t_L g2503 ( 
.A(n_2491),
.B(n_2454),
.Y(n_2503)
);

OAI21xp5_ASAP7_75t_L g2504 ( 
.A1(n_2493),
.A2(n_2459),
.B(n_2473),
.Y(n_2504)
);

NOR2x1_ASAP7_75t_L g2505 ( 
.A(n_2491),
.B(n_2471),
.Y(n_2505)
);

AND2x2_ASAP7_75t_L g2506 ( 
.A(n_2491),
.B(n_2468),
.Y(n_2506)
);

OR2x2_ASAP7_75t_L g2507 ( 
.A(n_2483),
.B(n_2461),
.Y(n_2507)
);

INVxp67_ASAP7_75t_L g2508 ( 
.A(n_2486),
.Y(n_2508)
);

INVx1_ASAP7_75t_L g2509 ( 
.A(n_2486),
.Y(n_2509)
);

NAND2xp5_ASAP7_75t_L g2510 ( 
.A(n_2489),
.B(n_2473),
.Y(n_2510)
);

NOR2xp33_ASAP7_75t_SL g2511 ( 
.A(n_2494),
.B(n_2416),
.Y(n_2511)
);

AND2x2_ASAP7_75t_L g2512 ( 
.A(n_2494),
.B(n_2468),
.Y(n_2512)
);

INVx1_ASAP7_75t_L g2513 ( 
.A(n_2483),
.Y(n_2513)
);

NAND2xp5_ASAP7_75t_L g2514 ( 
.A(n_2513),
.B(n_2488),
.Y(n_2514)
);

AOI21xp5_ASAP7_75t_L g2515 ( 
.A1(n_2504),
.A2(n_2494),
.B(n_2469),
.Y(n_2515)
);

OR2x2_ASAP7_75t_L g2516 ( 
.A(n_2507),
.B(n_2495),
.Y(n_2516)
);

NOR2x1_ASAP7_75t_L g2517 ( 
.A(n_2505),
.B(n_2484),
.Y(n_2517)
);

OR2x2_ASAP7_75t_L g2518 ( 
.A(n_2507),
.B(n_2495),
.Y(n_2518)
);

NAND2xp5_ASAP7_75t_L g2519 ( 
.A(n_2513),
.B(n_2488),
.Y(n_2519)
);

INVx1_ASAP7_75t_L g2520 ( 
.A(n_2509),
.Y(n_2520)
);

NOR2xp33_ASAP7_75t_L g2521 ( 
.A(n_2496),
.B(n_2464),
.Y(n_2521)
);

INVx1_ASAP7_75t_L g2522 ( 
.A(n_2509),
.Y(n_2522)
);

NAND2xp5_ASAP7_75t_L g2523 ( 
.A(n_2508),
.B(n_2495),
.Y(n_2523)
);

AND2x2_ASAP7_75t_L g2524 ( 
.A(n_2502),
.B(n_2480),
.Y(n_2524)
);

INVx1_ASAP7_75t_L g2525 ( 
.A(n_2502),
.Y(n_2525)
);

AND2x2_ASAP7_75t_SL g2526 ( 
.A(n_2511),
.B(n_2452),
.Y(n_2526)
);

AND2x2_ASAP7_75t_L g2527 ( 
.A(n_2503),
.B(n_2480),
.Y(n_2527)
);

INVx1_ASAP7_75t_L g2528 ( 
.A(n_2503),
.Y(n_2528)
);

AOI22xp5_ASAP7_75t_L g2529 ( 
.A1(n_2521),
.A2(n_2505),
.B1(n_2497),
.B2(n_2499),
.Y(n_2529)
);

OR2x2_ASAP7_75t_L g2530 ( 
.A(n_2528),
.B(n_2510),
.Y(n_2530)
);

INVxp67_ASAP7_75t_L g2531 ( 
.A(n_2523),
.Y(n_2531)
);

NAND2xp5_ASAP7_75t_L g2532 ( 
.A(n_2525),
.B(n_2497),
.Y(n_2532)
);

OR2x2_ASAP7_75t_L g2533 ( 
.A(n_2523),
.B(n_2499),
.Y(n_2533)
);

INVx1_ASAP7_75t_SL g2534 ( 
.A(n_2516),
.Y(n_2534)
);

OAI31xp33_ASAP7_75t_L g2535 ( 
.A1(n_2515),
.A2(n_2512),
.A3(n_2506),
.B(n_2469),
.Y(n_2535)
);

AOI22xp33_ASAP7_75t_L g2536 ( 
.A1(n_2526),
.A2(n_2518),
.B1(n_2517),
.B2(n_2524),
.Y(n_2536)
);

INVx1_ASAP7_75t_L g2537 ( 
.A(n_2514),
.Y(n_2537)
);

NAND2xp5_ASAP7_75t_L g2538 ( 
.A(n_2527),
.B(n_2506),
.Y(n_2538)
);

NOR2xp33_ASAP7_75t_L g2539 ( 
.A(n_2520),
.B(n_2512),
.Y(n_2539)
);

OAI21xp5_ASAP7_75t_L g2540 ( 
.A1(n_2522),
.A2(n_2484),
.B(n_2475),
.Y(n_2540)
);

NAND2xp5_ASAP7_75t_SL g2541 ( 
.A(n_2514),
.B(n_2484),
.Y(n_2541)
);

OAI322xp33_ASAP7_75t_L g2542 ( 
.A1(n_2519),
.A2(n_2465),
.A3(n_2475),
.B1(n_2500),
.B2(n_2498),
.C1(n_2501),
.C2(n_2481),
.Y(n_2542)
);

OAI22xp5_ASAP7_75t_L g2543 ( 
.A1(n_2536),
.A2(n_2519),
.B1(n_2484),
.B2(n_2465),
.Y(n_2543)
);

AOI222xp33_ASAP7_75t_L g2544 ( 
.A1(n_2531),
.A2(n_2534),
.B1(n_2537),
.B2(n_2541),
.C1(n_2532),
.C2(n_2540),
.Y(n_2544)
);

AOI221x1_ASAP7_75t_L g2545 ( 
.A1(n_2539),
.A2(n_2538),
.B1(n_2531),
.B2(n_2535),
.C(n_2529),
.Y(n_2545)
);

AOI32xp33_ASAP7_75t_L g2546 ( 
.A1(n_2533),
.A2(n_2481),
.A3(n_2482),
.B1(n_2485),
.B2(n_2501),
.Y(n_2546)
);

AOI22xp5_ASAP7_75t_L g2547 ( 
.A1(n_2530),
.A2(n_2482),
.B1(n_2485),
.B2(n_2498),
.Y(n_2547)
);

AND2x2_ASAP7_75t_L g2548 ( 
.A(n_2542),
.B(n_2489),
.Y(n_2548)
);

NAND2xp5_ASAP7_75t_L g2549 ( 
.A(n_2534),
.B(n_2500),
.Y(n_2549)
);

INVx1_ASAP7_75t_SL g2550 ( 
.A(n_2534),
.Y(n_2550)
);

INVx2_ASAP7_75t_L g2551 ( 
.A(n_2534),
.Y(n_2551)
);

AOI22xp5_ASAP7_75t_L g2552 ( 
.A1(n_2534),
.A2(n_2436),
.B1(n_2285),
.B2(n_2490),
.Y(n_2552)
);

INVxp67_ASAP7_75t_L g2553 ( 
.A(n_2534),
.Y(n_2553)
);

INVx1_ASAP7_75t_SL g2554 ( 
.A(n_2534),
.Y(n_2554)
);

NAND3xp33_ASAP7_75t_SL g2555 ( 
.A(n_2534),
.B(n_2436),
.C(n_2367),
.Y(n_2555)
);

AOI21xp5_ASAP7_75t_L g2556 ( 
.A1(n_2534),
.A2(n_2490),
.B(n_2476),
.Y(n_2556)
);

OR2x2_ASAP7_75t_L g2557 ( 
.A(n_2534),
.B(n_2462),
.Y(n_2557)
);

INVx2_ASAP7_75t_SL g2558 ( 
.A(n_2551),
.Y(n_2558)
);

NOR2xp33_ASAP7_75t_L g2559 ( 
.A(n_2550),
.B(n_2490),
.Y(n_2559)
);

INVx2_ASAP7_75t_L g2560 ( 
.A(n_2554),
.Y(n_2560)
);

OAI21xp33_ASAP7_75t_SL g2561 ( 
.A1(n_2544),
.A2(n_2458),
.B(n_2467),
.Y(n_2561)
);

OAI22xp33_ASAP7_75t_L g2562 ( 
.A1(n_2552),
.A2(n_2478),
.B1(n_2453),
.B2(n_2451),
.Y(n_2562)
);

OAI21xp33_ASAP7_75t_L g2563 ( 
.A1(n_2553),
.A2(n_2367),
.B(n_2462),
.Y(n_2563)
);

OAI21xp33_ASAP7_75t_L g2564 ( 
.A1(n_2543),
.A2(n_2549),
.B(n_2548),
.Y(n_2564)
);

INVx1_ASAP7_75t_L g2565 ( 
.A(n_2557),
.Y(n_2565)
);

BUFx3_ASAP7_75t_L g2566 ( 
.A(n_2547),
.Y(n_2566)
);

AOI22xp5_ASAP7_75t_L g2567 ( 
.A1(n_2555),
.A2(n_2474),
.B1(n_2467),
.B2(n_2472),
.Y(n_2567)
);

NOR3xp33_ASAP7_75t_L g2568 ( 
.A(n_2556),
.B(n_2380),
.C(n_2292),
.Y(n_2568)
);

INVx2_ASAP7_75t_L g2569 ( 
.A(n_2546),
.Y(n_2569)
);

AOI22xp5_ASAP7_75t_L g2570 ( 
.A1(n_2545),
.A2(n_2474),
.B1(n_2472),
.B2(n_2443),
.Y(n_2570)
);

XNOR2xp5_ASAP7_75t_L g2571 ( 
.A(n_2550),
.B(n_2380),
.Y(n_2571)
);

AND2x2_ASAP7_75t_SL g2572 ( 
.A(n_2560),
.B(n_2478),
.Y(n_2572)
);

NOR3xp33_ASAP7_75t_L g2573 ( 
.A(n_2558),
.B(n_2325),
.C(n_2352),
.Y(n_2573)
);

AOI21xp5_ASAP7_75t_L g2574 ( 
.A1(n_2564),
.A2(n_2458),
.B(n_2352),
.Y(n_2574)
);

NAND2xp5_ASAP7_75t_SL g2575 ( 
.A(n_2569),
.B(n_2561),
.Y(n_2575)
);

HB1xp67_ASAP7_75t_L g2576 ( 
.A(n_2559),
.Y(n_2576)
);

NAND4xp75_ASAP7_75t_L g2577 ( 
.A(n_2565),
.B(n_2386),
.C(n_2451),
.D(n_2453),
.Y(n_2577)
);

INVx1_ASAP7_75t_L g2578 ( 
.A(n_2565),
.Y(n_2578)
);

INVx1_ASAP7_75t_L g2579 ( 
.A(n_2566),
.Y(n_2579)
);

NOR2x1_ASAP7_75t_L g2580 ( 
.A(n_2571),
.B(n_2477),
.Y(n_2580)
);

NAND2xp5_ASAP7_75t_L g2581 ( 
.A(n_2563),
.B(n_2456),
.Y(n_2581)
);

OAI22xp33_ASAP7_75t_L g2582 ( 
.A1(n_2570),
.A2(n_2456),
.B1(n_2288),
.B2(n_2477),
.Y(n_2582)
);

NOR3xp33_ASAP7_75t_L g2583 ( 
.A(n_2568),
.B(n_2383),
.C(n_2382),
.Y(n_2583)
);

NAND2xp5_ASAP7_75t_L g2584 ( 
.A(n_2579),
.B(n_2562),
.Y(n_2584)
);

AOI22xp5_ASAP7_75t_L g2585 ( 
.A1(n_2573),
.A2(n_2567),
.B1(n_2288),
.B2(n_2383),
.Y(n_2585)
);

O2A1O1Ixp33_ASAP7_75t_L g2586 ( 
.A1(n_2575),
.A2(n_2578),
.B(n_2576),
.C(n_2581),
.Y(n_2586)
);

AOI221xp5_ASAP7_75t_L g2587 ( 
.A1(n_2574),
.A2(n_2357),
.B1(n_2342),
.B2(n_2343),
.C(n_2479),
.Y(n_2587)
);

OAI22xp5_ASAP7_75t_L g2588 ( 
.A1(n_2580),
.A2(n_2457),
.B1(n_2479),
.B2(n_2288),
.Y(n_2588)
);

NAND4xp25_ASAP7_75t_SL g2589 ( 
.A(n_2583),
.B(n_2449),
.C(n_2442),
.D(n_2440),
.Y(n_2589)
);

INVxp67_ASAP7_75t_L g2590 ( 
.A(n_2572),
.Y(n_2590)
);

AOI211x1_ASAP7_75t_SL g2591 ( 
.A1(n_2582),
.A2(n_2479),
.B(n_2384),
.C(n_2359),
.Y(n_2591)
);

AOI211xp5_ASAP7_75t_L g2592 ( 
.A1(n_2577),
.A2(n_2382),
.B(n_2443),
.C(n_2357),
.Y(n_2592)
);

OAI21xp33_ASAP7_75t_L g2593 ( 
.A1(n_2579),
.A2(n_2449),
.B(n_2375),
.Y(n_2593)
);

AOI322xp5_ASAP7_75t_L g2594 ( 
.A1(n_2584),
.A2(n_2443),
.A3(n_2440),
.B1(n_2441),
.B2(n_2400),
.C1(n_2348),
.C2(n_2390),
.Y(n_2594)
);

AOI221xp5_ASAP7_75t_L g2595 ( 
.A1(n_2586),
.A2(n_2343),
.B1(n_2346),
.B2(n_2428),
.C(n_2425),
.Y(n_2595)
);

AOI221x1_ASAP7_75t_SL g2596 ( 
.A1(n_2592),
.A2(n_2590),
.B1(n_2593),
.B2(n_2588),
.C(n_2591),
.Y(n_2596)
);

INVxp67_ASAP7_75t_SL g2597 ( 
.A(n_2585),
.Y(n_2597)
);

OAI211xp5_ASAP7_75t_SL g2598 ( 
.A1(n_2587),
.A2(n_2379),
.B(n_2213),
.C(n_2348),
.Y(n_2598)
);

INVxp33_ASAP7_75t_SL g2599 ( 
.A(n_2589),
.Y(n_2599)
);

OR2x2_ASAP7_75t_L g2600 ( 
.A(n_2584),
.B(n_2423),
.Y(n_2600)
);

OAI211xp5_ASAP7_75t_SL g2601 ( 
.A1(n_2586),
.A2(n_2379),
.B(n_2348),
.C(n_2362),
.Y(n_2601)
);

AOI221xp5_ASAP7_75t_L g2602 ( 
.A1(n_2586),
.A2(n_2346),
.B1(n_2424),
.B2(n_2428),
.C(n_2425),
.Y(n_2602)
);

AND2x2_ASAP7_75t_L g2603 ( 
.A(n_2585),
.B(n_2390),
.Y(n_2603)
);

AOI221xp5_ASAP7_75t_L g2604 ( 
.A1(n_2586),
.A2(n_2424),
.B1(n_2359),
.B2(n_2362),
.C(n_2361),
.Y(n_2604)
);

AND4x2_ASAP7_75t_L g2605 ( 
.A(n_2586),
.B(n_2390),
.C(n_2318),
.D(n_2392),
.Y(n_2605)
);

OAI21xp5_ASAP7_75t_L g2606 ( 
.A1(n_2597),
.A2(n_2382),
.B(n_2224),
.Y(n_2606)
);

INVx2_ASAP7_75t_L g2607 ( 
.A(n_2600),
.Y(n_2607)
);

OR2x2_ASAP7_75t_L g2608 ( 
.A(n_2603),
.B(n_2423),
.Y(n_2608)
);

AND3x4_ASAP7_75t_L g2609 ( 
.A(n_2599),
.B(n_2400),
.C(n_2441),
.Y(n_2609)
);

NOR3xp33_ASAP7_75t_L g2610 ( 
.A(n_2601),
.B(n_2339),
.C(n_2379),
.Y(n_2610)
);

INVx1_ASAP7_75t_SL g2611 ( 
.A(n_2596),
.Y(n_2611)
);

HB1xp67_ASAP7_75t_L g2612 ( 
.A(n_2602),
.Y(n_2612)
);

XNOR2xp5_ASAP7_75t_L g2613 ( 
.A(n_2595),
.B(n_2360),
.Y(n_2613)
);

INVx1_ASAP7_75t_L g2614 ( 
.A(n_2598),
.Y(n_2614)
);

XOR2xp5_ASAP7_75t_L g2615 ( 
.A(n_2605),
.B(n_2377),
.Y(n_2615)
);

INVx1_ASAP7_75t_L g2616 ( 
.A(n_2604),
.Y(n_2616)
);

AOI22xp5_ASAP7_75t_L g2617 ( 
.A1(n_2594),
.A2(n_2379),
.B1(n_2359),
.B2(n_2324),
.Y(n_2617)
);

INVx2_ASAP7_75t_L g2618 ( 
.A(n_2600),
.Y(n_2618)
);

AOI22xp5_ASAP7_75t_L g2619 ( 
.A1(n_2611),
.A2(n_2379),
.B1(n_2384),
.B2(n_2441),
.Y(n_2619)
);

NOR3xp33_ASAP7_75t_L g2620 ( 
.A(n_2607),
.B(n_2354),
.C(n_2384),
.Y(n_2620)
);

OR2x2_ASAP7_75t_L g2621 ( 
.A(n_2618),
.B(n_2381),
.Y(n_2621)
);

OAI221xp5_ASAP7_75t_SL g2622 ( 
.A1(n_2614),
.A2(n_2390),
.B1(n_2348),
.B2(n_2437),
.C(n_2378),
.Y(n_2622)
);

NAND2xp5_ASAP7_75t_L g2623 ( 
.A(n_2615),
.B(n_2381),
.Y(n_2623)
);

AND2x2_ASAP7_75t_L g2624 ( 
.A(n_2612),
.B(n_2608),
.Y(n_2624)
);

NAND3xp33_ASAP7_75t_L g2625 ( 
.A(n_2616),
.B(n_2005),
.C(n_2008),
.Y(n_2625)
);

NAND3xp33_ASAP7_75t_SL g2626 ( 
.A(n_2616),
.B(n_2353),
.C(n_2376),
.Y(n_2626)
);

OAI322xp33_ASAP7_75t_L g2627 ( 
.A1(n_2613),
.A2(n_2378),
.A3(n_2376),
.B1(n_2381),
.B2(n_2355),
.C1(n_2356),
.C2(n_2353),
.Y(n_2627)
);

AOI22xp5_ASAP7_75t_L g2628 ( 
.A1(n_2609),
.A2(n_2441),
.B1(n_2363),
.B2(n_2364),
.Y(n_2628)
);

NAND3xp33_ASAP7_75t_L g2629 ( 
.A(n_2610),
.B(n_2005),
.C(n_2008),
.Y(n_2629)
);

OR2x2_ASAP7_75t_L g2630 ( 
.A(n_2625),
.B(n_2617),
.Y(n_2630)
);

AO22x2_ASAP7_75t_L g2631 ( 
.A1(n_2624),
.A2(n_2606),
.B1(n_2356),
.B2(n_2355),
.Y(n_2631)
);

INVx3_ASAP7_75t_L g2632 ( 
.A(n_2621),
.Y(n_2632)
);

AND2x4_ASAP7_75t_L g2633 ( 
.A(n_2620),
.B(n_2377),
.Y(n_2633)
);

OAI21xp5_ASAP7_75t_L g2634 ( 
.A1(n_2619),
.A2(n_2360),
.B(n_2372),
.Y(n_2634)
);

OAI22xp5_ASAP7_75t_SL g2635 ( 
.A1(n_2623),
.A2(n_2353),
.B1(n_2334),
.B2(n_2354),
.Y(n_2635)
);

AND2x2_ASAP7_75t_L g2636 ( 
.A(n_2628),
.B(n_2394),
.Y(n_2636)
);

INVx1_ASAP7_75t_L g2637 ( 
.A(n_2626),
.Y(n_2637)
);

INVx2_ASAP7_75t_L g2638 ( 
.A(n_2630),
.Y(n_2638)
);

AOI22xp5_ASAP7_75t_L g2639 ( 
.A1(n_2632),
.A2(n_2629),
.B1(n_2627),
.B2(n_2622),
.Y(n_2639)
);

AOI22xp5_ASAP7_75t_L g2640 ( 
.A1(n_2637),
.A2(n_2635),
.B1(n_2633),
.B2(n_2636),
.Y(n_2640)
);

AO22x2_ASAP7_75t_L g2641 ( 
.A1(n_2636),
.A2(n_2354),
.B1(n_2363),
.B2(n_2364),
.Y(n_2641)
);

AO22x2_ASAP7_75t_L g2642 ( 
.A1(n_2631),
.A2(n_2354),
.B1(n_2392),
.B2(n_2394),
.Y(n_2642)
);

AOI22xp5_ASAP7_75t_L g2643 ( 
.A1(n_2634),
.A2(n_2354),
.B1(n_2336),
.B2(n_2334),
.Y(n_2643)
);

HB1xp67_ASAP7_75t_L g2644 ( 
.A(n_2638),
.Y(n_2644)
);

OAI22xp5_ASAP7_75t_SL g2645 ( 
.A1(n_2640),
.A2(n_2353),
.B1(n_2334),
.B2(n_2026),
.Y(n_2645)
);

NOR2x1p5_ASAP7_75t_L g2646 ( 
.A(n_2639),
.B(n_2334),
.Y(n_2646)
);

OAI22xp5_ASAP7_75t_L g2647 ( 
.A1(n_2641),
.A2(n_2334),
.B1(n_2175),
.B2(n_2337),
.Y(n_2647)
);

AO22x2_ASAP7_75t_L g2648 ( 
.A1(n_2647),
.A2(n_2643),
.B1(n_2642),
.B2(n_2366),
.Y(n_2648)
);

HB1xp67_ASAP7_75t_L g2649 ( 
.A(n_2644),
.Y(n_2649)
);

AOI22xp5_ASAP7_75t_SL g2650 ( 
.A1(n_2649),
.A2(n_2646),
.B1(n_2645),
.B2(n_2334),
.Y(n_2650)
);

AOI22xp33_ASAP7_75t_L g2651 ( 
.A1(n_2650),
.A2(n_2648),
.B1(n_2334),
.B2(n_2336),
.Y(n_2651)
);

OAI21xp5_ASAP7_75t_SL g2652 ( 
.A1(n_2651),
.A2(n_2008),
.B(n_2009),
.Y(n_2652)
);

OAI21xp5_ASAP7_75t_L g2653 ( 
.A1(n_2651),
.A2(n_2372),
.B(n_2207),
.Y(n_2653)
);

XNOR2xp5_ASAP7_75t_L g2654 ( 
.A(n_2653),
.B(n_2335),
.Y(n_2654)
);

HB1xp67_ASAP7_75t_L g2655 ( 
.A(n_2652),
.Y(n_2655)
);

AOI221xp5_ASAP7_75t_L g2656 ( 
.A1(n_2655),
.A2(n_2351),
.B1(n_2349),
.B2(n_2350),
.C(n_2340),
.Y(n_2656)
);

AOI211xp5_ASAP7_75t_L g2657 ( 
.A1(n_2656),
.A2(n_2654),
.B(n_2340),
.C(n_2337),
.Y(n_2657)
);


endmodule