module fake_jpeg_2584_n_700 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_700);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_700;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_696;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_686;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_678;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_699;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_672;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_688;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_689;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_698;
wire n_195;
wire n_450;
wire n_557;
wire n_681;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_694;
wire n_692;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_668;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_682;
wire n_305;
wire n_161;
wire n_441;
wire n_697;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_679;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_691;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_615;
wire n_598;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_676;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_670;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_683;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_690;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_693;
wire n_674;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_684;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_680;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_695;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_687;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_673;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_665;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_677;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_671;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_669;
wire n_524;
wire n_402;
wire n_563;
wire n_685;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_675;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx4_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_17),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_14),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_0),
.Y(n_31)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_16),
.Y(n_33)
);

BUFx16f_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

BUFx10_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_16),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_15),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_19),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_10),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

CKINVDCx14_ASAP7_75t_R g44 ( 
.A(n_18),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_8),
.Y(n_45)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_10),
.Y(n_46)
);

INVx13_ASAP7_75t_L g47 ( 
.A(n_13),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_1),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_17),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_7),
.Y(n_51)
);

BUFx16f_ASAP7_75t_L g52 ( 
.A(n_14),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_13),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_0),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_3),
.Y(n_55)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_3),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_13),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_14),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_52),
.Y(n_59)
);

INVx1_ASAP7_75t_SL g193 ( 
.A(n_59),
.Y(n_193)
);

INVx2_ASAP7_75t_SL g60 ( 
.A(n_34),
.Y(n_60)
);

INVx2_ASAP7_75t_SL g137 ( 
.A(n_60),
.Y(n_137)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_52),
.Y(n_61)
);

INVx4_ASAP7_75t_SL g230 ( 
.A(n_61),
.Y(n_230)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_52),
.Y(n_62)
);

INVx2_ASAP7_75t_SL g231 ( 
.A(n_62),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_44),
.B(n_19),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_63),
.B(n_80),
.Y(n_177)
);

OR2x2_ASAP7_75t_L g64 ( 
.A(n_20),
.B(n_19),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_64),
.B(n_87),
.Y(n_144)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_57),
.Y(n_65)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_65),
.Y(n_135)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_66),
.Y(n_136)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_34),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g149 ( 
.A(n_67),
.Y(n_149)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_68),
.Y(n_171)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_69),
.Y(n_151)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_20),
.Y(n_70)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_70),
.Y(n_143)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_71),
.Y(n_154)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_57),
.Y(n_72)
);

INVx5_ASAP7_75t_L g142 ( 
.A(n_72),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_24),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_73),
.Y(n_145)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_20),
.Y(n_74)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_74),
.Y(n_155)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_34),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g168 ( 
.A(n_75),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_24),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_76),
.Y(n_158)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_20),
.Y(n_77)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_77),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_24),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_78),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_34),
.A2(n_19),
.B1(n_18),
.B2(n_17),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_79),
.A2(n_100),
.B1(n_132),
.B2(n_31),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_44),
.B(n_18),
.Y(n_80)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_24),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_81),
.Y(n_186)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_57),
.Y(n_82)
);

INVx5_ASAP7_75t_L g152 ( 
.A(n_82),
.Y(n_152)
);

BUFx12_ASAP7_75t_L g83 ( 
.A(n_52),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g213 ( 
.A(n_83),
.Y(n_213)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_43),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_84),
.Y(n_188)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_34),
.Y(n_85)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_85),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_43),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_86),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_21),
.B(n_18),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_56),
.Y(n_88)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_88),
.Y(n_161)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_57),
.Y(n_89)
);

INVx5_ASAP7_75t_L g198 ( 
.A(n_89),
.Y(n_198)
);

BUFx12f_ASAP7_75t_L g90 ( 
.A(n_52),
.Y(n_90)
);

INVx8_ASAP7_75t_L g166 ( 
.A(n_90),
.Y(n_166)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_57),
.Y(n_91)
);

INVx5_ASAP7_75t_L g210 ( 
.A(n_91),
.Y(n_210)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_57),
.Y(n_92)
);

INVx3_ASAP7_75t_SL g187 ( 
.A(n_92),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_21),
.B(n_17),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_93),
.B(n_108),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_43),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_94),
.Y(n_200)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_57),
.Y(n_95)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_95),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_43),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_96),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_53),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_97),
.Y(n_217)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_22),
.Y(n_98)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_98),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_53),
.Y(n_99)
);

INVx6_ASAP7_75t_L g159 ( 
.A(n_99),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_53),
.A2(n_16),
.B1(n_12),
.B2(n_2),
.Y(n_100)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_53),
.Y(n_101)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_101),
.Y(n_164)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_26),
.Y(n_102)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_102),
.Y(n_146)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_22),
.Y(n_103)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_103),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_22),
.Y(n_104)
);

INVx6_ASAP7_75t_L g182 ( 
.A(n_104),
.Y(n_182)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_56),
.Y(n_105)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_105),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_22),
.Y(n_106)
);

INVx6_ASAP7_75t_L g195 ( 
.A(n_106),
.Y(n_195)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_27),
.Y(n_107)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_107),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_23),
.B(n_12),
.Y(n_108)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_27),
.Y(n_109)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_109),
.Y(n_190)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_27),
.Y(n_110)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_110),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_27),
.Y(n_111)
);

INVx6_ASAP7_75t_L g206 ( 
.A(n_111),
.Y(n_206)
);

INVx11_ASAP7_75t_L g112 ( 
.A(n_47),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_112),
.Y(n_169)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_56),
.Y(n_113)
);

HB1xp67_ASAP7_75t_L g141 ( 
.A(n_113),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_21),
.B(n_0),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_114),
.B(n_116),
.Y(n_232)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_56),
.Y(n_115)
);

HB1xp67_ASAP7_75t_L g162 ( 
.A(n_115),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_25),
.B(n_0),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_25),
.B(n_33),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_117),
.B(n_118),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_25),
.B(n_11),
.Y(n_118)
);

BUFx12f_ASAP7_75t_L g119 ( 
.A(n_39),
.Y(n_119)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_119),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_39),
.Y(n_120)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_120),
.Y(n_175)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_39),
.Y(n_121)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_121),
.Y(n_180)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_39),
.Y(n_122)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_122),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_48),
.B(n_0),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_123),
.B(n_31),
.Y(n_148)
);

INVx5_ASAP7_75t_L g124 ( 
.A(n_48),
.Y(n_124)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_124),
.Y(n_216)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_26),
.Y(n_125)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_125),
.Y(n_222)
);

INVx11_ASAP7_75t_L g126 ( 
.A(n_47),
.Y(n_126)
);

INVxp67_ASAP7_75t_SL g209 ( 
.A(n_126),
.Y(n_209)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_48),
.Y(n_127)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_127),
.Y(n_185)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_26),
.Y(n_128)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_128),
.Y(n_229)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_29),
.Y(n_129)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_129),
.Y(n_179)
);

INVx13_ASAP7_75t_L g130 ( 
.A(n_47),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_130),
.Y(n_203)
);

INVx6_ASAP7_75t_L g131 ( 
.A(n_48),
.Y(n_131)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_131),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_33),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_29),
.Y(n_133)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_133),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_134),
.A2(n_183),
.B1(n_192),
.B2(n_199),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_60),
.A2(n_32),
.B1(n_40),
.B2(n_28),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_147),
.A2(n_150),
.B1(n_173),
.B2(n_178),
.Y(n_260)
);

AND2x2_ASAP7_75t_L g258 ( 
.A(n_148),
.B(n_1),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_102),
.A2(n_32),
.B1(n_40),
.B2(n_28),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_123),
.B(n_37),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_157),
.B(n_172),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_67),
.B(n_37),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_125),
.A2(n_32),
.B1(n_40),
.B2(n_28),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_64),
.B(n_37),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_174),
.B(n_176),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_59),
.B(n_41),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_128),
.A2(n_32),
.B1(n_40),
.B2(n_28),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_81),
.A2(n_33),
.B1(n_38),
.B2(n_41),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_133),
.Y(n_184)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_184),
.Y(n_245)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_98),
.Y(n_189)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_189),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_84),
.A2(n_38),
.B1(n_41),
.B2(n_50),
.Y(n_192)
);

OR2x2_ASAP7_75t_L g197 ( 
.A(n_130),
.B(n_29),
.Y(n_197)
);

NAND3xp33_ASAP7_75t_L g269 ( 
.A(n_197),
.B(n_221),
.C(n_2),
.Y(n_269)
);

OAI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_104),
.A2(n_31),
.B1(n_55),
.B2(n_23),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_59),
.B(n_38),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g298 ( 
.A(n_201),
.B(n_202),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_61),
.B(n_50),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_61),
.A2(n_90),
.B1(n_112),
.B2(n_126),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_205),
.A2(n_224),
.B1(n_228),
.B2(n_36),
.Y(n_278)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_107),
.Y(n_207)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_207),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_90),
.B(n_50),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_211),
.B(n_220),
.Y(n_237)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_131),
.Y(n_212)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_212),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_103),
.B(n_23),
.Y(n_214)
);

OR2x2_ASAP7_75t_L g293 ( 
.A(n_214),
.B(n_219),
.Y(n_293)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_65),
.Y(n_215)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_215),
.Y(n_264)
);

OAI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_106),
.A2(n_55),
.B1(n_42),
.B2(n_45),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_218),
.A2(n_30),
.B1(n_51),
.B2(n_54),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_73),
.A2(n_49),
.B1(n_55),
.B2(n_42),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_119),
.B(n_49),
.Y(n_220)
);

AND2x2_ASAP7_75t_L g221 ( 
.A(n_119),
.B(n_45),
.Y(n_221)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_101),
.Y(n_223)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_223),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_L g224 ( 
.A1(n_111),
.A2(n_45),
.B1(n_42),
.B2(n_49),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_72),
.B(n_54),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_225),
.B(n_233),
.Y(n_250)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_120),
.Y(n_227)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_227),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_82),
.A2(n_54),
.B1(n_51),
.B2(n_30),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_89),
.B(n_95),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_91),
.Y(n_234)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_234),
.Y(n_274)
);

INVx4_ASAP7_75t_L g236 ( 
.A(n_231),
.Y(n_236)
);

INVx4_ASAP7_75t_L g361 ( 
.A(n_236),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_232),
.B(n_92),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_238),
.B(n_268),
.Y(n_351)
);

AOI22xp33_ASAP7_75t_L g240 ( 
.A1(n_199),
.A2(n_99),
.B1(n_97),
.B2(n_96),
.Y(n_240)
);

OAI22xp33_ASAP7_75t_SL g324 ( 
.A1(n_240),
.A2(n_170),
.B1(n_204),
.B2(n_200),
.Y(n_324)
);

INVx6_ASAP7_75t_L g242 ( 
.A(n_145),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g326 ( 
.A(n_242),
.Y(n_326)
);

INVx6_ASAP7_75t_L g244 ( 
.A(n_145),
.Y(n_244)
);

INVx3_ASAP7_75t_L g332 ( 
.A(n_244),
.Y(n_332)
);

INVx3_ASAP7_75t_L g246 ( 
.A(n_193),
.Y(n_246)
);

INVxp67_ASAP7_75t_SL g385 ( 
.A(n_246),
.Y(n_385)
);

INVx3_ASAP7_75t_L g249 ( 
.A(n_193),
.Y(n_249)
);

INVx3_ASAP7_75t_L g364 ( 
.A(n_249),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_251),
.A2(n_261),
.B1(n_284),
.B2(n_286),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_218),
.A2(n_94),
.B1(n_86),
.B2(n_78),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g352 ( 
.A1(n_252),
.A2(n_282),
.B1(n_288),
.B2(n_320),
.Y(n_352)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_194),
.Y(n_254)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_254),
.Y(n_323)
);

INVx4_ASAP7_75t_L g255 ( 
.A(n_231),
.Y(n_255)
);

INVx3_ASAP7_75t_L g381 ( 
.A(n_255),
.Y(n_381)
);

AOI22xp33_ASAP7_75t_SL g256 ( 
.A1(n_221),
.A2(n_51),
.B1(n_30),
.B2(n_47),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g329 ( 
.A(n_256),
.Y(n_329)
);

INVx5_ASAP7_75t_L g257 ( 
.A(n_166),
.Y(n_257)
);

BUFx3_ASAP7_75t_L g341 ( 
.A(n_257),
.Y(n_341)
);

AND2x2_ASAP7_75t_L g343 ( 
.A(n_258),
.B(n_269),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_140),
.B(n_1),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_259),
.B(n_265),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_224),
.A2(n_76),
.B1(n_79),
.B2(n_36),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_164),
.Y(n_262)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_262),
.Y(n_331)
);

INVx5_ASAP7_75t_L g263 ( 
.A(n_166),
.Y(n_263)
);

INVx1_ASAP7_75t_SL g360 ( 
.A(n_263),
.Y(n_360)
);

CKINVDCx16_ASAP7_75t_R g265 ( 
.A(n_197),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_161),
.Y(n_266)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_266),
.Y(n_346)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_165),
.Y(n_267)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_267),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_226),
.B(n_1),
.Y(n_268)
);

INVx4_ASAP7_75t_L g270 ( 
.A(n_137),
.Y(n_270)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_270),
.Y(n_363)
);

AOI22xp33_ASAP7_75t_SL g271 ( 
.A1(n_144),
.A2(n_26),
.B1(n_36),
.B2(n_35),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g340 ( 
.A(n_271),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_177),
.B(n_2),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_272),
.B(n_285),
.Y(n_365)
);

INVx3_ASAP7_75t_L g273 ( 
.A(n_135),
.Y(n_273)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_273),
.Y(n_369)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_180),
.Y(n_275)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_275),
.Y(n_327)
);

AOI22xp33_ASAP7_75t_SL g276 ( 
.A1(n_196),
.A2(n_36),
.B1(n_35),
.B2(n_58),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_SL g325 ( 
.A1(n_276),
.A2(n_278),
.B1(n_300),
.B2(n_317),
.Y(n_325)
);

INVx3_ASAP7_75t_L g279 ( 
.A(n_135),
.Y(n_279)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_279),
.Y(n_330)
);

AND2x2_ASAP7_75t_L g280 ( 
.A(n_137),
.B(n_2),
.Y(n_280)
);

AND2x2_ASAP7_75t_L g354 ( 
.A(n_280),
.B(n_283),
.Y(n_354)
);

A2O1A1Ixp33_ASAP7_75t_L g281 ( 
.A1(n_203),
.A2(n_83),
.B(n_36),
.C(n_35),
.Y(n_281)
);

AOI31xp33_ASAP7_75t_L g336 ( 
.A1(n_281),
.A2(n_213),
.A3(n_168),
.B(n_187),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_175),
.A2(n_36),
.B1(n_83),
.B2(n_58),
.Y(n_282)
);

AND2x2_ASAP7_75t_L g283 ( 
.A(n_179),
.B(n_3),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_228),
.A2(n_36),
.B1(n_58),
.B2(n_6),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_143),
.B(n_4),
.Y(n_285)
);

OAI22xp33_ASAP7_75t_L g286 ( 
.A1(n_150),
.A2(n_58),
.B1(n_5),
.B2(n_6),
.Y(n_286)
);

INVx5_ASAP7_75t_L g287 ( 
.A(n_149),
.Y(n_287)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_287),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_173),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_181),
.Y(n_289)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_289),
.Y(n_337)
);

INVxp67_ASAP7_75t_L g290 ( 
.A(n_209),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_290),
.B(n_291),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_155),
.B(n_4),
.Y(n_291)
);

INVx3_ASAP7_75t_L g292 ( 
.A(n_142),
.Y(n_292)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_292),
.Y(n_342)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_167),
.Y(n_294)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_294),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_136),
.B(n_4),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_295),
.B(n_297),
.Y(n_374)
);

INVx2_ASAP7_75t_SL g296 ( 
.A(n_149),
.Y(n_296)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_296),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_151),
.B(n_5),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_208),
.B(n_5),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_299),
.B(n_304),
.Y(n_375)
);

AOI22xp33_ASAP7_75t_SL g300 ( 
.A1(n_146),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_185),
.Y(n_301)
);

AND2x2_ASAP7_75t_L g358 ( 
.A(n_301),
.B(n_303),
.Y(n_358)
);

BUFx2_ASAP7_75t_L g302 ( 
.A(n_187),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_302),
.Y(n_376)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_141),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_154),
.B(n_7),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_205),
.A2(n_147),
.B(n_178),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g373 ( 
.A1(n_305),
.A2(n_310),
.B(n_163),
.Y(n_373)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_162),
.Y(n_306)
);

AND2x2_ASAP7_75t_L g362 ( 
.A(n_306),
.B(n_307),
.Y(n_362)
);

INVx3_ASAP7_75t_L g307 ( 
.A(n_142),
.Y(n_307)
);

INVx3_ASAP7_75t_L g308 ( 
.A(n_152),
.Y(n_308)
);

AND2x2_ASAP7_75t_L g380 ( 
.A(n_308),
.B(n_309),
.Y(n_380)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_175),
.Y(n_309)
);

O2A1O1Ixp33_ASAP7_75t_L g310 ( 
.A1(n_209),
.A2(n_7),
.B(n_8),
.C(n_9),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_171),
.B(n_7),
.Y(n_311)
);

AND2x2_ASAP7_75t_L g384 ( 
.A(n_311),
.B(n_313),
.Y(n_384)
);

INVxp67_ASAP7_75t_L g312 ( 
.A(n_146),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_312),
.Y(n_377)
);

CKINVDCx16_ASAP7_75t_R g313 ( 
.A(n_230),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_139),
.Y(n_314)
);

OR2x2_ASAP7_75t_L g370 ( 
.A(n_314),
.B(n_315),
.Y(n_370)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_139),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_222),
.B(n_9),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_316),
.B(n_169),
.Y(n_333)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_156),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_156),
.Y(n_318)
);

AOI22xp33_ASAP7_75t_SL g334 ( 
.A1(n_318),
.A2(n_321),
.B1(n_322),
.B2(n_230),
.Y(n_334)
);

OAI22xp33_ASAP7_75t_SL g319 ( 
.A1(n_186),
.A2(n_9),
.B1(n_11),
.B2(n_188),
.Y(n_319)
);

AOI22xp33_ASAP7_75t_L g359 ( 
.A1(n_319),
.A2(n_191),
.B1(n_204),
.B2(n_158),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_186),
.A2(n_9),
.B1(n_11),
.B2(n_188),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_159),
.Y(n_321)
);

INVx3_ASAP7_75t_L g322 ( 
.A(n_152),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_324),
.A2(n_338),
.B1(n_344),
.B2(n_356),
.Y(n_395)
);

NAND2x1p5_ASAP7_75t_L g328 ( 
.A(n_258),
.B(n_229),
.Y(n_328)
);

OAI21xp33_ASAP7_75t_L g390 ( 
.A1(n_328),
.A2(n_333),
.B(n_336),
.Y(n_390)
);

INVxp67_ASAP7_75t_L g411 ( 
.A(n_334),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_235),
.A2(n_206),
.B1(n_182),
.B2(n_195),
.Y(n_338)
);

OAI32xp33_ASAP7_75t_L g339 ( 
.A1(n_243),
.A2(n_229),
.A3(n_222),
.B1(n_153),
.B2(n_160),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_339),
.B(n_345),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_235),
.A2(n_182),
.B1(n_195),
.B2(n_206),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_283),
.B(n_138),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_283),
.B(n_138),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_349),
.B(n_355),
.Y(n_415)
);

INVx6_ASAP7_75t_L g353 ( 
.A(n_242),
.Y(n_353)
);

INVx4_ASAP7_75t_L g391 ( 
.A(n_353),
.Y(n_391)
);

OAI32xp33_ASAP7_75t_L g355 ( 
.A1(n_258),
.A2(n_153),
.A3(n_216),
.B1(n_160),
.B2(n_190),
.Y(n_355)
);

OAI22xp33_ASAP7_75t_L g356 ( 
.A1(n_252),
.A2(n_159),
.B1(n_217),
.B2(n_158),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_311),
.B(n_213),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_357),
.B(n_368),
.Y(n_429)
);

OAI22xp33_ASAP7_75t_SL g396 ( 
.A1(n_359),
.A2(n_366),
.B1(n_379),
.B2(n_282),
.Y(n_396)
);

AOI22xp33_ASAP7_75t_L g366 ( 
.A1(n_260),
.A2(n_216),
.B1(n_217),
.B2(n_191),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_250),
.B(n_210),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_237),
.B(n_210),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_372),
.B(n_257),
.Y(n_432)
);

INVx1_ASAP7_75t_SL g418 ( 
.A(n_373),
.Y(n_418)
);

INVx6_ASAP7_75t_L g378 ( 
.A(n_244),
.Y(n_378)
);

INVx4_ASAP7_75t_L g392 ( 
.A(n_378),
.Y(n_392)
);

AOI22xp33_ASAP7_75t_L g379 ( 
.A1(n_305),
.A2(n_170),
.B1(n_200),
.B2(n_190),
.Y(n_379)
);

OAI21xp5_ASAP7_75t_SL g382 ( 
.A1(n_293),
.A2(n_198),
.B(n_163),
.Y(n_382)
);

AOI21xp5_ASAP7_75t_SL g410 ( 
.A1(n_382),
.A2(n_290),
.B(n_302),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_L g386 ( 
.A1(n_293),
.A2(n_198),
.B1(n_168),
.B2(n_11),
.Y(n_386)
);

AO21x2_ASAP7_75t_L g420 ( 
.A1(n_386),
.A2(n_310),
.B(n_309),
.Y(n_420)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_380),
.Y(n_387)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_387),
.Y(n_471)
);

OAI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_367),
.A2(n_251),
.B1(n_261),
.B2(n_320),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_388),
.A2(n_426),
.B1(n_433),
.B2(n_437),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_377),
.B(n_277),
.Y(n_389)
);

OAI21xp33_ASAP7_75t_L g446 ( 
.A1(n_389),
.A2(n_402),
.B(n_432),
.Y(n_446)
);

HB1xp67_ASAP7_75t_L g393 ( 
.A(n_330),
.Y(n_393)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_393),
.Y(n_473)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_380),
.Y(n_394)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_394),
.Y(n_479)
);

AOI22xp5_ASAP7_75t_SL g469 ( 
.A1(n_396),
.A2(n_335),
.B1(n_376),
.B2(n_383),
.Y(n_469)
);

AOI21xp5_ASAP7_75t_L g397 ( 
.A1(n_373),
.A2(n_281),
.B(n_286),
.Y(n_397)
);

AOI21xp5_ASAP7_75t_L g458 ( 
.A1(n_397),
.A2(n_424),
.B(n_360),
.Y(n_458)
);

AOI22xp33_ASAP7_75t_SL g398 ( 
.A1(n_340),
.A2(n_273),
.B1(n_308),
.B2(n_307),
.Y(n_398)
);

INVxp67_ASAP7_75t_L g445 ( 
.A(n_398),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_358),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_399),
.B(n_403),
.Y(n_461)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_353),
.Y(n_400)
);

INVxp67_ASAP7_75t_L g457 ( 
.A(n_400),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_377),
.B(n_298),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_358),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_338),
.A2(n_321),
.B1(n_280),
.B2(n_245),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_L g440 ( 
.A1(n_404),
.A2(n_408),
.B1(n_370),
.B2(n_349),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_358),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_405),
.B(n_406),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_SL g406 ( 
.A(n_368),
.B(n_280),
.Y(n_406)
);

XOR2xp5_ASAP7_75t_L g407 ( 
.A(n_357),
.B(n_274),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_407),
.B(n_414),
.C(n_431),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_344),
.A2(n_367),
.B1(n_352),
.B2(n_356),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_370),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_409),
.B(n_425),
.Y(n_462)
);

OAI21xp5_ASAP7_75t_SL g456 ( 
.A1(n_410),
.A2(n_422),
.B(n_428),
.Y(n_456)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_380),
.Y(n_412)
);

INVxp67_ASAP7_75t_L g464 ( 
.A(n_412),
.Y(n_464)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_347),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_SL g451 ( 
.A(n_413),
.B(n_416),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_384),
.B(n_372),
.C(n_351),
.Y(n_414)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_347),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_327),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_SL g460 ( 
.A(n_417),
.B(n_419),
.Y(n_460)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_327),
.Y(n_419)
);

OAI22xp33_ASAP7_75t_SL g463 ( 
.A1(n_420),
.A2(n_409),
.B1(n_435),
.B2(n_397),
.Y(n_463)
);

XNOR2xp5_ASAP7_75t_SL g421 ( 
.A(n_384),
.B(n_253),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_SL g477 ( 
.A(n_421),
.B(n_275),
.Y(n_477)
);

AOI21xp5_ASAP7_75t_SL g422 ( 
.A1(n_329),
.A2(n_303),
.B(n_248),
.Y(n_422)
);

BUFx5_ASAP7_75t_L g423 ( 
.A(n_369),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_423),
.Y(n_442)
);

AOI21xp5_ASAP7_75t_L g424 ( 
.A1(n_382),
.A2(n_270),
.B(n_255),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_SL g425 ( 
.A(n_354),
.B(n_266),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_SL g426 ( 
.A1(n_325),
.A2(n_254),
.B1(n_262),
.B2(n_239),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_378),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_427),
.B(n_430),
.Y(n_467)
);

AOI22xp33_ASAP7_75t_SL g428 ( 
.A1(n_340),
.A2(n_279),
.B1(n_292),
.B2(n_322),
.Y(n_428)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_332),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_L g431 ( 
.A(n_384),
.B(n_264),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_L g433 ( 
.A1(n_352),
.A2(n_239),
.B1(n_241),
.B2(n_267),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_371),
.B(n_247),
.Y(n_434)
);

BUFx24_ASAP7_75t_SL g475 ( 
.A(n_434),
.Y(n_475)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_370),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_435),
.B(n_436),
.Y(n_478)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_337),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_L g437 ( 
.A1(n_386),
.A2(n_241),
.B1(n_301),
.B2(n_289),
.Y(n_437)
);

XOR2xp5_ASAP7_75t_SL g438 ( 
.A(n_429),
.B(n_354),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_L g481 ( 
.A(n_438),
.B(n_477),
.Y(n_481)
);

AOI22xp33_ASAP7_75t_L g505 ( 
.A1(n_440),
.A2(n_463),
.B1(n_480),
.B2(n_363),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_429),
.B(n_354),
.C(n_328),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_443),
.B(n_444),
.C(n_468),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_407),
.B(n_328),
.C(n_329),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_432),
.Y(n_447)
);

CKINVDCx14_ASAP7_75t_R g502 ( 
.A(n_447),
.Y(n_502)
);

OAI22xp5_ASAP7_75t_L g448 ( 
.A1(n_408),
.A2(n_345),
.B1(n_375),
.B2(n_336),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_L g486 ( 
.A1(n_448),
.A2(n_469),
.B1(n_420),
.B2(n_410),
.Y(n_486)
);

AOI22xp5_ASAP7_75t_L g450 ( 
.A1(n_388),
.A2(n_333),
.B1(n_350),
.B2(n_339),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_SL g494 ( 
.A1(n_450),
.A2(n_453),
.B1(n_454),
.B2(n_465),
.Y(n_494)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_402),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_452),
.B(n_389),
.Y(n_485)
);

AOI22xp5_ASAP7_75t_L g453 ( 
.A1(n_415),
.A2(n_355),
.B1(n_343),
.B2(n_374),
.Y(n_453)
);

AOI22xp5_ASAP7_75t_L g454 ( 
.A1(n_415),
.A2(n_343),
.B1(n_365),
.B2(n_332),
.Y(n_454)
);

OAI21xp5_ASAP7_75t_L g455 ( 
.A1(n_418),
.A2(n_343),
.B(n_362),
.Y(n_455)
);

OAI21xp5_ASAP7_75t_SL g501 ( 
.A1(n_455),
.A2(n_458),
.B(n_472),
.Y(n_501)
);

XNOR2x1_ASAP7_75t_L g459 ( 
.A(n_421),
.B(n_362),
.Y(n_459)
);

XOR2xp5_ASAP7_75t_L g484 ( 
.A(n_459),
.B(n_425),
.Y(n_484)
);

AOI22xp5_ASAP7_75t_L g465 ( 
.A1(n_401),
.A2(n_330),
.B1(n_342),
.B2(n_369),
.Y(n_465)
);

AOI22xp5_ASAP7_75t_L g466 ( 
.A1(n_401),
.A2(n_342),
.B1(n_362),
.B2(n_360),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_SL g516 ( 
.A1(n_466),
.A2(n_474),
.B1(n_391),
.B2(n_331),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_414),
.B(n_431),
.C(n_406),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_418),
.B(n_337),
.C(n_383),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_470),
.B(n_394),
.C(n_387),
.Y(n_488)
);

OAI21xp5_ASAP7_75t_L g472 ( 
.A1(n_390),
.A2(n_385),
.B(n_376),
.Y(n_472)
);

AOI22xp5_ASAP7_75t_L g474 ( 
.A1(n_433),
.A2(n_326),
.B1(n_335),
.B2(n_341),
.Y(n_474)
);

OAI22xp5_ASAP7_75t_SL g476 ( 
.A1(n_420),
.A2(n_395),
.B1(n_404),
.B2(n_403),
.Y(n_476)
);

AOI22xp5_ASAP7_75t_L g490 ( 
.A1(n_476),
.A2(n_420),
.B1(n_399),
.B2(n_426),
.Y(n_490)
);

OAI22xp33_ASAP7_75t_SL g480 ( 
.A1(n_420),
.A2(n_341),
.B1(n_326),
.B2(n_381),
.Y(n_480)
);

CKINVDCx20_ASAP7_75t_R g482 ( 
.A(n_460),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_482),
.B(n_485),
.Y(n_533)
);

MAJx2_ASAP7_75t_L g525 ( 
.A(n_484),
.B(n_439),
.C(n_444),
.Y(n_525)
);

OAI22xp5_ASAP7_75t_L g558 ( 
.A1(n_486),
.A2(n_487),
.B1(n_490),
.B2(n_491),
.Y(n_558)
);

OAI22xp5_ASAP7_75t_L g487 ( 
.A1(n_447),
.A2(n_420),
.B1(n_395),
.B2(n_405),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g536 ( 
.A(n_488),
.B(n_500),
.C(n_510),
.Y(n_536)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_460),
.Y(n_489)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_489),
.Y(n_527)
);

AOI22xp5_ASAP7_75t_L g491 ( 
.A1(n_476),
.A2(n_424),
.B1(n_411),
.B2(n_437),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_451),
.Y(n_492)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_492),
.Y(n_532)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_451),
.Y(n_493)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_493),
.Y(n_540)
);

OAI22xp5_ASAP7_75t_L g495 ( 
.A1(n_466),
.A2(n_411),
.B1(n_412),
.B2(n_422),
.Y(n_495)
);

AOI22xp5_ASAP7_75t_L g523 ( 
.A1(n_495),
.A2(n_517),
.B1(n_480),
.B2(n_441),
.Y(n_523)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_478),
.Y(n_496)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_496),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_SL g497 ( 
.A(n_446),
.B(n_436),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_497),
.B(n_507),
.Y(n_554)
);

AOI22xp5_ASAP7_75t_L g498 ( 
.A1(n_440),
.A2(n_416),
.B1(n_413),
.B2(n_419),
.Y(n_498)
);

OAI22xp5_ASAP7_75t_SL g537 ( 
.A1(n_498),
.A2(n_504),
.B1(n_515),
.B2(n_474),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_478),
.B(n_417),
.Y(n_499)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_499),
.Y(n_545)
);

XNOR2xp5_ASAP7_75t_L g500 ( 
.A(n_468),
.B(n_346),
.Y(n_500)
);

AOI21xp5_ASAP7_75t_L g503 ( 
.A1(n_458),
.A2(n_364),
.B(n_430),
.Y(n_503)
);

AOI21xp5_ASAP7_75t_L g522 ( 
.A1(n_503),
.A2(n_512),
.B(n_456),
.Y(n_522)
);

AOI22xp5_ASAP7_75t_L g504 ( 
.A1(n_463),
.A2(n_400),
.B1(n_427),
.B2(n_392),
.Y(n_504)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_505),
.Y(n_549)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_473),
.Y(n_506)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_506),
.Y(n_551)
);

INVx1_ASAP7_75t_SL g507 ( 
.A(n_472),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_473),
.Y(n_508)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_508),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_471),
.B(n_392),
.Y(n_509)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_509),
.Y(n_559)
);

XOR2xp5_ASAP7_75t_L g510 ( 
.A(n_439),
.B(n_348),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_467),
.Y(n_511)
);

INVxp67_ASAP7_75t_L g539 ( 
.A(n_511),
.Y(n_539)
);

AOI21xp5_ASAP7_75t_L g512 ( 
.A1(n_456),
.A2(n_364),
.B(n_381),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_439),
.B(n_348),
.C(n_346),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g547 ( 
.A(n_513),
.B(n_470),
.C(n_464),
.Y(n_547)
);

CKINVDCx20_ASAP7_75t_R g514 ( 
.A(n_467),
.Y(n_514)
);

CKINVDCx20_ASAP7_75t_R g541 ( 
.A(n_514),
.Y(n_541)
);

AOI22xp5_ASAP7_75t_L g515 ( 
.A1(n_465),
.A2(n_391),
.B1(n_326),
.B2(n_363),
.Y(n_515)
);

AND2x2_ASAP7_75t_L g526 ( 
.A(n_516),
.B(n_519),
.Y(n_526)
);

OAI22xp5_ASAP7_75t_L g517 ( 
.A1(n_441),
.A2(n_323),
.B1(n_331),
.B2(n_263),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_SL g518 ( 
.A(n_452),
.B(n_361),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_SL g530 ( 
.A(n_518),
.B(n_461),
.Y(n_530)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_471),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_479),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_520),
.B(n_462),
.Y(n_535)
);

CKINVDCx20_ASAP7_75t_R g521 ( 
.A(n_457),
.Y(n_521)
);

CKINVDCx20_ASAP7_75t_R g543 ( 
.A(n_521),
.Y(n_543)
);

HB1xp67_ASAP7_75t_L g580 ( 
.A(n_522),
.Y(n_580)
);

OAI22xp5_ASAP7_75t_SL g563 ( 
.A1(n_523),
.A2(n_552),
.B1(n_482),
.B2(n_490),
.Y(n_563)
);

XNOR2xp5_ASAP7_75t_L g524 ( 
.A(n_510),
.B(n_468),
.Y(n_524)
);

XOR2xp5_ASAP7_75t_L g593 ( 
.A(n_524),
.B(n_528),
.Y(n_593)
);

MAJx2_ASAP7_75t_L g581 ( 
.A(n_525),
.B(n_438),
.C(n_477),
.Y(n_581)
);

XNOR2xp5_ASAP7_75t_L g528 ( 
.A(n_483),
.B(n_443),
.Y(n_528)
);

AO22x1_ASAP7_75t_SL g529 ( 
.A1(n_486),
.A2(n_448),
.B1(n_479),
.B2(n_469),
.Y(n_529)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_529),
.Y(n_578)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_530),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_SL g531 ( 
.A(n_485),
.B(n_475),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_SL g592 ( 
.A(n_531),
.B(n_544),
.Y(n_592)
);

XNOR2xp5_ASAP7_75t_L g534 ( 
.A(n_483),
.B(n_500),
.Y(n_534)
);

XNOR2xp5_ASAP7_75t_L g590 ( 
.A(n_534),
.B(n_540),
.Y(n_590)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_535),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_537),
.B(n_546),
.Y(n_570)
);

AOI21xp5_ASAP7_75t_L g538 ( 
.A1(n_501),
.A2(n_512),
.B(n_503),
.Y(n_538)
);

NOR3xp33_ASAP7_75t_L g562 ( 
.A(n_538),
.B(n_556),
.C(n_507),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_SL g544 ( 
.A(n_513),
.B(n_454),
.Y(n_544)
);

CKINVDCx20_ASAP7_75t_R g546 ( 
.A(n_502),
.Y(n_546)
);

MAJIxp5_ASAP7_75t_L g561 ( 
.A(n_547),
.B(n_557),
.C(n_560),
.Y(n_561)
);

CKINVDCx20_ASAP7_75t_R g548 ( 
.A(n_499),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_548),
.B(n_533),
.Y(n_571)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_497),
.B(n_453),
.Y(n_550)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_550),
.Y(n_573)
);

AOI22xp5_ASAP7_75t_L g552 ( 
.A1(n_487),
.A2(n_450),
.B1(n_461),
.B2(n_449),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_L g553 ( 
.A(n_488),
.B(n_442),
.Y(n_553)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_553),
.Y(n_574)
);

AOI21xp5_ASAP7_75t_L g556 ( 
.A1(n_501),
.A2(n_445),
.B(n_455),
.Y(n_556)
);

MAJIxp5_ASAP7_75t_L g557 ( 
.A(n_484),
.B(n_444),
.C(n_443),
.Y(n_557)
);

MAJIxp5_ASAP7_75t_L g560 ( 
.A(n_481),
.B(n_477),
.C(n_459),
.Y(n_560)
);

O2A1O1Ixp33_ASAP7_75t_SL g611 ( 
.A1(n_562),
.A2(n_556),
.B(n_529),
.C(n_549),
.Y(n_611)
);

AOI22xp5_ASAP7_75t_L g603 ( 
.A1(n_563),
.A2(n_566),
.B1(n_567),
.B2(n_569),
.Y(n_603)
);

MAJIxp5_ASAP7_75t_L g564 ( 
.A(n_528),
.B(n_470),
.C(n_481),
.Y(n_564)
);

MAJIxp5_ASAP7_75t_L g607 ( 
.A(n_564),
.B(n_583),
.C(n_585),
.Y(n_607)
);

XNOR2x2_ASAP7_75t_SL g565 ( 
.A(n_533),
.B(n_496),
.Y(n_565)
);

XNOR2xp5_ASAP7_75t_L g594 ( 
.A(n_565),
.B(n_542),
.Y(n_594)
);

AOI22xp5_ASAP7_75t_L g566 ( 
.A1(n_558),
.A2(n_494),
.B1(n_514),
.B2(n_498),
.Y(n_566)
);

OAI22xp5_ASAP7_75t_SL g567 ( 
.A1(n_552),
.A2(n_548),
.B1(n_541),
.B2(n_545),
.Y(n_567)
);

AOI22xp5_ASAP7_75t_L g569 ( 
.A1(n_541),
.A2(n_494),
.B1(n_495),
.B2(n_493),
.Y(n_569)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_571),
.Y(n_596)
);

NOR2xp33_ASAP7_75t_L g575 ( 
.A(n_546),
.B(n_521),
.Y(n_575)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_575),
.Y(n_598)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_527),
.Y(n_576)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_576),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_L g577 ( 
.A(n_543),
.B(n_492),
.Y(n_577)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_577),
.Y(n_605)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_527),
.Y(n_579)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_579),
.Y(n_606)
);

XOR2xp5_ASAP7_75t_L g604 ( 
.A(n_581),
.B(n_584),
.Y(n_604)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_532),
.Y(n_582)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_582),
.Y(n_613)
);

MAJIxp5_ASAP7_75t_L g583 ( 
.A(n_534),
.B(n_438),
.C(n_489),
.Y(n_583)
);

XNOR2xp5_ASAP7_75t_SL g584 ( 
.A(n_525),
.B(n_459),
.Y(n_584)
);

MAJIxp5_ASAP7_75t_L g585 ( 
.A(n_536),
.B(n_449),
.C(n_462),
.Y(n_585)
);

XNOR2xp5_ASAP7_75t_SL g586 ( 
.A(n_524),
.B(n_491),
.Y(n_586)
);

XOR2xp5_ASAP7_75t_L g610 ( 
.A(n_586),
.B(n_588),
.Y(n_610)
);

MAJx2_ASAP7_75t_L g587 ( 
.A(n_557),
.B(n_560),
.C(n_536),
.Y(n_587)
);

MAJIxp5_ASAP7_75t_SL g599 ( 
.A(n_587),
.B(n_540),
.C(n_542),
.Y(n_599)
);

XNOR2xp5_ASAP7_75t_SL g588 ( 
.A(n_547),
.B(n_554),
.Y(n_588)
);

MAJIxp5_ASAP7_75t_L g589 ( 
.A(n_532),
.B(n_511),
.C(n_519),
.Y(n_589)
);

MAJIxp5_ASAP7_75t_L g617 ( 
.A(n_589),
.B(n_590),
.C(n_506),
.Y(n_617)
);

OAI22xp5_ASAP7_75t_SL g591 ( 
.A1(n_545),
.A2(n_504),
.B1(n_469),
.B2(n_520),
.Y(n_591)
);

AOI22xp5_ASAP7_75t_L g609 ( 
.A1(n_591),
.A2(n_537),
.B1(n_523),
.B2(n_526),
.Y(n_609)
);

AO21x1_ASAP7_75t_L g623 ( 
.A1(n_594),
.A2(n_601),
.B(n_569),
.Y(n_623)
);

AOI22xp5_ASAP7_75t_SL g595 ( 
.A1(n_563),
.A2(n_539),
.B1(n_549),
.B2(n_554),
.Y(n_595)
);

OAI22xp5_ASAP7_75t_L g625 ( 
.A1(n_595),
.A2(n_609),
.B1(n_611),
.B2(n_614),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_567),
.B(n_543),
.Y(n_597)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_597),
.Y(n_628)
);

XNOR2xp5_ASAP7_75t_L g621 ( 
.A(n_599),
.B(n_608),
.Y(n_621)
);

OAI21xp5_ASAP7_75t_SL g601 ( 
.A1(n_570),
.A2(n_538),
.B(n_522),
.Y(n_601)
);

NOR2xp33_ASAP7_75t_L g602 ( 
.A(n_574),
.B(n_539),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_602),
.B(n_616),
.Y(n_640)
);

XNOR2xp5_ASAP7_75t_L g608 ( 
.A(n_585),
.B(n_529),
.Y(n_608)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_565),
.Y(n_612)
);

INVx1_ASAP7_75t_SL g637 ( 
.A(n_612),
.Y(n_637)
);

AOI22xp5_ASAP7_75t_L g614 ( 
.A1(n_578),
.A2(n_559),
.B1(n_526),
.B2(n_516),
.Y(n_614)
);

XOR2xp5_ASAP7_75t_L g615 ( 
.A(n_593),
.B(n_559),
.Y(n_615)
);

XOR2xp5_ASAP7_75t_L g627 ( 
.A(n_615),
.B(n_619),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_571),
.B(n_555),
.Y(n_616)
);

XNOR2xp5_ASAP7_75t_L g626 ( 
.A(n_617),
.B(n_583),
.Y(n_626)
);

MAJIxp5_ASAP7_75t_L g618 ( 
.A(n_593),
.B(n_555),
.C(n_526),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_SL g624 ( 
.A(n_618),
.B(n_590),
.Y(n_624)
);

XOR2xp5_ASAP7_75t_L g619 ( 
.A(n_586),
.B(n_509),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_L g620 ( 
.A(n_568),
.B(n_573),
.Y(n_620)
);

OAI21x1_ASAP7_75t_L g622 ( 
.A1(n_620),
.A2(n_592),
.B(n_572),
.Y(n_622)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_622),
.Y(n_648)
);

OR2x2_ASAP7_75t_L g651 ( 
.A(n_623),
.B(n_604),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_SL g643 ( 
.A(n_624),
.B(n_626),
.Y(n_643)
);

AOI22xp5_ASAP7_75t_L g629 ( 
.A1(n_596),
.A2(n_570),
.B1(n_578),
.B2(n_566),
.Y(n_629)
);

AOI22xp5_ASAP7_75t_L g647 ( 
.A1(n_629),
.A2(n_603),
.B1(n_609),
.B2(n_614),
.Y(n_647)
);

AOI22xp5_ASAP7_75t_SL g630 ( 
.A1(n_597),
.A2(n_580),
.B1(n_612),
.B2(n_616),
.Y(n_630)
);

XNOR2xp5_ASAP7_75t_L g649 ( 
.A(n_630),
.B(n_634),
.Y(n_649)
);

MAJIxp5_ASAP7_75t_L g631 ( 
.A(n_607),
.B(n_561),
.C(n_587),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_SL g654 ( 
.A(n_631),
.B(n_632),
.Y(n_654)
);

MAJIxp5_ASAP7_75t_L g632 ( 
.A(n_607),
.B(n_561),
.C(n_588),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_SL g633 ( 
.A(n_598),
.B(n_589),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_SL g656 ( 
.A(n_633),
.B(n_635),
.Y(n_656)
);

AOI22xp5_ASAP7_75t_SL g634 ( 
.A1(n_611),
.A2(n_591),
.B1(n_584),
.B2(n_581),
.Y(n_634)
);

MAJIxp5_ASAP7_75t_L g635 ( 
.A(n_615),
.B(n_564),
.C(n_508),
.Y(n_635)
);

AND2x2_ASAP7_75t_L g636 ( 
.A(n_618),
.B(n_517),
.Y(n_636)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_636),
.Y(n_652)
);

CKINVDCx16_ASAP7_75t_R g638 ( 
.A(n_595),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_SL g659 ( 
.A(n_638),
.B(n_642),
.Y(n_659)
);

NOR2xp67_ASAP7_75t_SL g639 ( 
.A(n_608),
.B(n_551),
.Y(n_639)
);

AOI21xp5_ASAP7_75t_L g646 ( 
.A1(n_639),
.A2(n_594),
.B(n_601),
.Y(n_646)
);

XNOR2xp5_ASAP7_75t_L g641 ( 
.A(n_599),
.B(n_515),
.Y(n_641)
);

NOR2xp33_ASAP7_75t_L g653 ( 
.A(n_641),
.B(n_613),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_SL g642 ( 
.A(n_605),
.B(n_551),
.Y(n_642)
);

MAJIxp5_ASAP7_75t_L g644 ( 
.A(n_635),
.B(n_617),
.C(n_610),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_644),
.B(n_645),
.Y(n_662)
);

MAJIxp5_ASAP7_75t_L g645 ( 
.A(n_631),
.B(n_610),
.C(n_619),
.Y(n_645)
);

OR2x2_ASAP7_75t_L g672 ( 
.A(n_646),
.B(n_650),
.Y(n_672)
);

INVxp67_ASAP7_75t_L g667 ( 
.A(n_647),
.Y(n_667)
);

AOI21xp5_ASAP7_75t_L g650 ( 
.A1(n_623),
.A2(n_603),
.B(n_604),
.Y(n_650)
);

OAI21x1_ASAP7_75t_L g663 ( 
.A1(n_651),
.A2(n_646),
.B(n_650),
.Y(n_663)
);

AOI22xp33_ASAP7_75t_SL g666 ( 
.A1(n_653),
.A2(n_637),
.B1(n_625),
.B2(n_636),
.Y(n_666)
);

AOI22xp5_ASAP7_75t_L g655 ( 
.A1(n_628),
.A2(n_606),
.B1(n_600),
.B2(n_442),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_655),
.B(n_660),
.Y(n_665)
);

XOR2xp5_ASAP7_75t_L g657 ( 
.A(n_627),
.B(n_423),
.Y(n_657)
);

XOR2xp5_ASAP7_75t_L g664 ( 
.A(n_657),
.B(n_658),
.Y(n_664)
);

XNOR2xp5_ASAP7_75t_SL g658 ( 
.A(n_621),
.B(n_246),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_SL g660 ( 
.A(n_632),
.B(n_323),
.Y(n_660)
);

CKINVDCx16_ASAP7_75t_R g661 ( 
.A(n_640),
.Y(n_661)
);

NOR2xp33_ASAP7_75t_L g669 ( 
.A(n_661),
.B(n_637),
.Y(n_669)
);

NAND2x1_ASAP7_75t_L g681 ( 
.A(n_663),
.B(n_658),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_666),
.B(n_669),
.Y(n_683)
);

XOR2xp5_ASAP7_75t_L g668 ( 
.A(n_644),
.B(n_626),
.Y(n_668)
);

XOR2xp5_ASAP7_75t_L g684 ( 
.A(n_668),
.B(n_670),
.Y(n_684)
);

MAJIxp5_ASAP7_75t_L g670 ( 
.A(n_654),
.B(n_636),
.C(n_621),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_670),
.B(n_671),
.Y(n_685)
);

NOR2xp33_ASAP7_75t_SL g671 ( 
.A(n_643),
.B(n_641),
.Y(n_671)
);

AOI21xp5_ASAP7_75t_L g673 ( 
.A1(n_648),
.A2(n_627),
.B(n_629),
.Y(n_673)
);

OR2x2_ASAP7_75t_L g680 ( 
.A(n_673),
.B(n_674),
.Y(n_680)
);

AOI22xp5_ASAP7_75t_SL g674 ( 
.A1(n_652),
.A2(n_659),
.B1(n_649),
.B2(n_651),
.Y(n_674)
);

OAI21xp5_ASAP7_75t_L g675 ( 
.A1(n_652),
.A2(n_630),
.B(n_634),
.Y(n_675)
);

AOI21xp5_ASAP7_75t_L g678 ( 
.A1(n_675),
.A2(n_647),
.B(n_657),
.Y(n_678)
);

NOR2xp33_ASAP7_75t_SL g676 ( 
.A(n_662),
.B(n_656),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_SL g690 ( 
.A(n_676),
.B(n_679),
.Y(n_690)
);

OAI21xp5_ASAP7_75t_L g677 ( 
.A1(n_672),
.A2(n_645),
.B(n_649),
.Y(n_677)
);

OR2x2_ASAP7_75t_L g687 ( 
.A(n_677),
.B(n_678),
.Y(n_687)
);

NOR2xp33_ASAP7_75t_SL g679 ( 
.A(n_668),
.B(n_655),
.Y(n_679)
);

OAI21xp5_ASAP7_75t_L g691 ( 
.A1(n_681),
.A2(n_682),
.B(n_674),
.Y(n_691)
);

AOI21xp5_ASAP7_75t_L g682 ( 
.A1(n_672),
.A2(n_361),
.B(n_296),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_684),
.B(n_667),
.Y(n_688)
);

AOI21xp5_ASAP7_75t_SL g686 ( 
.A1(n_683),
.A2(n_675),
.B(n_665),
.Y(n_686)
);

OAI21xp5_ASAP7_75t_L g694 ( 
.A1(n_686),
.A2(n_680),
.B(n_684),
.Y(n_694)
);

AND2x2_ASAP7_75t_L g693 ( 
.A(n_688),
.B(n_689),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_685),
.B(n_667),
.Y(n_689)
);

AO21x1_ASAP7_75t_L g692 ( 
.A1(n_691),
.A2(n_680),
.B(n_681),
.Y(n_692)
);

AOI21xp5_ASAP7_75t_L g695 ( 
.A1(n_692),
.A2(n_694),
.B(n_687),
.Y(n_695)
);

MAJIxp5_ASAP7_75t_L g697 ( 
.A(n_695),
.B(n_696),
.C(n_664),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_693),
.B(n_690),
.Y(n_696)
);

OAI21xp5_ASAP7_75t_L g698 ( 
.A1(n_697),
.A2(n_664),
.B(n_236),
.Y(n_698)
);

A2O1A1Ixp33_ASAP7_75t_SL g699 ( 
.A1(n_698),
.A2(n_287),
.B(n_249),
.C(n_312),
.Y(n_699)
);

MAJIxp5_ASAP7_75t_L g700 ( 
.A(n_699),
.B(n_9),
.C(n_11),
.Y(n_700)
);


endmodule