module fake_ariane_1144_n_1223 (n_83, n_8, n_56, n_60, n_160, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_158, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_52, n_157, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1223);

input n_83;
input n_8;
input n_56;
input n_60;
input n_160;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_158;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_52;
input n_157;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1223;

wire n_295;
wire n_356;
wire n_556;
wire n_170;
wire n_190;
wire n_698;
wire n_1127;
wire n_1072;
wire n_695;
wire n_913;
wire n_180;
wire n_730;
wire n_386;
wire n_516;
wire n_307;
wire n_589;
wire n_332;
wire n_1008;
wire n_581;
wire n_294;
wire n_1020;
wire n_1209;
wire n_1137;
wire n_646;
wire n_1174;
wire n_197;
wire n_640;
wire n_463;
wire n_1024;
wire n_830;
wire n_176;
wire n_691;
wire n_1214;
wire n_404;
wire n_172;
wire n_943;
wire n_1118;
wire n_678;
wire n_1058;
wire n_651;
wire n_987;
wire n_936;
wire n_347;
wire n_423;
wire n_1042;
wire n_961;
wire n_183;
wire n_469;
wire n_1046;
wire n_479;
wire n_726;
wire n_603;
wire n_1123;
wire n_878;
wire n_373;
wire n_299;
wire n_836;
wire n_541;
wire n_499;
wire n_1169;
wire n_789;
wire n_788;
wire n_850;
wire n_908;
wire n_771;
wire n_1036;
wire n_564;
wire n_610;
wire n_205;
wire n_752;
wire n_1029;
wire n_341;
wire n_1187;
wire n_985;
wire n_245;
wire n_421;
wire n_549;
wire n_760;
wire n_522;
wire n_319;
wire n_591;
wire n_906;
wire n_690;
wire n_1180;
wire n_416;
wire n_969;
wire n_283;
wire n_1109;
wire n_919;
wire n_525;
wire n_187;
wire n_806;
wire n_367;
wire n_1111;
wire n_970;
wire n_713;
wire n_649;
wire n_598;
wire n_345;
wire n_374;
wire n_318;
wire n_817;
wire n_643;
wire n_679;
wire n_244;
wire n_226;
wire n_924;
wire n_927;
wire n_781;
wire n_220;
wire n_261;
wire n_1095;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_189;
wire n_717;
wire n_819;
wire n_286;
wire n_443;
wire n_586;
wire n_864;
wire n_952;
wire n_1096;
wire n_686;
wire n_605;
wire n_776;
wire n_424;
wire n_528;
wire n_584;
wire n_1154;
wire n_1166;
wire n_387;
wire n_1200;
wire n_406;
wire n_826;
wire n_1130;
wire n_524;
wire n_391;
wire n_349;
wire n_634;
wire n_756;
wire n_466;
wire n_940;
wire n_1016;
wire n_346;
wire n_1138;
wire n_214;
wire n_1149;
wire n_764;
wire n_979;
wire n_348;
wire n_552;
wire n_1077;
wire n_462;
wire n_1196;
wire n_607;
wire n_670;
wire n_897;
wire n_956;
wire n_949;
wire n_410;
wire n_1181;
wire n_379;
wire n_445;
wire n_515;
wire n_807;
wire n_765;
wire n_1131;
wire n_264;
wire n_891;
wire n_737;
wire n_885;
wire n_198;
wire n_232;
wire n_441;
wire n_568;
wire n_1032;
wire n_1217;
wire n_385;
wire n_637;
wire n_917;
wire n_1208;
wire n_327;
wire n_1088;
wire n_766;
wire n_372;
wire n_1177;
wire n_377;
wire n_396;
wire n_802;
wire n_631;
wire n_399;
wire n_1167;
wire n_1170;
wire n_1151;
wire n_554;
wire n_960;
wire n_520;
wire n_980;
wire n_870;
wire n_714;
wire n_905;
wire n_279;
wire n_958;
wire n_702;
wire n_945;
wire n_790;
wire n_857;
wire n_207;
wire n_898;
wire n_363;
wire n_720;
wire n_968;
wire n_1067;
wire n_354;
wire n_813;
wire n_926;
wire n_725;
wire n_419;
wire n_1009;
wire n_230;
wire n_270;
wire n_194;
wire n_1064;
wire n_633;
wire n_900;
wire n_1133;
wire n_883;
wire n_338;
wire n_1163;
wire n_995;
wire n_285;
wire n_1093;
wire n_473;
wire n_186;
wire n_801;
wire n_1184;
wire n_202;
wire n_193;
wire n_733;
wire n_761;
wire n_818;
wire n_500;
wire n_665;
wire n_336;
wire n_731;
wire n_754;
wire n_779;
wire n_871;
wire n_315;
wire n_903;
wire n_1073;
wire n_594;
wire n_1173;
wire n_311;
wire n_239;
wire n_402;
wire n_1068;
wire n_1052;
wire n_272;
wire n_829;
wire n_1198;
wire n_1062;
wire n_668;
wire n_339;
wire n_738;
wire n_758;
wire n_833;
wire n_672;
wire n_487;
wire n_740;
wire n_879;
wire n_1117;
wire n_167;
wire n_422;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_597;
wire n_816;
wire n_1018;
wire n_855;
wire n_1047;
wire n_259;
wire n_835;
wire n_808;
wire n_953;
wire n_446;
wire n_553;
wire n_1076;
wire n_753;
wire n_1050;
wire n_566;
wire n_814;
wire n_578;
wire n_701;
wire n_1003;
wire n_1125;
wire n_625;
wire n_405;
wire n_557;
wire n_169;
wire n_1201;
wire n_1107;
wire n_173;
wire n_858;
wire n_645;
wire n_989;
wire n_242;
wire n_331;
wire n_309;
wire n_320;
wire n_559;
wire n_1134;
wire n_1185;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_1035;
wire n_1141;
wire n_350;
wire n_291;
wire n_822;
wire n_1143;
wire n_381;
wire n_344;
wire n_840;
wire n_721;
wire n_433;
wire n_481;
wire n_600;
wire n_426;
wire n_795;
wire n_1053;
wire n_1084;
wire n_398;
wire n_210;
wire n_1090;
wire n_200;
wire n_529;
wire n_502;
wire n_166;
wire n_253;
wire n_561;
wire n_770;
wire n_218;
wire n_821;
wire n_839;
wire n_928;
wire n_1099;
wire n_271;
wire n_1153;
wire n_507;
wire n_486;
wire n_465;
wire n_901;
wire n_759;
wire n_247;
wire n_569;
wire n_567;
wire n_825;
wire n_732;
wire n_1103;
wire n_1145;
wire n_971;
wire n_240;
wire n_369;
wire n_1192;
wire n_224;
wire n_787;
wire n_894;
wire n_1105;
wire n_547;
wire n_1195;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_1172;
wire n_222;
wire n_478;
wire n_703;
wire n_1207;
wire n_748;
wire n_1212;
wire n_786;
wire n_510;
wire n_1061;
wire n_1045;
wire n_831;
wire n_256;
wire n_868;
wire n_326;
wire n_681;
wire n_778;
wire n_227;
wire n_1160;
wire n_874;
wire n_188;
wire n_323;
wire n_550;
wire n_1023;
wire n_997;
wire n_635;
wire n_707;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_694;
wire n_884;
wire n_1116;
wire n_983;
wire n_282;
wire n_328;
wire n_368;
wire n_1113;
wire n_1034;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_248;
wire n_277;
wire n_467;
wire n_1085;
wire n_1152;
wire n_432;
wire n_545;
wire n_1015;
wire n_1162;
wire n_536;
wire n_644;
wire n_293;
wire n_823;
wire n_921;
wire n_620;
wire n_1197;
wire n_228;
wire n_325;
wire n_276;
wire n_1074;
wire n_688;
wire n_859;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_1098;
wire n_693;
wire n_863;
wire n_1165;
wire n_303;
wire n_671;
wire n_442;
wire n_777;
wire n_929;
wire n_168;
wire n_352;
wire n_538;
wire n_206;
wire n_920;
wire n_899;
wire n_576;
wire n_843;
wire n_1080;
wire n_511;
wire n_1086;
wire n_611;
wire n_1092;
wire n_365;
wire n_455;
wire n_429;
wire n_238;
wire n_654;
wire n_588;
wire n_1013;
wire n_986;
wire n_1104;
wire n_638;
wire n_334;
wire n_192;
wire n_1128;
wire n_729;
wire n_887;
wire n_661;
wire n_488;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_1122;
wire n_1205;
wire n_300;
wire n_533;
wire n_904;
wire n_505;
wire n_163;
wire n_869;
wire n_846;
wire n_1132;
wire n_390;
wire n_1156;
wire n_498;
wire n_501;
wire n_438;
wire n_1059;
wire n_314;
wire n_684;
wire n_1120;
wire n_440;
wire n_1202;
wire n_627;
wire n_1039;
wire n_1188;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_1150;
wire n_233;
wire n_728;
wire n_977;
wire n_388;
wire n_449;
wire n_333;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_957;
wire n_1216;
wire n_512;
wire n_715;
wire n_889;
wire n_1066;
wire n_935;
wire n_579;
wire n_1218;
wire n_844;
wire n_1012;
wire n_459;
wire n_685;
wire n_221;
wire n_321;
wire n_911;
wire n_1136;
wire n_361;
wire n_458;
wire n_1190;
wire n_1144;
wire n_383;
wire n_623;
wire n_838;
wire n_1213;
wire n_237;
wire n_780;
wire n_861;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_877;
wire n_1021;
wire n_1065;
wire n_453;
wire n_1119;
wire n_734;
wire n_491;
wire n_810;
wire n_181;
wire n_723;
wire n_1142;
wire n_617;
wire n_616;
wire n_658;
wire n_705;
wire n_630;
wire n_1140;
wire n_570;
wire n_1055;
wire n_260;
wire n_362;
wire n_543;
wire n_942;
wire n_310;
wire n_709;
wire n_601;
wire n_683;
wire n_236;
wire n_565;
wire n_1089;
wire n_281;
wire n_628;
wire n_809;
wire n_461;
wire n_1121;
wire n_490;
wire n_262;
wire n_209;
wire n_743;
wire n_1194;
wire n_225;
wire n_907;
wire n_235;
wire n_1006;
wire n_881;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_1019;
wire n_297;
wire n_962;
wire n_662;
wire n_641;
wire n_1005;
wire n_503;
wire n_941;
wire n_1112;
wire n_700;
wire n_1159;
wire n_910;
wire n_1210;
wire n_290;
wire n_527;
wire n_741;
wire n_772;
wire n_747;
wire n_847;
wire n_939;
wire n_1135;
wire n_371;
wire n_845;
wire n_888;
wire n_199;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_217;
wire n_1114;
wire n_676;
wire n_178;
wire n_708;
wire n_551;
wire n_308;
wire n_417;
wire n_201;
wire n_1038;
wire n_572;
wire n_343;
wire n_1199;
wire n_865;
wire n_1222;
wire n_1041;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_993;
wire n_380;
wire n_948;
wire n_582;
wire n_284;
wire n_922;
wire n_1004;
wire n_448;
wire n_593;
wire n_755;
wire n_1097;
wire n_1219;
wire n_710;
wire n_860;
wire n_249;
wire n_534;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_609;
wire n_851;
wire n_1043;
wire n_278;
wire n_255;
wire n_560;
wire n_450;
wire n_890;
wire n_257;
wire n_1193;
wire n_842;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_1022;
wire n_1033;
wire n_896;
wire n_409;
wire n_171;
wire n_947;
wire n_930;
wire n_519;
wire n_902;
wire n_384;
wire n_1031;
wire n_1179;
wire n_468;
wire n_1056;
wire n_853;
wire n_526;
wire n_742;
wire n_716;
wire n_1081;
wire n_182;
wire n_696;
wire n_1040;
wire n_674;
wire n_482;
wire n_316;
wire n_196;
wire n_1158;
wire n_798;
wire n_769;
wire n_820;
wire n_577;
wire n_407;
wire n_774;
wire n_872;
wire n_933;
wire n_916;
wire n_254;
wire n_596;
wire n_954;
wire n_912;
wire n_1168;
wire n_476;
wire n_460;
wire n_219;
wire n_832;
wire n_535;
wire n_231;
wire n_366;
wire n_744;
wire n_762;
wire n_656;
wire n_1157;
wire n_555;
wire n_492;
wire n_234;
wire n_574;
wire n_848;
wire n_804;
wire n_280;
wire n_982;
wire n_915;
wire n_215;
wire n_252;
wire n_664;
wire n_629;
wire n_1075;
wire n_454;
wire n_966;
wire n_992;
wire n_298;
wire n_955;
wire n_532;
wire n_415;
wire n_794;
wire n_1182;
wire n_763;
wire n_655;
wire n_540;
wire n_544;
wire n_216;
wire n_692;
wire n_1186;
wire n_599;
wire n_768;
wire n_1091;
wire n_514;
wire n_418;
wire n_984;
wire n_537;
wire n_1063;
wire n_223;
wire n_403;
wire n_750;
wire n_991;
wire n_834;
wire n_389;
wire n_1007;
wire n_800;
wire n_657;
wire n_513;
wire n_837;
wire n_288;
wire n_179;
wire n_812;
wire n_1126;
wire n_395;
wire n_621;
wire n_1178;
wire n_195;
wire n_606;
wire n_1026;
wire n_951;
wire n_938;
wire n_213;
wire n_862;
wire n_304;
wire n_895;
wire n_659;
wire n_583;
wire n_509;
wire n_1014;
wire n_724;
wire n_306;
wire n_666;
wire n_1000;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_1206;
wire n_378;
wire n_203;
wire n_436;
wire n_946;
wire n_757;
wire n_375;
wire n_324;
wire n_1030;
wire n_1146;
wire n_1100;
wire n_1171;
wire n_585;
wire n_875;
wire n_669;
wire n_785;
wire n_827;
wire n_931;
wire n_1203;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_697;
wire n_622;
wire n_967;
wire n_998;
wire n_999;
wire n_1083;
wire n_472;
wire n_937;
wire n_296;
wire n_265;
wire n_746;
wire n_208;
wire n_456;
wire n_292;
wire n_880;
wire n_793;
wire n_852;
wire n_1079;
wire n_174;
wire n_275;
wire n_704;
wire n_1060;
wire n_1175;
wire n_1044;
wire n_1148;
wire n_204;
wire n_751;
wire n_615;
wire n_1027;
wire n_1070;
wire n_996;
wire n_521;
wire n_1211;
wire n_963;
wire n_873;
wire n_1082;
wire n_1139;
wire n_496;
wire n_739;
wire n_1028;
wire n_342;
wire n_866;
wire n_517;
wire n_925;
wire n_246;
wire n_1221;
wire n_530;
wire n_1094;
wire n_792;
wire n_1001;
wire n_1115;
wire n_824;
wire n_428;
wire n_1002;
wire n_358;
wire n_580;
wire n_1051;
wire n_892;
wire n_608;
wire n_959;
wire n_494;
wire n_719;
wire n_434;
wire n_263;
wire n_360;
wire n_1102;
wire n_975;
wire n_1101;
wire n_1129;
wire n_563;
wire n_229;
wire n_394;
wire n_923;
wire n_1189;
wire n_1124;
wire n_250;
wire n_932;
wire n_1183;
wire n_773;
wire n_165;
wire n_1037;
wire n_981;
wire n_1010;
wire n_882;
wire n_990;
wire n_1110;
wire n_317;
wire n_867;
wire n_243;
wire n_803;
wire n_329;
wire n_718;
wire n_185;
wire n_340;
wire n_944;
wire n_749;
wire n_1204;
wire n_994;
wire n_289;
wire n_548;
wire n_542;
wire n_815;
wire n_973;
wire n_523;
wire n_1078;
wire n_268;
wire n_972;
wire n_470;
wire n_266;
wire n_457;
wire n_1087;
wire n_164;
wire n_632;
wire n_184;
wire n_177;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_782;
wire n_856;
wire n_425;
wire n_1161;
wire n_431;
wire n_1176;
wire n_811;
wire n_1054;
wire n_508;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1155;
wire n_1191;
wire n_1071;
wire n_484;
wire n_712;
wire n_411;
wire n_849;
wire n_909;
wire n_976;
wire n_353;
wire n_736;
wire n_767;
wire n_1025;
wire n_1164;
wire n_1215;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_964;
wire n_1057;
wire n_382;
wire n_191;
wire n_797;
wire n_489;
wire n_480;
wire n_978;
wire n_211;
wire n_642;
wire n_1011;
wire n_408;
wire n_828;
wire n_595;
wire n_322;
wire n_251;
wire n_974;
wire n_506;
wire n_893;
wire n_602;
wire n_799;
wire n_558;
wire n_1147;
wire n_592;
wire n_397;
wire n_854;
wire n_841;
wire n_471;
wire n_351;
wire n_886;
wire n_965;
wire n_393;
wire n_1069;
wire n_474;
wire n_653;
wire n_359;
wire n_573;
wire n_796;
wire n_805;
wire n_934;
wire n_531;
wire n_783;
wire n_1220;
wire n_675;

INVx2_ASAP7_75t_L g163 ( 
.A(n_138),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_30),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_100),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_115),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_143),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_111),
.Y(n_168)
);

BUFx10_ASAP7_75t_L g169 ( 
.A(n_80),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_15),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_22),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_83),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_12),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_157),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_75),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_123),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_37),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_125),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_147),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_2),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_27),
.Y(n_181)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_37),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_62),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_82),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_2),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_160),
.Y(n_186)
);

INVx1_ASAP7_75t_SL g187 ( 
.A(n_90),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_150),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_49),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_128),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_32),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_86),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_110),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_59),
.Y(n_194)
);

CKINVDCx14_ASAP7_75t_R g195 ( 
.A(n_146),
.Y(n_195)
);

INVx1_ASAP7_75t_SL g196 ( 
.A(n_104),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_8),
.Y(n_197)
);

INVx2_ASAP7_75t_SL g198 ( 
.A(n_108),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_144),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_15),
.Y(n_200)
);

HB1xp67_ASAP7_75t_L g201 ( 
.A(n_162),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_12),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_152),
.Y(n_203)
);

INVx1_ASAP7_75t_SL g204 ( 
.A(n_158),
.Y(n_204)
);

INVx2_ASAP7_75t_SL g205 ( 
.A(n_41),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_49),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_159),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_76),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_51),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_0),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_13),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_50),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_148),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_7),
.Y(n_214)
);

BUFx10_ASAP7_75t_L g215 ( 
.A(n_63),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_18),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_117),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_20),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_153),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_120),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_27),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_81),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_10),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_106),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_73),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_47),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_95),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_118),
.Y(n_228)
);

INVx1_ASAP7_75t_SL g229 ( 
.A(n_136),
.Y(n_229)
);

BUFx3_ASAP7_75t_L g230 ( 
.A(n_103),
.Y(n_230)
);

INVx2_ASAP7_75t_SL g231 ( 
.A(n_135),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_44),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_45),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_55),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_10),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_91),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_40),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_11),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_161),
.Y(n_239)
);

INVx2_ASAP7_75t_SL g240 ( 
.A(n_156),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_154),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_122),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_132),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_99),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_151),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_145),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_142),
.Y(n_247)
);

INVx1_ASAP7_75t_SL g248 ( 
.A(n_47),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_43),
.Y(n_249)
);

INVx1_ASAP7_75t_SL g250 ( 
.A(n_14),
.Y(n_250)
);

INVx1_ASAP7_75t_SL g251 ( 
.A(n_68),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_70),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_72),
.Y(n_253)
);

BUFx10_ASAP7_75t_L g254 ( 
.A(n_94),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_89),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_9),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_107),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_1),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_1),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_78),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_55),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_53),
.Y(n_262)
);

INVx1_ASAP7_75t_SL g263 ( 
.A(n_109),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_149),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_21),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_40),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_77),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_131),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_28),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_3),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_137),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_155),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_43),
.Y(n_273)
);

BUFx5_ASAP7_75t_L g274 ( 
.A(n_18),
.Y(n_274)
);

CKINVDCx16_ASAP7_75t_R g275 ( 
.A(n_19),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_141),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_85),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_121),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_24),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_139),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_114),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_140),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_14),
.Y(n_283)
);

INVxp67_ASAP7_75t_SL g284 ( 
.A(n_283),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_274),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_274),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_274),
.Y(n_287)
);

CKINVDCx16_ASAP7_75t_R g288 ( 
.A(n_275),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_274),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_169),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_168),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_169),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_222),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_274),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_274),
.Y(n_295)
);

HB1xp67_ASAP7_75t_L g296 ( 
.A(n_170),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_205),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_169),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_274),
.Y(n_299)
);

BUFx3_ASAP7_75t_L g300 ( 
.A(n_230),
.Y(n_300)
);

BUFx3_ASAP7_75t_L g301 ( 
.A(n_230),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_247),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_215),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_272),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_274),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_164),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_195),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_164),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_215),
.Y(n_309)
);

BUFx2_ASAP7_75t_L g310 ( 
.A(n_170),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g311 ( 
.A(n_205),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_164),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_201),
.B(n_0),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_215),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_254),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_254),
.Y(n_316)
);

BUFx10_ASAP7_75t_L g317 ( 
.A(n_164),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_180),
.Y(n_318)
);

BUFx3_ASAP7_75t_L g319 ( 
.A(n_172),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_254),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_175),
.B(n_3),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_165),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_178),
.B(n_4),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_181),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_164),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_171),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_185),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_212),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_165),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_171),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_183),
.B(n_4),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_214),
.Y(n_332)
);

INVxp67_ASAP7_75t_L g333 ( 
.A(n_221),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_223),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_232),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_249),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_173),
.Y(n_337)
);

INVxp33_ASAP7_75t_L g338 ( 
.A(n_259),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_186),
.B(n_5),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_193),
.B(n_5),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_265),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_269),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_173),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_270),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_182),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_177),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_237),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_166),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_177),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_256),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_237),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_182),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_189),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_166),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_256),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_189),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_208),
.B(n_6),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_167),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_220),
.B(n_6),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_262),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_SL g361 ( 
.A(n_198),
.B(n_7),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_167),
.Y(n_362)
);

INVxp67_ASAP7_75t_SL g363 ( 
.A(n_237),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_237),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_262),
.Y(n_365)
);

INVxp67_ASAP7_75t_L g366 ( 
.A(n_258),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_237),
.Y(n_367)
);

INVxp67_ASAP7_75t_SL g368 ( 
.A(n_283),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_258),
.Y(n_369)
);

BUFx3_ASAP7_75t_L g370 ( 
.A(n_227),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_283),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_283),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_176),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_176),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_285),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_285),
.Y(n_376)
);

HB1xp67_ASAP7_75t_L g377 ( 
.A(n_310),
.Y(n_377)
);

AND2x2_ASAP7_75t_L g378 ( 
.A(n_319),
.B(n_283),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_299),
.Y(n_379)
);

CKINVDCx8_ASAP7_75t_R g380 ( 
.A(n_288),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_290),
.B(n_179),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_299),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_305),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_286),
.Y(n_384)
);

AND2x2_ASAP7_75t_L g385 ( 
.A(n_319),
.B(n_198),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_284),
.B(n_239),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_305),
.Y(n_387)
);

HB1xp67_ASAP7_75t_L g388 ( 
.A(n_310),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_363),
.B(n_245),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_306),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_287),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_289),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_306),
.Y(n_393)
);

BUFx6f_ASAP7_75t_L g394 ( 
.A(n_294),
.Y(n_394)
);

INVxp67_ASAP7_75t_L g395 ( 
.A(n_296),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_295),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_308),
.Y(n_397)
);

AND2x4_ASAP7_75t_L g398 ( 
.A(n_370),
.B(n_231),
.Y(n_398)
);

AND2x4_ASAP7_75t_L g399 ( 
.A(n_370),
.B(n_231),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_308),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_312),
.Y(n_401)
);

INVx3_ASAP7_75t_L g402 ( 
.A(n_317),
.Y(n_402)
);

INVxp67_ASAP7_75t_L g403 ( 
.A(n_300),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_326),
.A2(n_248),
.B1(n_250),
.B2(n_261),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_312),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_325),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_368),
.B(n_257),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_325),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_347),
.Y(n_409)
);

BUFx6f_ASAP7_75t_L g410 ( 
.A(n_347),
.Y(n_410)
);

BUFx6f_ASAP7_75t_L g411 ( 
.A(n_351),
.Y(n_411)
);

HB1xp67_ASAP7_75t_L g412 ( 
.A(n_330),
.Y(n_412)
);

INVxp67_ASAP7_75t_L g413 ( 
.A(n_300),
.Y(n_413)
);

INVx4_ASAP7_75t_L g414 ( 
.A(n_317),
.Y(n_414)
);

AND2x4_ASAP7_75t_L g415 ( 
.A(n_301),
.B(n_240),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_291),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_351),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_364),
.Y(n_418)
);

INVxp33_ASAP7_75t_L g419 ( 
.A(n_338),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_364),
.Y(n_420)
);

HB1xp67_ASAP7_75t_L g421 ( 
.A(n_337),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_371),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_301),
.B(n_260),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_SL g424 ( 
.A(n_290),
.B(n_179),
.Y(n_424)
);

BUFx6f_ASAP7_75t_L g425 ( 
.A(n_371),
.Y(n_425)
);

BUFx6f_ASAP7_75t_L g426 ( 
.A(n_372),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_372),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_367),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_317),
.B(n_264),
.Y(n_429)
);

AND2x4_ASAP7_75t_L g430 ( 
.A(n_318),
.B(n_240),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_292),
.B(n_252),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_345),
.Y(n_432)
);

BUFx6f_ASAP7_75t_L g433 ( 
.A(n_323),
.Y(n_433)
);

INVx5_ASAP7_75t_L g434 ( 
.A(n_321),
.Y(n_434)
);

AND2x6_ASAP7_75t_L g435 ( 
.A(n_331),
.B(n_163),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_352),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_353),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_356),
.Y(n_438)
);

BUFx6f_ASAP7_75t_L g439 ( 
.A(n_359),
.Y(n_439)
);

INVx3_ASAP7_75t_L g440 ( 
.A(n_360),
.Y(n_440)
);

OAI21x1_ASAP7_75t_L g441 ( 
.A1(n_361),
.A2(n_241),
.B(n_163),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_324),
.B(n_267),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_365),
.Y(n_443)
);

INVx6_ASAP7_75t_L g444 ( 
.A(n_339),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_384),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_384),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_384),
.Y(n_447)
);

BUFx3_ASAP7_75t_L g448 ( 
.A(n_375),
.Y(n_448)
);

NOR3xp33_ASAP7_75t_L g449 ( 
.A(n_395),
.B(n_313),
.C(n_340),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_385),
.B(n_292),
.Y(n_450)
);

INVx2_ASAP7_75t_SL g451 ( 
.A(n_444),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_391),
.Y(n_452)
);

INVx3_ASAP7_75t_L g453 ( 
.A(n_394),
.Y(n_453)
);

OR2x2_ASAP7_75t_L g454 ( 
.A(n_419),
.B(n_366),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_391),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_391),
.Y(n_456)
);

AOI22xp33_ASAP7_75t_L g457 ( 
.A1(n_435),
.A2(n_357),
.B1(n_298),
.B2(n_309),
.Y(n_457)
);

BUFx2_ASAP7_75t_L g458 ( 
.A(n_377),
.Y(n_458)
);

AOI22xp33_ASAP7_75t_L g459 ( 
.A1(n_435),
.A2(n_298),
.B1(n_309),
.B2(n_303),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_392),
.Y(n_460)
);

AOI22xp5_ASAP7_75t_L g461 ( 
.A1(n_435),
.A2(n_343),
.B1(n_349),
.B2(n_346),
.Y(n_461)
);

INVxp33_ASAP7_75t_SL g462 ( 
.A(n_412),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_375),
.B(n_303),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_392),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_392),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_SL g466 ( 
.A(n_403),
.B(n_322),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_385),
.B(n_402),
.Y(n_467)
);

BUFx10_ASAP7_75t_L g468 ( 
.A(n_444),
.Y(n_468)
);

INVx2_ASAP7_75t_SL g469 ( 
.A(n_444),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_444),
.B(n_322),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_396),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_396),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_396),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_390),
.Y(n_474)
);

INVx1_ASAP7_75t_SL g475 ( 
.A(n_416),
.Y(n_475)
);

AND2x2_ASAP7_75t_L g476 ( 
.A(n_385),
.B(n_430),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_390),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_393),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_376),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_376),
.Y(n_480)
);

INVx2_ASAP7_75t_SL g481 ( 
.A(n_444),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_393),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_400),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_400),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_SL g485 ( 
.A(n_403),
.B(n_329),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_401),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_402),
.B(n_314),
.Y(n_487)
);

INVx6_ASAP7_75t_L g488 ( 
.A(n_414),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_379),
.B(n_314),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_401),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_379),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_413),
.B(n_329),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_SL g493 ( 
.A(n_380),
.B(n_315),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_402),
.B(n_315),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_382),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_413),
.B(n_348),
.Y(n_496)
);

AOI22xp33_ASAP7_75t_L g497 ( 
.A1(n_435),
.A2(n_316),
.B1(n_320),
.B2(n_369),
.Y(n_497)
);

INVx3_ASAP7_75t_L g498 ( 
.A(n_394),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_405),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_382),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_405),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_383),
.Y(n_502)
);

INVx4_ASAP7_75t_L g503 ( 
.A(n_402),
.Y(n_503)
);

CKINVDCx20_ASAP7_75t_R g504 ( 
.A(n_380),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_406),
.Y(n_505)
);

AOI22xp5_ASAP7_75t_L g506 ( 
.A1(n_435),
.A2(n_404),
.B1(n_350),
.B2(n_355),
.Y(n_506)
);

BUFx4f_ASAP7_75t_L g507 ( 
.A(n_433),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_SL g508 ( 
.A(n_381),
.B(n_348),
.Y(n_508)
);

BUFx3_ASAP7_75t_L g509 ( 
.A(n_383),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_SL g510 ( 
.A(n_424),
.B(n_354),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_406),
.Y(n_511)
);

INVx4_ASAP7_75t_L g512 ( 
.A(n_414),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_409),
.Y(n_513)
);

INVxp33_ASAP7_75t_SL g514 ( 
.A(n_412),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_387),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_470),
.B(n_433),
.Y(n_516)
);

INVx3_ASAP7_75t_L g517 ( 
.A(n_448),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_467),
.B(n_451),
.Y(n_518)
);

A2O1A1Ixp33_ASAP7_75t_L g519 ( 
.A1(n_476),
.A2(n_404),
.B(n_441),
.C(n_442),
.Y(n_519)
);

BUFx3_ASAP7_75t_L g520 ( 
.A(n_448),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_474),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_474),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_450),
.B(n_433),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_477),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_455),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_477),
.Y(n_526)
);

INVx2_ASAP7_75t_SL g527 ( 
.A(n_454),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_451),
.B(n_433),
.Y(n_528)
);

OAI22xp5_ASAP7_75t_L g529 ( 
.A1(n_469),
.A2(n_433),
.B1(n_439),
.B2(n_395),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_SL g530 ( 
.A(n_468),
.B(n_469),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_SL g531 ( 
.A(n_468),
.B(n_433),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_SL g532 ( 
.A(n_468),
.B(n_433),
.Y(n_532)
);

BUFx6f_ASAP7_75t_L g533 ( 
.A(n_448),
.Y(n_533)
);

INVx3_ASAP7_75t_L g534 ( 
.A(n_509),
.Y(n_534)
);

OR2x2_ASAP7_75t_L g535 ( 
.A(n_458),
.B(n_377),
.Y(n_535)
);

BUFx6f_ASAP7_75t_L g536 ( 
.A(n_509),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_481),
.B(n_439),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_481),
.B(n_439),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_L g539 ( 
.A(n_463),
.B(n_439),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_476),
.B(n_439),
.Y(n_540)
);

OAI22xp5_ASAP7_75t_L g541 ( 
.A1(n_463),
.A2(n_439),
.B1(n_434),
.B2(n_388),
.Y(n_541)
);

NAND3xp33_ASAP7_75t_L g542 ( 
.A(n_492),
.B(n_358),
.C(n_354),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_489),
.B(n_439),
.Y(n_543)
);

INVxp67_ASAP7_75t_L g544 ( 
.A(n_454),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_478),
.Y(n_545)
);

AND2x4_ASAP7_75t_L g546 ( 
.A(n_489),
.B(n_430),
.Y(n_546)
);

INVx5_ASAP7_75t_L g547 ( 
.A(n_488),
.Y(n_547)
);

BUFx5_ASAP7_75t_L g548 ( 
.A(n_468),
.Y(n_548)
);

AOI22xp5_ASAP7_75t_L g549 ( 
.A1(n_449),
.A2(n_435),
.B1(n_431),
.B2(n_362),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_487),
.B(n_388),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_496),
.B(n_398),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_494),
.B(n_398),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_503),
.B(n_398),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_SL g554 ( 
.A(n_507),
.B(n_434),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_478),
.Y(n_555)
);

NOR2x1_ASAP7_75t_R g556 ( 
.A(n_458),
.B(n_358),
.Y(n_556)
);

AND2x2_ASAP7_75t_L g557 ( 
.A(n_475),
.B(n_316),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_503),
.B(n_398),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_503),
.B(n_398),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_SL g560 ( 
.A(n_475),
.B(n_380),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_503),
.B(n_399),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_482),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_509),
.B(n_399),
.Y(n_563)
);

NOR2xp67_ASAP7_75t_L g564 ( 
.A(n_506),
.B(n_320),
.Y(n_564)
);

INVxp67_ASAP7_75t_L g565 ( 
.A(n_493),
.Y(n_565)
);

HB1xp67_ASAP7_75t_L g566 ( 
.A(n_462),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_459),
.B(n_399),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_482),
.Y(n_568)
);

INVx3_ASAP7_75t_L g569 ( 
.A(n_479),
.Y(n_569)
);

OAI22xp33_ASAP7_75t_L g570 ( 
.A1(n_506),
.A2(n_362),
.B1(n_374),
.B2(n_373),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_L g571 ( 
.A(n_508),
.B(n_414),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_457),
.B(n_399),
.Y(n_572)
);

AND2x2_ASAP7_75t_L g573 ( 
.A(n_493),
.B(n_373),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_483),
.Y(n_574)
);

NAND2xp33_ASAP7_75t_L g575 ( 
.A(n_479),
.B(n_435),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_510),
.B(n_414),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_512),
.B(n_399),
.Y(n_577)
);

INVx2_ASAP7_75t_SL g578 ( 
.A(n_466),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_512),
.B(n_415),
.Y(n_579)
);

NOR2xp33_ASAP7_75t_L g580 ( 
.A(n_485),
.B(n_374),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_512),
.B(n_415),
.Y(n_581)
);

HB1xp67_ASAP7_75t_L g582 ( 
.A(n_514),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_L g583 ( 
.A(n_497),
.B(n_479),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_483),
.Y(n_584)
);

NOR2xp67_ASAP7_75t_L g585 ( 
.A(n_461),
.B(n_297),
.Y(n_585)
);

OR2x2_ASAP7_75t_L g586 ( 
.A(n_461),
.B(n_421),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_455),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_512),
.B(n_415),
.Y(n_588)
);

BUFx3_ASAP7_75t_L g589 ( 
.A(n_504),
.Y(n_589)
);

INVx2_ASAP7_75t_SL g590 ( 
.A(n_484),
.Y(n_590)
);

INVxp67_ASAP7_75t_L g591 ( 
.A(n_484),
.Y(n_591)
);

AOI22xp33_ASAP7_75t_L g592 ( 
.A1(n_480),
.A2(n_435),
.B1(n_434),
.B2(n_430),
.Y(n_592)
);

AOI22xp33_ASAP7_75t_L g593 ( 
.A1(n_480),
.A2(n_435),
.B1(n_434),
.B2(n_430),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_486),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_SL g595 ( 
.A(n_507),
.B(n_434),
.Y(n_595)
);

NAND2x1p5_ASAP7_75t_L g596 ( 
.A(n_507),
.B(n_440),
.Y(n_596)
);

NOR2xp33_ASAP7_75t_L g597 ( 
.A(n_480),
.B(n_386),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_491),
.B(n_415),
.Y(n_598)
);

AND2x2_ASAP7_75t_L g599 ( 
.A(n_491),
.B(n_421),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_486),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_490),
.Y(n_601)
);

OR2x2_ASAP7_75t_L g602 ( 
.A(n_445),
.B(n_423),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_SL g603 ( 
.A(n_507),
.B(n_434),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_490),
.Y(n_604)
);

INVxp67_ASAP7_75t_L g605 ( 
.A(n_499),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_455),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_491),
.B(n_415),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_495),
.B(n_500),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_495),
.B(n_429),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_495),
.B(n_429),
.Y(n_610)
);

OAI22xp5_ASAP7_75t_SL g611 ( 
.A1(n_499),
.A2(n_293),
.B1(n_304),
.B2(n_302),
.Y(n_611)
);

BUFx2_ASAP7_75t_L g612 ( 
.A(n_453),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_500),
.B(n_378),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_546),
.B(n_430),
.Y(n_614)
);

O2A1O1Ixp33_ASAP7_75t_L g615 ( 
.A1(n_540),
.A2(n_502),
.B(n_515),
.C(n_500),
.Y(n_615)
);

AOI21xp5_ASAP7_75t_L g616 ( 
.A1(n_516),
.A2(n_515),
.B(n_502),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_L g617 ( 
.A(n_550),
.B(n_502),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_569),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_546),
.B(n_515),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_521),
.Y(n_620)
);

AND2x2_ASAP7_75t_L g621 ( 
.A(n_544),
.B(n_311),
.Y(n_621)
);

AOI21xp5_ASAP7_75t_L g622 ( 
.A1(n_516),
.A2(n_498),
.B(n_453),
.Y(n_622)
);

O2A1O1Ixp33_ASAP7_75t_L g623 ( 
.A1(n_570),
.A2(n_501),
.B(n_511),
.C(n_505),
.Y(n_623)
);

AOI21xp5_ASAP7_75t_L g624 ( 
.A1(n_575),
.A2(n_498),
.B(n_453),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_SL g625 ( 
.A(n_548),
.B(n_434),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_546),
.B(n_423),
.Y(n_626)
);

BUFx12f_ASAP7_75t_L g627 ( 
.A(n_527),
.Y(n_627)
);

AND2x2_ASAP7_75t_L g628 ( 
.A(n_566),
.B(n_333),
.Y(n_628)
);

AOI21xp5_ASAP7_75t_L g629 ( 
.A1(n_528),
.A2(n_498),
.B(n_453),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_SL g630 ( 
.A(n_548),
.B(n_533),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_L g631 ( 
.A(n_550),
.B(n_498),
.Y(n_631)
);

OAI21xp5_ASAP7_75t_L g632 ( 
.A1(n_539),
.A2(n_446),
.B(n_445),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_591),
.B(n_378),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_605),
.B(n_378),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_SL g635 ( 
.A(n_548),
.B(n_434),
.Y(n_635)
);

AOI21xp5_ASAP7_75t_L g636 ( 
.A1(n_537),
.A2(n_538),
.B(n_532),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_539),
.B(n_446),
.Y(n_637)
);

BUFx6f_ASAP7_75t_L g638 ( 
.A(n_533),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_522),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_L g640 ( 
.A(n_565),
.B(n_501),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_543),
.B(n_551),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_SL g642 ( 
.A(n_548),
.B(n_447),
.Y(n_642)
);

AND2x2_ASAP7_75t_SL g643 ( 
.A(n_583),
.B(n_241),
.Y(n_643)
);

AND2x2_ASAP7_75t_L g644 ( 
.A(n_582),
.B(n_442),
.Y(n_644)
);

AOI21xp5_ASAP7_75t_L g645 ( 
.A1(n_531),
.A2(n_511),
.B(n_505),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_569),
.Y(n_646)
);

NOR2xp33_ASAP7_75t_L g647 ( 
.A(n_573),
.B(n_513),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_543),
.B(n_597),
.Y(n_648)
);

AOI21xp5_ASAP7_75t_L g649 ( 
.A1(n_531),
.A2(n_513),
.B(n_452),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_597),
.B(n_447),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_SL g651 ( 
.A(n_548),
.B(n_452),
.Y(n_651)
);

AND2x2_ASAP7_75t_L g652 ( 
.A(n_557),
.B(n_443),
.Y(n_652)
);

AOI22xp5_ASAP7_75t_L g653 ( 
.A1(n_580),
.A2(n_488),
.B1(n_460),
.B2(n_464),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_590),
.B(n_456),
.Y(n_654)
);

AOI22xp5_ASAP7_75t_L g655 ( 
.A1(n_580),
.A2(n_488),
.B1(n_460),
.B2(n_464),
.Y(n_655)
);

AOI21xp5_ASAP7_75t_L g656 ( 
.A1(n_532),
.A2(n_471),
.B(n_456),
.Y(n_656)
);

AOI21xp5_ASAP7_75t_L g657 ( 
.A1(n_518),
.A2(n_608),
.B(n_547),
.Y(n_657)
);

NOR2xp33_ASAP7_75t_L g658 ( 
.A(n_578),
.B(n_542),
.Y(n_658)
);

OAI21xp5_ASAP7_75t_L g659 ( 
.A1(n_523),
.A2(n_472),
.B(n_471),
.Y(n_659)
);

INVx2_ASAP7_75t_SL g660 ( 
.A(n_589),
.Y(n_660)
);

NAND3xp33_ASAP7_75t_L g661 ( 
.A(n_535),
.B(n_473),
.C(n_472),
.Y(n_661)
);

AND2x4_ASAP7_75t_L g662 ( 
.A(n_599),
.B(n_443),
.Y(n_662)
);

INVx3_ASAP7_75t_L g663 ( 
.A(n_520),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_523),
.B(n_473),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_525),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_SL g666 ( 
.A(n_548),
.B(n_465),
.Y(n_666)
);

AOI21xp5_ASAP7_75t_L g667 ( 
.A1(n_547),
.A2(n_465),
.B(n_387),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_525),
.Y(n_668)
);

OAI21xp5_ASAP7_75t_L g669 ( 
.A1(n_553),
.A2(n_465),
.B(n_441),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_609),
.B(n_386),
.Y(n_670)
);

NAND2x1_ASAP7_75t_L g671 ( 
.A(n_517),
.B(n_488),
.Y(n_671)
);

BUFx6f_ASAP7_75t_L g672 ( 
.A(n_533),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_SL g673 ( 
.A(n_533),
.B(n_394),
.Y(n_673)
);

INVx5_ASAP7_75t_L g674 ( 
.A(n_536),
.Y(n_674)
);

AOI21xp5_ASAP7_75t_L g675 ( 
.A1(n_547),
.A2(n_488),
.B(n_441),
.Y(n_675)
);

AOI21xp5_ASAP7_75t_L g676 ( 
.A1(n_547),
.A2(n_394),
.B(n_389),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_587),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_610),
.B(n_389),
.Y(n_678)
);

A2O1A1Ixp33_ASAP7_75t_L g679 ( 
.A1(n_583),
.A2(n_407),
.B(n_440),
.C(n_174),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_602),
.B(n_524),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_587),
.Y(n_681)
);

AOI21xp5_ASAP7_75t_L g682 ( 
.A1(n_558),
.A2(n_394),
.B(n_407),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_526),
.B(n_440),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_611),
.Y(n_684)
);

AOI22xp33_ASAP7_75t_L g685 ( 
.A1(n_572),
.A2(n_438),
.B1(n_437),
.B2(n_436),
.Y(n_685)
);

AOI21xp5_ASAP7_75t_L g686 ( 
.A1(n_559),
.A2(n_394),
.B(n_253),
.Y(n_686)
);

A2O1A1Ixp33_ASAP7_75t_L g687 ( 
.A1(n_545),
.A2(n_440),
.B(n_438),
.C(n_437),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_555),
.B(n_307),
.Y(n_688)
);

NOR2xp33_ASAP7_75t_L g689 ( 
.A(n_586),
.B(n_394),
.Y(n_689)
);

BUFx6f_ASAP7_75t_L g690 ( 
.A(n_536),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_562),
.Y(n_691)
);

NOR3xp33_ASAP7_75t_L g692 ( 
.A(n_556),
.B(n_261),
.C(n_194),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_606),
.Y(n_693)
);

AOI21xp5_ASAP7_75t_L g694 ( 
.A1(n_561),
.A2(n_253),
.B(n_252),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_606),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_568),
.B(n_432),
.Y(n_696)
);

OAI22xp5_ASAP7_75t_L g697 ( 
.A1(n_517),
.A2(n_211),
.B1(n_266),
.B2(n_273),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_574),
.B(n_432),
.Y(n_698)
);

NAND3xp33_ASAP7_75t_SL g699 ( 
.A(n_549),
.B(n_197),
.C(n_191),
.Y(n_699)
);

A2O1A1Ixp33_ASAP7_75t_L g700 ( 
.A1(n_584),
.A2(n_438),
.B(n_437),
.C(n_436),
.Y(n_700)
);

INVx3_ASAP7_75t_L g701 ( 
.A(n_520),
.Y(n_701)
);

A2O1A1Ixp33_ASAP7_75t_L g702 ( 
.A1(n_594),
.A2(n_436),
.B(n_432),
.C(n_335),
.Y(n_702)
);

CKINVDCx10_ASAP7_75t_R g703 ( 
.A(n_589),
.Y(n_703)
);

NOR2xp33_ASAP7_75t_L g704 ( 
.A(n_534),
.B(n_200),
.Y(n_704)
);

NOR2xp33_ASAP7_75t_L g705 ( 
.A(n_534),
.B(n_202),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_600),
.Y(n_706)
);

HB1xp67_ASAP7_75t_L g707 ( 
.A(n_585),
.Y(n_707)
);

AOI21xp5_ASAP7_75t_L g708 ( 
.A1(n_552),
.A2(n_280),
.B(n_255),
.Y(n_708)
);

OAI21xp5_ASAP7_75t_L g709 ( 
.A1(n_613),
.A2(n_417),
.B(n_409),
.Y(n_709)
);

BUFx12f_ASAP7_75t_L g710 ( 
.A(n_627),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_665),
.Y(n_711)
);

AOI21x1_ASAP7_75t_L g712 ( 
.A1(n_641),
.A2(n_530),
.B(n_554),
.Y(n_712)
);

AOI21xp5_ASAP7_75t_L g713 ( 
.A1(n_648),
.A2(n_577),
.B(n_579),
.Y(n_713)
);

INVx5_ASAP7_75t_L g714 ( 
.A(n_638),
.Y(n_714)
);

AOI21xp5_ASAP7_75t_L g715 ( 
.A1(n_650),
.A2(n_588),
.B(n_581),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_SL g716 ( 
.A(n_643),
.B(n_536),
.Y(n_716)
);

AOI21xp5_ASAP7_75t_L g717 ( 
.A1(n_637),
.A2(n_530),
.B(n_554),
.Y(n_717)
);

AOI21xp5_ASAP7_75t_L g718 ( 
.A1(n_664),
.A2(n_603),
.B(n_595),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_617),
.B(n_564),
.Y(n_719)
);

OAI22xp5_ASAP7_75t_L g720 ( 
.A1(n_617),
.A2(n_604),
.B1(n_601),
.B2(n_563),
.Y(n_720)
);

NOR2xp33_ASAP7_75t_L g721 ( 
.A(n_644),
.B(n_560),
.Y(n_721)
);

AOI21xp5_ASAP7_75t_L g722 ( 
.A1(n_675),
.A2(n_603),
.B(n_595),
.Y(n_722)
);

O2A1O1Ixp33_ASAP7_75t_L g723 ( 
.A1(n_647),
.A2(n_541),
.B(n_529),
.C(n_571),
.Y(n_723)
);

INVx1_ASAP7_75t_SL g724 ( 
.A(n_703),
.Y(n_724)
);

AND2x2_ASAP7_75t_L g725 ( 
.A(n_628),
.B(n_327),
.Y(n_725)
);

NOR2xp33_ASAP7_75t_L g726 ( 
.A(n_647),
.B(n_571),
.Y(n_726)
);

NOR2xp33_ASAP7_75t_L g727 ( 
.A(n_688),
.B(n_576),
.Y(n_727)
);

AOI21xp5_ASAP7_75t_L g728 ( 
.A1(n_616),
.A2(n_607),
.B(n_598),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_662),
.B(n_576),
.Y(n_729)
);

INVx5_ASAP7_75t_L g730 ( 
.A(n_638),
.Y(n_730)
);

OR2x2_ASAP7_75t_L g731 ( 
.A(n_621),
.B(n_519),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_662),
.B(n_536),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_620),
.Y(n_733)
);

INVx3_ASAP7_75t_L g734 ( 
.A(n_638),
.Y(n_734)
);

O2A1O1Ixp5_ASAP7_75t_L g735 ( 
.A1(n_679),
.A2(n_519),
.B(n_567),
.C(n_417),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_652),
.B(n_612),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_680),
.B(n_592),
.Y(n_737)
);

INVx4_ASAP7_75t_L g738 ( 
.A(n_674),
.Y(n_738)
);

AOI21xp5_ASAP7_75t_L g739 ( 
.A1(n_666),
.A2(n_596),
.B(n_593),
.Y(n_739)
);

A2O1A1Ixp33_ASAP7_75t_L g740 ( 
.A1(n_640),
.A2(n_593),
.B(n_592),
.C(n_268),
.Y(n_740)
);

AND2x2_ASAP7_75t_L g741 ( 
.A(n_684),
.B(n_328),
.Y(n_741)
);

OAI22xp5_ASAP7_75t_L g742 ( 
.A1(n_631),
.A2(n_596),
.B1(n_238),
.B2(n_279),
.Y(n_742)
);

HB1xp67_ASAP7_75t_L g743 ( 
.A(n_619),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_640),
.B(n_332),
.Y(n_744)
);

BUFx3_ASAP7_75t_L g745 ( 
.A(n_660),
.Y(n_745)
);

BUFx12f_ASAP7_75t_L g746 ( 
.A(n_638),
.Y(n_746)
);

AOI21xp5_ASAP7_75t_L g747 ( 
.A1(n_666),
.A2(n_196),
.B(n_187),
.Y(n_747)
);

A2O1A1Ixp33_ASAP7_75t_L g748 ( 
.A1(n_631),
.A2(n_420),
.B(n_428),
.C(n_334),
.Y(n_748)
);

NOR3xp33_ASAP7_75t_SL g749 ( 
.A(n_699),
.B(n_209),
.C(n_206),
.Y(n_749)
);

OAI22xp5_ASAP7_75t_L g750 ( 
.A1(n_643),
.A2(n_235),
.B1(n_234),
.B2(n_210),
.Y(n_750)
);

OAI21xp33_ASAP7_75t_L g751 ( 
.A1(n_704),
.A2(n_218),
.B(n_216),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_689),
.B(n_336),
.Y(n_752)
);

A2O1A1Ixp33_ASAP7_75t_L g753 ( 
.A1(n_623),
.A2(n_420),
.B(n_428),
.C(n_344),
.Y(n_753)
);

A2O1A1Ixp33_ASAP7_75t_L g754 ( 
.A1(n_658),
.A2(n_341),
.B(n_342),
.C(n_397),
.Y(n_754)
);

NAND2x1_ASAP7_75t_L g755 ( 
.A(n_663),
.B(n_410),
.Y(n_755)
);

AO21x1_ASAP7_75t_L g756 ( 
.A1(n_659),
.A2(n_408),
.B(n_397),
.Y(n_756)
);

BUFx2_ASAP7_75t_SL g757 ( 
.A(n_674),
.Y(n_757)
);

INVxp67_ASAP7_75t_L g758 ( 
.A(n_689),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_668),
.Y(n_759)
);

BUFx6f_ASAP7_75t_L g760 ( 
.A(n_672),
.Y(n_760)
);

BUFx2_ASAP7_75t_L g761 ( 
.A(n_707),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_670),
.B(n_226),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_639),
.Y(n_763)
);

O2A1O1Ixp33_ASAP7_75t_L g764 ( 
.A1(n_658),
.A2(n_427),
.B(n_422),
.C(n_418),
.Y(n_764)
);

O2A1O1Ixp33_ASAP7_75t_L g765 ( 
.A1(n_633),
.A2(n_427),
.B(n_422),
.C(n_418),
.Y(n_765)
);

A2O1A1Ixp33_ASAP7_75t_L g766 ( 
.A1(n_704),
.A2(n_427),
.B(n_397),
.C(n_408),
.Y(n_766)
);

O2A1O1Ixp33_ASAP7_75t_L g767 ( 
.A1(n_634),
.A2(n_422),
.B(n_418),
.C(n_408),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_678),
.B(n_233),
.Y(n_768)
);

AOI21xp5_ASAP7_75t_L g769 ( 
.A1(n_657),
.A2(n_229),
.B(n_204),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_SL g770 ( 
.A(n_672),
.B(n_410),
.Y(n_770)
);

A2O1A1Ixp33_ASAP7_75t_L g771 ( 
.A1(n_705),
.A2(n_263),
.B(n_251),
.C(n_281),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_691),
.Y(n_772)
);

OR2x2_ASAP7_75t_L g773 ( 
.A(n_697),
.B(n_410),
.Y(n_773)
);

O2A1O1Ixp33_ASAP7_75t_L g774 ( 
.A1(n_705),
.A2(n_8),
.B(n_9),
.C(n_11),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_733),
.Y(n_775)
);

AOI21xp5_ASAP7_75t_L g776 ( 
.A1(n_726),
.A2(n_635),
.B(n_625),
.Y(n_776)
);

AO32x2_ASAP7_75t_L g777 ( 
.A1(n_720),
.A2(n_742),
.A3(n_750),
.B1(n_756),
.B2(n_731),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_725),
.B(n_706),
.Y(n_778)
);

INVx8_ASAP7_75t_L g779 ( 
.A(n_746),
.Y(n_779)
);

AOI21xp5_ASAP7_75t_L g780 ( 
.A1(n_726),
.A2(n_635),
.B(n_625),
.Y(n_780)
);

OAI21x1_ASAP7_75t_L g781 ( 
.A1(n_722),
.A2(n_669),
.B(n_636),
.Y(n_781)
);

OAI21xp5_ASAP7_75t_L g782 ( 
.A1(n_727),
.A2(n_661),
.B(n_655),
.Y(n_782)
);

O2A1O1Ixp5_ASAP7_75t_L g783 ( 
.A1(n_727),
.A2(n_630),
.B(n_642),
.C(n_651),
.Y(n_783)
);

OAI21x1_ASAP7_75t_L g784 ( 
.A1(n_728),
.A2(n_632),
.B(n_649),
.Y(n_784)
);

OAI21x1_ASAP7_75t_L g785 ( 
.A1(n_735),
.A2(n_656),
.B(n_645),
.Y(n_785)
);

AOI21xp5_ASAP7_75t_L g786 ( 
.A1(n_713),
.A2(n_651),
.B(n_642),
.Y(n_786)
);

AOI21xp5_ASAP7_75t_L g787 ( 
.A1(n_715),
.A2(n_630),
.B(n_622),
.Y(n_787)
);

AO31x2_ASAP7_75t_L g788 ( 
.A1(n_718),
.A2(n_687),
.A3(n_700),
.B(n_702),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_721),
.B(n_626),
.Y(n_789)
);

OAI21x1_ASAP7_75t_L g790 ( 
.A1(n_735),
.A2(n_629),
.B(n_615),
.Y(n_790)
);

A2O1A1Ixp33_ASAP7_75t_L g791 ( 
.A1(n_723),
.A2(n_614),
.B(n_653),
.C(n_682),
.Y(n_791)
);

AOI22xp33_ASAP7_75t_L g792 ( 
.A1(n_721),
.A2(n_695),
.B1(n_681),
.B2(n_693),
.Y(n_792)
);

INVx3_ASAP7_75t_L g793 ( 
.A(n_738),
.Y(n_793)
);

OR2x2_ASAP7_75t_L g794 ( 
.A(n_736),
.B(n_654),
.Y(n_794)
);

OAI21x1_ASAP7_75t_L g795 ( 
.A1(n_717),
.A2(n_624),
.B(n_667),
.Y(n_795)
);

OAI21x1_ASAP7_75t_L g796 ( 
.A1(n_712),
.A2(n_673),
.B(n_709),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_744),
.B(n_692),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_711),
.Y(n_798)
);

AND2x2_ASAP7_75t_L g799 ( 
.A(n_741),
.B(n_663),
.Y(n_799)
);

BUFx8_ASAP7_75t_L g800 ( 
.A(n_710),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_763),
.Y(n_801)
);

AOI21xp5_ASAP7_75t_L g802 ( 
.A1(n_739),
.A2(n_671),
.B(n_729),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_SL g803 ( 
.A(n_758),
.B(n_672),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_772),
.Y(n_804)
);

INVxp67_ASAP7_75t_L g805 ( 
.A(n_761),
.Y(n_805)
);

OAI21x1_ASAP7_75t_L g806 ( 
.A1(n_765),
.A2(n_673),
.B(n_685),
.Y(n_806)
);

AOI21x1_ASAP7_75t_L g807 ( 
.A1(n_716),
.A2(n_686),
.B(n_696),
.Y(n_807)
);

BUFx8_ASAP7_75t_L g808 ( 
.A(n_760),
.Y(n_808)
);

O2A1O1Ixp33_ASAP7_75t_SL g809 ( 
.A1(n_774),
.A2(n_687),
.B(n_700),
.C(n_702),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_762),
.B(n_768),
.Y(n_810)
);

O2A1O1Ixp33_ASAP7_75t_L g811 ( 
.A1(n_771),
.A2(n_708),
.B(n_683),
.C(n_698),
.Y(n_811)
);

HB1xp67_ASAP7_75t_L g812 ( 
.A(n_743),
.Y(n_812)
);

INVxp67_ASAP7_75t_SL g813 ( 
.A(n_743),
.Y(n_813)
);

AND2x4_ASAP7_75t_L g814 ( 
.A(n_714),
.B(n_674),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_719),
.B(n_701),
.Y(n_815)
);

O2A1O1Ixp33_ASAP7_75t_L g816 ( 
.A1(n_751),
.A2(n_694),
.B(n_646),
.C(n_618),
.Y(n_816)
);

OAI21x1_ASAP7_75t_L g817 ( 
.A1(n_767),
.A2(n_676),
.B(n_685),
.Y(n_817)
);

CKINVDCx11_ASAP7_75t_R g818 ( 
.A(n_724),
.Y(n_818)
);

OAI21xp5_ASAP7_75t_L g819 ( 
.A1(n_758),
.A2(n_701),
.B(n_677),
.Y(n_819)
);

CKINVDCx20_ASAP7_75t_R g820 ( 
.A(n_745),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_759),
.Y(n_821)
);

CKINVDCx20_ASAP7_75t_R g822 ( 
.A(n_749),
.Y(n_822)
);

AND2x2_ASAP7_75t_L g823 ( 
.A(n_732),
.B(n_13),
.Y(n_823)
);

OAI21x1_ASAP7_75t_L g824 ( 
.A1(n_770),
.A2(n_674),
.B(n_672),
.Y(n_824)
);

AOI21xp5_ASAP7_75t_L g825 ( 
.A1(n_770),
.A2(n_690),
.B(n_282),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_754),
.Y(n_826)
);

AND2x4_ASAP7_75t_L g827 ( 
.A(n_714),
.B(n_690),
.Y(n_827)
);

INVx4_ASAP7_75t_L g828 ( 
.A(n_714),
.Y(n_828)
);

OA22x2_ASAP7_75t_L g829 ( 
.A1(n_737),
.A2(n_282),
.B1(n_281),
.B2(n_280),
.Y(n_829)
);

CKINVDCx5p33_ASAP7_75t_R g830 ( 
.A(n_800),
.Y(n_830)
);

INVx6_ASAP7_75t_L g831 ( 
.A(n_808),
.Y(n_831)
);

AOI22xp33_ASAP7_75t_SL g832 ( 
.A1(n_829),
.A2(n_752),
.B1(n_769),
.B2(n_747),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_778),
.B(n_789),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_775),
.Y(n_834)
);

AOI22xp5_ASAP7_75t_L g835 ( 
.A1(n_822),
.A2(n_716),
.B1(n_749),
.B2(n_740),
.Y(n_835)
);

CKINVDCx20_ASAP7_75t_R g836 ( 
.A(n_818),
.Y(n_836)
);

BUFx12f_ASAP7_75t_L g837 ( 
.A(n_818),
.Y(n_837)
);

AOI22xp33_ASAP7_75t_L g838 ( 
.A1(n_829),
.A2(n_773),
.B1(n_690),
.B2(n_411),
.Y(n_838)
);

CKINVDCx11_ASAP7_75t_R g839 ( 
.A(n_820),
.Y(n_839)
);

CKINVDCx20_ASAP7_75t_R g840 ( 
.A(n_800),
.Y(n_840)
);

AND2x2_ASAP7_75t_L g841 ( 
.A(n_799),
.B(n_16),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_801),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_798),
.Y(n_843)
);

BUFx12f_ASAP7_75t_L g844 ( 
.A(n_800),
.Y(n_844)
);

AOI22xp33_ASAP7_75t_L g845 ( 
.A1(n_810),
.A2(n_690),
.B1(n_425),
.B2(n_426),
.Y(n_845)
);

AOI22xp33_ASAP7_75t_L g846 ( 
.A1(n_782),
.A2(n_411),
.B1(n_425),
.B2(n_426),
.Y(n_846)
);

OAI22xp33_ASAP7_75t_L g847 ( 
.A1(n_797),
.A2(n_730),
.B1(n_714),
.B2(n_738),
.Y(n_847)
);

OAI22xp5_ASAP7_75t_L g848 ( 
.A1(n_805),
.A2(n_748),
.B1(n_753),
.B2(n_734),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_804),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_794),
.B(n_734),
.Y(n_850)
);

AOI22xp33_ASAP7_75t_L g851 ( 
.A1(n_822),
.A2(n_410),
.B1(n_411),
.B2(n_425),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_821),
.Y(n_852)
);

BUFx4f_ASAP7_75t_SL g853 ( 
.A(n_820),
.Y(n_853)
);

INVx2_ASAP7_75t_L g854 ( 
.A(n_798),
.Y(n_854)
);

AOI22xp33_ASAP7_75t_L g855 ( 
.A1(n_826),
.A2(n_410),
.B1(n_411),
.B2(n_425),
.Y(n_855)
);

AOI22xp33_ASAP7_75t_L g856 ( 
.A1(n_812),
.A2(n_410),
.B1(n_411),
.B2(n_425),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_812),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_813),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_823),
.B(n_730),
.Y(n_859)
);

CKINVDCx11_ASAP7_75t_R g860 ( 
.A(n_779),
.Y(n_860)
);

OAI22xp5_ASAP7_75t_L g861 ( 
.A1(n_791),
.A2(n_730),
.B1(n_755),
.B2(n_757),
.Y(n_861)
);

BUFx10_ASAP7_75t_L g862 ( 
.A(n_814),
.Y(n_862)
);

INVx2_ASAP7_75t_SL g863 ( 
.A(n_779),
.Y(n_863)
);

OAI22xp33_ASAP7_75t_L g864 ( 
.A1(n_815),
.A2(n_730),
.B1(n_760),
.B2(n_255),
.Y(n_864)
);

AOI22xp33_ASAP7_75t_L g865 ( 
.A1(n_792),
.A2(n_410),
.B1(n_426),
.B2(n_425),
.Y(n_865)
);

CKINVDCx6p67_ASAP7_75t_R g866 ( 
.A(n_779),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_803),
.Y(n_867)
);

INVx3_ASAP7_75t_SL g868 ( 
.A(n_827),
.Y(n_868)
);

INVx6_ASAP7_75t_L g869 ( 
.A(n_808),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_803),
.Y(n_870)
);

OAI22xp5_ASAP7_75t_L g871 ( 
.A1(n_791),
.A2(n_776),
.B1(n_780),
.B2(n_792),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_808),
.B(n_760),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_819),
.Y(n_873)
);

BUFx6f_ASAP7_75t_L g874 ( 
.A(n_814),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_827),
.B(n_760),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_796),
.Y(n_876)
);

AOI22xp33_ASAP7_75t_SL g877 ( 
.A1(n_777),
.A2(n_199),
.B1(n_184),
.B2(n_228),
.Y(n_877)
);

CKINVDCx5p33_ASAP7_75t_R g878 ( 
.A(n_827),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_788),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_788),
.Y(n_880)
);

AOI22xp33_ASAP7_75t_L g881 ( 
.A1(n_802),
.A2(n_411),
.B1(n_426),
.B2(n_425),
.Y(n_881)
);

INVx4_ASAP7_75t_L g882 ( 
.A(n_814),
.Y(n_882)
);

CKINVDCx5p33_ASAP7_75t_R g883 ( 
.A(n_793),
.Y(n_883)
);

AOI22xp5_ASAP7_75t_L g884 ( 
.A1(n_828),
.A2(n_236),
.B1(n_190),
.B2(n_192),
.Y(n_884)
);

OAI22xp5_ASAP7_75t_L g885 ( 
.A1(n_811),
.A2(n_766),
.B1(n_764),
.B2(n_243),
.Y(n_885)
);

AOI22xp33_ASAP7_75t_SL g886 ( 
.A1(n_777),
.A2(n_199),
.B1(n_188),
.B2(n_278),
.Y(n_886)
);

OAI22xp33_ASAP7_75t_L g887 ( 
.A1(n_828),
.A2(n_225),
.B1(n_203),
.B2(n_277),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_879),
.Y(n_888)
);

INVx2_ASAP7_75t_L g889 ( 
.A(n_876),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_880),
.Y(n_890)
);

BUFx2_ASAP7_75t_L g891 ( 
.A(n_876),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_880),
.Y(n_892)
);

OAI21x1_ASAP7_75t_L g893 ( 
.A1(n_871),
.A2(n_781),
.B(n_790),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_834),
.Y(n_894)
);

AND2x2_ASAP7_75t_L g895 ( 
.A(n_857),
.B(n_777),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_867),
.Y(n_896)
);

OAI21x1_ASAP7_75t_L g897 ( 
.A1(n_881),
.A2(n_790),
.B(n_784),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_843),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_842),
.Y(n_899)
);

INVx3_ASAP7_75t_L g900 ( 
.A(n_870),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_843),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_849),
.Y(n_902)
);

AO31x2_ASAP7_75t_L g903 ( 
.A1(n_873),
.A2(n_787),
.A3(n_786),
.B(n_777),
.Y(n_903)
);

HB1xp67_ASAP7_75t_L g904 ( 
.A(n_858),
.Y(n_904)
);

HB1xp67_ASAP7_75t_L g905 ( 
.A(n_850),
.Y(n_905)
);

OR2x2_ASAP7_75t_L g906 ( 
.A(n_833),
.B(n_788),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_854),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_854),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_852),
.Y(n_909)
);

INVx1_ASAP7_75t_SL g910 ( 
.A(n_859),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_877),
.B(n_788),
.Y(n_911)
);

OA21x2_ASAP7_75t_L g912 ( 
.A1(n_881),
.A2(n_785),
.B(n_784),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_874),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_886),
.B(n_793),
.Y(n_914)
);

AND2x4_ASAP7_75t_L g915 ( 
.A(n_874),
.B(n_824),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_875),
.Y(n_916)
);

BUFx6f_ASAP7_75t_L g917 ( 
.A(n_874),
.Y(n_917)
);

HB1xp67_ASAP7_75t_L g918 ( 
.A(n_848),
.Y(n_918)
);

AO31x2_ASAP7_75t_L g919 ( 
.A1(n_861),
.A2(n_825),
.A3(n_809),
.B(n_783),
.Y(n_919)
);

NOR2x1p5_ASAP7_75t_L g920 ( 
.A(n_844),
.B(n_807),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_847),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_874),
.Y(n_922)
);

INVx2_ASAP7_75t_L g923 ( 
.A(n_862),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_832),
.Y(n_924)
);

BUFx2_ASAP7_75t_L g925 ( 
.A(n_883),
.Y(n_925)
);

OR2x2_ASAP7_75t_L g926 ( 
.A(n_905),
.B(n_841),
.Y(n_926)
);

AO32x2_ASAP7_75t_L g927 ( 
.A1(n_905),
.A2(n_904),
.A3(n_910),
.B1(n_895),
.B2(n_906),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_904),
.Y(n_928)
);

NOR2x1_ASAP7_75t_SL g929 ( 
.A(n_917),
.B(n_844),
.Y(n_929)
);

AOI21xp5_ASAP7_75t_SL g930 ( 
.A1(n_920),
.A2(n_882),
.B(n_872),
.Y(n_930)
);

NOR2xp33_ASAP7_75t_L g931 ( 
.A(n_918),
.B(n_835),
.Y(n_931)
);

OR2x6_ASAP7_75t_L g932 ( 
.A(n_920),
.B(n_831),
.Y(n_932)
);

NOR2x1_ASAP7_75t_SL g933 ( 
.A(n_917),
.B(n_837),
.Y(n_933)
);

AND2x2_ASAP7_75t_L g934 ( 
.A(n_895),
.B(n_838),
.Y(n_934)
);

AOI22xp33_ASAP7_75t_L g935 ( 
.A1(n_918),
.A2(n_838),
.B1(n_851),
.B2(n_865),
.Y(n_935)
);

AND2x2_ASAP7_75t_L g936 ( 
.A(n_895),
.B(n_882),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_910),
.B(n_846),
.Y(n_937)
);

OR2x2_ASAP7_75t_L g938 ( 
.A(n_906),
.B(n_868),
.Y(n_938)
);

OAI21xp5_ASAP7_75t_L g939 ( 
.A1(n_924),
.A2(n_884),
.B(n_846),
.Y(n_939)
);

AND2x4_ASAP7_75t_L g940 ( 
.A(n_915),
.B(n_878),
.Y(n_940)
);

AND2x2_ASAP7_75t_L g941 ( 
.A(n_925),
.B(n_868),
.Y(n_941)
);

NOR2xp33_ASAP7_75t_L g942 ( 
.A(n_925),
.B(n_837),
.Y(n_942)
);

NOR2xp33_ASAP7_75t_L g943 ( 
.A(n_925),
.B(n_900),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_894),
.B(n_845),
.Y(n_944)
);

AND2x2_ASAP7_75t_L g945 ( 
.A(n_894),
.B(n_817),
.Y(n_945)
);

HB1xp67_ASAP7_75t_L g946 ( 
.A(n_900),
.Y(n_946)
);

OR2x2_ASAP7_75t_L g947 ( 
.A(n_906),
.B(n_863),
.Y(n_947)
);

AND2x2_ASAP7_75t_L g948 ( 
.A(n_917),
.B(n_839),
.Y(n_948)
);

OR2x2_ASAP7_75t_L g949 ( 
.A(n_916),
.B(n_845),
.Y(n_949)
);

AO32x1_ASAP7_75t_L g950 ( 
.A1(n_924),
.A2(n_885),
.A3(n_809),
.B1(n_865),
.B2(n_855),
.Y(n_950)
);

OR2x2_ASAP7_75t_L g951 ( 
.A(n_916),
.B(n_866),
.Y(n_951)
);

AOI221x1_ASAP7_75t_SL g952 ( 
.A1(n_924),
.A2(n_16),
.B1(n_17),
.B2(n_19),
.C(n_20),
.Y(n_952)
);

NAND4xp25_ASAP7_75t_L g953 ( 
.A(n_894),
.B(n_899),
.C(n_902),
.D(n_900),
.Y(n_953)
);

AND2x2_ASAP7_75t_L g954 ( 
.A(n_899),
.B(n_902),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_899),
.Y(n_955)
);

AOI22xp5_ASAP7_75t_L g956 ( 
.A1(n_921),
.A2(n_851),
.B1(n_864),
.B2(n_840),
.Y(n_956)
);

OR2x6_ASAP7_75t_L g957 ( 
.A(n_915),
.B(n_831),
.Y(n_957)
);

A2O1A1Ixp33_ASAP7_75t_L g958 ( 
.A1(n_911),
.A2(n_816),
.B(n_855),
.C(n_817),
.Y(n_958)
);

AND2x2_ASAP7_75t_L g959 ( 
.A(n_902),
.B(n_795),
.Y(n_959)
);

INVx3_ASAP7_75t_L g960 ( 
.A(n_900),
.Y(n_960)
);

AOI221xp5_ASAP7_75t_L g961 ( 
.A1(n_911),
.A2(n_887),
.B1(n_199),
.B2(n_244),
.C(n_207),
.Y(n_961)
);

AO21x2_ASAP7_75t_L g962 ( 
.A1(n_914),
.A2(n_806),
.B(n_856),
.Y(n_962)
);

OAI22xp5_ASAP7_75t_L g963 ( 
.A1(n_914),
.A2(n_869),
.B1(n_831),
.B2(n_853),
.Y(n_963)
);

AO21x2_ASAP7_75t_L g964 ( 
.A1(n_889),
.A2(n_856),
.B(n_862),
.Y(n_964)
);

INVx4_ASAP7_75t_L g965 ( 
.A(n_917),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_954),
.Y(n_966)
);

AOI221xp5_ASAP7_75t_L g967 ( 
.A1(n_952),
.A2(n_909),
.B1(n_896),
.B2(n_888),
.C(n_921),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_928),
.B(n_896),
.Y(n_968)
);

INVxp67_ASAP7_75t_L g969 ( 
.A(n_943),
.Y(n_969)
);

AND2x2_ASAP7_75t_L g970 ( 
.A(n_936),
.B(n_900),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_954),
.B(n_955),
.Y(n_971)
);

AND2x2_ASAP7_75t_L g972 ( 
.A(n_936),
.B(n_909),
.Y(n_972)
);

BUFx2_ASAP7_75t_L g973 ( 
.A(n_946),
.Y(n_973)
);

BUFx2_ASAP7_75t_L g974 ( 
.A(n_960),
.Y(n_974)
);

AND2x2_ASAP7_75t_L g975 ( 
.A(n_943),
.B(n_909),
.Y(n_975)
);

AND2x4_ASAP7_75t_L g976 ( 
.A(n_940),
.B(n_915),
.Y(n_976)
);

AND2x2_ASAP7_75t_L g977 ( 
.A(n_927),
.B(n_891),
.Y(n_977)
);

AOI22xp33_ASAP7_75t_L g978 ( 
.A1(n_931),
.A2(n_921),
.B1(n_888),
.B2(n_890),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_927),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_927),
.Y(n_980)
);

AND2x2_ASAP7_75t_SL g981 ( 
.A(n_940),
.B(n_917),
.Y(n_981)
);

OR2x2_ASAP7_75t_L g982 ( 
.A(n_926),
.B(n_888),
.Y(n_982)
);

AOI22xp33_ASAP7_75t_SL g983 ( 
.A1(n_931),
.A2(n_836),
.B1(n_869),
.B2(n_912),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_927),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_953),
.Y(n_985)
);

AND2x2_ASAP7_75t_L g986 ( 
.A(n_960),
.B(n_891),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_959),
.Y(n_987)
);

AND2x2_ASAP7_75t_L g988 ( 
.A(n_960),
.B(n_891),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_959),
.Y(n_989)
);

AOI22xp5_ASAP7_75t_L g990 ( 
.A1(n_935),
.A2(n_869),
.B1(n_839),
.B2(n_922),
.Y(n_990)
);

NAND2x1p5_ASAP7_75t_L g991 ( 
.A(n_981),
.B(n_965),
.Y(n_991)
);

AOI22xp33_ASAP7_75t_L g992 ( 
.A1(n_983),
.A2(n_939),
.B1(n_934),
.B2(n_961),
.Y(n_992)
);

AOI221xp5_ASAP7_75t_L g993 ( 
.A1(n_967),
.A2(n_934),
.B1(n_935),
.B2(n_958),
.C(n_956),
.Y(n_993)
);

AOI21xp5_ASAP7_75t_L g994 ( 
.A1(n_983),
.A2(n_950),
.B(n_958),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_966),
.Y(n_995)
);

AND2x2_ASAP7_75t_L g996 ( 
.A(n_981),
.B(n_948),
.Y(n_996)
);

INVx2_ASAP7_75t_L g997 ( 
.A(n_977),
.Y(n_997)
);

INVxp67_ASAP7_75t_L g998 ( 
.A(n_985),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_979),
.B(n_945),
.Y(n_999)
);

INVx2_ASAP7_75t_L g1000 ( 
.A(n_977),
.Y(n_1000)
);

AOI221xp5_ASAP7_75t_L g1001 ( 
.A1(n_967),
.A2(n_937),
.B1(n_944),
.B2(n_963),
.C(n_945),
.Y(n_1001)
);

AND2x2_ASAP7_75t_L g1002 ( 
.A(n_981),
.B(n_965),
.Y(n_1002)
);

INVx4_ASAP7_75t_L g1003 ( 
.A(n_976),
.Y(n_1003)
);

HB1xp67_ASAP7_75t_L g1004 ( 
.A(n_985),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_966),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_968),
.Y(n_1006)
);

INVxp67_ASAP7_75t_SL g1007 ( 
.A(n_979),
.Y(n_1007)
);

INVx2_ASAP7_75t_L g1008 ( 
.A(n_987),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_968),
.Y(n_1009)
);

INVxp67_ASAP7_75t_SL g1010 ( 
.A(n_980),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_987),
.Y(n_1011)
);

INVx2_ASAP7_75t_L g1012 ( 
.A(n_1008),
.Y(n_1012)
);

AND2x4_ASAP7_75t_L g1013 ( 
.A(n_1003),
.B(n_976),
.Y(n_1013)
);

INVx2_ASAP7_75t_L g1014 ( 
.A(n_1008),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_995),
.Y(n_1015)
);

AND2x2_ASAP7_75t_L g1016 ( 
.A(n_1003),
.B(n_969),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_995),
.Y(n_1017)
);

INVx2_ASAP7_75t_L g1018 ( 
.A(n_1008),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_998),
.B(n_975),
.Y(n_1019)
);

NOR3xp33_ASAP7_75t_SL g1020 ( 
.A(n_1001),
.B(n_830),
.C(n_942),
.Y(n_1020)
);

INVx2_ASAP7_75t_L g1021 ( 
.A(n_997),
.Y(n_1021)
);

AND2x2_ASAP7_75t_L g1022 ( 
.A(n_1003),
.B(n_972),
.Y(n_1022)
);

OR2x2_ASAP7_75t_L g1023 ( 
.A(n_1019),
.B(n_998),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_1015),
.Y(n_1024)
);

AND2x4_ASAP7_75t_L g1025 ( 
.A(n_1013),
.B(n_1003),
.Y(n_1025)
);

INVx2_ASAP7_75t_L g1026 ( 
.A(n_1021),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_1015),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_1017),
.Y(n_1028)
);

AND2x2_ASAP7_75t_L g1029 ( 
.A(n_1016),
.B(n_1004),
.Y(n_1029)
);

AND2x2_ASAP7_75t_L g1030 ( 
.A(n_1029),
.B(n_1016),
.Y(n_1030)
);

OR2x2_ASAP7_75t_L g1031 ( 
.A(n_1023),
.B(n_999),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_1029),
.B(n_1001),
.Y(n_1032)
);

HB1xp67_ASAP7_75t_L g1033 ( 
.A(n_1023),
.Y(n_1033)
);

HB1xp67_ASAP7_75t_L g1034 ( 
.A(n_1033),
.Y(n_1034)
);

INVx2_ASAP7_75t_L g1035 ( 
.A(n_1030),
.Y(n_1035)
);

AOI21xp33_ASAP7_75t_L g1036 ( 
.A1(n_1032),
.A2(n_1026),
.B(n_1024),
.Y(n_1036)
);

OAI22xp5_ASAP7_75t_L g1037 ( 
.A1(n_1031),
.A2(n_1020),
.B1(n_993),
.B2(n_992),
.Y(n_1037)
);

AND2x2_ASAP7_75t_L g1038 ( 
.A(n_1030),
.B(n_1025),
.Y(n_1038)
);

OAI22xp5_ASAP7_75t_L g1039 ( 
.A1(n_1032),
.A2(n_993),
.B1(n_1025),
.B2(n_994),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_1033),
.B(n_1028),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_1033),
.Y(n_1041)
);

NAND2xp33_ASAP7_75t_SL g1042 ( 
.A(n_1032),
.B(n_1025),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_1033),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_1033),
.B(n_1024),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_SL g1045 ( 
.A(n_1034),
.B(n_1027),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_SL g1046 ( 
.A(n_1034),
.B(n_1027),
.Y(n_1046)
);

OAI21xp33_ASAP7_75t_L g1047 ( 
.A1(n_1035),
.A2(n_994),
.B(n_1007),
.Y(n_1047)
);

INVxp67_ASAP7_75t_SL g1048 ( 
.A(n_1041),
.Y(n_1048)
);

AND2x2_ASAP7_75t_L g1049 ( 
.A(n_1038),
.B(n_1013),
.Y(n_1049)
);

AOI21xp33_ASAP7_75t_L g1050 ( 
.A1(n_1039),
.A2(n_1026),
.B(n_1010),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_1035),
.B(n_1043),
.Y(n_1051)
);

OAI22xp33_ASAP7_75t_L g1052 ( 
.A1(n_1037),
.A2(n_980),
.B1(n_984),
.B2(n_990),
.Y(n_1052)
);

INVx2_ASAP7_75t_L g1053 ( 
.A(n_1044),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_1040),
.Y(n_1054)
);

INVx2_ASAP7_75t_L g1055 ( 
.A(n_1036),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_1042),
.B(n_1007),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_1034),
.Y(n_1057)
);

OAI211xp5_ASAP7_75t_L g1058 ( 
.A1(n_1042),
.A2(n_860),
.B(n_942),
.C(n_1010),
.Y(n_1058)
);

OAI221xp5_ASAP7_75t_L g1059 ( 
.A1(n_1039),
.A2(n_984),
.B1(n_990),
.B2(n_1021),
.C(n_997),
.Y(n_1059)
);

OAI31xp33_ASAP7_75t_L g1060 ( 
.A1(n_1039),
.A2(n_997),
.A3(n_1000),
.B(n_1014),
.Y(n_1060)
);

OAI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_1047),
.A2(n_1014),
.B(n_1012),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_1057),
.Y(n_1062)
);

OAI22xp5_ASAP7_75t_L g1063 ( 
.A1(n_1056),
.A2(n_1013),
.B1(n_991),
.B2(n_1017),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_1048),
.Y(n_1064)
);

XNOR2x1_ASAP7_75t_L g1065 ( 
.A(n_1055),
.B(n_932),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_1053),
.B(n_1055),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_1051),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_1045),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_1053),
.B(n_1006),
.Y(n_1069)
);

AO22x2_ASAP7_75t_L g1070 ( 
.A1(n_1054),
.A2(n_1018),
.B1(n_1012),
.B2(n_1000),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_1045),
.B(n_1006),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_1046),
.B(n_1009),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_1046),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_1049),
.Y(n_1074)
);

AOI321xp33_ASAP7_75t_L g1075 ( 
.A1(n_1052),
.A2(n_978),
.A3(n_1000),
.B1(n_1018),
.B2(n_999),
.C(n_951),
.Y(n_1075)
);

AND2x2_ASAP7_75t_L g1076 ( 
.A(n_1049),
.B(n_1058),
.Y(n_1076)
);

INVxp67_ASAP7_75t_L g1077 ( 
.A(n_1059),
.Y(n_1077)
);

OAI22xp5_ASAP7_75t_SL g1078 ( 
.A1(n_1050),
.A2(n_991),
.B1(n_932),
.B2(n_1009),
.Y(n_1078)
);

OR2x2_ASAP7_75t_L g1079 ( 
.A(n_1060),
.B(n_1005),
.Y(n_1079)
);

NAND3xp33_ASAP7_75t_L g1080 ( 
.A(n_1068),
.B(n_1022),
.C(n_947),
.Y(n_1080)
);

NOR2xp33_ASAP7_75t_SL g1081 ( 
.A(n_1074),
.B(n_991),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_1064),
.Y(n_1082)
);

AOI221xp5_ASAP7_75t_L g1083 ( 
.A1(n_1066),
.A2(n_1011),
.B1(n_962),
.B2(n_1005),
.C(n_982),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_1067),
.B(n_1022),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_1073),
.B(n_975),
.Y(n_1085)
);

NOR3xp33_ASAP7_75t_L g1086 ( 
.A(n_1062),
.B(n_982),
.C(n_1002),
.Y(n_1086)
);

OAI22xp33_ASAP7_75t_L g1087 ( 
.A1(n_1077),
.A2(n_1079),
.B1(n_1061),
.B2(n_1072),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_SL g1088 ( 
.A(n_1076),
.B(n_991),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_1069),
.Y(n_1089)
);

INVxp67_ASAP7_75t_L g1090 ( 
.A(n_1065),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_1071),
.B(n_1011),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_1070),
.Y(n_1092)
);

NOR4xp25_ASAP7_75t_L g1093 ( 
.A(n_1075),
.B(n_1002),
.C(n_996),
.D(n_971),
.Y(n_1093)
);

AOI222xp33_ASAP7_75t_L g1094 ( 
.A1(n_1070),
.A2(n_950),
.B1(n_933),
.B2(n_929),
.C1(n_199),
.C2(n_996),
.Y(n_1094)
);

AOI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_1078),
.A2(n_950),
.B(n_930),
.Y(n_1095)
);

AOI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_1078),
.A2(n_950),
.B(n_971),
.Y(n_1096)
);

AOI221x1_ASAP7_75t_L g1097 ( 
.A1(n_1082),
.A2(n_1063),
.B1(n_21),
.B2(n_22),
.C(n_23),
.Y(n_1097)
);

NAND5xp2_ASAP7_75t_L g1098 ( 
.A(n_1089),
.B(n_1081),
.C(n_1084),
.D(n_1090),
.E(n_1092),
.Y(n_1098)
);

AOI221xp5_ASAP7_75t_L g1099 ( 
.A1(n_1087),
.A2(n_962),
.B1(n_989),
.B2(n_972),
.C(n_964),
.Y(n_1099)
);

AOI21xp5_ASAP7_75t_L g1100 ( 
.A1(n_1088),
.A2(n_941),
.B(n_932),
.Y(n_1100)
);

BUFx3_ASAP7_75t_L g1101 ( 
.A(n_1085),
.Y(n_1101)
);

OAI221xp5_ASAP7_75t_L g1102 ( 
.A1(n_1093),
.A2(n_1096),
.B1(n_1095),
.B2(n_1094),
.C(n_1083),
.Y(n_1102)
);

NOR2xp33_ASAP7_75t_R g1103 ( 
.A(n_1091),
.B(n_17),
.Y(n_1103)
);

AOI21xp33_ASAP7_75t_L g1104 ( 
.A1(n_1080),
.A2(n_949),
.B(n_217),
.Y(n_1104)
);

AOI22xp5_ASAP7_75t_L g1105 ( 
.A1(n_1086),
.A2(n_932),
.B1(n_976),
.B2(n_940),
.Y(n_1105)
);

OAI221xp5_ASAP7_75t_SL g1106 ( 
.A1(n_1093),
.A2(n_989),
.B1(n_957),
.B2(n_938),
.C(n_970),
.Y(n_1106)
);

AOI222xp33_ASAP7_75t_L g1107 ( 
.A1(n_1092),
.A2(n_199),
.B1(n_973),
.B2(n_893),
.C1(n_224),
.C2(n_219),
.Y(n_1107)
);

NOR2xp33_ASAP7_75t_R g1108 ( 
.A(n_1082),
.B(n_23),
.Y(n_1108)
);

O2A1O1Ixp33_ASAP7_75t_L g1109 ( 
.A1(n_1087),
.A2(n_24),
.B(n_25),
.C(n_26),
.Y(n_1109)
);

AOI211xp5_ASAP7_75t_L g1110 ( 
.A1(n_1087),
.A2(n_976),
.B(n_988),
.C(n_986),
.Y(n_1110)
);

NOR2xp33_ASAP7_75t_SL g1111 ( 
.A(n_1082),
.B(n_973),
.Y(n_1111)
);

O2A1O1Ixp5_ASAP7_75t_SL g1112 ( 
.A1(n_1082),
.A2(n_25),
.B(n_26),
.C(n_28),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_1092),
.Y(n_1113)
);

NOR2xp33_ASAP7_75t_R g1114 ( 
.A(n_1082),
.B(n_29),
.Y(n_1114)
);

O2A1O1Ixp33_ASAP7_75t_L g1115 ( 
.A1(n_1087),
.A2(n_29),
.B(n_30),
.C(n_31),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_1092),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_1089),
.B(n_974),
.Y(n_1117)
);

A2O1A1Ixp33_ASAP7_75t_L g1118 ( 
.A1(n_1096),
.A2(n_893),
.B(n_897),
.C(n_970),
.Y(n_1118)
);

AOI21xp33_ASAP7_75t_L g1119 ( 
.A1(n_1082),
.A2(n_31),
.B(n_32),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_1089),
.B(n_974),
.Y(n_1120)
);

OAI311xp33_ASAP7_75t_L g1121 ( 
.A1(n_1102),
.A2(n_33),
.A3(n_34),
.B1(n_35),
.C1(n_36),
.Y(n_1121)
);

AOI221xp5_ASAP7_75t_L g1122 ( 
.A1(n_1113),
.A2(n_276),
.B1(n_242),
.B2(n_246),
.C(n_271),
.Y(n_1122)
);

NOR3xp33_ASAP7_75t_L g1123 ( 
.A(n_1098),
.B(n_213),
.C(n_34),
.Y(n_1123)
);

OAI211xp5_ASAP7_75t_L g1124 ( 
.A1(n_1097),
.A2(n_965),
.B(n_35),
.C(n_36),
.Y(n_1124)
);

NAND4xp25_ASAP7_75t_L g1125 ( 
.A(n_1101),
.B(n_986),
.C(n_988),
.D(n_39),
.Y(n_1125)
);

OAI22xp33_ASAP7_75t_L g1126 ( 
.A1(n_1116),
.A2(n_957),
.B1(n_923),
.B2(n_917),
.Y(n_1126)
);

AOI211x1_ASAP7_75t_SL g1127 ( 
.A1(n_1117),
.A2(n_33),
.B(n_38),
.C(n_39),
.Y(n_1127)
);

A2O1A1Ixp33_ASAP7_75t_L g1128 ( 
.A1(n_1109),
.A2(n_893),
.B(n_897),
.C(n_42),
.Y(n_1128)
);

AOI321xp33_ASAP7_75t_L g1129 ( 
.A1(n_1106),
.A2(n_922),
.A3(n_913),
.B1(n_923),
.B2(n_915),
.C(n_889),
.Y(n_1129)
);

A2O1A1Ixp33_ASAP7_75t_L g1130 ( 
.A1(n_1115),
.A2(n_897),
.B(n_41),
.C(n_42),
.Y(n_1130)
);

AOI221xp5_ASAP7_75t_L g1131 ( 
.A1(n_1104),
.A2(n_964),
.B1(n_44),
.B2(n_45),
.C(n_46),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_1108),
.Y(n_1132)
);

INVx2_ASAP7_75t_L g1133 ( 
.A(n_1120),
.Y(n_1133)
);

OAI221xp5_ASAP7_75t_L g1134 ( 
.A1(n_1118),
.A2(n_1099),
.B1(n_1111),
.B2(n_1107),
.C(n_1119),
.Y(n_1134)
);

AOI21xp5_ASAP7_75t_L g1135 ( 
.A1(n_1119),
.A2(n_38),
.B(n_46),
.Y(n_1135)
);

AOI221xp5_ASAP7_75t_L g1136 ( 
.A1(n_1114),
.A2(n_48),
.B1(n_50),
.B2(n_51),
.C(n_52),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_1103),
.B(n_48),
.Y(n_1137)
);

XNOR2x1_ASAP7_75t_L g1138 ( 
.A(n_1112),
.B(n_52),
.Y(n_1138)
);

OAI311xp33_ASAP7_75t_L g1139 ( 
.A1(n_1110),
.A2(n_53),
.A3(n_54),
.B1(n_56),
.C1(n_57),
.Y(n_1139)
);

AOI221xp5_ASAP7_75t_SL g1140 ( 
.A1(n_1100),
.A2(n_54),
.B1(n_56),
.B2(n_57),
.C(n_58),
.Y(n_1140)
);

AOI221xp5_ASAP7_75t_L g1141 ( 
.A1(n_1105),
.A2(n_58),
.B1(n_59),
.B2(n_60),
.C(n_61),
.Y(n_1141)
);

NAND3xp33_ASAP7_75t_SL g1142 ( 
.A(n_1109),
.B(n_60),
.C(n_61),
.Y(n_1142)
);

OAI21xp5_ASAP7_75t_L g1143 ( 
.A1(n_1109),
.A2(n_912),
.B(n_923),
.Y(n_1143)
);

INVx1_ASAP7_75t_SL g1144 ( 
.A(n_1108),
.Y(n_1144)
);

NOR2x1_ASAP7_75t_L g1145 ( 
.A(n_1138),
.B(n_957),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_1137),
.Y(n_1146)
);

NAND4xp75_ASAP7_75t_L g1147 ( 
.A(n_1132),
.B(n_923),
.C(n_912),
.D(n_913),
.Y(n_1147)
);

NAND2x1p5_ASAP7_75t_SL g1148 ( 
.A(n_1133),
.B(n_913),
.Y(n_1148)
);

XOR2xp5_ASAP7_75t_L g1149 ( 
.A(n_1127),
.B(n_64),
.Y(n_1149)
);

AND2x2_ASAP7_75t_L g1150 ( 
.A(n_1123),
.B(n_957),
.Y(n_1150)
);

NAND4xp75_ASAP7_75t_L g1151 ( 
.A(n_1140),
.B(n_1135),
.C(n_1136),
.D(n_1122),
.Y(n_1151)
);

OR2x2_ASAP7_75t_L g1152 ( 
.A(n_1125),
.B(n_903),
.Y(n_1152)
);

OR2x2_ASAP7_75t_L g1153 ( 
.A(n_1124),
.B(n_1144),
.Y(n_1153)
);

NAND4xp75_ASAP7_75t_L g1154 ( 
.A(n_1141),
.B(n_912),
.C(n_66),
.D(n_67),
.Y(n_1154)
);

AND2x4_ASAP7_75t_L g1155 ( 
.A(n_1128),
.B(n_917),
.Y(n_1155)
);

INVx2_ASAP7_75t_L g1156 ( 
.A(n_1134),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_1142),
.Y(n_1157)
);

INVx3_ASAP7_75t_L g1158 ( 
.A(n_1139),
.Y(n_1158)
);

OR2x2_ASAP7_75t_L g1159 ( 
.A(n_1130),
.B(n_903),
.Y(n_1159)
);

XOR2xp5_ASAP7_75t_L g1160 ( 
.A(n_1121),
.B(n_65),
.Y(n_1160)
);

NAND4xp75_ASAP7_75t_L g1161 ( 
.A(n_1143),
.B(n_912),
.C(n_922),
.D(n_913),
.Y(n_1161)
);

AND2x2_ASAP7_75t_L g1162 ( 
.A(n_1143),
.B(n_903),
.Y(n_1162)
);

OR2x2_ASAP7_75t_L g1163 ( 
.A(n_1126),
.B(n_903),
.Y(n_1163)
);

OR2x2_ASAP7_75t_L g1164 ( 
.A(n_1129),
.B(n_903),
.Y(n_1164)
);

NAND3xp33_ASAP7_75t_SL g1165 ( 
.A(n_1131),
.B(n_922),
.C(n_889),
.Y(n_1165)
);

NAND4xp75_ASAP7_75t_L g1166 ( 
.A(n_1132),
.B(n_912),
.C(n_71),
.D(n_74),
.Y(n_1166)
);

AOI22xp5_ASAP7_75t_L g1167 ( 
.A1(n_1123),
.A2(n_917),
.B1(n_915),
.B2(n_889),
.Y(n_1167)
);

NOR3xp33_ASAP7_75t_L g1168 ( 
.A(n_1156),
.B(n_69),
.C(n_79),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_SL g1169 ( 
.A(n_1158),
.B(n_917),
.Y(n_1169)
);

AOI22xp5_ASAP7_75t_L g1170 ( 
.A1(n_1146),
.A2(n_915),
.B1(n_908),
.B2(n_907),
.Y(n_1170)
);

NOR3xp33_ASAP7_75t_SL g1171 ( 
.A(n_1151),
.B(n_84),
.C(n_87),
.Y(n_1171)
);

OR2x2_ASAP7_75t_L g1172 ( 
.A(n_1153),
.B(n_903),
.Y(n_1172)
);

NAND4xp75_ASAP7_75t_L g1173 ( 
.A(n_1157),
.B(n_88),
.C(n_92),
.D(n_93),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_1149),
.Y(n_1174)
);

OR2x6_ASAP7_75t_L g1175 ( 
.A(n_1151),
.B(n_426),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_1160),
.Y(n_1176)
);

INVx2_ASAP7_75t_L g1177 ( 
.A(n_1148),
.Y(n_1177)
);

NOR3xp33_ASAP7_75t_L g1178 ( 
.A(n_1145),
.B(n_1165),
.C(n_1154),
.Y(n_1178)
);

BUFx2_ASAP7_75t_L g1179 ( 
.A(n_1155),
.Y(n_1179)
);

OAI22xp5_ASAP7_75t_L g1180 ( 
.A1(n_1152),
.A2(n_890),
.B1(n_892),
.B2(n_907),
.Y(n_1180)
);

OAI21xp5_ASAP7_75t_L g1181 ( 
.A1(n_1154),
.A2(n_890),
.B(n_892),
.Y(n_1181)
);

AOI21xp5_ASAP7_75t_L g1182 ( 
.A1(n_1159),
.A2(n_426),
.B(n_411),
.Y(n_1182)
);

XNOR2x1_ASAP7_75t_L g1183 ( 
.A(n_1176),
.B(n_1150),
.Y(n_1183)
);

INVx2_ASAP7_75t_SL g1184 ( 
.A(n_1179),
.Y(n_1184)
);

AOI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_1169),
.A2(n_1174),
.B(n_1177),
.Y(n_1185)
);

XNOR2xp5_ASAP7_75t_L g1186 ( 
.A(n_1171),
.B(n_1166),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_1175),
.Y(n_1187)
);

NAND3xp33_ASAP7_75t_SL g1188 ( 
.A(n_1168),
.B(n_1167),
.C(n_1164),
.Y(n_1188)
);

OAI22x1_ASAP7_75t_L g1189 ( 
.A1(n_1172),
.A2(n_1163),
.B1(n_1162),
.B2(n_1147),
.Y(n_1189)
);

NOR2xp33_ASAP7_75t_L g1190 ( 
.A(n_1175),
.B(n_1161),
.Y(n_1190)
);

INVx4_ASAP7_75t_L g1191 ( 
.A(n_1178),
.Y(n_1191)
);

NOR2xp67_ASAP7_75t_SL g1192 ( 
.A(n_1173),
.B(n_426),
.Y(n_1192)
);

AO22x2_ASAP7_75t_L g1193 ( 
.A1(n_1180),
.A2(n_96),
.B1(n_97),
.B2(n_98),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_1182),
.B(n_903),
.Y(n_1194)
);

AOI22xp5_ASAP7_75t_L g1195 ( 
.A1(n_1170),
.A2(n_908),
.B1(n_907),
.B2(n_901),
.Y(n_1195)
);

BUFx2_ASAP7_75t_L g1196 ( 
.A(n_1181),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_1175),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_1184),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_1183),
.Y(n_1199)
);

AOI22xp5_ASAP7_75t_L g1200 ( 
.A1(n_1185),
.A2(n_908),
.B1(n_901),
.B2(n_898),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1196),
.Y(n_1201)
);

NAND4xp25_ASAP7_75t_L g1202 ( 
.A(n_1191),
.B(n_101),
.C(n_102),
.D(n_105),
.Y(n_1202)
);

AOI22xp5_ASAP7_75t_L g1203 ( 
.A1(n_1188),
.A2(n_901),
.B1(n_898),
.B2(n_892),
.Y(n_1203)
);

AOI22xp5_ASAP7_75t_L g1204 ( 
.A1(n_1189),
.A2(n_901),
.B1(n_898),
.B2(n_919),
.Y(n_1204)
);

AOI22xp5_ASAP7_75t_L g1205 ( 
.A1(n_1190),
.A2(n_898),
.B1(n_919),
.B2(n_903),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_1187),
.Y(n_1206)
);

OAI22xp5_ASAP7_75t_L g1207 ( 
.A1(n_1186),
.A2(n_919),
.B1(n_903),
.B2(n_116),
.Y(n_1207)
);

INVx2_ASAP7_75t_L g1208 ( 
.A(n_1198),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_1199),
.B(n_1197),
.Y(n_1209)
);

INVx2_ASAP7_75t_L g1210 ( 
.A(n_1201),
.Y(n_1210)
);

INVx2_ASAP7_75t_L g1211 ( 
.A(n_1206),
.Y(n_1211)
);

XOR2xp5_ASAP7_75t_L g1212 ( 
.A(n_1202),
.B(n_1193),
.Y(n_1212)
);

OAI22xp5_ASAP7_75t_L g1213 ( 
.A1(n_1204),
.A2(n_1194),
.B1(n_1195),
.B2(n_1193),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_1212),
.B(n_1210),
.Y(n_1214)
);

OAI22xp5_ASAP7_75t_SL g1215 ( 
.A1(n_1208),
.A2(n_1207),
.B1(n_1192),
.B2(n_1200),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_1211),
.Y(n_1216)
);

OAI21xp5_ASAP7_75t_L g1217 ( 
.A1(n_1209),
.A2(n_1203),
.B(n_1205),
.Y(n_1217)
);

XNOR2xp5_ASAP7_75t_L g1218 ( 
.A(n_1214),
.B(n_1213),
.Y(n_1218)
);

OAI22xp5_ASAP7_75t_L g1219 ( 
.A1(n_1218),
.A2(n_1216),
.B1(n_1215),
.B2(n_1217),
.Y(n_1219)
);

OAI21xp33_ASAP7_75t_L g1220 ( 
.A1(n_1219),
.A2(n_112),
.B(n_113),
.Y(n_1220)
);

XNOR2x1_ASAP7_75t_L g1221 ( 
.A(n_1220),
.B(n_119),
.Y(n_1221)
);

AOI221xp5_ASAP7_75t_L g1222 ( 
.A1(n_1221),
.A2(n_124),
.B1(n_126),
.B2(n_127),
.C(n_129),
.Y(n_1222)
);

AOI211xp5_ASAP7_75t_L g1223 ( 
.A1(n_1222),
.A2(n_130),
.B(n_133),
.C(n_134),
.Y(n_1223)
);


endmodule