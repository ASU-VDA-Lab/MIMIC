module fake_jpeg_29839_n_71 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_71);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_71;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_40;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_62;
wire n_31;
wire n_56;
wire n_67;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;
wire n_70;
wire n_66;

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_19),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_15),
.B(n_24),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVx2_ASAP7_75t_SL g30 ( 
.A(n_17),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_31),
.A2(n_30),
.B1(n_32),
.B2(n_29),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_33),
.A2(n_39),
.B1(n_3),
.B2(n_4),
.Y(n_45)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_31),
.Y(n_34)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_32),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_35),
.B(n_27),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_26),
.B(n_0),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_36),
.B(n_4),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_28),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_37),
.B(n_38),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_30),
.B(n_0),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_L g39 ( 
.A1(n_26),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_35),
.A2(n_29),
.B1(n_27),
.B2(n_14),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_40),
.A2(n_45),
.B1(n_6),
.B2(n_8),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_43),
.B(n_44),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_36),
.B(n_2),
.Y(n_44)
);

XNOR2xp5_ASAP7_75t_L g58 ( 
.A(n_47),
.B(n_6),
.Y(n_58)
);

XNOR2xp5_ASAP7_75t_SL g49 ( 
.A(n_41),
.B(n_16),
.Y(n_49)
);

XNOR2xp5_ASAP7_75t_SL g60 ( 
.A(n_49),
.B(n_18),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_48),
.B(n_5),
.Y(n_50)
);

XNOR2xp5_ASAP7_75t_SL g61 ( 
.A(n_50),
.B(n_58),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_40),
.B(n_5),
.Y(n_51)
);

OAI21xp5_ASAP7_75t_L g63 ( 
.A1(n_51),
.A2(n_57),
.B(n_20),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_53),
.A2(n_10),
.B1(n_11),
.B2(n_13),
.Y(n_59)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_56),
.Y(n_62)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_59),
.A2(n_63),
.B1(n_55),
.B2(n_54),
.Y(n_66)
);

XNOR2xp5_ASAP7_75t_L g65 ( 
.A(n_60),
.B(n_64),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_L g64 ( 
.A1(n_54),
.A2(n_21),
.B(n_22),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_66),
.A2(n_67),
.B1(n_52),
.B2(n_49),
.Y(n_68)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_62),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_68),
.B(n_61),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_SL g70 ( 
.A1(n_69),
.A2(n_60),
.B(n_65),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_70),
.A2(n_65),
.B1(n_23),
.B2(n_25),
.Y(n_71)
);


endmodule