module fake_netlist_1_911_n_579 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_73, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_71, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_72, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_579);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_73;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_71;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_72;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_579;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_540;
wire n_563;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_554;
wire n_447;
wire n_171;
wire n_567;
wire n_196;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_446;
wire n_342;
wire n_423;
wire n_370;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_260;
wire n_78;
wire n_539;
wire n_201;
wire n_197;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_409;
wire n_363;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_75;
wire n_376;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_497;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_74;
wire n_561;
wire n_335;
wire n_272;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_99;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g74 ( .A(n_66), .Y(n_74) );
INVx1_ASAP7_75t_L g75 ( .A(n_45), .Y(n_75) );
INVx1_ASAP7_75t_L g76 ( .A(n_64), .Y(n_76) );
INVx1_ASAP7_75t_L g77 ( .A(n_1), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_8), .Y(n_78) );
INVxp67_ASAP7_75t_SL g79 ( .A(n_60), .Y(n_79) );
INVxp67_ASAP7_75t_SL g80 ( .A(n_36), .Y(n_80) );
CKINVDCx5p33_ASAP7_75t_R g81 ( .A(n_29), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_15), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_35), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_43), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_5), .Y(n_85) );
CKINVDCx5p33_ASAP7_75t_R g86 ( .A(n_22), .Y(n_86) );
HB1xp67_ASAP7_75t_L g87 ( .A(n_21), .Y(n_87) );
INVx2_ASAP7_75t_L g88 ( .A(n_12), .Y(n_88) );
CKINVDCx5p33_ASAP7_75t_R g89 ( .A(n_27), .Y(n_89) );
INVx2_ASAP7_75t_L g90 ( .A(n_48), .Y(n_90) );
CKINVDCx16_ASAP7_75t_R g91 ( .A(n_39), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_10), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_61), .Y(n_93) );
OR2x2_ASAP7_75t_L g94 ( .A(n_19), .B(n_68), .Y(n_94) );
CKINVDCx5p33_ASAP7_75t_R g95 ( .A(n_72), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_73), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_41), .Y(n_97) );
BUFx6f_ASAP7_75t_L g98 ( .A(n_69), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_5), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_55), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_20), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_2), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_21), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_3), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_20), .Y(n_105) );
INVx2_ASAP7_75t_L g106 ( .A(n_67), .Y(n_106) );
INVxp67_ASAP7_75t_SL g107 ( .A(n_49), .Y(n_107) );
CKINVDCx14_ASAP7_75t_R g108 ( .A(n_59), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_3), .Y(n_109) );
CKINVDCx5p33_ASAP7_75t_R g110 ( .A(n_4), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_34), .Y(n_111) );
INVxp33_ASAP7_75t_SL g112 ( .A(n_30), .Y(n_112) );
CKINVDCx20_ASAP7_75t_R g113 ( .A(n_54), .Y(n_113) );
INVxp33_ASAP7_75t_L g114 ( .A(n_53), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_2), .Y(n_115) );
HB1xp67_ASAP7_75t_L g116 ( .A(n_42), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_22), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_12), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_33), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_25), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_28), .Y(n_121) );
INVxp33_ASAP7_75t_SL g122 ( .A(n_71), .Y(n_122) );
NAND2xp5_ASAP7_75t_SL g123 ( .A(n_98), .B(n_0), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_74), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_116), .Y(n_125) );
AND2x6_ASAP7_75t_L g126 ( .A(n_74), .B(n_37), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_75), .Y(n_127) );
BUFx2_ASAP7_75t_L g128 ( .A(n_87), .Y(n_128) );
OA21x2_ASAP7_75t_L g129 ( .A1(n_75), .A2(n_32), .B(n_65), .Y(n_129) );
AOI22xp5_ASAP7_75t_L g130 ( .A1(n_91), .A2(n_0), .B1(n_1), .B2(n_4), .Y(n_130) );
OA21x2_ASAP7_75t_L g131 ( .A1(n_76), .A2(n_96), .B(n_121), .Y(n_131) );
OAI22xp5_ASAP7_75t_L g132 ( .A1(n_77), .A2(n_6), .B1(n_7), .B2(n_8), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_76), .Y(n_133) );
BUFx2_ASAP7_75t_L g134 ( .A(n_86), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_83), .Y(n_135) );
INVx2_ASAP7_75t_L g136 ( .A(n_90), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_83), .Y(n_137) );
BUFx6f_ASAP7_75t_L g138 ( .A(n_98), .Y(n_138) );
CKINVDCx5p33_ASAP7_75t_R g139 ( .A(n_108), .Y(n_139) );
CKINVDCx5p33_ASAP7_75t_R g140 ( .A(n_113), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g141 ( .A(n_101), .B(n_6), .Y(n_141) );
BUFx6f_ASAP7_75t_L g142 ( .A(n_98), .Y(n_142) );
CKINVDCx5p33_ASAP7_75t_R g143 ( .A(n_110), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_88), .Y(n_144) );
INVxp67_ASAP7_75t_L g145 ( .A(n_102), .Y(n_145) );
NOR2xp33_ASAP7_75t_L g146 ( .A(n_84), .B(n_7), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_88), .Y(n_147) );
CKINVDCx5p33_ASAP7_75t_R g148 ( .A(n_122), .Y(n_148) );
CKINVDCx5p33_ASAP7_75t_R g149 ( .A(n_112), .Y(n_149) );
AND2x2_ASAP7_75t_L g150 ( .A(n_114), .B(n_9), .Y(n_150) );
CKINVDCx5p33_ASAP7_75t_R g151 ( .A(n_81), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_77), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_78), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_78), .Y(n_154) );
INVx2_ASAP7_75t_L g155 ( .A(n_90), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_84), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_106), .B(n_9), .Y(n_157) );
BUFx2_ASAP7_75t_L g158 ( .A(n_94), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_93), .Y(n_159) );
AND2x4_ASAP7_75t_L g160 ( .A(n_82), .B(n_10), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_82), .Y(n_161) );
NOR2xp33_ASAP7_75t_R g162 ( .A(n_89), .B(n_44), .Y(n_162) );
BUFx6f_ASAP7_75t_L g163 ( .A(n_98), .Y(n_163) );
INVx1_ASAP7_75t_L g164 ( .A(n_85), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_85), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_93), .Y(n_166) );
NOR2xp33_ASAP7_75t_L g167 ( .A(n_125), .B(n_106), .Y(n_167) );
NOR2xp33_ASAP7_75t_SL g168 ( .A(n_139), .B(n_94), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_160), .Y(n_169) );
NOR2xp33_ASAP7_75t_L g170 ( .A(n_158), .B(n_121), .Y(n_170) );
CKINVDCx16_ASAP7_75t_R g171 ( .A(n_134), .Y(n_171) );
BUFx3_ASAP7_75t_L g172 ( .A(n_126), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_158), .B(n_95), .Y(n_173) );
AND2x4_ASAP7_75t_L g174 ( .A(n_160), .B(n_104), .Y(n_174) );
INVx2_ASAP7_75t_L g175 ( .A(n_138), .Y(n_175) );
NAND2xp5_ASAP7_75t_SL g176 ( .A(n_139), .B(n_120), .Y(n_176) );
INVx5_ASAP7_75t_L g177 ( .A(n_126), .Y(n_177) );
INVx2_ASAP7_75t_L g178 ( .A(n_138), .Y(n_178) );
BUFx6f_ASAP7_75t_L g179 ( .A(n_138), .Y(n_179) );
AND2x2_ASAP7_75t_L g180 ( .A(n_128), .B(n_104), .Y(n_180) );
NOR2x1p5_ASAP7_75t_L g181 ( .A(n_140), .B(n_103), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_160), .Y(n_182) );
NOR2xp33_ASAP7_75t_L g183 ( .A(n_148), .B(n_120), .Y(n_183) );
OR2x6_ASAP7_75t_L g184 ( .A(n_132), .B(n_103), .Y(n_184) );
INVx4_ASAP7_75t_L g185 ( .A(n_126), .Y(n_185) );
BUFx3_ASAP7_75t_L g186 ( .A(n_126), .Y(n_186) );
OAI22xp5_ASAP7_75t_L g187 ( .A1(n_128), .A2(n_143), .B1(n_149), .B2(n_148), .Y(n_187) );
INVx2_ASAP7_75t_L g188 ( .A(n_138), .Y(n_188) );
INVx2_ASAP7_75t_L g189 ( .A(n_138), .Y(n_189) );
INVx3_ASAP7_75t_L g190 ( .A(n_160), .Y(n_190) );
AND2x2_ASAP7_75t_L g191 ( .A(n_145), .B(n_92), .Y(n_191) );
INVx8_ASAP7_75t_L g192 ( .A(n_126), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_131), .Y(n_193) );
INVx2_ASAP7_75t_L g194 ( .A(n_142), .Y(n_194) );
INVx3_ASAP7_75t_L g195 ( .A(n_136), .Y(n_195) );
INVx1_ASAP7_75t_L g196 ( .A(n_131), .Y(n_196) );
NAND2xp5_ASAP7_75t_SL g197 ( .A(n_151), .B(n_119), .Y(n_197) );
HB1xp67_ASAP7_75t_L g198 ( .A(n_134), .Y(n_198) );
BUFx6f_ASAP7_75t_L g199 ( .A(n_142), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_131), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_131), .Y(n_201) );
AO22x2_ASAP7_75t_L g202 ( .A1(n_124), .A2(n_119), .B1(n_96), .B2(n_97), .Y(n_202) );
BUFx6f_ASAP7_75t_L g203 ( .A(n_142), .Y(n_203) );
BUFx2_ASAP7_75t_L g204 ( .A(n_143), .Y(n_204) );
AND2x4_ASAP7_75t_L g205 ( .A(n_124), .B(n_118), .Y(n_205) );
INVx1_ASAP7_75t_L g206 ( .A(n_136), .Y(n_206) );
INVx2_ASAP7_75t_SL g207 ( .A(n_150), .Y(n_207) );
INVx3_ASAP7_75t_L g208 ( .A(n_155), .Y(n_208) );
AND2x6_ASAP7_75t_L g209 ( .A(n_150), .B(n_100), .Y(n_209) );
AND2x4_ASAP7_75t_L g210 ( .A(n_166), .B(n_118), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_152), .Y(n_211) );
AND2x4_ASAP7_75t_L g212 ( .A(n_127), .B(n_117), .Y(n_212) );
AND2x4_ASAP7_75t_L g213 ( .A(n_127), .B(n_133), .Y(n_213) );
AND2x4_ASAP7_75t_L g214 ( .A(n_166), .B(n_117), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_133), .B(n_97), .Y(n_215) );
INVx2_ASAP7_75t_SL g216 ( .A(n_135), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_155), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_153), .Y(n_218) );
NOR2xp33_ASAP7_75t_L g219 ( .A(n_149), .B(n_100), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_135), .Y(n_220) );
AND2x4_ASAP7_75t_L g221 ( .A(n_137), .B(n_115), .Y(n_221) );
NOR3xp33_ASAP7_75t_L g222 ( .A(n_130), .B(n_115), .C(n_92), .Y(n_222) );
BUFx3_ASAP7_75t_L g223 ( .A(n_126), .Y(n_223) );
NAND3xp33_ASAP7_75t_L g224 ( .A(n_146), .B(n_99), .C(n_109), .Y(n_224) );
INVxp67_ASAP7_75t_L g225 ( .A(n_151), .Y(n_225) );
AND2x2_ASAP7_75t_L g226 ( .A(n_154), .B(n_99), .Y(n_226) );
NOR2xp33_ASAP7_75t_L g227 ( .A(n_161), .B(n_111), .Y(n_227) );
INVx6_ASAP7_75t_L g228 ( .A(n_126), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_137), .B(n_111), .Y(n_229) );
BUFx2_ASAP7_75t_L g230 ( .A(n_198), .Y(n_230) );
NAND2xp5_ASAP7_75t_SL g231 ( .A(n_185), .B(n_162), .Y(n_231) );
AOI22xp5_ASAP7_75t_L g232 ( .A1(n_202), .A2(n_156), .B1(n_159), .B2(n_165), .Y(n_232) );
NAND2xp5_ASAP7_75t_SL g233 ( .A(n_185), .B(n_141), .Y(n_233) );
OAI22xp5_ASAP7_75t_L g234 ( .A1(n_184), .A2(n_156), .B1(n_159), .B2(n_164), .Y(n_234) );
AOI22xp33_ASAP7_75t_L g235 ( .A1(n_209), .A2(n_157), .B1(n_105), .B2(n_109), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_213), .Y(n_236) );
INVx2_ASAP7_75t_L g237 ( .A(n_193), .Y(n_237) );
CKINVDCx5p33_ASAP7_75t_R g238 ( .A(n_171), .Y(n_238) );
NAND2xp5_ASAP7_75t_SL g239 ( .A(n_185), .B(n_105), .Y(n_239) );
INVx2_ASAP7_75t_L g240 ( .A(n_193), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_213), .B(n_79), .Y(n_241) );
INVx2_ASAP7_75t_L g242 ( .A(n_196), .Y(n_242) );
INVx3_ASAP7_75t_L g243 ( .A(n_190), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_213), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_216), .B(n_80), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_216), .B(n_147), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_220), .B(n_107), .Y(n_247) );
AOI22xp33_ASAP7_75t_L g248 ( .A1(n_209), .A2(n_123), .B1(n_144), .B2(n_129), .Y(n_248) );
NAND2xp33_ASAP7_75t_R g249 ( .A(n_204), .B(n_140), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_207), .B(n_129), .Y(n_250) );
NOR2xp67_ASAP7_75t_L g251 ( .A(n_190), .B(n_50), .Y(n_251) );
NAND2xp5_ASAP7_75t_SL g252 ( .A(n_177), .B(n_98), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_220), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_190), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_169), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_207), .B(n_129), .Y(n_256) );
OAI221xp5_ASAP7_75t_L g257 ( .A1(n_222), .A2(n_129), .B1(n_98), .B2(n_163), .C(n_142), .Y(n_257) );
BUFx3_ASAP7_75t_L g258 ( .A(n_192), .Y(n_258) );
INVx3_ASAP7_75t_L g259 ( .A(n_195), .Y(n_259) );
BUFx3_ASAP7_75t_L g260 ( .A(n_192), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_173), .B(n_163), .Y(n_261) );
CKINVDCx5p33_ASAP7_75t_R g262 ( .A(n_204), .Y(n_262) );
AOI22xp33_ASAP7_75t_L g263 ( .A1(n_209), .A2(n_163), .B1(n_142), .B2(n_14), .Y(n_263) );
INVxp67_ASAP7_75t_L g264 ( .A(n_168), .Y(n_264) );
INVx2_ASAP7_75t_SL g265 ( .A(n_192), .Y(n_265) );
AND2x2_ASAP7_75t_L g266 ( .A(n_191), .B(n_11), .Y(n_266) );
INVx2_ASAP7_75t_L g267 ( .A(n_196), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_169), .Y(n_268) );
BUFx3_ASAP7_75t_L g269 ( .A(n_192), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_182), .Y(n_270) );
AND2x4_ASAP7_75t_L g271 ( .A(n_174), .B(n_11), .Y(n_271) );
BUFx3_ASAP7_75t_L g272 ( .A(n_172), .Y(n_272) );
BUFx3_ASAP7_75t_L g273 ( .A(n_172), .Y(n_273) );
NOR2xp33_ASAP7_75t_L g274 ( .A(n_176), .B(n_46), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_182), .Y(n_275) );
INVx2_ASAP7_75t_L g276 ( .A(n_200), .Y(n_276) );
INVx2_ASAP7_75t_L g277 ( .A(n_200), .Y(n_277) );
INVx2_ASAP7_75t_L g278 ( .A(n_201), .Y(n_278) );
BUFx12f_ASAP7_75t_L g279 ( .A(n_209), .Y(n_279) );
CKINVDCx5p33_ASAP7_75t_R g280 ( .A(n_187), .Y(n_280) );
NOR2xp33_ASAP7_75t_L g281 ( .A(n_170), .B(n_47), .Y(n_281) );
OR2x6_ASAP7_75t_L g282 ( .A(n_202), .B(n_163), .Y(n_282) );
INVx2_ASAP7_75t_L g283 ( .A(n_201), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_211), .B(n_163), .Y(n_284) );
INVx2_ASAP7_75t_L g285 ( .A(n_206), .Y(n_285) );
INVx3_ASAP7_75t_L g286 ( .A(n_195), .Y(n_286) );
NOR2xp33_ASAP7_75t_L g287 ( .A(n_183), .B(n_219), .Y(n_287) );
INVx2_ASAP7_75t_L g288 ( .A(n_206), .Y(n_288) );
BUFx4f_ASAP7_75t_L g289 ( .A(n_228), .Y(n_289) );
NAND3xp33_ASAP7_75t_L g290 ( .A(n_224), .B(n_13), .C(n_14), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_217), .Y(n_291) );
INVx2_ASAP7_75t_L g292 ( .A(n_217), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_202), .Y(n_293) );
INVx3_ASAP7_75t_L g294 ( .A(n_195), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_205), .B(n_13), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_202), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_236), .Y(n_297) );
OAI22xp5_ASAP7_75t_L g298 ( .A1(n_282), .A2(n_174), .B1(n_228), .B2(n_225), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_236), .Y(n_299) );
HB1xp67_ASAP7_75t_L g300 ( .A(n_282), .Y(n_300) );
CKINVDCx20_ASAP7_75t_R g301 ( .A(n_262), .Y(n_301) );
AOI21xp5_ASAP7_75t_L g302 ( .A1(n_250), .A2(n_223), .B(n_186), .Y(n_302) );
AOI22xp5_ASAP7_75t_SL g303 ( .A1(n_238), .A2(n_209), .B1(n_180), .B2(n_191), .Y(n_303) );
INVx2_ASAP7_75t_SL g304 ( .A(n_230), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_244), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_287), .B(n_209), .Y(n_306) );
INVx3_ASAP7_75t_L g307 ( .A(n_279), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_244), .B(n_210), .Y(n_308) );
AOI22xp5_ASAP7_75t_L g309 ( .A1(n_271), .A2(n_181), .B1(n_180), .B2(n_197), .Y(n_309) );
CKINVDCx5p33_ASAP7_75t_R g310 ( .A(n_249), .Y(n_310) );
AOI21xp5_ASAP7_75t_L g311 ( .A1(n_256), .A2(n_223), .B(n_186), .Y(n_311) );
AND2x4_ASAP7_75t_L g312 ( .A(n_271), .B(n_226), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_266), .B(n_214), .Y(n_313) );
INVx3_ASAP7_75t_L g314 ( .A(n_279), .Y(n_314) );
AOI21xp5_ASAP7_75t_L g315 ( .A1(n_237), .A2(n_177), .B(n_174), .Y(n_315) );
OR2x6_ASAP7_75t_L g316 ( .A(n_279), .B(n_184), .Y(n_316) );
BUFx6f_ASAP7_75t_L g317 ( .A(n_258), .Y(n_317) );
AND2x2_ASAP7_75t_L g318 ( .A(n_230), .B(n_184), .Y(n_318) );
AOI22xp33_ASAP7_75t_L g319 ( .A1(n_293), .A2(n_205), .B1(n_212), .B2(n_214), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_243), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_243), .Y(n_321) );
O2A1O1Ixp33_ASAP7_75t_L g322 ( .A1(n_234), .A2(n_184), .B(n_229), .C(n_215), .Y(n_322) );
AND2x4_ASAP7_75t_L g323 ( .A(n_271), .B(n_221), .Y(n_323) );
AOI22xp33_ASAP7_75t_L g324 ( .A1(n_293), .A2(n_214), .B1(n_210), .B2(n_212), .Y(n_324) );
INVx4_ASAP7_75t_L g325 ( .A(n_282), .Y(n_325) );
NAND2xp5_ASAP7_75t_SL g326 ( .A(n_296), .B(n_177), .Y(n_326) );
OR2x2_ASAP7_75t_L g327 ( .A(n_280), .B(n_226), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_243), .Y(n_328) );
INVx3_ASAP7_75t_SL g329 ( .A(n_271), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_243), .Y(n_330) );
AND2x2_ASAP7_75t_L g331 ( .A(n_266), .B(n_210), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_241), .B(n_212), .Y(n_332) );
AND2x2_ASAP7_75t_L g333 ( .A(n_264), .B(n_221), .Y(n_333) );
AOI21xp5_ASAP7_75t_L g334 ( .A1(n_237), .A2(n_177), .B(n_218), .Y(n_334) );
BUFx6f_ASAP7_75t_L g335 ( .A(n_258), .Y(n_335) );
CKINVDCx20_ASAP7_75t_R g336 ( .A(n_234), .Y(n_336) );
HB1xp67_ASAP7_75t_L g337 ( .A(n_282), .Y(n_337) );
CKINVDCx5p33_ASAP7_75t_R g338 ( .A(n_232), .Y(n_338) );
INVx2_ASAP7_75t_L g339 ( .A(n_237), .Y(n_339) );
OAI22xp33_ASAP7_75t_L g340 ( .A1(n_282), .A2(n_208), .B1(n_221), .B2(n_205), .Y(n_340) );
AND2x4_ASAP7_75t_L g341 ( .A(n_258), .B(n_167), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_246), .Y(n_342) );
AO32x2_ASAP7_75t_L g343 ( .A1(n_257), .A2(n_208), .A3(n_227), .B1(n_228), .B2(n_177), .Y(n_343) );
INVx6_ASAP7_75t_L g344 ( .A(n_260), .Y(n_344) );
INVx1_ASAP7_75t_SL g345 ( .A(n_241), .Y(n_345) );
CKINVDCx20_ASAP7_75t_R g346 ( .A(n_232), .Y(n_346) );
INVxp67_ASAP7_75t_L g347 ( .A(n_245), .Y(n_347) );
OR2x6_ASAP7_75t_SL g348 ( .A(n_295), .B(n_15), .Y(n_348) );
BUFx3_ASAP7_75t_L g349 ( .A(n_285), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_339), .Y(n_350) );
AOI221xp5_ASAP7_75t_L g351 ( .A1(n_322), .A2(n_247), .B1(n_235), .B2(n_296), .C(n_270), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_347), .B(n_255), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_339), .Y(n_353) );
INVx2_ASAP7_75t_L g354 ( .A(n_349), .Y(n_354) );
OA21x2_ASAP7_75t_L g355 ( .A1(n_302), .A2(n_248), .B(n_251), .Y(n_355) );
OAI22xp5_ASAP7_75t_L g356 ( .A1(n_340), .A2(n_253), .B1(n_242), .B2(n_278), .Y(n_356) );
CKINVDCx16_ASAP7_75t_R g357 ( .A(n_301), .Y(n_357) );
INVx2_ASAP7_75t_L g358 ( .A(n_349), .Y(n_358) );
OAI221xp5_ASAP7_75t_L g359 ( .A1(n_309), .A2(n_247), .B1(n_245), .B2(n_268), .C(n_275), .Y(n_359) );
AOI22xp33_ASAP7_75t_L g360 ( .A1(n_336), .A2(n_275), .B1(n_255), .B2(n_268), .Y(n_360) );
OR2x6_ASAP7_75t_L g361 ( .A(n_323), .B(n_240), .Y(n_361) );
INVx2_ASAP7_75t_L g362 ( .A(n_297), .Y(n_362) );
INVx2_ASAP7_75t_L g363 ( .A(n_299), .Y(n_363) );
CKINVDCx8_ASAP7_75t_R g364 ( .A(n_316), .Y(n_364) );
INVxp67_ASAP7_75t_SL g365 ( .A(n_340), .Y(n_365) );
CKINVDCx5p33_ASAP7_75t_R g366 ( .A(n_301), .Y(n_366) );
INVxp67_ASAP7_75t_L g367 ( .A(n_304), .Y(n_367) );
AO21x2_ASAP7_75t_L g368 ( .A1(n_306), .A2(n_251), .B(n_290), .Y(n_368) );
AOI22xp33_ASAP7_75t_L g369 ( .A1(n_336), .A2(n_270), .B1(n_254), .B2(n_253), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_305), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_342), .Y(n_371) );
CKINVDCx5p33_ASAP7_75t_R g372 ( .A(n_310), .Y(n_372) );
AOI221x1_ASAP7_75t_L g373 ( .A1(n_298), .A2(n_290), .B1(n_281), .B2(n_261), .C(n_274), .Y(n_373) );
INVxp33_ASAP7_75t_L g374 ( .A(n_303), .Y(n_374) );
NAND2x1p5_ASAP7_75t_L g375 ( .A(n_325), .B(n_283), .Y(n_375) );
OAI21x1_ASAP7_75t_L g376 ( .A1(n_311), .A2(n_283), .B(n_242), .Y(n_376) );
OR2x6_ASAP7_75t_L g377 ( .A(n_323), .B(n_283), .Y(n_377) );
AOI22xp5_ASAP7_75t_L g378 ( .A1(n_346), .A2(n_254), .B1(n_292), .B2(n_285), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_308), .Y(n_379) );
AOI22xp5_ASAP7_75t_L g380 ( .A1(n_346), .A2(n_285), .B1(n_292), .B2(n_288), .Y(n_380) );
BUFx12f_ASAP7_75t_L g381 ( .A(n_316), .Y(n_381) );
AOI221x1_ASAP7_75t_L g382 ( .A1(n_356), .A2(n_325), .B1(n_313), .B2(n_323), .C(n_312), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_371), .Y(n_383) );
BUFx8_ASAP7_75t_L g384 ( .A(n_381), .Y(n_384) );
AND2x2_ASAP7_75t_L g385 ( .A(n_371), .B(n_312), .Y(n_385) );
OAI21xp33_ASAP7_75t_L g386 ( .A1(n_380), .A2(n_327), .B(n_333), .Y(n_386) );
NAND2x1_ASAP7_75t_L g387 ( .A(n_350), .B(n_288), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_360), .B(n_345), .Y(n_388) );
OAI22xp5_ASAP7_75t_L g389 ( .A1(n_380), .A2(n_338), .B1(n_329), .B2(n_319), .Y(n_389) );
OAI221xp5_ASAP7_75t_L g390 ( .A1(n_369), .A2(n_318), .B1(n_319), .B2(n_324), .C(n_316), .Y(n_390) );
INVx4_ASAP7_75t_L g391 ( .A(n_361), .Y(n_391) );
OAI22xp33_ASAP7_75t_L g392 ( .A1(n_378), .A2(n_348), .B1(n_300), .B2(n_337), .Y(n_392) );
OAI211xp5_ASAP7_75t_L g393 ( .A1(n_364), .A2(n_332), .B(n_324), .C(n_331), .Y(n_393) );
NAND3xp33_ASAP7_75t_L g394 ( .A(n_373), .B(n_263), .C(n_284), .Y(n_394) );
AOI22xp33_ASAP7_75t_L g395 ( .A1(n_374), .A2(n_341), .B1(n_300), .B2(n_337), .Y(n_395) );
OA21x2_ASAP7_75t_L g396 ( .A1(n_376), .A2(n_284), .B(n_334), .Y(n_396) );
AOI22xp33_ASAP7_75t_SL g397 ( .A1(n_365), .A2(n_341), .B1(n_307), .B2(n_314), .Y(n_397) );
BUFx2_ASAP7_75t_L g398 ( .A(n_361), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_370), .Y(n_399) );
INVx1_ASAP7_75t_SL g400 ( .A(n_366), .Y(n_400) );
AOI22xp33_ASAP7_75t_L g401 ( .A1(n_359), .A2(n_307), .B1(n_314), .B2(n_294), .Y(n_401) );
OAI221xp5_ASAP7_75t_L g402 ( .A1(n_378), .A2(n_320), .B1(n_330), .B2(n_328), .C(n_321), .Y(n_402) );
OAI21x1_ASAP7_75t_L g403 ( .A1(n_376), .A2(n_326), .B(n_315), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_370), .Y(n_404) );
OAI22xp5_ASAP7_75t_L g405 ( .A1(n_361), .A2(n_288), .B1(n_292), .B2(n_291), .Y(n_405) );
OAI22xp5_ASAP7_75t_L g406 ( .A1(n_361), .A2(n_291), .B1(n_276), .B2(n_277), .Y(n_406) );
A2O1A1Ixp33_ASAP7_75t_L g407 ( .A1(n_351), .A2(n_267), .B(n_242), .C(n_240), .Y(n_407) );
OAI22xp33_ASAP7_75t_L g408 ( .A1(n_357), .A2(n_344), .B1(n_317), .B2(n_335), .Y(n_408) );
INVx2_ASAP7_75t_L g409 ( .A(n_350), .Y(n_409) );
NAND2x1p5_ASAP7_75t_L g410 ( .A(n_353), .B(n_317), .Y(n_410) );
AND4x1_ASAP7_75t_L g411 ( .A(n_382), .B(n_364), .C(n_357), .D(n_373), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_409), .Y(n_412) );
OR2x6_ASAP7_75t_L g413 ( .A(n_391), .B(n_361), .Y(n_413) );
AND2x4_ASAP7_75t_L g414 ( .A(n_391), .B(n_353), .Y(n_414) );
NAND4xp25_ASAP7_75t_SL g415 ( .A(n_393), .B(n_381), .C(n_352), .D(n_379), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_409), .Y(n_416) );
AOI22xp33_ASAP7_75t_L g417 ( .A1(n_386), .A2(n_379), .B1(n_362), .B2(n_363), .Y(n_417) );
INVx2_ASAP7_75t_L g418 ( .A(n_396), .Y(n_418) );
AND2x2_ASAP7_75t_L g419 ( .A(n_399), .B(n_362), .Y(n_419) );
OA21x2_ASAP7_75t_L g420 ( .A1(n_382), .A2(n_363), .B(n_362), .Y(n_420) );
AOI221xp5_ASAP7_75t_L g421 ( .A1(n_392), .A2(n_367), .B1(n_363), .B2(n_372), .C(n_208), .Y(n_421) );
INVx2_ASAP7_75t_L g422 ( .A(n_396), .Y(n_422) );
INVx2_ASAP7_75t_SL g423 ( .A(n_391), .Y(n_423) );
AOI21xp5_ASAP7_75t_L g424 ( .A1(n_407), .A2(n_355), .B(n_377), .Y(n_424) );
OR2x2_ASAP7_75t_L g425 ( .A(n_404), .B(n_377), .Y(n_425) );
AOI33xp33_ASAP7_75t_L g426 ( .A1(n_400), .A2(n_16), .A3(n_17), .B1(n_18), .B2(n_19), .B3(n_23), .Y(n_426) );
OAI22xp5_ASAP7_75t_L g427 ( .A1(n_389), .A2(n_377), .B1(n_375), .B2(n_358), .Y(n_427) );
BUFx2_ASAP7_75t_L g428 ( .A(n_398), .Y(n_428) );
OAI211xp5_ASAP7_75t_L g429 ( .A1(n_397), .A2(n_286), .B(n_259), .C(n_294), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_383), .Y(n_430) );
INVx2_ASAP7_75t_L g431 ( .A(n_403), .Y(n_431) );
OAI22xp5_ASAP7_75t_L g432 ( .A1(n_390), .A2(n_377), .B1(n_375), .B2(n_358), .Y(n_432) );
AO21x2_ASAP7_75t_L g433 ( .A1(n_394), .A2(n_368), .B(n_354), .Y(n_433) );
NOR2x2_ASAP7_75t_L g434 ( .A(n_384), .B(n_377), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_387), .Y(n_435) );
AND2x2_ASAP7_75t_L g436 ( .A(n_385), .B(n_354), .Y(n_436) );
BUFx3_ASAP7_75t_L g437 ( .A(n_387), .Y(n_437) );
OAI21x1_ASAP7_75t_L g438 ( .A1(n_403), .A2(n_355), .B(n_375), .Y(n_438) );
NAND3xp33_ASAP7_75t_L g439 ( .A(n_401), .B(n_355), .C(n_326), .Y(n_439) );
OAI31xp33_ASAP7_75t_L g440 ( .A1(n_388), .A2(n_259), .A3(n_286), .B(n_294), .Y(n_440) );
AND2x2_ASAP7_75t_L g441 ( .A(n_385), .B(n_368), .Y(n_441) );
AOI221xp5_ASAP7_75t_L g442 ( .A1(n_395), .A2(n_259), .B1(n_286), .B2(n_294), .C(n_239), .Y(n_442) );
AO21x2_ASAP7_75t_L g443 ( .A1(n_407), .A2(n_368), .B(n_355), .Y(n_443) );
BUFx10_ASAP7_75t_L g444 ( .A(n_384), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_412), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_416), .Y(n_446) );
OAI31xp33_ASAP7_75t_L g447 ( .A1(n_415), .A2(n_408), .A3(n_405), .B(n_402), .Y(n_447) );
OR2x2_ASAP7_75t_L g448 ( .A(n_428), .B(n_410), .Y(n_448) );
AND2x4_ASAP7_75t_L g449 ( .A(n_441), .B(n_56), .Y(n_449) );
AOI31xp67_ASAP7_75t_L g450 ( .A1(n_418), .A2(n_175), .A3(n_178), .B(n_188), .Y(n_450) );
AND2x2_ASAP7_75t_L g451 ( .A(n_441), .B(n_410), .Y(n_451) );
BUFx2_ASAP7_75t_L g452 ( .A(n_437), .Y(n_452) );
AND2x2_ASAP7_75t_SL g453 ( .A(n_428), .B(n_406), .Y(n_453) );
AND2x4_ASAP7_75t_L g454 ( .A(n_435), .B(n_58), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_418), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_430), .B(n_384), .Y(n_456) );
OAI211xp5_ASAP7_75t_L g457 ( .A1(n_421), .A2(n_286), .B(n_259), .C(n_252), .Y(n_457) );
AOI221xp5_ASAP7_75t_L g458 ( .A1(n_421), .A2(n_233), .B1(n_188), .B2(n_175), .C(n_189), .Y(n_458) );
AOI22xp33_ASAP7_75t_L g459 ( .A1(n_415), .A2(n_335), .B1(n_317), .B2(n_344), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_422), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_419), .B(n_16), .Y(n_461) );
AND2x4_ASAP7_75t_L g462 ( .A(n_435), .B(n_57), .Y(n_462) );
AOI221xp5_ASAP7_75t_L g463 ( .A1(n_432), .A2(n_189), .B1(n_194), .B2(n_178), .C(n_179), .Y(n_463) );
INVx2_ASAP7_75t_L g464 ( .A(n_422), .Y(n_464) );
OAI31xp33_ASAP7_75t_L g465 ( .A1(n_429), .A2(n_231), .A3(n_240), .B(n_267), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_422), .Y(n_466) );
AND2x2_ASAP7_75t_L g467 ( .A(n_419), .B(n_343), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_436), .B(n_343), .Y(n_468) );
AND2x2_ASAP7_75t_L g469 ( .A(n_436), .B(n_343), .Y(n_469) );
AOI22xp33_ASAP7_75t_L g470 ( .A1(n_427), .A2(n_432), .B1(n_413), .B2(n_440), .Y(n_470) );
OAI33xp33_ASAP7_75t_L g471 ( .A1(n_427), .A2(n_17), .A3(n_18), .B1(n_23), .B2(n_194), .B3(n_267), .Y(n_471) );
AND2x4_ASAP7_75t_L g472 ( .A(n_437), .B(n_24), .Y(n_472) );
AOI211xp5_ASAP7_75t_L g473 ( .A1(n_429), .A2(n_335), .B(n_317), .C(n_277), .Y(n_473) );
AND2x2_ASAP7_75t_L g474 ( .A(n_414), .B(n_26), .Y(n_474) );
AND2x2_ASAP7_75t_L g475 ( .A(n_414), .B(n_31), .Y(n_475) );
OR2x6_ASAP7_75t_L g476 ( .A(n_413), .B(n_335), .Y(n_476) );
INVx2_ASAP7_75t_L g477 ( .A(n_431), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_420), .Y(n_478) );
INVx2_ASAP7_75t_L g479 ( .A(n_431), .Y(n_479) );
NAND2x1p5_ASAP7_75t_L g480 ( .A(n_437), .B(n_278), .Y(n_480) );
INVx2_ASAP7_75t_L g481 ( .A(n_431), .Y(n_481) );
BUFx3_ASAP7_75t_L g482 ( .A(n_414), .Y(n_482) );
CKINVDCx5p33_ASAP7_75t_R g483 ( .A(n_456), .Y(n_483) );
AOI21xp5_ASAP7_75t_L g484 ( .A1(n_473), .A2(n_424), .B(n_440), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_445), .Y(n_485) );
OR2x2_ASAP7_75t_L g486 ( .A(n_446), .B(n_425), .Y(n_486) );
OAI33xp33_ASAP7_75t_L g487 ( .A1(n_461), .A2(n_425), .A3(n_426), .B1(n_439), .B2(n_411), .B3(n_444), .Y(n_487) );
AND2x4_ASAP7_75t_L g488 ( .A(n_482), .B(n_423), .Y(n_488) );
OR2x6_ASAP7_75t_L g489 ( .A(n_452), .B(n_413), .Y(n_489) );
CKINVDCx8_ASAP7_75t_R g490 ( .A(n_449), .Y(n_490) );
OR2x2_ASAP7_75t_L g491 ( .A(n_451), .B(n_413), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_455), .Y(n_492) );
NOR2xp33_ASAP7_75t_SL g493 ( .A(n_453), .B(n_444), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_455), .Y(n_494) );
NAND2xp33_ASAP7_75t_SL g495 ( .A(n_474), .B(n_434), .Y(n_495) );
AOI21xp5_ASAP7_75t_L g496 ( .A1(n_473), .A2(n_424), .B(n_438), .Y(n_496) );
NAND2xp33_ASAP7_75t_R g497 ( .A(n_452), .B(n_444), .Y(n_497) );
AND2x2_ASAP7_75t_L g498 ( .A(n_482), .B(n_413), .Y(n_498) );
AO21x1_ASAP7_75t_L g499 ( .A1(n_447), .A2(n_411), .B(n_438), .Y(n_499) );
NAND2xp33_ASAP7_75t_R g500 ( .A(n_472), .B(n_413), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_460), .Y(n_501) );
OR2x2_ASAP7_75t_L g502 ( .A(n_448), .B(n_420), .Y(n_502) );
INVx2_ASAP7_75t_L g503 ( .A(n_466), .Y(n_503) );
NAND2xp33_ASAP7_75t_SL g504 ( .A(n_474), .B(n_417), .Y(n_504) );
AND3x2_ASAP7_75t_L g505 ( .A(n_475), .B(n_442), .C(n_439), .Y(n_505) );
AND2x4_ASAP7_75t_L g506 ( .A(n_449), .B(n_438), .Y(n_506) );
AOI22xp33_ASAP7_75t_L g507 ( .A1(n_470), .A2(n_442), .B1(n_443), .B2(n_433), .Y(n_507) );
CKINVDCx14_ASAP7_75t_R g508 ( .A(n_475), .Y(n_508) );
OR2x2_ASAP7_75t_L g509 ( .A(n_464), .B(n_38), .Y(n_509) );
NAND3xp33_ASAP7_75t_L g510 ( .A(n_459), .B(n_199), .C(n_203), .Y(n_510) );
NOR2xp33_ASAP7_75t_R g511 ( .A(n_453), .B(n_40), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_467), .B(n_276), .Y(n_512) );
AOI22xp5_ASAP7_75t_L g513 ( .A1(n_493), .A2(n_453), .B1(n_471), .B2(n_468), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_485), .B(n_478), .Y(n_514) );
AOI211x1_ASAP7_75t_L g515 ( .A1(n_499), .A2(n_457), .B(n_478), .C(n_469), .Y(n_515) );
OAI22xp5_ASAP7_75t_L g516 ( .A1(n_490), .A2(n_472), .B1(n_454), .B2(n_462), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_508), .B(n_481), .Y(n_517) );
O2A1O1Ixp33_ASAP7_75t_L g518 ( .A1(n_487), .A2(n_454), .B(n_462), .C(n_472), .Y(n_518) );
AOI22xp5_ASAP7_75t_L g519 ( .A1(n_493), .A2(n_462), .B1(n_454), .B2(n_472), .Y(n_519) );
OAI22xp33_ASAP7_75t_L g520 ( .A1(n_500), .A2(n_476), .B1(n_480), .B2(n_454), .Y(n_520) );
AOI221xp5_ASAP7_75t_L g521 ( .A1(n_487), .A2(n_462), .B1(n_463), .B2(n_477), .C(n_479), .Y(n_521) );
HB1xp67_ASAP7_75t_L g522 ( .A(n_497), .Y(n_522) );
NOR2xp33_ASAP7_75t_L g523 ( .A(n_483), .B(n_476), .Y(n_523) );
A2O1A1Ixp33_ASAP7_75t_L g524 ( .A1(n_495), .A2(n_465), .B(n_479), .C(n_458), .Y(n_524) );
NOR2xp33_ASAP7_75t_L g525 ( .A(n_491), .B(n_476), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_486), .B(n_476), .Y(n_526) );
AOI22xp33_ASAP7_75t_L g527 ( .A1(n_504), .A2(n_476), .B1(n_480), .B2(n_344), .Y(n_527) );
NOR2x2_ASAP7_75t_L g528 ( .A(n_489), .B(n_511), .Y(n_528) );
OR4x1_ASAP7_75t_L g529 ( .A(n_492), .B(n_450), .C(n_51), .D(n_52), .Y(n_529) );
INVxp67_ASAP7_75t_L g530 ( .A(n_488), .Y(n_530) );
NAND2xp5_ASAP7_75t_SL g531 ( .A(n_488), .B(n_278), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_494), .Y(n_532) );
AO22x2_ASAP7_75t_L g533 ( .A1(n_502), .A2(n_62), .B1(n_63), .B2(n_70), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_501), .Y(n_534) );
AOI32xp33_ASAP7_75t_L g535 ( .A1(n_506), .A2(n_260), .A3(n_269), .B1(n_265), .B2(n_272), .Y(n_535) );
INVx2_ASAP7_75t_L g536 ( .A(n_503), .Y(n_536) );
OAI22xp5_ASAP7_75t_L g537 ( .A1(n_489), .A2(n_228), .B1(n_269), .B2(n_260), .Y(n_537) );
OAI21xp5_ASAP7_75t_L g538 ( .A1(n_518), .A2(n_484), .B(n_510), .Y(n_538) );
AOI31xp33_ASAP7_75t_L g539 ( .A1(n_522), .A2(n_507), .A3(n_498), .B(n_496), .Y(n_539) );
AO22x1_ASAP7_75t_L g540 ( .A1(n_516), .A2(n_505), .B1(n_489), .B2(n_512), .Y(n_540) );
AND3x2_ASAP7_75t_L g541 ( .A(n_523), .B(n_505), .C(n_509), .Y(n_541) );
AND2x2_ASAP7_75t_L g542 ( .A(n_536), .B(n_179), .Y(n_542) );
NOR2x1_ASAP7_75t_L g543 ( .A(n_516), .B(n_520), .Y(n_543) );
AOI221xp5_ASAP7_75t_L g544 ( .A1(n_515), .A2(n_199), .B1(n_203), .B2(n_272), .C(n_273), .Y(n_544) );
AOI222xp33_ASAP7_75t_L g545 ( .A1(n_530), .A2(n_199), .B1(n_203), .B2(n_272), .C1(n_273), .C2(n_289), .Y(n_545) );
AOI21xp5_ASAP7_75t_SL g546 ( .A1(n_519), .A2(n_269), .B(n_265), .Y(n_546) );
XOR2x2_ASAP7_75t_L g547 ( .A(n_517), .B(n_273), .Y(n_547) );
INVx1_ASAP7_75t_SL g548 ( .A(n_528), .Y(n_548) );
NAND2x1p5_ASAP7_75t_L g549 ( .A(n_531), .B(n_289), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_532), .B(n_289), .Y(n_550) );
OAI21xp33_ASAP7_75t_L g551 ( .A1(n_513), .A2(n_533), .B(n_527), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_534), .Y(n_552) );
OAI221xp5_ASAP7_75t_L g553 ( .A1(n_524), .A2(n_535), .B1(n_521), .B2(n_525), .C(n_526), .Y(n_553) );
NOR2xp33_ASAP7_75t_L g554 ( .A(n_548), .B(n_514), .Y(n_554) );
OAI211xp5_ASAP7_75t_SL g555 ( .A1(n_551), .A2(n_537), .B(n_533), .C(n_529), .Y(n_555) );
XNOR2xp5_ASAP7_75t_L g556 ( .A(n_543), .B(n_537), .Y(n_556) );
AOI31xp33_ASAP7_75t_L g557 ( .A1(n_543), .A2(n_538), .A3(n_553), .B(n_540), .Y(n_557) );
NOR2x1_ASAP7_75t_L g558 ( .A(n_546), .B(n_539), .Y(n_558) );
OAI21x1_ASAP7_75t_SL g559 ( .A1(n_540), .A2(n_552), .B(n_544), .Y(n_559) );
NOR2xp33_ASAP7_75t_R g560 ( .A(n_541), .B(n_546), .Y(n_560) );
NAND2xp5_ASAP7_75t_SL g561 ( .A(n_557), .B(n_547), .Y(n_561) );
NAND4xp25_ASAP7_75t_L g562 ( .A(n_554), .B(n_545), .C(n_550), .D(n_542), .Y(n_562) );
AND3x2_ASAP7_75t_L g563 ( .A(n_560), .B(n_549), .C(n_559), .Y(n_563) );
INVxp67_ASAP7_75t_L g564 ( .A(n_554), .Y(n_564) );
NOR3xp33_ASAP7_75t_L g565 ( .A(n_557), .B(n_555), .C(n_551), .Y(n_565) );
NOR2x1_ASAP7_75t_L g566 ( .A(n_557), .B(n_558), .Y(n_566) );
OAI22xp5_ASAP7_75t_L g567 ( .A1(n_557), .A2(n_543), .B1(n_556), .B2(n_548), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_565), .B(n_567), .Y(n_568) );
AND2x4_ASAP7_75t_L g569 ( .A(n_566), .B(n_563), .Y(n_569) );
INVx1_ASAP7_75t_SL g570 ( .A(n_563), .Y(n_570) );
AND2x4_ASAP7_75t_L g571 ( .A(n_564), .B(n_561), .Y(n_571) );
BUFx2_ASAP7_75t_L g572 ( .A(n_569), .Y(n_572) );
NOR2x1p5_ASAP7_75t_L g573 ( .A(n_569), .B(n_562), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_571), .Y(n_574) );
HB1xp67_ASAP7_75t_L g575 ( .A(n_574), .Y(n_575) );
INVxp67_ASAP7_75t_L g576 ( .A(n_572), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_575), .Y(n_577) );
AOI22xp5_ASAP7_75t_L g578 ( .A1(n_577), .A2(n_573), .B1(n_568), .B2(n_572), .Y(n_578) );
AOI21xp5_ASAP7_75t_L g579 ( .A1(n_578), .A2(n_576), .B(n_570), .Y(n_579) );
endmodule