module real_aes_17216_n_344 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_64, n_254, n_207, n_10, n_83, n_181, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_239, n_100, n_54, n_112, n_319, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_184, n_28, n_202, n_56, n_34, n_98, n_121, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_304, n_311, n_324, n_25, n_278, n_236, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_323, n_199, n_142, n_223, n_67, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_58, n_165, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_193, n_293, n_162, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_60, n_233, n_290, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_340, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_344);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_184;
input n_28;
input n_202;
input n_56;
input n_34;
input n_98;
input n_121;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_304;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_323;
input n_199;
input n_142;
input n_223;
input n_67;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_58;
input n_165;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_193;
input n_293;
input n_162;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_60;
input n_233;
input n_290;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_340;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_344;
wire n_476;
wire n_887;
wire n_599;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_1797;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_1641;
wire n_503;
wire n_1781;
wire n_1762;
wire n_1591;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_1621;
wire n_1729;
wire n_1737;
wire n_761;
wire n_421;
wire n_919;
wire n_1217;
wire n_1423;
wire n_1034;
wire n_549;
wire n_571;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_1730;
wire n_1744;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1835;
wire n_1468;
wire n_1713;
wire n_870;
wire n_1248;
wire n_1602;
wire n_548;
wire n_1859;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_1520;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_1379;
wire n_400;
wire n_1597;
wire n_1845;
wire n_1415;
wire n_1160;
wire n_1849;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_1687;
wire n_553;
wire n_1805;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1382;
wire n_1225;
wire n_875;
wire n_1199;
wire n_951;
wire n_1441;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1833;
wire n_1477;
wire n_595;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_1599;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_1688;
wire n_956;
wire n_1242;
wire n_1537;
wire n_874;
wire n_796;
wire n_1126;
wire n_383;
wire n_1607;
wire n_455;
wire n_1771;
wire n_1809;
wire n_682;
wire n_1745;
wire n_1820;
wire n_812;
wire n_817;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1639;
wire n_1224;
wire n_1694;
wire n_688;
wire n_1042;
wire n_1588;
wire n_363;
wire n_1317;
wire n_417;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1731;
wire n_1589;
wire n_947;
wire n_970;
wire n_1677;
wire n_1149;
wire n_368;
wire n_527;
wire n_1676;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1346;
wire n_1383;
wire n_1675;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_805;
wire n_1600;
wire n_619;
wire n_1284;
wire n_1095;
wire n_1250;
wire n_360;
wire n_1583;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_488;
wire n_501;
wire n_1380;
wire n_1658;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1502;
wire n_404;
wire n_1073;
wire n_1301;
wire n_728;
wire n_1632;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1768;
wire n_1243;
wire n_1846;
wire n_1003;
wire n_346;
wire n_749;
wire n_914;
wire n_1837;
wire n_1286;
wire n_494;
wire n_1661;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1813;
wire n_1628;
wire n_1587;
wire n_1821;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_1825;
wire n_1615;
wire n_1763;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_1714;
wire n_420;
wire n_1666;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_1814;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1510;
wire n_1495;
wire n_1727;
wire n_712;
wire n_422;
wire n_861;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_1742;
wire n_724;
wire n_1648;
wire n_440;
wire n_1231;
wire n_1305;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_1793;
wire n_837;
wire n_1349;
wire n_1708;
wire n_1445;
wire n_1631;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_1751;
wire n_1765;
wire n_1538;
wire n_652;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_1787;
wire n_424;
wire n_877;
wire n_802;
wire n_1488;
wire n_1572;
wire n_1514;
wire n_480;
wire n_1652;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1657;
wire n_1616;
wire n_1828;
wire n_1860;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_635;
wire n_792;
wire n_1392;
wire n_1542;
wire n_665;
wire n_667;
wire n_991;
wire n_1712;
wire n_1556;
wire n_580;
wire n_1004;
wire n_1370;
wire n_1417;
wire n_1703;
wire n_1717;
wire n_1723;
wire n_979;
wire n_445;
wire n_596;
wire n_1740;
wire n_1197;
wire n_657;
wire n_1260;
wire n_355;
wire n_1606;
wire n_1129;
wire n_1760;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_1629;
wire n_1618;
wire n_461;
wire n_1770;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_1750;
wire n_1852;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_1830;
wire n_1594;
wire n_537;
wire n_1767;
wire n_1651;
wire n_560;
wire n_1094;
wire n_1776;
wire n_1719;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1613;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_948;
wire n_399;
wire n_700;
wire n_1499;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1635;
wire n_1518;
wire n_1702;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1577;
wire n_1839;
wire n_1642;
wire n_1406;
wire n_550;
wire n_966;
wire n_1568;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1612;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_1611;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_1665;
wire n_535;
wire n_882;
wire n_1210;
wire n_1741;
wire n_1456;
wire n_746;
wire n_656;
wire n_1614;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_1653;
wire n_529;
wire n_504;
wire n_973;
wire n_1853;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_1668;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1769;
wire n_1812;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_1680;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_1854;
wire n_617;
wire n_602;
wire n_402;
wire n_733;
wire n_1404;
wire n_658;
wire n_676;
wire n_1856;
wire n_531;
wire n_1848;
wire n_1031;
wire n_1394;
wire n_807;
wire n_1011;
wire n_416;
wire n_1567;
wire n_895;
wire n_1569;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_1626;
wire n_645;
wire n_1145;
wire n_1529;
wire n_557;
wire n_1681;
wire n_1620;
wire n_985;
wire n_777;
wire n_1659;
wire n_910;
wire n_642;
wire n_613;
wire n_1773;
wire n_1125;
wire n_1347;
wire n_1655;
wire n_1766;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_1623;
wire n_735;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1716;
wire n_1232;
wire n_471;
wire n_1857;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_1580;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1634;
wire n_1353;
wire n_1002;
wire n_1165;
wire n_1551;
wire n_1667;
wire n_1058;
wire n_1216;
wire n_662;
wire n_1862;
wire n_850;
wire n_720;
wire n_354;
wire n_1026;
wire n_1756;
wire n_1803;
wire n_492;
wire n_407;
wire n_1023;
wire n_419;
wire n_730;
wire n_1699;
wire n_1794;
wire n_1748;
wire n_643;
wire n_1403;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_1513;
wire n_1194;
wire n_389;
wire n_1609;
wire n_1462;
wire n_701;
wire n_809;
wire n_1532;
wire n_679;
wire n_520;
wire n_926;
wire n_1643;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1784;
wire n_1548;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_1409;
wire n_753;
wire n_1188;
wire n_623;
wire n_1474;
wire n_1032;
wire n_721;
wire n_1431;
wire n_1806;
wire n_1829;
wire n_1133;
wire n_1775;
wire n_1593;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1732;
wire n_1162;
wire n_1463;
wire n_762;
wire n_1524;
wire n_1298;
wire n_442;
wire n_1633;
wire n_740;
wire n_1686;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_1807;
wire n_459;
wire n_1172;
wire n_998;
wire n_1689;
wire n_1625;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1733;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1783;
wire n_1759;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_1578;
wire n_473;
wire n_1779;
wire n_967;
wire n_1709;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_1840;
wire n_968;
wire n_710;
wire n_1040;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_1795;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1451;
wire n_1069;
wire n_842;
wire n_1788;
wire n_798;
wire n_1700;
wire n_668;
wire n_862;
wire n_869;
wire n_1816;
wire n_1811;
wire n_1066;
wire n_1377;
wire n_800;
wire n_1175;
wire n_1170;
wire n_778;
wire n_522;
wire n_1475;
wire n_943;
wire n_977;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1734;
wire n_1333;
wire n_577;
wire n_1610;
wire n_759;
wire n_1235;
wire n_900;
wire n_841;
wire n_1724;
wire n_1218;
wire n_736;
wire n_1706;
wire n_766;
wire n_1113;
wire n_1268;
wire n_852;
wire n_1695;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_1778;
wire n_865;
wire n_1644;
wire n_1736;
wire n_1707;
wire n_856;
wire n_594;
wire n_1146;
wire n_1685;
wire n_1810;
wire n_1435;
wire n_1800;
wire n_374;
wire n_932;
wire n_958;
wire n_1755;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_1540;
wire n_519;
wire n_1116;
wire n_709;
wire n_1834;
wire n_388;
wire n_1470;
wire n_816;
wire n_625;
wire n_953;
wire n_1565;
wire n_1373;
wire n_1558;
wire n_716;
wire n_1683;
wire n_356;
wire n_584;
wire n_896;
wire n_1817;
wire n_1722;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_1638;
wire n_370;
wire n_1663;
wire n_352;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_1168;
wire n_1598;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1850;
wire n_1332;
wire n_1263;
wire n_1411;
wire n_1115;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_1726;
wire n_1827;
wire n_1656;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_1555;
wire n_664;
wire n_367;
wire n_1017;
wire n_936;
wire n_581;
wire n_1215;
wire n_582;
wire n_641;
wire n_1738;
wire n_940;
wire n_745;
wire n_1608;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1743;
wire n_1752;
wire n_1792;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_1560;
wire n_1223;
wire n_405;
wire n_621;
wire n_1012;
wire n_1414;
wire n_1241;
wire n_1671;
wire n_502;
wire n_434;
wire n_769;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1669;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1670;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1660;
wire n_1060;
wire n_1154;
wire n_1786;
wire n_361;
wire n_632;
wire n_1344;
wire n_1450;
wire n_1603;
wire n_1720;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_1764;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_902;
wire n_1749;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_1832;
wire n_366;
wire n_727;
wire n_1083;
wire n_397;
wire n_1855;
wire n_1056;
wire n_1592;
wire n_1605;
wire n_1802;
wire n_663;
wire n_588;
wire n_1682;
wire n_1698;
wire n_1448;
wire n_707;
wire n_915;
wire n_1785;
wire n_1774;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1782;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1798;
wire n_1038;
wire n_1085;
wire n_1838;
wire n_845;
wire n_1673;
wire n_1619;
wire n_1127;
wire n_1718;
wire n_484;
wire n_893;
wire n_1068;
wire n_747;
wire n_1672;
wire n_1753;
wire n_1244;
wire n_1581;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_1772;
wire n_653;
wire n_1725;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1696;
wire n_1355;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_1693;
wire n_1791;
wire n_418;
wire n_771;
wire n_524;
wire n_1378;
wire n_1496;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1824;
wire n_1270;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_1761;
wire n_863;
wire n_525;
wire n_1226;
wire n_1617;
wire n_1790;
wire n_644;
wire n_1150;
wire n_1861;
wire n_1341;
wire n_833;
wire n_1229;
wire n_1690;
wire n_929;
wire n_1143;
wire n_1190;
wire n_1728;
wire n_543;
wire n_1710;
wire n_585;
wire n_465;
wire n_719;
wire n_1343;
wire n_1457;
wire n_1604;
wire n_1156;
wire n_988;
wire n_1757;
wire n_1466;
wire n_921;
wire n_1396;
wire n_1799;
wire n_640;
wire n_1176;
wire n_1691;
wire n_1721;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_1804;
wire n_1480;
wire n_1101;
wire n_1251;
wire n_1076;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1715;
wire n_1407;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1704;
wire n_1844;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1590;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_1841;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1292;
wire n_1192;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_1789;
wire n_987;
wire n_1596;
wire n_362;
wire n_1065;
wire n_1064;
wire n_540;
wire n_1075;
wire n_1822;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_1777;
wire n_458;
wire n_444;
wire n_1200;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_1819;
wire n_1674;
wire n_376;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_460;
wire n_1679;
wire n_1595;
wire n_1735;
wire n_666;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1847;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1622;
wire n_1381;
wire n_1582;
wire n_1747;
wire n_573;
wire n_1099;
wire n_1654;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_1541;
wire n_408;
wire n_1754;
wire n_372;
wire n_578;
wire n_892;
wire n_938;
wire n_774;
wire n_559;
wire n_1049;
wire n_466;
wire n_1277;
wire n_1584;
wire n_984;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_1851;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_532;
wire n_1025;
wire n_1826;
wire n_1836;
wire n_924;
wire n_1264;
wire n_1858;
wire n_1527;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_1678;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1637;
wire n_1290;
wire n_1318;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_1519;
wire n_425;
wire n_1650;
wire n_879;
wire n_1640;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_1818;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1780;
wire n_1823;
wire n_1547;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_1843;
wire n_410;
wire n_1684;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1356;
wire n_1646;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1249;
wire n_1416;
wire n_387;
wire n_1239;
wire n_1796;
wire n_1662;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_1801;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_1252;
wire n_430;
wire n_1647;
wire n_1132;
wire n_1649;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_851;
wire n_470;
wire n_1155;
wire n_934;
wire n_1636;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1808;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_1481;
wire n_907;
wire n_1430;
wire n_1758;
wire n_1005;
wire n_1312;
wire n_1697;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1842;
wire n_1536;
wire n_1746;
wire n_1711;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1601;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_1573;
wire n_1130;
wire n_794;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1624;
wire n_1253;
wire n_1183;
wire n_1831;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_1300;
wire n_575;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1701;
wire n_1664;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1815;
wire n_1412;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1739;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_483;
wire n_1630;
wire n_394;
wire n_1280;
wire n_1352;
wire n_729;
wire n_1323;
wire n_703;
wire n_1369;
wire n_1097;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_348;
wire n_1528;
wire n_603;
wire n_1692;
wire n_1288;
wire n_868;
wire n_1705;
wire n_1024;
wire n_1144;
wire n_1627;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_1645;
wire n_429;
AOI22xp33_ASAP7_75t_L g1205 ( .A1(n_0), .A2(n_267), .B1(n_664), .B2(n_668), .Y(n_1205) );
AOI22xp33_ASAP7_75t_L g1217 ( .A1(n_0), .A2(n_232), .B1(n_467), .B2(n_1218), .Y(n_1217) );
INVx1_ASAP7_75t_L g825 ( .A(n_1), .Y(n_825) );
INVx1_ASAP7_75t_L g1772 ( .A(n_2), .Y(n_1772) );
AO22x1_ASAP7_75t_L g1792 ( .A1(n_2), .A2(n_207), .B1(n_686), .B2(n_692), .Y(n_1792) );
AND2x2_ASAP7_75t_L g446 ( .A(n_3), .B(n_447), .Y(n_446) );
AND2x2_ASAP7_75t_L g477 ( .A(n_3), .B(n_237), .Y(n_477) );
NOR2xp33_ASAP7_75t_L g517 ( .A(n_3), .B(n_518), .Y(n_517) );
INVx1_ASAP7_75t_L g527 ( .A(n_3), .Y(n_527) );
INVx1_ASAP7_75t_L g1779 ( .A(n_4), .Y(n_1779) );
AOI22xp33_ASAP7_75t_L g1791 ( .A1(n_4), .A2(n_119), .B1(n_512), .B2(n_1064), .Y(n_1791) );
INVx1_ASAP7_75t_L g1831 ( .A(n_5), .Y(n_1831) );
OAI22xp5_ASAP7_75t_L g1843 ( .A1(n_5), .A2(n_83), .B1(n_372), .B2(n_1844), .Y(n_1843) );
OAI22xp5_ASAP7_75t_L g1361 ( .A1(n_6), .A2(n_257), .B1(n_1362), .B2(n_1365), .Y(n_1361) );
OAI22xp33_ASAP7_75t_L g1397 ( .A1(n_6), .A2(n_257), .B1(n_1398), .B2(n_1401), .Y(n_1397) );
INVx1_ASAP7_75t_L g655 ( .A(n_7), .Y(n_655) );
OAI221xp5_ASAP7_75t_L g700 ( .A1(n_7), .A2(n_136), .B1(n_701), .B2(n_705), .C(n_710), .Y(n_700) );
INVx1_ASAP7_75t_L g755 ( .A(n_8), .Y(n_755) );
INVx1_ASAP7_75t_L g1171 ( .A(n_9), .Y(n_1171) );
INVx1_ASAP7_75t_L g1820 ( .A(n_10), .Y(n_1820) );
INVx1_ASAP7_75t_L g1044 ( .A(n_11), .Y(n_1044) );
OA222x2_ASAP7_75t_L g1057 ( .A1(n_11), .A2(n_138), .B1(n_164), .B2(n_488), .C1(n_624), .C2(n_1058), .Y(n_1057) );
INVxp67_ASAP7_75t_SL g1158 ( .A(n_12), .Y(n_1158) );
AOI22xp33_ASAP7_75t_L g1186 ( .A1(n_12), .A2(n_113), .B1(n_660), .B2(n_850), .Y(n_1186) );
INVx1_ASAP7_75t_L g1156 ( .A(n_13), .Y(n_1156) );
AOI22xp33_ASAP7_75t_L g1187 ( .A1(n_13), .A2(n_154), .B1(n_403), .B2(n_1188), .Y(n_1187) );
AOI22xp33_ASAP7_75t_SL g1206 ( .A1(n_14), .A2(n_194), .B1(n_412), .B2(n_661), .Y(n_1206) );
AOI221xp5_ASAP7_75t_L g1216 ( .A1(n_14), .A2(n_110), .B1(n_511), .B2(n_819), .C(n_1064), .Y(n_1216) );
OAI221xp5_ASAP7_75t_L g371 ( .A1(n_15), .A2(n_334), .B1(n_372), .B2(n_377), .C(n_383), .Y(n_371) );
OAI21xp33_ASAP7_75t_SL g487 ( .A1(n_15), .A2(n_488), .B(n_491), .Y(n_487) );
INVx1_ASAP7_75t_L g1354 ( .A(n_16), .Y(n_1354) );
AOI22xp33_ASAP7_75t_L g996 ( .A1(n_17), .A2(n_73), .B1(n_551), .B2(n_997), .Y(n_996) );
AOI221xp5_ASAP7_75t_L g1015 ( .A1(n_17), .A2(n_303), .B1(n_934), .B2(n_1016), .C(n_1017), .Y(n_1015) );
INVx2_ASAP7_75t_L g367 ( .A(n_18), .Y(n_367) );
INVx1_ASAP7_75t_L g824 ( .A(n_19), .Y(n_824) );
OAI322xp33_ASAP7_75t_L g828 ( .A1(n_19), .A2(n_829), .A3(n_835), .B1(n_837), .B2(n_844), .C1(n_851), .C2(n_856), .Y(n_828) );
AOI22xp33_ASAP7_75t_L g1168 ( .A1(n_20), .A2(n_154), .B1(n_467), .B2(n_719), .Y(n_1168) );
AOI22xp5_ASAP7_75t_L g1189 ( .A1(n_20), .A2(n_302), .B1(n_1188), .B2(n_1190), .Y(n_1189) );
AOI22xp5_ASAP7_75t_L g1589 ( .A1(n_21), .A2(n_26), .B1(n_1535), .B2(n_1543), .Y(n_1589) );
CKINVDCx5p33_ASAP7_75t_R g1296 ( .A(n_22), .Y(n_1296) );
AOI22xp33_ASAP7_75t_L g1036 ( .A1(n_23), .A2(n_167), .B1(n_1034), .B2(n_1037), .Y(n_1036) );
INVxp67_ASAP7_75t_SL g1076 ( .A(n_23), .Y(n_1076) );
INVx1_ASAP7_75t_L g1320 ( .A(n_24), .Y(n_1320) );
AOI221xp5_ASAP7_75t_L g815 ( .A1(n_25), .A2(n_224), .B1(n_689), .B2(n_816), .C(n_818), .Y(n_815) );
INVx1_ASAP7_75t_L g842 ( .A(n_25), .Y(n_842) );
OAI22xp33_ASAP7_75t_L g416 ( .A1(n_27), .A2(n_277), .B1(n_417), .B2(n_420), .Y(n_416) );
INVx1_ASAP7_75t_L g481 ( .A(n_27), .Y(n_481) );
INVx1_ASAP7_75t_L g930 ( .A(n_28), .Y(n_930) );
OAI211xp5_ASAP7_75t_L g1349 ( .A1(n_29), .A2(n_774), .B(n_1350), .C(n_1353), .Y(n_1349) );
INVx1_ASAP7_75t_L g1396 ( .A(n_29), .Y(n_1396) );
CKINVDCx5p33_ASAP7_75t_R g984 ( .A(n_30), .Y(n_984) );
OAI22xp5_ASAP7_75t_L g756 ( .A1(n_31), .A2(n_309), .B1(n_417), .B2(n_420), .Y(n_756) );
INVxp67_ASAP7_75t_SL g758 ( .A(n_31), .Y(n_758) );
INVx1_ASAP7_75t_L g1246 ( .A(n_32), .Y(n_1246) );
AOI221xp5_ASAP7_75t_L g1261 ( .A1(n_32), .A2(n_133), .B1(n_551), .B2(n_1262), .C(n_1264), .Y(n_1261) );
INVx1_ASAP7_75t_L g595 ( .A(n_33), .Y(n_595) );
AOI221x1_ASAP7_75t_SL g601 ( .A1(n_33), .A2(n_185), .B1(n_467), .B2(n_602), .C(n_606), .Y(n_601) );
INVx1_ASAP7_75t_L g1329 ( .A(n_34), .Y(n_1329) );
HB1xp67_ASAP7_75t_L g1523 ( .A(n_35), .Y(n_1523) );
AND2x2_ASAP7_75t_L g1536 ( .A(n_35), .B(n_1521), .Y(n_1536) );
AOI22xp33_ASAP7_75t_L g1669 ( .A1(n_36), .A2(n_174), .B1(n_1543), .B2(n_1564), .Y(n_1669) );
AOI22xp33_ASAP7_75t_L g1107 ( .A1(n_37), .A2(n_214), .B1(n_1041), .B2(n_1108), .Y(n_1107) );
AOI22xp5_ASAP7_75t_L g1138 ( .A1(n_37), .A2(n_289), .B1(n_939), .B2(n_1139), .Y(n_1138) );
AOI22xp33_ASAP7_75t_L g820 ( .A1(n_38), .A2(n_288), .B1(n_617), .B2(n_821), .Y(n_820) );
INVxp67_ASAP7_75t_L g833 ( .A(n_38), .Y(n_833) );
INVx1_ASAP7_75t_L g586 ( .A(n_39), .Y(n_586) );
AOI22xp33_ASAP7_75t_L g616 ( .A1(n_39), .A2(n_168), .B1(n_512), .B2(n_617), .Y(n_616) );
INVx1_ASAP7_75t_L g790 ( .A(n_40), .Y(n_790) );
OAI211xp5_ASAP7_75t_SL g926 ( .A1(n_41), .A2(n_927), .B(n_929), .C(n_932), .Y(n_926) );
OAI22xp5_ASAP7_75t_L g975 ( .A1(n_41), .A2(n_265), .B1(n_645), .B2(n_859), .Y(n_975) );
INVx1_ASAP7_75t_L g744 ( .A(n_42), .Y(n_744) );
AOI22xp33_ASAP7_75t_L g803 ( .A1(n_43), .A2(n_285), .B1(n_617), .B2(n_804), .Y(n_803) );
AOI22xp33_ASAP7_75t_L g849 ( .A1(n_43), .A2(n_224), .B1(n_660), .B2(n_850), .Y(n_849) );
INVx1_ASAP7_75t_L g1253 ( .A(n_44), .Y(n_1253) );
OAI22xp33_ASAP7_75t_L g1259 ( .A1(n_44), .A2(n_56), .B1(n_372), .B2(n_377), .Y(n_1259) );
AOI22xp33_ASAP7_75t_L g1204 ( .A1(n_45), .A2(n_232), .B1(n_664), .B2(n_668), .Y(n_1204) );
AOI221xp5_ASAP7_75t_L g1213 ( .A1(n_45), .A2(n_267), .B1(n_533), .B2(n_535), .C(n_715), .Y(n_1213) );
OAI22xp5_ASAP7_75t_L g1464 ( .A1(n_46), .A2(n_1465), .B1(n_1466), .B2(n_1467), .Y(n_1464) );
INVx1_ASAP7_75t_L g1465 ( .A(n_46), .Y(n_1465) );
CKINVDCx5p33_ASAP7_75t_R g583 ( .A(n_47), .Y(n_583) );
AOI22xp33_ASAP7_75t_SL g1032 ( .A1(n_48), .A2(n_264), .B1(n_1033), .B2(n_1034), .Y(n_1032) );
INVxp67_ASAP7_75t_SL g1066 ( .A(n_48), .Y(n_1066) );
INVxp67_ASAP7_75t_SL g1161 ( .A(n_49), .Y(n_1161) );
AOI22xp33_ASAP7_75t_SL g1191 ( .A1(n_49), .A2(n_89), .B1(n_660), .B2(n_850), .Y(n_1191) );
INVx1_ASAP7_75t_L g885 ( .A(n_50), .Y(n_885) );
OAI22xp5_ASAP7_75t_L g1283 ( .A1(n_51), .A2(n_396), .B1(n_1284), .B2(n_1287), .Y(n_1283) );
INVx1_ASAP7_75t_L g1301 ( .A(n_51), .Y(n_1301) );
CKINVDCx5p33_ASAP7_75t_R g1198 ( .A(n_52), .Y(n_1198) );
INVx1_ASAP7_75t_L g882 ( .A(n_53), .Y(n_882) );
AOI221xp5_ASAP7_75t_L g910 ( .A1(n_53), .A2(n_254), .B1(n_535), .B2(n_911), .C(n_912), .Y(n_910) );
OAI221xp5_ASAP7_75t_L g940 ( .A1(n_54), .A2(n_112), .B1(n_706), .B2(n_941), .C(n_942), .Y(n_940) );
OAI22xp33_ASAP7_75t_L g968 ( .A1(n_54), .A2(n_112), .B1(n_969), .B2(n_971), .Y(n_968) );
AOI22xp33_ASAP7_75t_L g1486 ( .A1(n_55), .A2(n_177), .B1(n_467), .B2(n_720), .Y(n_1486) );
INVx1_ASAP7_75t_L g1511 ( .A(n_55), .Y(n_1511) );
OAI221xp5_ASAP7_75t_L g1249 ( .A1(n_56), .A2(n_294), .B1(n_491), .B2(n_620), .C(n_622), .Y(n_1249) );
INVx1_ASAP7_75t_L g730 ( .A(n_57), .Y(n_730) );
AOI22xp33_ASAP7_75t_SL g947 ( .A1(n_58), .A2(n_240), .B1(n_948), .B2(n_949), .Y(n_947) );
AOI22xp33_ASAP7_75t_L g959 ( .A1(n_58), .A2(n_337), .B1(n_660), .B2(n_681), .Y(n_959) );
AOI22xp5_ASAP7_75t_L g1562 ( .A1(n_59), .A2(n_192), .B1(n_1535), .B2(n_1540), .Y(n_1562) );
AOI22xp5_ASAP7_75t_L g1550 ( .A1(n_60), .A2(n_323), .B1(n_1543), .B2(n_1551), .Y(n_1550) );
BUFx6f_ASAP7_75t_L g452 ( .A(n_61), .Y(n_452) );
AOI21xp5_ASAP7_75t_L g735 ( .A1(n_62), .A2(n_660), .B(n_736), .Y(n_735) );
INVxp67_ASAP7_75t_SL g768 ( .A(n_62), .Y(n_768) );
INVx1_ASAP7_75t_L g1208 ( .A(n_63), .Y(n_1208) );
CKINVDCx5p33_ASAP7_75t_R g1241 ( .A(n_64), .Y(n_1241) );
INVx1_ASAP7_75t_L g1290 ( .A(n_65), .Y(n_1290) );
AOI22xp33_ASAP7_75t_L g1310 ( .A1(n_65), .A2(n_69), .B1(n_686), .B2(n_720), .Y(n_1310) );
AOI22xp5_ASAP7_75t_L g1563 ( .A1(n_66), .A2(n_301), .B1(n_1543), .B2(n_1564), .Y(n_1563) );
AOI22xp5_ASAP7_75t_L g1569 ( .A1(n_67), .A2(n_121), .B1(n_1535), .B2(n_1540), .Y(n_1569) );
AOI22xp33_ASAP7_75t_L g1488 ( .A1(n_68), .A2(n_206), .B1(n_719), .B2(n_1131), .Y(n_1488) );
INVx1_ASAP7_75t_L g1506 ( .A(n_68), .Y(n_1506) );
AOI221xp5_ASAP7_75t_L g1278 ( .A1(n_69), .A2(n_328), .B1(n_751), .B2(n_1188), .C(n_1279), .Y(n_1278) );
INVxp67_ASAP7_75t_SL g1251 ( .A(n_70), .Y(n_1251) );
OAI22xp5_ASAP7_75t_L g1266 ( .A1(n_70), .A2(n_396), .B1(n_1267), .B2(n_1268), .Y(n_1266) );
OAI221xp5_ASAP7_75t_L g731 ( .A1(n_71), .A2(n_238), .B1(n_372), .B2(n_377), .C(n_383), .Y(n_731) );
OAI221xp5_ASAP7_75t_L g781 ( .A1(n_71), .A2(n_309), .B1(n_491), .B2(n_620), .C(n_622), .Y(n_781) );
OAI22xp5_ASAP7_75t_L g886 ( .A1(n_72), .A2(n_275), .B1(n_389), .B2(n_396), .Y(n_886) );
INVxp67_ASAP7_75t_SL g891 ( .A(n_72), .Y(n_891) );
AOI22xp33_ASAP7_75t_SL g1013 ( .A1(n_73), .A2(n_137), .B1(n_805), .B2(n_938), .Y(n_1013) );
AOI21xp33_ASAP7_75t_L g423 ( .A1(n_74), .A2(n_424), .B(n_427), .Y(n_423) );
AOI221xp5_ASAP7_75t_L g531 ( .A1(n_74), .A2(n_101), .B1(n_532), .B2(n_534), .C(n_536), .Y(n_531) );
INVx1_ASAP7_75t_L g1087 ( .A(n_75), .Y(n_1087) );
CKINVDCx5p33_ASAP7_75t_R g860 ( .A(n_76), .Y(n_860) );
INVx1_ASAP7_75t_L g811 ( .A(n_77), .Y(n_811) );
OAI211xp5_ASAP7_75t_L g861 ( .A1(n_77), .A2(n_862), .B(n_863), .C(n_866), .Y(n_861) );
CKINVDCx5p33_ASAP7_75t_R g1096 ( .A(n_78), .Y(n_1096) );
INVx1_ASAP7_75t_L g1255 ( .A(n_79), .Y(n_1255) );
OAI222xp33_ASAP7_75t_L g1258 ( .A1(n_79), .A2(n_283), .B1(n_294), .B2(n_393), .C1(n_580), .C2(n_843), .Y(n_1258) );
AOI21xp33_ASAP7_75t_L g945 ( .A1(n_80), .A2(n_497), .B(n_946), .Y(n_945) );
INVx1_ASAP7_75t_L g955 ( .A(n_80), .Y(n_955) );
XOR2x2_ASAP7_75t_L g353 ( .A(n_81), .B(n_354), .Y(n_353) );
AOI22xp33_ASAP7_75t_L g1439 ( .A1(n_82), .A2(n_305), .B1(n_874), .B2(n_1440), .Y(n_1439) );
AOI221xp5_ASAP7_75t_L g1447 ( .A1(n_82), .A2(n_325), .B1(n_497), .B2(n_819), .C(n_1448), .Y(n_1447) );
INVx1_ASAP7_75t_L g1825 ( .A(n_83), .Y(n_1825) );
AOI22xp5_ASAP7_75t_L g1554 ( .A1(n_84), .A2(n_336), .B1(n_1535), .B2(n_1540), .Y(n_1554) );
OAI221xp5_ASAP7_75t_L g1470 ( .A1(n_85), .A2(n_118), .B1(n_1067), .B2(n_1471), .C(n_1472), .Y(n_1470) );
INVx1_ASAP7_75t_L g1493 ( .A(n_85), .Y(n_1493) );
AOI22xp33_ASAP7_75t_SL g671 ( .A1(n_86), .A2(n_342), .B1(n_660), .B2(n_661), .Y(n_671) );
AOI221xp5_ASAP7_75t_L g688 ( .A1(n_86), .A2(n_190), .B1(n_602), .B2(n_689), .C(n_690), .Y(n_688) );
CKINVDCx5p33_ASAP7_75t_R g1178 ( .A(n_87), .Y(n_1178) );
XOR2xp5_ASAP7_75t_L g1194 ( .A(n_88), .B(n_1195), .Y(n_1194) );
AOI221xp5_ASAP7_75t_L g1167 ( .A1(n_89), .A2(n_113), .B1(n_497), .B2(n_901), .C(n_936), .Y(n_1167) );
INVx1_ASAP7_75t_L g1474 ( .A(n_90), .Y(n_1474) );
OAI221xp5_ASAP7_75t_SL g1498 ( .A1(n_90), .A2(n_116), .B1(n_375), .B2(n_565), .C(n_876), .Y(n_1498) );
OAI22xp5_ASAP7_75t_L g388 ( .A1(n_91), .A2(n_199), .B1(n_389), .B2(n_396), .Y(n_388) );
INVxp67_ASAP7_75t_SL g519 ( .A(n_91), .Y(n_519) );
AOI22xp5_ASAP7_75t_SL g1555 ( .A1(n_92), .A2(n_204), .B1(n_1543), .B2(n_1551), .Y(n_1555) );
INVx1_ASAP7_75t_L g1221 ( .A(n_93), .Y(n_1221) );
AOI221xp5_ASAP7_75t_L g1039 ( .A1(n_94), .A2(n_108), .B1(n_736), .B2(n_1040), .C(n_1041), .Y(n_1039) );
AOI22xp33_ASAP7_75t_SL g1077 ( .A1(n_94), .A2(n_264), .B1(n_720), .B2(n_939), .Y(n_1077) );
AOI222xp33_ASAP7_75t_L g428 ( .A1(n_95), .A2(n_142), .B1(n_324), .B2(n_398), .C1(n_429), .C2(n_431), .Y(n_428) );
INVx1_ASAP7_75t_L g539 ( .A(n_95), .Y(n_539) );
CKINVDCx5p33_ASAP7_75t_R g1242 ( .A(n_96), .Y(n_1242) );
INVx1_ASAP7_75t_L g878 ( .A(n_97), .Y(n_878) );
AOI221xp5_ASAP7_75t_L g900 ( .A1(n_97), .A2(n_183), .B1(n_901), .B2(n_903), .C(n_905), .Y(n_900) );
OAI22xp33_ASAP7_75t_L g1297 ( .A1(n_98), .A2(n_139), .B1(n_372), .B2(n_377), .Y(n_1297) );
OAI22xp5_ASAP7_75t_L g1311 ( .A1(n_98), .A2(n_281), .B1(n_620), .B2(n_622), .Y(n_1311) );
CKINVDCx5p33_ASAP7_75t_R g1247 ( .A(n_99), .Y(n_1247) );
OAI221xp5_ASAP7_75t_L g1419 ( .A1(n_100), .A2(n_220), .B1(n_1193), .B2(n_1420), .C(n_1421), .Y(n_1419) );
OAI211xp5_ASAP7_75t_L g1445 ( .A1(n_100), .A2(n_701), .B(n_1446), .C(n_1449), .Y(n_1445) );
AOI221xp5_ASAP7_75t_L g400 ( .A1(n_101), .A2(n_213), .B1(n_401), .B2(n_404), .C(n_408), .Y(n_400) );
XNOR2xp5_ASAP7_75t_L g1815 ( .A(n_102), .B(n_1816), .Y(n_1815) );
INVx1_ASAP7_75t_L g1521 ( .A(n_103), .Y(n_1521) );
INVx1_ASAP7_75t_L g1286 ( .A(n_104), .Y(n_1286) );
AOI22xp33_ASAP7_75t_L g1306 ( .A1(n_104), .A2(n_328), .B1(n_467), .B2(n_720), .Y(n_1306) );
INVx1_ASAP7_75t_L g1252 ( .A(n_105), .Y(n_1252) );
INVx1_ASAP7_75t_L g370 ( .A(n_106), .Y(n_370) );
OAI21xp33_ASAP7_75t_L g461 ( .A1(n_106), .A2(n_462), .B(n_471), .Y(n_461) );
AOI221xp5_ASAP7_75t_L g1487 ( .A1(n_107), .A2(n_144), .B1(n_602), .B2(n_689), .C(n_936), .Y(n_1487) );
INVx1_ASAP7_75t_L g1502 ( .A(n_107), .Y(n_1502) );
AOI221xp5_ASAP7_75t_L g1063 ( .A1(n_108), .A2(n_149), .B1(n_689), .B2(n_1064), .C(n_1065), .Y(n_1063) );
OAI22xp5_ASAP7_75t_L g1443 ( .A1(n_109), .A2(n_250), .B1(n_794), .B2(n_859), .Y(n_1443) );
AOI22xp33_ASAP7_75t_L g1201 ( .A1(n_110), .A2(n_236), .B1(n_1202), .B2(n_1203), .Y(n_1201) );
INVx1_ASAP7_75t_L g1323 ( .A(n_111), .Y(n_1323) );
AOI22xp5_ASAP7_75t_L g1557 ( .A1(n_114), .A2(n_312), .B1(n_1540), .B2(n_1551), .Y(n_1557) );
OAI222xp33_ASAP7_75t_L g1784 ( .A1(n_115), .A2(n_320), .B1(n_372), .B2(n_377), .C1(n_1048), .C2(n_1785), .Y(n_1784) );
INVx1_ASAP7_75t_L g1795 ( .A(n_115), .Y(n_1795) );
INVx1_ASAP7_75t_L g1481 ( .A(n_116), .Y(n_1481) );
INVx1_ASAP7_75t_L g555 ( .A(n_117), .Y(n_555) );
OAI22xp5_ASAP7_75t_L g619 ( .A1(n_117), .A2(n_234), .B1(n_620), .B2(n_622), .Y(n_619) );
INVx1_ASAP7_75t_L g1491 ( .A(n_118), .Y(n_1491) );
INVx1_ASAP7_75t_L g1777 ( .A(n_119), .Y(n_1777) );
AOI22xp33_ASAP7_75t_L g937 ( .A1(n_120), .A2(n_228), .B1(n_938), .B2(n_939), .Y(n_937) );
INVx1_ASAP7_75t_L g958 ( .A(n_120), .Y(n_958) );
XOR2x2_ASAP7_75t_L g634 ( .A(n_121), .B(n_635), .Y(n_634) );
AOI22xp5_ASAP7_75t_L g1083 ( .A1(n_122), .A2(n_1084), .B1(n_1085), .B2(n_1146), .Y(n_1083) );
INVx1_ASAP7_75t_L g1146 ( .A(n_122), .Y(n_1146) );
INVx1_ASAP7_75t_L g1478 ( .A(n_123), .Y(n_1478) );
OAI21xp33_ASAP7_75t_L g1496 ( .A1(n_123), .A2(n_639), .B(n_1497), .Y(n_1496) );
CKINVDCx5p33_ASAP7_75t_R g985 ( .A(n_124), .Y(n_985) );
CKINVDCx5p33_ASAP7_75t_R g1281 ( .A(n_125), .Y(n_1281) );
AOI22xp33_ASAP7_75t_SL g1829 ( .A1(n_126), .A2(n_242), .B1(n_719), .B2(n_939), .Y(n_1829) );
AOI221xp5_ASAP7_75t_L g1849 ( .A1(n_126), .A2(n_322), .B1(n_660), .B2(n_736), .C(n_1040), .Y(n_1849) );
OAI22xp33_ASAP7_75t_L g1368 ( .A1(n_127), .A2(n_308), .B1(n_1369), .B2(n_1373), .Y(n_1368) );
OAI22xp5_ASAP7_75t_L g1380 ( .A1(n_127), .A2(n_308), .B1(n_1381), .B2(n_1382), .Y(n_1380) );
INVx1_ASAP7_75t_L g808 ( .A(n_128), .Y(n_808) );
CKINVDCx5p33_ASAP7_75t_R g643 ( .A(n_129), .Y(n_643) );
OAI211xp5_ASAP7_75t_SL g1164 ( .A1(n_130), .A2(n_1165), .B(n_1166), .C(n_1169), .Y(n_1164) );
INVx1_ASAP7_75t_L g1184 ( .A(n_130), .Y(n_1184) );
AOI22xp33_ASAP7_75t_SL g992 ( .A1(n_131), .A2(n_291), .B1(n_993), .B2(n_995), .Y(n_992) );
AOI22xp33_ASAP7_75t_L g1018 ( .A1(n_131), .A2(n_280), .B1(n_805), .B2(n_938), .Y(n_1018) );
OAI222xp33_ASAP7_75t_L g1153 ( .A1(n_132), .A2(n_259), .B1(n_706), .B2(n_941), .C1(n_1154), .C2(n_1157), .Y(n_1153) );
INVx1_ASAP7_75t_L g1181 ( .A(n_132), .Y(n_1181) );
INVx1_ASAP7_75t_L g1232 ( .A(n_133), .Y(n_1232) );
INVx1_ASAP7_75t_L g1432 ( .A(n_134), .Y(n_1432) );
XNOR2x1_ASAP7_75t_L g1149 ( .A(n_135), .B(n_1150), .Y(n_1149) );
INVx1_ASAP7_75t_L g652 ( .A(n_136), .Y(n_652) );
AOI22xp33_ASAP7_75t_L g998 ( .A1(n_137), .A2(n_303), .B1(n_431), .B2(n_999), .Y(n_998) );
INVx1_ASAP7_75t_L g1054 ( .A(n_138), .Y(n_1054) );
INVx1_ASAP7_75t_L g1302 ( .A(n_139), .Y(n_1302) );
AOI221xp5_ASAP7_75t_SL g1485 ( .A1(n_140), .A2(n_300), .B1(n_602), .B2(n_689), .C(n_715), .Y(n_1485) );
INVx1_ASAP7_75t_L g1508 ( .A(n_140), .Y(n_1508) );
CKINVDCx5p33_ASAP7_75t_R g1483 ( .A(n_141), .Y(n_1483) );
INVx1_ASAP7_75t_L g504 ( .A(n_142), .Y(n_504) );
AOI221xp5_ASAP7_75t_L g798 ( .A1(n_143), .A2(n_198), .B1(n_511), .B2(n_799), .C(n_802), .Y(n_798) );
INVxp67_ASAP7_75t_L g830 ( .A(n_143), .Y(n_830) );
INVx1_ASAP7_75t_L g1512 ( .A(n_144), .Y(n_1512) );
AOI22xp33_ASAP7_75t_L g663 ( .A1(n_145), .A2(n_293), .B1(n_664), .B2(n_666), .Y(n_663) );
AOI22xp33_ASAP7_75t_L g691 ( .A1(n_145), .A2(n_251), .B1(n_692), .B2(n_693), .Y(n_691) );
AOI221xp5_ASAP7_75t_L g933 ( .A1(n_146), .A2(n_337), .B1(n_934), .B2(n_935), .C(n_936), .Y(n_933) );
AOI22xp33_ASAP7_75t_L g964 ( .A1(n_146), .A2(n_240), .B1(n_660), .B2(n_965), .Y(n_964) );
INVxp67_ASAP7_75t_SL g1424 ( .A(n_147), .Y(n_1424) );
AOI221xp5_ASAP7_75t_L g1458 ( .A1(n_147), .A2(n_239), .B1(n_535), .B2(n_715), .C(n_1448), .Y(n_1458) );
CKINVDCx5p33_ASAP7_75t_R g573 ( .A(n_148), .Y(n_573) );
AOI221xp5_ASAP7_75t_L g1035 ( .A1(n_149), .A2(n_173), .B1(n_748), .B2(n_850), .C(n_997), .Y(n_1035) );
AOI221xp5_ASAP7_75t_L g879 ( .A1(n_150), .A2(n_183), .B1(n_551), .B2(n_880), .C(n_881), .Y(n_879) );
INVx1_ASAP7_75t_L g916 ( .A(n_150), .Y(n_916) );
INVxp67_ASAP7_75t_SL g1091 ( .A(n_151), .Y(n_1091) );
OAI221xp5_ASAP7_75t_L g1109 ( .A1(n_151), .A2(n_383), .B1(n_389), .B2(n_1110), .C(n_1115), .Y(n_1109) );
AOI21xp5_ASAP7_75t_L g1104 ( .A1(n_152), .A2(n_748), .B(n_1105), .Y(n_1104) );
INVx1_ASAP7_75t_L g1128 ( .A(n_152), .Y(n_1128) );
INVx1_ASAP7_75t_L g1114 ( .A(n_153), .Y(n_1114) );
AOI22xp33_ASAP7_75t_SL g1130 ( .A1(n_153), .A2(n_214), .B1(n_692), .B2(n_1131), .Y(n_1130) );
AOI22xp33_ASAP7_75t_L g750 ( .A1(n_155), .A2(n_339), .B1(n_398), .B2(n_751), .Y(n_750) );
INVxp67_ASAP7_75t_SL g778 ( .A(n_155), .Y(n_778) );
INVx1_ASAP7_75t_L g1197 ( .A(n_156), .Y(n_1197) );
INVx1_ASAP7_75t_L g1774 ( .A(n_157), .Y(n_1774) );
AOI22xp33_ASAP7_75t_L g1800 ( .A1(n_157), .A2(n_249), .B1(n_692), .B2(n_939), .Y(n_1800) );
INVx1_ASAP7_75t_L g1292 ( .A(n_158), .Y(n_1292) );
INVx1_ASAP7_75t_L g1442 ( .A(n_159), .Y(n_1442) );
INVx1_ASAP7_75t_L g734 ( .A(n_160), .Y(n_734) );
INVx1_ASAP7_75t_L g1666 ( .A(n_161), .Y(n_1666) );
AOI22xp5_ASAP7_75t_SL g1568 ( .A1(n_162), .A2(n_169), .B1(n_1543), .B2(n_1551), .Y(n_1568) );
INVx1_ASAP7_75t_L g1357 ( .A(n_163), .Y(n_1357) );
OAI211xp5_ASAP7_75t_L g1385 ( .A1(n_163), .A2(n_1333), .B(n_1386), .C(n_1388), .Y(n_1385) );
OAI221xp5_ASAP7_75t_L g1049 ( .A1(n_164), .A2(n_166), .B1(n_587), .B2(n_1050), .C(n_1051), .Y(n_1049) );
INVx1_ASAP7_75t_L g1170 ( .A(n_165), .Y(n_1170) );
INVxp67_ASAP7_75t_SL g1060 ( .A(n_166), .Y(n_1060) );
INVxp33_ASAP7_75t_SL g1068 ( .A(n_167), .Y(n_1068) );
INVx1_ASAP7_75t_L g578 ( .A(n_168), .Y(n_578) );
INVx2_ASAP7_75t_L g1538 ( .A(n_170), .Y(n_1538) );
AND2x2_ASAP7_75t_L g1541 ( .A(n_170), .B(n_1539), .Y(n_1541) );
AND2x2_ASAP7_75t_L g1546 ( .A(n_170), .B(n_290), .Y(n_1546) );
XNOR2xp5_ASAP7_75t_L g923 ( .A(n_171), .B(n_924), .Y(n_923) );
AOI22xp5_ASAP7_75t_SL g1588 ( .A1(n_171), .A2(n_241), .B1(n_1540), .B2(n_1545), .Y(n_1588) );
INVx1_ASAP7_75t_L g1209 ( .A(n_172), .Y(n_1209) );
INVx1_ASAP7_75t_L g1074 ( .A(n_173), .Y(n_1074) );
OAI21xp33_ASAP7_75t_L g1822 ( .A1(n_175), .A2(n_624), .B(n_1823), .Y(n_1822) );
OAI221xp5_ASAP7_75t_L g1852 ( .A1(n_175), .A2(n_274), .B1(n_961), .B2(n_1853), .C(n_1854), .Y(n_1852) );
AOI22xp5_ASAP7_75t_L g1542 ( .A1(n_176), .A2(n_306), .B1(n_1543), .B2(n_1545), .Y(n_1542) );
INVx1_ASAP7_75t_L g1501 ( .A(n_177), .Y(n_1501) );
AOI22xp5_ASAP7_75t_L g1549 ( .A1(n_178), .A2(n_246), .B1(n_1535), .B2(n_1540), .Y(n_1549) );
INVx1_ASAP7_75t_L g742 ( .A(n_179), .Y(n_742) );
INVx1_ASAP7_75t_L g1805 ( .A(n_180), .Y(n_1805) );
OAI221xp5_ASAP7_75t_L g887 ( .A1(n_181), .A2(n_268), .B1(n_372), .B2(n_377), .C(n_383), .Y(n_887) );
INVx1_ASAP7_75t_L g921 ( .A(n_181), .Y(n_921) );
INVx1_ASAP7_75t_L g1321 ( .A(n_182), .Y(n_1321) );
CKINVDCx5p33_ASAP7_75t_R g570 ( .A(n_184), .Y(n_570) );
INVx1_ASAP7_75t_L g581 ( .A(n_185), .Y(n_581) );
AOI22xp5_ASAP7_75t_L g1558 ( .A1(n_186), .A2(n_269), .B1(n_1535), .B2(n_1543), .Y(n_1558) );
CKINVDCx5p33_ASAP7_75t_R g989 ( .A(n_187), .Y(n_989) );
CKINVDCx5p33_ASAP7_75t_R g1776 ( .A(n_188), .Y(n_1776) );
INVx1_ASAP7_75t_L g1053 ( .A(n_189), .Y(n_1053) );
OAI22xp5_ASAP7_75t_L g1080 ( .A1(n_189), .A2(n_227), .B1(n_474), .B2(n_483), .Y(n_1080) );
AOI22xp33_ASAP7_75t_L g659 ( .A1(n_190), .A2(n_200), .B1(n_660), .B2(n_661), .Y(n_659) );
CKINVDCx5p33_ASAP7_75t_R g1117 ( .A(n_191), .Y(n_1117) );
AOI22xp33_ASAP7_75t_SL g1828 ( .A1(n_193), .A2(n_310), .B1(n_604), .B2(n_911), .Y(n_1828) );
AOI221xp5_ASAP7_75t_L g1848 ( .A1(n_193), .A2(n_221), .B1(n_664), .B2(n_748), .C(n_1040), .Y(n_1848) );
AOI22xp33_ASAP7_75t_L g1214 ( .A1(n_194), .A2(n_236), .B1(n_719), .B2(n_939), .Y(n_1214) );
AOI22xp33_ASAP7_75t_SL g1001 ( .A1(n_195), .A2(n_280), .B1(n_978), .B2(n_995), .Y(n_1001) );
AOI221xp5_ASAP7_75t_L g1008 ( .A1(n_195), .A2(n_291), .B1(n_534), .B2(n_819), .C(n_1009), .Y(n_1008) );
INVx2_ASAP7_75t_L g369 ( .A(n_196), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_196), .B(n_367), .Y(n_392) );
INVx1_ASAP7_75t_L g434 ( .A(n_196), .Y(n_434) );
INVx1_ASAP7_75t_L g974 ( .A(n_197), .Y(n_974) );
INVxp67_ASAP7_75t_L g847 ( .A(n_198), .Y(n_847) );
INVxp67_ASAP7_75t_SL g439 ( .A(n_199), .Y(n_439) );
AOI22xp33_ASAP7_75t_L g718 ( .A1(n_200), .A2(n_342), .B1(n_693), .B2(n_719), .Y(n_718) );
XOR2xp5_ASAP7_75t_L g543 ( .A(n_201), .B(n_544), .Y(n_543) );
INVx1_ASAP7_75t_L g1782 ( .A(n_202), .Y(n_1782) );
NAND2xp33_ASAP7_75t_SL g1801 ( .A(n_202), .B(n_512), .Y(n_1801) );
INVx1_ASAP7_75t_L g1226 ( .A(n_203), .Y(n_1226) );
OAI22xp33_ASAP7_75t_L g556 ( .A1(n_205), .A2(n_299), .B1(n_557), .B2(n_558), .Y(n_556) );
INVx1_ASAP7_75t_L g629 ( .A(n_205), .Y(n_629) );
INVx1_ASAP7_75t_L g1509 ( .A(n_206), .Y(n_1509) );
AOI21xp5_ASAP7_75t_L g1783 ( .A1(n_207), .A2(n_433), .B(n_751), .Y(n_1783) );
INVx1_ASAP7_75t_L g1803 ( .A(n_208), .Y(n_1803) );
CKINVDCx5p33_ASAP7_75t_R g1005 ( .A(n_209), .Y(n_1005) );
AOI22xp33_ASAP7_75t_L g1834 ( .A1(n_210), .A2(n_321), .B1(n_719), .B2(n_1835), .Y(n_1834) );
AOI22xp33_ASAP7_75t_L g1847 ( .A1(n_210), .A2(n_242), .B1(n_660), .B2(n_1188), .Y(n_1847) );
OAI22xp5_ASAP7_75t_L g644 ( .A1(n_211), .A2(n_292), .B1(n_645), .B2(n_647), .Y(n_644) );
OAI211xp5_ASAP7_75t_L g683 ( .A1(n_211), .A2(n_684), .B(n_687), .C(n_695), .Y(n_683) );
BUFx3_ASAP7_75t_L g361 ( .A(n_212), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_213), .B(n_496), .Y(n_495) );
INVx1_ASAP7_75t_L g410 ( .A(n_215), .Y(n_410) );
OAI21xp5_ASAP7_75t_SL g1022 ( .A1(n_216), .A2(n_794), .B(n_1023), .Y(n_1022) );
OAI221xp5_ASAP7_75t_L g1293 ( .A1(n_217), .A2(n_281), .B1(n_1103), .B2(n_1294), .C(n_1295), .Y(n_1293) );
OAI211xp5_ASAP7_75t_L g1299 ( .A1(n_217), .A2(n_893), .B(n_1300), .C(n_1303), .Y(n_1299) );
INVx1_ASAP7_75t_L g1824 ( .A(n_218), .Y(n_1824) );
CKINVDCx5p33_ASAP7_75t_R g1280 ( .A(n_219), .Y(n_1280) );
OAI221xp5_ASAP7_75t_SL g1450 ( .A1(n_220), .A2(n_316), .B1(n_1451), .B2(n_1453), .C(n_1454), .Y(n_1450) );
AOI22xp33_ASAP7_75t_L g1837 ( .A1(n_221), .A2(n_322), .B1(n_1016), .B2(n_1838), .Y(n_1837) );
OAI21xp5_ASAP7_75t_L g1172 ( .A1(n_222), .A2(n_645), .B(n_1173), .Y(n_1172) );
AOI22xp5_ASAP7_75t_L g1534 ( .A1(n_223), .A2(n_266), .B1(n_1535), .B2(n_1540), .Y(n_1534) );
INVx1_ASAP7_75t_L g1767 ( .A(n_225), .Y(n_1767) );
NOR2xp33_ASAP7_75t_L g1769 ( .A(n_225), .B(n_389), .Y(n_1769) );
OAI22xp33_ASAP7_75t_L g672 ( .A1(n_226), .A2(n_335), .B1(n_673), .B2(n_677), .Y(n_672) );
INVx1_ASAP7_75t_L g696 ( .A(n_226), .Y(n_696) );
INVx1_ASAP7_75t_L g1043 ( .A(n_227), .Y(n_1043) );
INVx1_ASAP7_75t_L g963 ( .A(n_228), .Y(n_963) );
INVx1_ASAP7_75t_L g754 ( .A(n_229), .Y(n_754) );
CKINVDCx5p33_ASAP7_75t_R g1090 ( .A(n_230), .Y(n_1090) );
CKINVDCx5p33_ASAP7_75t_R g1237 ( .A(n_231), .Y(n_1237) );
AOI22xp33_ASAP7_75t_L g667 ( .A1(n_233), .A2(n_251), .B1(n_664), .B2(n_668), .Y(n_667) );
INVx1_ASAP7_75t_L g711 ( .A(n_233), .Y(n_711) );
OAI221xp5_ASAP7_75t_L g564 ( .A1(n_234), .A2(n_256), .B1(n_375), .B2(n_565), .C(n_566), .Y(n_564) );
INVx1_ASAP7_75t_L g931 ( .A(n_235), .Y(n_931) );
INVx1_ASAP7_75t_L g447 ( .A(n_237), .Y(n_447) );
BUFx3_ASAP7_75t_L g518 ( .A(n_237), .Y(n_518) );
INVxp67_ASAP7_75t_SL g785 ( .A(n_238), .Y(n_785) );
INVx1_ASAP7_75t_L g1435 ( .A(n_239), .Y(n_1435) );
NOR2xp33_ASAP7_75t_L g1142 ( .A(n_243), .B(n_1143), .Y(n_1142) );
CKINVDCx5p33_ASAP7_75t_R g591 ( .A(n_244), .Y(n_591) );
OAI322xp33_ASAP7_75t_SL g1422 ( .A1(n_245), .A2(n_673), .A3(n_1330), .B1(n_1423), .B2(n_1427), .C1(n_1429), .C2(n_1434), .Y(n_1422) );
OAI22xp33_ASAP7_75t_SL g1459 ( .A1(n_245), .A2(n_250), .B1(n_1165), .B2(n_1460), .Y(n_1459) );
CKINVDCx5p33_ASAP7_75t_R g1473 ( .A(n_247), .Y(n_1473) );
INVx1_ASAP7_75t_L g1098 ( .A(n_248), .Y(n_1098) );
INVx1_ASAP7_75t_L g1780 ( .A(n_249), .Y(n_1780) );
CKINVDCx5p33_ASAP7_75t_R g1288 ( .A(n_252), .Y(n_1288) );
AOI221xp5_ASAP7_75t_L g873 ( .A1(n_253), .A2(n_319), .B1(n_551), .B2(n_874), .C(n_875), .Y(n_873) );
INVx1_ASAP7_75t_L g906 ( .A(n_253), .Y(n_906) );
INVx1_ASAP7_75t_L g877 ( .A(n_254), .Y(n_877) );
INVx1_ASAP7_75t_L g1438 ( .A(n_255), .Y(n_1438) );
OA222x2_ASAP7_75t_L g623 ( .A1(n_256), .A2(n_271), .B1(n_326), .B2(n_462), .C1(n_488), .C2(n_624), .Y(n_623) );
INVx1_ASAP7_75t_L g1332 ( .A(n_258), .Y(n_1332) );
INVx1_ASAP7_75t_L g1182 ( .A(n_259), .Y(n_1182) );
XOR2xp5_ASAP7_75t_L g868 ( .A(n_260), .B(n_869), .Y(n_868) );
OAI21xp5_ASAP7_75t_L g1222 ( .A1(n_261), .A2(n_794), .B(n_1223), .Y(n_1222) );
INVx1_ASAP7_75t_L g413 ( .A(n_262), .Y(n_413) );
CKINVDCx5p33_ASAP7_75t_R g1113 ( .A(n_263), .Y(n_1113) );
OAI22xp5_ASAP7_75t_SL g1413 ( .A1(n_266), .A2(n_1414), .B1(n_1415), .B2(n_1461), .Y(n_1413) );
INVx1_ASAP7_75t_L g1461 ( .A(n_266), .Y(n_1461) );
AOI22xp5_ASAP7_75t_L g1514 ( .A1(n_266), .A2(n_1414), .B1(n_1415), .B2(n_1461), .Y(n_1514) );
INVxp67_ASAP7_75t_SL g896 ( .A(n_268), .Y(n_896) );
INVx1_ASAP7_75t_L g364 ( .A(n_270), .Y(n_364) );
INVx1_ASAP7_75t_L g382 ( .A(n_270), .Y(n_382) );
INVx1_ASAP7_75t_L g561 ( .A(n_271), .Y(n_561) );
CKINVDCx5p33_ASAP7_75t_R g1235 ( .A(n_272), .Y(n_1235) );
INVx1_ASAP7_75t_L g1832 ( .A(n_273), .Y(n_1832) );
INVxp67_ASAP7_75t_SL g1857 ( .A(n_274), .Y(n_1857) );
INVx1_ASAP7_75t_L g899 ( .A(n_275), .Y(n_899) );
OAI22xp5_ASAP7_75t_L g872 ( .A1(n_276), .A2(n_313), .B1(n_417), .B2(n_420), .Y(n_872) );
INVx1_ASAP7_75t_L g897 ( .A(n_276), .Y(n_897) );
INVxp67_ASAP7_75t_SL g455 ( .A(n_277), .Y(n_455) );
AOI21xp33_ASAP7_75t_L g747 ( .A1(n_278), .A2(n_559), .B(n_748), .Y(n_747) );
INVxp67_ASAP7_75t_L g771 ( .A(n_278), .Y(n_771) );
INVx1_ASAP7_75t_L g1328 ( .A(n_279), .Y(n_1328) );
INVx1_ASAP7_75t_L g1052 ( .A(n_282), .Y(n_1052) );
NOR2xp33_ASAP7_75t_L g1055 ( .A(n_282), .B(n_760), .Y(n_1055) );
INVx1_ASAP7_75t_L g1271 ( .A(n_283), .Y(n_1271) );
CKINVDCx5p33_ASAP7_75t_R g1006 ( .A(n_284), .Y(n_1006) );
INVxp33_ASAP7_75t_L g838 ( .A(n_285), .Y(n_838) );
CKINVDCx5p33_ASAP7_75t_R g943 ( .A(n_286), .Y(n_943) );
CKINVDCx5p33_ASAP7_75t_R g1766 ( .A(n_287), .Y(n_1766) );
INVx1_ASAP7_75t_L g848 ( .A(n_288), .Y(n_848) );
INVx1_ASAP7_75t_L g1118 ( .A(n_289), .Y(n_1118) );
INVx1_ASAP7_75t_L g1539 ( .A(n_290), .Y(n_1539) );
AND2x2_ASAP7_75t_L g1544 ( .A(n_290), .B(n_1538), .Y(n_1544) );
AOI21xp33_ASAP7_75t_L g714 ( .A1(n_293), .A2(n_602), .B(n_715), .Y(n_714) );
INVx1_ASAP7_75t_L g1325 ( .A(n_295), .Y(n_1325) );
INVx1_ASAP7_75t_L g1668 ( .A(n_296), .Y(n_1668) );
CKINVDCx16_ASAP7_75t_R g1786 ( .A(n_297), .Y(n_1786) );
XOR2x2_ASAP7_75t_L g726 ( .A(n_298), .B(n_727), .Y(n_726) );
INVx1_ASAP7_75t_L g628 ( .A(n_299), .Y(n_628) );
INVx1_ASAP7_75t_L g1504 ( .A(n_300), .Y(n_1504) );
INVx1_ASAP7_75t_L g1155 ( .A(n_302), .Y(n_1155) );
INVx1_ASAP7_75t_L g1220 ( .A(n_304), .Y(n_1220) );
INVxp67_ASAP7_75t_SL g1457 ( .A(n_305), .Y(n_1457) );
INVx1_ASAP7_75t_L g1099 ( .A(n_307), .Y(n_1099) );
OAI221xp5_ASAP7_75t_L g1132 ( .A1(n_307), .A2(n_488), .B1(n_610), .B2(n_1133), .C(n_1141), .Y(n_1132) );
AOI22xp33_ASAP7_75t_L g1850 ( .A1(n_310), .A2(n_321), .B1(n_1188), .B2(n_1190), .Y(n_1850) );
INVx1_ASAP7_75t_L g814 ( .A(n_311), .Y(n_814) );
INVxp67_ASAP7_75t_SL g919 ( .A(n_313), .Y(n_919) );
BUFx6f_ASAP7_75t_L g450 ( .A(n_314), .Y(n_450) );
INVx1_ASAP7_75t_L g739 ( .A(n_315), .Y(n_739) );
INVxp67_ASAP7_75t_SL g1417 ( .A(n_316), .Y(n_1417) );
CKINVDCx5p33_ASAP7_75t_R g988 ( .A(n_317), .Y(n_988) );
CKINVDCx5p33_ASAP7_75t_R g1285 ( .A(n_318), .Y(n_1285) );
INVx1_ASAP7_75t_L g913 ( .A(n_319), .Y(n_913) );
NOR2xp33_ASAP7_75t_R g1796 ( .A(n_320), .B(n_488), .Y(n_1796) );
INVx1_ASAP7_75t_L g1762 ( .A(n_323), .Y(n_1762) );
AOI22xp33_ASAP7_75t_L g1809 ( .A1(n_323), .A2(n_1810), .B1(n_1814), .B2(n_1858), .Y(n_1809) );
AOI21xp33_ASAP7_75t_L g510 ( .A1(n_324), .A2(n_511), .B(n_514), .Y(n_510) );
INVx1_ASAP7_75t_L g1433 ( .A(n_325), .Y(n_1433) );
INVx1_ASAP7_75t_L g552 ( .A(n_326), .Y(n_552) );
CKINVDCx5p33_ASAP7_75t_R g1233 ( .A(n_327), .Y(n_1233) );
INVx1_ASAP7_75t_L g1081 ( .A(n_329), .Y(n_1081) );
XOR2xp5_ASAP7_75t_L g981 ( .A(n_330), .B(n_982), .Y(n_981) );
INVx2_ASAP7_75t_L g437 ( .A(n_331), .Y(n_437) );
INVx1_ASAP7_75t_L g444 ( .A(n_331), .Y(n_444) );
INVx1_ASAP7_75t_L g466 ( .A(n_331), .Y(n_466) );
XOR2x2_ASAP7_75t_L g1314 ( .A(n_332), .B(n_1315), .Y(n_1314) );
INVx1_ASAP7_75t_L g883 ( .A(n_333), .Y(n_883) );
INVx1_ASAP7_75t_L g472 ( .A(n_334), .Y(n_472) );
INVx1_ASAP7_75t_L g698 ( .A(n_335), .Y(n_698) );
INVx1_ASAP7_75t_L g1274 ( .A(n_336), .Y(n_1274) );
CKINVDCx5p33_ASAP7_75t_R g1101 ( .A(n_338), .Y(n_1101) );
INVxp67_ASAP7_75t_SL g766 ( .A(n_339), .Y(n_766) );
CKINVDCx5p33_ASAP7_75t_R g795 ( .A(n_340), .Y(n_795) );
INVx1_ASAP7_75t_L g1334 ( .A(n_341), .Y(n_1334) );
INVx1_ASAP7_75t_L g1426 ( .A(n_343), .Y(n_1426) );
AOI21xp5_ASAP7_75t_L g344 ( .A1(n_345), .A2(n_1515), .B(n_1527), .Y(n_344) );
XNOR2xp5_ASAP7_75t_L g345 ( .A(n_346), .B(n_1410), .Y(n_345) );
OAI22xp5_ASAP7_75t_L g346 ( .A1(n_347), .A2(n_348), .B1(n_1314), .B2(n_1409), .Y(n_346) );
INVx2_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
AOI22x1_ASAP7_75t_L g348 ( .A1(n_349), .A2(n_350), .B1(n_979), .B2(n_1312), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
XOR2x2_ASAP7_75t_L g350 ( .A(n_351), .B(n_788), .Y(n_350) );
OAI22xp5_ASAP7_75t_L g351 ( .A1(n_352), .A2(n_631), .B1(n_632), .B2(n_787), .Y(n_351) );
INVx1_ASAP7_75t_L g787 ( .A(n_352), .Y(n_787) );
AOI22xp5_ASAP7_75t_L g352 ( .A1(n_353), .A2(n_541), .B1(n_542), .B2(n_630), .Y(n_352) );
INVx2_ASAP7_75t_L g630 ( .A(n_353), .Y(n_630) );
NOR2x1_ASAP7_75t_L g354 ( .A(n_355), .B(n_453), .Y(n_354) );
A2O1A1Ixp33_ASAP7_75t_L g355 ( .A1(n_356), .A2(n_399), .B(n_435), .C(n_438), .Y(n_355) );
AOI211xp5_ASAP7_75t_SL g356 ( .A1(n_357), .A2(n_370), .B(n_371), .C(n_388), .Y(n_356) );
AOI211xp5_ASAP7_75t_L g729 ( .A1(n_357), .A2(n_730), .B(n_731), .C(n_732), .Y(n_729) );
AOI211xp5_ASAP7_75t_SL g884 ( .A1(n_357), .A2(n_885), .B(n_886), .C(n_887), .Y(n_884) );
AOI22xp33_ASAP7_75t_L g1046 ( .A1(n_357), .A2(n_1047), .B1(n_1049), .B2(n_1054), .Y(n_1046) );
AOI221xp5_ASAP7_75t_L g1257 ( .A1(n_357), .A2(n_548), .B1(n_1252), .B2(n_1258), .C(n_1259), .Y(n_1257) );
AOI221xp5_ASAP7_75t_L g1291 ( .A1(n_357), .A2(n_548), .B1(n_1292), .B2(n_1293), .C(n_1297), .Y(n_1291) );
INVx2_ASAP7_75t_L g1856 ( .A(n_357), .Y(n_1856) );
INVx2_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
OR2x2_ASAP7_75t_L g647 ( .A(n_358), .B(n_648), .Y(n_647) );
OR2x6_ASAP7_75t_L g859 ( .A(n_358), .B(n_648), .Y(n_859) );
NAND2x1p5_ASAP7_75t_L g358 ( .A(n_359), .B(n_365), .Y(n_358) );
BUFx3_ASAP7_75t_L g412 ( .A(n_359), .Y(n_412) );
AND2x2_ASAP7_75t_L g418 ( .A(n_359), .B(n_419), .Y(n_418) );
INVx8_ASAP7_75t_L g563 ( .A(n_359), .Y(n_563) );
BUFx3_ASAP7_75t_L g751 ( .A(n_359), .Y(n_751) );
HB1xp67_ASAP7_75t_L g1202 ( .A(n_359), .Y(n_1202) );
AND2x4_ASAP7_75t_L g359 ( .A(n_360), .B(n_362), .Y(n_359) );
AND2x4_ASAP7_75t_L g394 ( .A(n_360), .B(n_395), .Y(n_394) );
INVx2_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
BUFx6f_ASAP7_75t_L g376 ( .A(n_361), .Y(n_376) );
AND2x4_ASAP7_75t_L g422 ( .A(n_361), .B(n_381), .Y(n_422) );
OR2x2_ASAP7_75t_L g430 ( .A(n_361), .B(n_363), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_361), .B(n_382), .Y(n_576) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVxp67_ASAP7_75t_L g395 ( .A(n_364), .Y(n_395) );
AND2x6_ASAP7_75t_L g373 ( .A(n_365), .B(n_374), .Y(n_373) );
AND2x2_ASAP7_75t_L g378 ( .A(n_365), .B(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g387 ( .A(n_365), .Y(n_387) );
AND2x4_ASAP7_75t_L g654 ( .A(n_365), .B(n_522), .Y(n_654) );
AND2x4_ASAP7_75t_L g365 ( .A(n_366), .B(n_368), .Y(n_365) );
NAND2x1p5_ASAP7_75t_L g433 ( .A(n_366), .B(n_434), .Y(n_433) );
NAND3x1_ASAP7_75t_L g854 ( .A(n_366), .B(n_434), .C(n_855), .Y(n_854) );
OR2x4_ASAP7_75t_L g1381 ( .A(n_366), .B(n_430), .Y(n_1381) );
INVx1_ASAP7_75t_L g1384 ( .A(n_366), .Y(n_1384) );
AND2x4_ASAP7_75t_L g1387 ( .A(n_366), .B(n_422), .Y(n_1387) );
OR2x6_ASAP7_75t_L g1402 ( .A(n_366), .B(n_575), .Y(n_1402) );
INVx3_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
BUFx3_ASAP7_75t_L g415 ( .A(n_367), .Y(n_415) );
NAND2xp33_ASAP7_75t_SL g749 ( .A(n_367), .B(n_369), .Y(n_749) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
AND2x2_ASAP7_75t_L g414 ( .A(n_369), .B(n_415), .Y(n_414) );
AND3x4_ASAP7_75t_L g662 ( .A(n_369), .B(n_415), .C(n_436), .Y(n_662) );
HB1xp67_ASAP7_75t_L g1406 ( .A(n_369), .Y(n_1406) );
INVx4_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
AOI221xp5_ASAP7_75t_L g1042 ( .A1(n_373), .A2(n_378), .B1(n_1043), .B2(n_1044), .C(n_1045), .Y(n_1042) );
AOI22xp33_ASAP7_75t_L g1097 ( .A1(n_373), .A2(n_378), .B1(n_1098), .B2(n_1099), .Y(n_1097) );
AND2x2_ASAP7_75t_L g653 ( .A(n_374), .B(n_654), .Y(n_653) );
NAND2x1_ASAP7_75t_L g865 ( .A(n_374), .B(n_654), .Y(n_865) );
AND2x4_ASAP7_75t_SL g970 ( .A(n_374), .B(n_654), .Y(n_970) );
INVx3_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx2_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
NAND2x1p5_ASAP7_75t_L g385 ( .A(n_376), .B(n_386), .Y(n_385) );
AND2x4_ASAP7_75t_L g398 ( .A(n_376), .B(n_380), .Y(n_398) );
BUFx2_ASAP7_75t_L g1392 ( .A(n_376), .Y(n_1392) );
INVx2_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
HB1xp67_ASAP7_75t_L g1845 ( .A(n_378), .Y(n_1845) );
INVx1_ASAP7_75t_L g565 ( .A(n_379), .Y(n_565) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx2_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g386 ( .A(n_382), .Y(n_386) );
CKINVDCx5p33_ASAP7_75t_R g1045 ( .A(n_383), .Y(n_1045) );
OAI221xp5_ASAP7_75t_L g1770 ( .A1(n_383), .A2(n_1771), .B1(n_1775), .B2(n_1778), .C(n_1781), .Y(n_1770) );
OR2x6_ASAP7_75t_L g383 ( .A(n_384), .B(n_387), .Y(n_383) );
INVx1_ASAP7_75t_L g426 ( .A(n_384), .Y(n_426) );
OAI221xp5_ASAP7_75t_L g1284 ( .A1(n_384), .A2(n_432), .B1(n_841), .B2(n_1285), .C(n_1286), .Y(n_1284) );
OAI221xp5_ASAP7_75t_L g1775 ( .A1(n_384), .A2(n_414), .B1(n_1050), .B2(n_1776), .C(n_1777), .Y(n_1775) );
BUFx2_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
BUFx6f_ASAP7_75t_L g407 ( .A(n_385), .Y(n_407) );
BUFx3_ASAP7_75t_L g876 ( .A(n_385), .Y(n_876) );
BUFx2_ASAP7_75t_L g1395 ( .A(n_386), .Y(n_1395) );
INVx1_ASAP7_75t_L g567 ( .A(n_387), .Y(n_567) );
CKINVDCx5p33_ASAP7_75t_R g753 ( .A(n_389), .Y(n_753) );
OR2x6_ASAP7_75t_SL g389 ( .A(n_390), .B(n_393), .Y(n_389) );
INVx2_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
AND2x4_ASAP7_75t_L g397 ( .A(n_391), .B(n_398), .Y(n_397) );
HB1xp67_ASAP7_75t_L g549 ( .A(n_391), .Y(n_549) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
INVx1_ASAP7_75t_L g419 ( .A(n_392), .Y(n_419) );
OR2x2_ASAP7_75t_L g642 ( .A(n_392), .B(n_530), .Y(n_642) );
INVx1_ASAP7_75t_L g832 ( .A(n_393), .Y(n_832) );
INVx3_ASAP7_75t_L g1175 ( .A(n_393), .Y(n_1175) );
BUFx2_ASAP7_75t_L g1327 ( .A(n_393), .Y(n_1327) );
INVx2_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
BUFx6f_ASAP7_75t_L g403 ( .A(n_394), .Y(n_403) );
BUFx8_ASAP7_75t_L g431 ( .A(n_394), .Y(n_431) );
BUFx6f_ASAP7_75t_L g559 ( .A(n_394), .Y(n_559) );
INVx3_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
AOI221xp5_ASAP7_75t_L g752 ( .A1(n_397), .A2(n_753), .B1(n_754), .B2(n_755), .C(n_756), .Y(n_752) );
NAND2xp5_ASAP7_75t_L g1145 ( .A(n_397), .B(n_598), .Y(n_1145) );
INVx5_ASAP7_75t_L g409 ( .A(n_398), .Y(n_409) );
BUFx3_ASAP7_75t_L g551 ( .A(n_398), .Y(n_551) );
BUFx3_ASAP7_75t_L g999 ( .A(n_398), .Y(n_999) );
BUFx2_ASAP7_75t_L g1034 ( .A(n_398), .Y(n_1034) );
BUFx12f_ASAP7_75t_L g1188 ( .A(n_398), .Y(n_1188) );
NOR3xp33_ASAP7_75t_SL g399 ( .A(n_400), .B(n_416), .C(n_423), .Y(n_399) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
BUFx6f_ASAP7_75t_L g594 ( .A(n_403), .Y(n_594) );
BUFx6f_ASAP7_75t_L g846 ( .A(n_403), .Y(n_846) );
INVx2_ASAP7_75t_L g1282 ( .A(n_403), .Y(n_1282) );
INVx2_ASAP7_75t_L g1324 ( .A(n_403), .Y(n_1324) );
AND2x4_ASAP7_75t_L g1383 ( .A(n_403), .B(n_1384), .Y(n_1383) );
INVx2_ASAP7_75t_L g1853 ( .A(n_403), .Y(n_1853) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx2_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g579 ( .A(n_406), .Y(n_579) );
INVx1_ASAP7_75t_L g592 ( .A(n_406), .Y(n_592) );
INVx4_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
BUFx6f_ASAP7_75t_L g566 ( .A(n_407), .Y(n_566) );
OR2x2_ASAP7_75t_L g646 ( .A(n_407), .B(n_642), .Y(n_646) );
INVx3_ASAP7_75t_L g746 ( .A(n_407), .Y(n_746) );
OAI221xp5_ASAP7_75t_L g1279 ( .A1(n_407), .A2(n_414), .B1(n_1280), .B2(n_1281), .C(n_1282), .Y(n_1279) );
OAI221xp5_ASAP7_75t_L g408 ( .A1(n_409), .A2(n_410), .B1(n_411), .B2(n_413), .C(n_414), .Y(n_408) );
INVx2_ASAP7_75t_L g666 ( .A(n_409), .Y(n_666) );
INVx2_ASAP7_75t_R g668 ( .A(n_409), .Y(n_668) );
INVx1_ASAP7_75t_L g1108 ( .A(n_409), .Y(n_1108) );
OAI22xp5_ASAP7_75t_L g536 ( .A1(n_410), .A2(n_537), .B1(n_539), .B2(n_540), .Y(n_536) );
INVx2_ASAP7_75t_L g1033 ( .A(n_411), .Y(n_1033) );
INVx2_ASAP7_75t_SL g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g994 ( .A(n_412), .Y(n_994) );
NAND2xp5_ASAP7_75t_L g1295 ( .A(n_412), .B(n_1296), .Y(n_1295) );
OAI22xp5_ASAP7_75t_L g499 ( .A1(n_413), .A2(n_500), .B1(n_504), .B2(n_505), .Y(n_499) );
OAI221xp5_ASAP7_75t_L g590 ( .A1(n_414), .A2(n_591), .B1(n_592), .B2(n_593), .C(n_595), .Y(n_590) );
OAI221xp5_ASAP7_75t_L g875 ( .A1(n_414), .A2(n_558), .B1(n_876), .B2(n_877), .C(n_878), .Y(n_875) );
OAI221xp5_ASAP7_75t_L g1264 ( .A1(n_414), .A2(n_876), .B1(n_1237), .B2(n_1241), .C(n_1265), .Y(n_1264) );
INVx3_ASAP7_75t_L g1391 ( .A(n_415), .Y(n_1391) );
INVx2_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
AND2x2_ASAP7_75t_L g421 ( .A(n_419), .B(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx2_ASAP7_75t_L g554 ( .A(n_422), .Y(n_554) );
BUFx2_ASAP7_75t_L g661 ( .A(n_422), .Y(n_661) );
BUFx2_ASAP7_75t_L g681 ( .A(n_422), .Y(n_681) );
BUFx2_ASAP7_75t_L g850 ( .A(n_422), .Y(n_850) );
BUFx2_ASAP7_75t_L g995 ( .A(n_422), .Y(n_995) );
BUFx3_ASAP7_75t_L g1040 ( .A(n_422), .Y(n_1040) );
BUFx2_ASAP7_75t_L g1440 ( .A(n_422), .Y(n_1440) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_428), .B(n_432), .Y(n_427) );
INVx3_ASAP7_75t_L g585 ( .A(n_429), .Y(n_585) );
INVx2_ASAP7_75t_SL g674 ( .A(n_429), .Y(n_674) );
INVx2_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
BUFx3_ASAP7_75t_L g557 ( .A(n_430), .Y(n_557) );
BUFx3_ASAP7_75t_L g580 ( .A(n_430), .Y(n_580) );
BUFx4f_ASAP7_75t_L g841 ( .A(n_430), .Y(n_841) );
OR2x4_ASAP7_75t_L g1400 ( .A(n_430), .B(n_1384), .Y(n_1400) );
AND2x4_ASAP7_75t_L g678 ( .A(n_431), .B(n_679), .Y(n_678) );
INVx2_ASAP7_75t_SL g738 ( .A(n_431), .Y(n_738) );
INVx3_ASAP7_75t_L g954 ( .A(n_431), .Y(n_954) );
INVx3_ASAP7_75t_L g1106 ( .A(n_431), .Y(n_1106) );
INVx2_ASAP7_75t_SL g1116 ( .A(n_431), .Y(n_1116) );
OAI221xp5_ASAP7_75t_L g577 ( .A1(n_432), .A2(n_578), .B1(n_579), .B2(n_580), .C(n_581), .Y(n_577) );
INVx3_ASAP7_75t_L g736 ( .A(n_432), .Y(n_736) );
OAI221xp5_ASAP7_75t_L g881 ( .A1(n_432), .A2(n_841), .B1(n_876), .B2(n_882), .C(n_883), .Y(n_881) );
OAI221xp5_ASAP7_75t_L g1110 ( .A1(n_432), .A2(n_839), .B1(n_1111), .B2(n_1113), .C(n_1114), .Y(n_1110) );
OAI221xp5_ASAP7_75t_L g1267 ( .A1(n_432), .A2(n_557), .B1(n_876), .B2(n_1233), .C(n_1242), .Y(n_1267) );
INVx3_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
OR2x6_ASAP7_75t_L g670 ( .A(n_433), .B(n_516), .Y(n_670) );
OR2x2_ASAP7_75t_L g1513 ( .A(n_433), .B(n_516), .Y(n_1513) );
INVx2_ASAP7_75t_SL g435 ( .A(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g724 ( .A(n_436), .Y(n_724) );
OAI31xp33_ASAP7_75t_L g1768 ( .A1(n_436), .A2(n_1769), .A3(n_1770), .B(n_1784), .Y(n_1768) );
AOI22xp33_ASAP7_75t_SL g1840 ( .A1(n_436), .A2(n_892), .B1(n_1841), .B2(n_1857), .Y(n_1840) );
INVx2_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_437), .B(n_477), .Y(n_476) );
BUFx2_ASAP7_75t_L g516 ( .A(n_437), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_439), .B(n_440), .Y(n_438) );
AOI22xp33_ASAP7_75t_SL g627 ( .A1(n_440), .A2(n_456), .B1(n_628), .B2(n_629), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g786 ( .A(n_440), .B(n_754), .Y(n_786) );
INVx1_ASAP7_75t_L g893 ( .A(n_440), .Y(n_893) );
HB1xp67_ASAP7_75t_L g1061 ( .A(n_440), .Y(n_1061) );
AOI222xp33_ASAP7_75t_L g1086 ( .A1(n_440), .A2(n_456), .B1(n_1087), .B2(n_1088), .C1(n_1090), .C2(n_1091), .Y(n_1086) );
NAND2xp33_ASAP7_75t_SL g1270 ( .A(n_440), .B(n_1271), .Y(n_1270) );
AOI22xp33_ASAP7_75t_L g1765 ( .A1(n_440), .A2(n_456), .B1(n_1766), .B2(n_1767), .Y(n_1765) );
AND2x4_ASAP7_75t_L g440 ( .A(n_441), .B(n_445), .Y(n_440) );
AND2x4_ASAP7_75t_L g456 ( .A(n_441), .B(n_457), .Y(n_456) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
OR2x2_ASAP7_75t_L g483 ( .A(n_442), .B(n_484), .Y(n_483) );
OR2x2_ASAP7_75t_L g622 ( .A(n_442), .B(n_484), .Y(n_622) );
INVxp67_ASAP7_75t_L g648 ( .A(n_442), .Y(n_648) );
INVx1_ASAP7_75t_L g1378 ( .A(n_442), .Y(n_1378) );
BUFx2_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx2_ASAP7_75t_L g530 ( .A(n_443), .Y(n_530) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
AND2x2_ASAP7_75t_L g445 ( .A(n_446), .B(n_448), .Y(n_445) );
AND2x2_ASAP7_75t_L g457 ( .A(n_446), .B(n_458), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_446), .B(n_466), .Y(n_465) );
AND2x4_ASAP7_75t_L g685 ( .A(n_446), .B(n_686), .Y(n_685) );
AND2x4_ASAP7_75t_L g699 ( .A(n_446), .B(n_448), .Y(n_699) );
AND2x4_ASAP7_75t_SL g704 ( .A(n_446), .B(n_512), .Y(n_704) );
AND2x2_ASAP7_75t_L g928 ( .A(n_446), .B(n_467), .Y(n_928) );
BUFx2_ASAP7_75t_L g1475 ( .A(n_446), .Y(n_1475) );
HB1xp67_ASAP7_75t_L g1364 ( .A(n_447), .Y(n_1364) );
BUFx6f_ASAP7_75t_L g497 ( .A(n_448), .Y(n_497) );
INVx2_ASAP7_75t_L g801 ( .A(n_448), .Y(n_801) );
BUFx6f_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
BUFx3_ASAP7_75t_L g535 ( .A(n_449), .Y(n_535) );
INVx2_ASAP7_75t_L g605 ( .A(n_449), .Y(n_605) );
AND2x4_ASAP7_75t_L g1374 ( .A(n_449), .B(n_1364), .Y(n_1374) );
AND2x2_ASAP7_75t_L g449 ( .A(n_450), .B(n_451), .Y(n_449) );
INVx2_ASAP7_75t_L g459 ( .A(n_450), .Y(n_459) );
INVx2_ASAP7_75t_L g470 ( .A(n_450), .Y(n_470) );
INVx1_ASAP7_75t_L g486 ( .A(n_450), .Y(n_486) );
NAND2x1_ASAP7_75t_L g490 ( .A(n_450), .B(n_452), .Y(n_490) );
OR2x2_ASAP7_75t_L g503 ( .A(n_450), .B(n_452), .Y(n_503) );
AND2x2_ASAP7_75t_L g513 ( .A(n_450), .B(n_452), .Y(n_513) );
INVx2_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx1_ASAP7_75t_L g460 ( .A(n_452), .Y(n_460) );
AND2x2_ASAP7_75t_L g469 ( .A(n_452), .B(n_470), .Y(n_469) );
BUFx2_ASAP7_75t_L g480 ( .A(n_452), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_452), .B(n_470), .Y(n_509) );
OR2x2_ASAP7_75t_L g614 ( .A(n_452), .B(n_459), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_454), .B(n_494), .Y(n_453) );
AOI211xp5_ASAP7_75t_L g454 ( .A1(n_455), .A2(n_456), .B(n_461), .C(n_487), .Y(n_454) );
INVx3_ASAP7_75t_L g760 ( .A(n_456), .Y(n_760) );
NAND2xp5_ASAP7_75t_L g918 ( .A(n_456), .B(n_919), .Y(n_918) );
NAND2xp5_ASAP7_75t_L g1254 ( .A(n_456), .B(n_1255), .Y(n_1254) );
NAND2xp5_ASAP7_75t_L g1298 ( .A(n_456), .B(n_1296), .Y(n_1298) );
NAND2xp5_ASAP7_75t_L g1819 ( .A(n_456), .B(n_1820), .Y(n_1819) );
BUFx6f_ASAP7_75t_L g697 ( .A(n_457), .Y(n_697) );
INVx1_ASAP7_75t_L g810 ( .A(n_457), .Y(n_810) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_458), .B(n_477), .Y(n_524) );
INVx3_ASAP7_75t_L g618 ( .A(n_458), .Y(n_618) );
BUFx6f_ASAP7_75t_L g720 ( .A(n_458), .Y(n_720) );
AND2x2_ASAP7_75t_L g458 ( .A(n_459), .B(n_460), .Y(n_458) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
AOI222xp33_ASAP7_75t_L g782 ( .A1(n_463), .A2(n_520), .B1(n_730), .B2(n_755), .C1(n_783), .C2(n_785), .Y(n_782) );
AOI222xp33_ASAP7_75t_L g895 ( .A1(n_463), .A2(n_473), .B1(n_482), .B2(n_885), .C1(n_896), .C2(n_897), .Y(n_895) );
INVxp67_ASAP7_75t_L g1058 ( .A(n_463), .Y(n_1058) );
INVx1_ASAP7_75t_L g1089 ( .A(n_463), .Y(n_1089) );
AOI222xp33_ASAP7_75t_L g1250 ( .A1(n_463), .A2(n_520), .B1(n_783), .B2(n_1251), .C1(n_1252), .C2(n_1253), .Y(n_1250) );
AOI22xp33_ASAP7_75t_L g1823 ( .A1(n_463), .A2(n_783), .B1(n_1824), .B2(n_1825), .Y(n_1823) );
AND2x4_ASAP7_75t_L g463 ( .A(n_464), .B(n_467), .Y(n_463) );
AOI332xp33_ASAP7_75t_L g1300 ( .A1(n_464), .A2(n_467), .A3(n_521), .B1(n_523), .B2(n_783), .B3(n_1292), .C1(n_1301), .C2(n_1302), .Y(n_1300) );
INVx1_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
OR2x2_ASAP7_75t_L g488 ( .A(n_465), .B(n_489), .Y(n_488) );
OR2x2_ASAP7_75t_L g784 ( .A(n_465), .B(n_489), .Y(n_784) );
INVx1_ASAP7_75t_L g522 ( .A(n_466), .Y(n_522) );
INVx1_ASAP7_75t_L g855 ( .A(n_466), .Y(n_855) );
INVx3_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx1_ASAP7_75t_L g949 ( .A(n_468), .Y(n_949) );
INVx2_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
BUFx6f_ASAP7_75t_L g686 ( .A(n_469), .Y(n_686) );
BUFx3_ASAP7_75t_L g805 ( .A(n_469), .Y(n_805) );
BUFx3_ASAP7_75t_L g939 ( .A(n_469), .Y(n_939) );
AOI22xp5_ASAP7_75t_L g471 ( .A1(n_472), .A2(n_473), .B1(n_481), .B2(n_482), .Y(n_471) );
AOI22xp5_ASAP7_75t_L g1141 ( .A1(n_473), .A2(n_482), .B1(n_1096), .B2(n_1098), .Y(n_1141) );
AOI22xp33_ASAP7_75t_SL g1830 ( .A1(n_473), .A2(n_482), .B1(n_1831), .B2(n_1832), .Y(n_1830) );
INVx1_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
INVx2_ASAP7_75t_SL g621 ( .A(n_474), .Y(n_621) );
NAND2x2_ASAP7_75t_L g474 ( .A(n_475), .B(n_478), .Y(n_474) );
INVx1_ASAP7_75t_L g493 ( .A(n_475), .Y(n_493) );
INVx2_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_477), .B(n_485), .Y(n_484) );
AND2x6_ASAP7_75t_L g694 ( .A(n_477), .B(n_512), .Y(n_694) );
INVx1_ASAP7_75t_L g709 ( .A(n_477), .Y(n_709) );
AND2x2_ASAP7_75t_L g806 ( .A(n_477), .B(n_807), .Y(n_806) );
INVx2_ASAP7_75t_SL g478 ( .A(n_479), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
INVx1_ASAP7_75t_L g708 ( .A(n_480), .Y(n_708) );
BUFx2_ASAP7_75t_L g807 ( .A(n_480), .Y(n_807) );
AND2x4_ASAP7_75t_L g1355 ( .A(n_480), .B(n_1356), .Y(n_1355) );
INVx2_ASAP7_75t_SL g482 ( .A(n_483), .Y(n_482) );
AND2x4_ASAP7_75t_L g645 ( .A(n_483), .B(n_646), .Y(n_645) );
AND2x4_ASAP7_75t_L g794 ( .A(n_483), .B(n_646), .Y(n_794) );
INVx1_ASAP7_75t_L g1482 ( .A(n_484), .Y(n_1482) );
AND2x4_ASAP7_75t_L g1360 ( .A(n_485), .B(n_518), .Y(n_1360) );
INVx1_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
BUFx3_ASAP7_75t_L g608 ( .A(n_489), .Y(n_608) );
BUFx3_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
BUFx6f_ASAP7_75t_L g492 ( .A(n_490), .Y(n_492) );
OAI21xp5_ASAP7_75t_L g609 ( .A1(n_491), .A2(n_610), .B(n_611), .Y(n_609) );
CKINVDCx5p33_ASAP7_75t_R g922 ( .A(n_491), .Y(n_922) );
OAI21xp5_ASAP7_75t_L g1069 ( .A1(n_491), .A2(n_1070), .B(n_1078), .Y(n_1069) );
OAI21xp5_ASAP7_75t_SL g1120 ( .A1(n_491), .A2(n_1121), .B(n_1125), .Y(n_1120) );
OAI21xp5_ASAP7_75t_L g1797 ( .A1(n_491), .A2(n_779), .B(n_1798), .Y(n_1797) );
OR2x6_ASAP7_75t_L g491 ( .A(n_492), .B(n_493), .Y(n_491) );
INVx4_ASAP7_75t_L g713 ( .A(n_492), .Y(n_713) );
BUFx6f_ASAP7_75t_L g774 ( .A(n_492), .Y(n_774) );
BUFx4f_ASAP7_75t_L g944 ( .A(n_492), .Y(n_944) );
BUFx4f_ASAP7_75t_L g1129 ( .A(n_492), .Y(n_1129) );
BUFx4f_ASAP7_75t_L g1137 ( .A(n_492), .Y(n_1137) );
AOI322xp5_ASAP7_75t_L g494 ( .A1(n_495), .A2(n_498), .A3(n_510), .B1(n_519), .B2(n_520), .C1(n_525), .C2(n_531), .Y(n_494) );
BUFx3_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
INVx1_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
OAI22xp5_ASAP7_75t_L g1231 ( .A1(n_500), .A2(n_917), .B1(n_1232), .B2(n_1233), .Y(n_1231) );
BUFx4f_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
INVx1_ASAP7_75t_L g915 ( .A(n_501), .Y(n_915) );
INVxp67_ASAP7_75t_L g1245 ( .A(n_501), .Y(n_1245) );
OR2x6_ASAP7_75t_L g1363 ( .A(n_501), .B(n_1364), .Y(n_1363) );
OR2x6_ASAP7_75t_L g1371 ( .A(n_501), .B(n_1372), .Y(n_1371) );
INVx2_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
INVx3_ASAP7_75t_L g538 ( .A(n_502), .Y(n_538) );
BUFx4f_ASAP7_75t_L g908 ( .A(n_502), .Y(n_908) );
INVx3_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
INVx5_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
INVx6_ASAP7_75t_L g615 ( .A(n_506), .Y(n_615) );
BUFx6f_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
INVx2_ASAP7_75t_L g540 ( .A(n_507), .Y(n_540) );
INVx4_ASAP7_75t_L g909 ( .A(n_507), .Y(n_909) );
INVx2_ASAP7_75t_SL g917 ( .A(n_507), .Y(n_917) );
INVx1_ASAP7_75t_L g1163 ( .A(n_507), .Y(n_1163) );
INVx8_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
BUFx2_ASAP7_75t_L g769 ( .A(n_508), .Y(n_769) );
OR2x2_ASAP7_75t_L g1367 ( .A(n_508), .B(n_1356), .Y(n_1367) );
BUFx6f_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
AOI22xp33_ASAP7_75t_L g1472 ( .A1(n_511), .A2(n_805), .B1(n_1473), .B2(n_1474), .Y(n_1472) );
A2O1A1Ixp33_ASAP7_75t_L g1477 ( .A1(n_511), .A2(n_1139), .B(n_1478), .C(n_1479), .Y(n_1477) );
BUFx3_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
BUFx6f_ASAP7_75t_L g533 ( .A(n_512), .Y(n_533) );
BUFx3_ASAP7_75t_L g689 ( .A(n_512), .Y(n_689) );
INVx1_ASAP7_75t_L g902 ( .A(n_512), .Y(n_902) );
BUFx3_ASAP7_75t_L g911 ( .A(n_512), .Y(n_911) );
BUFx3_ASAP7_75t_L g934 ( .A(n_512), .Y(n_934) );
AND2x2_ASAP7_75t_L g1351 ( .A(n_512), .B(n_1352), .Y(n_1351) );
BUFx6f_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
INVx1_ASAP7_75t_L g1012 ( .A(n_513), .Y(n_1012) );
OAI33xp33_ASAP7_75t_L g1335 ( .A1(n_514), .A2(n_1336), .A3(n_1340), .B1(n_1342), .B2(n_1343), .B3(n_1345), .Y(n_1335) );
INVx2_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
HB1xp67_ASAP7_75t_L g600 ( .A(n_515), .Y(n_600) );
INVx2_ASAP7_75t_L g764 ( .A(n_515), .Y(n_764) );
AOI222xp33_ASAP7_75t_L g898 ( .A1(n_515), .A2(n_520), .B1(n_525), .B2(n_899), .C1(n_900), .C2(n_910), .Y(n_898) );
INVx2_ASAP7_75t_L g1079 ( .A(n_515), .Y(n_1079) );
INVx4_ASAP7_75t_L g1124 ( .A(n_515), .Y(n_1124) );
NAND2xp5_ASAP7_75t_L g1790 ( .A(n_515), .B(n_1791), .Y(n_1790) );
AOI31xp33_ASAP7_75t_L g1827 ( .A1(n_515), .A2(n_922), .A3(n_1828), .B(n_1829), .Y(n_1827) );
AND2x4_ASAP7_75t_L g515 ( .A(n_516), .B(n_517), .Y(n_515) );
INVx1_ASAP7_75t_L g598 ( .A(n_516), .Y(n_598) );
AND2x4_ASAP7_75t_L g526 ( .A(n_518), .B(n_527), .Y(n_526) );
INVx2_ASAP7_75t_L g717 ( .A(n_518), .Y(n_717) );
BUFx2_ASAP7_75t_L g1356 ( .A(n_518), .Y(n_1356) );
AND2x4_ASAP7_75t_L g520 ( .A(n_521), .B(n_523), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
OR2x2_ASAP7_75t_L g626 ( .A(n_522), .B(n_524), .Y(n_626) );
INVx1_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
CKINVDCx5p33_ASAP7_75t_R g610 ( .A(n_525), .Y(n_610) );
AOI211xp5_ASAP7_75t_L g1062 ( .A1(n_525), .A2(n_1063), .B(n_1069), .C(n_1080), .Y(n_1062) );
NAND3xp33_ASAP7_75t_L g1833 ( .A(n_525), .B(n_1834), .C(n_1837), .Y(n_1833) );
AND2x4_ASAP7_75t_L g525 ( .A(n_526), .B(n_528), .Y(n_525) );
INVx1_ASAP7_75t_SL g690 ( .A(n_526), .Y(n_690) );
AND2x2_ASAP7_75t_SL g780 ( .A(n_526), .B(n_530), .Y(n_780) );
INVx4_ASAP7_75t_L g819 ( .A(n_526), .Y(n_819) );
INVx4_ASAP7_75t_L g936 ( .A(n_526), .Y(n_936) );
NAND2xp5_ASAP7_75t_L g1307 ( .A(n_526), .B(n_528), .Y(n_1307) );
AND2x4_ASAP7_75t_L g716 ( .A(n_527), .B(n_717), .Y(n_716) );
INVx1_ASAP7_75t_L g1377 ( .A(n_527), .Y(n_1377) );
INVx1_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
OR2x2_ASAP7_75t_L g836 ( .A(n_530), .B(n_749), .Y(n_836) );
HB1xp67_ASAP7_75t_L g1408 ( .A(n_530), .Y(n_1408) );
BUFx2_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
BUFx2_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
INVx1_ASAP7_75t_L g904 ( .A(n_535), .Y(n_904) );
BUFx3_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
BUFx3_ASAP7_75t_L g607 ( .A(n_538), .Y(n_607) );
BUFx6f_ASAP7_75t_L g767 ( .A(n_538), .Y(n_767) );
INVx2_ASAP7_75t_SL g777 ( .A(n_538), .Y(n_777) );
INVx2_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
NAND4xp75_ASAP7_75t_L g544 ( .A(n_545), .B(n_599), .C(n_623), .D(n_627), .Y(n_544) );
OAI21x1_ASAP7_75t_L g545 ( .A1(n_546), .A2(n_568), .B(n_596), .Y(n_545) );
OAI21xp5_ASAP7_75t_L g546 ( .A1(n_547), .A2(n_550), .B(n_560), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
AOI22xp33_ASAP7_75t_L g1851 ( .A1(n_548), .A2(n_1824), .B1(n_1852), .B2(n_1855), .Y(n_1851) );
BUFx2_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
INVx1_ASAP7_75t_L g1048 ( .A(n_549), .Y(n_1048) );
AOI221xp5_ASAP7_75t_SL g550 ( .A1(n_551), .A2(n_552), .B1(n_553), .B2(n_555), .C(n_556), .Y(n_550) );
INVx1_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
INVx2_ASAP7_75t_L g965 ( .A(n_554), .Y(n_965) );
INVx2_ASAP7_75t_L g1203 ( .A(n_554), .Y(n_1203) );
INVx1_ASAP7_75t_L g1431 ( .A(n_557), .Y(n_1431) );
INVx2_ASAP7_75t_L g997 ( .A(n_558), .Y(n_997) );
INVx2_ASAP7_75t_SL g558 ( .A(n_559), .Y(n_558) );
HB1xp67_ASAP7_75t_L g572 ( .A(n_559), .Y(n_572) );
INVx5_ASAP7_75t_L g665 ( .A(n_559), .Y(n_665) );
INVx2_ASAP7_75t_SL g1038 ( .A(n_559), .Y(n_1038) );
INVx3_ASAP7_75t_L g1050 ( .A(n_559), .Y(n_1050) );
A2O1A1Ixp33_ASAP7_75t_L g560 ( .A1(n_561), .A2(n_562), .B(n_564), .C(n_567), .Y(n_560) );
AOI22xp33_ASAP7_75t_L g1854 ( .A1(n_562), .A2(n_681), .B1(n_1820), .B2(n_1832), .Y(n_1854) );
INVx3_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
INVx8_ASAP7_75t_L g660 ( .A(n_563), .Y(n_660) );
INVx2_ASAP7_75t_L g874 ( .A(n_563), .Y(n_874) );
INVx2_ASAP7_75t_L g978 ( .A(n_563), .Y(n_978) );
INVx2_ASAP7_75t_L g657 ( .A(n_565), .Y(n_657) );
OAI22xp33_ASAP7_75t_L g1319 ( .A1(n_566), .A2(n_839), .B1(n_1320), .B2(n_1321), .Y(n_1319) );
OAI22xp33_ASAP7_75t_L g1500 ( .A1(n_566), .A2(n_841), .B1(n_1501), .B2(n_1502), .Y(n_1500) );
OAI22xp5_ASAP7_75t_L g568 ( .A1(n_569), .A2(n_577), .B1(n_582), .B2(n_590), .Y(n_568) );
OAI22xp5_ASAP7_75t_L g569 ( .A1(n_570), .A2(n_571), .B1(n_573), .B2(n_574), .Y(n_569) );
OAI22xp5_ASAP7_75t_L g606 ( .A1(n_570), .A2(n_583), .B1(n_607), .B2(n_608), .Y(n_606) );
INVx1_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
OAI221xp5_ASAP7_75t_L g611 ( .A1(n_573), .A2(n_591), .B1(n_612), .B2(n_615), .C(n_616), .Y(n_611) );
OAI221xp5_ASAP7_75t_L g844 ( .A1(n_574), .A2(n_845), .B1(n_847), .B2(n_848), .C(n_849), .Y(n_844) );
OAI22xp5_ASAP7_75t_L g1423 ( .A1(n_574), .A2(n_1424), .B1(n_1425), .B2(n_1426), .Y(n_1423) );
OAI221xp5_ASAP7_75t_L g1434 ( .A1(n_574), .A2(n_1435), .B1(n_1436), .B2(n_1438), .C(n_1439), .Y(n_1434) );
BUFx3_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
INVx1_ASAP7_75t_L g589 ( .A(n_575), .Y(n_589) );
BUFx2_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
INVx1_ASAP7_75t_L g641 ( .A(n_576), .Y(n_641) );
OAI22xp5_ASAP7_75t_L g582 ( .A1(n_583), .A2(n_584), .B1(n_586), .B2(n_587), .Y(n_582) );
BUFx4f_ASAP7_75t_SL g584 ( .A(n_585), .Y(n_584) );
OAI21xp33_ASAP7_75t_L g957 ( .A1(n_587), .A2(n_958), .B(n_959), .Y(n_957) );
INVx3_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
BUFx2_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
INVx1_ASAP7_75t_L g1505 ( .A(n_589), .Y(n_1505) );
OAI21xp33_ASAP7_75t_L g733 ( .A1(n_592), .A2(n_734), .B(n_735), .Y(n_733) );
OAI221xp5_ASAP7_75t_L g960 ( .A1(n_593), .A2(n_943), .B1(n_961), .B2(n_963), .C(n_964), .Y(n_960) );
INVx2_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
INVx1_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
BUFx2_ASAP7_75t_L g889 ( .A(n_598), .Y(n_889) );
AOI21xp5_ASAP7_75t_SL g1468 ( .A1(n_598), .A2(n_1469), .B(n_1484), .Y(n_1468) );
AOI211x1_ASAP7_75t_L g599 ( .A1(n_600), .A2(n_601), .B(n_609), .C(n_619), .Y(n_599) );
INVx2_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
INVx2_ASAP7_75t_L g1016 ( .A(n_603), .Y(n_1016) );
INVx2_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
INVx1_ASAP7_75t_L g817 ( .A(n_604), .Y(n_817) );
INVx2_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
INVx2_ASAP7_75t_L g1064 ( .A(n_605), .Y(n_1064) );
INVx1_ASAP7_75t_L g1338 ( .A(n_607), .Y(n_1338) );
OAI22xp5_ASAP7_75t_L g770 ( .A1(n_608), .A2(n_612), .B1(n_739), .B2(n_771), .Y(n_770) );
OAI22xp5_ASAP7_75t_L g1238 ( .A1(n_608), .A2(n_1239), .B1(n_1241), .B2(n_1242), .Y(n_1238) );
INVx2_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
INVx2_ASAP7_75t_L g1799 ( .A(n_613), .Y(n_1799) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
BUFx2_ASAP7_75t_L g773 ( .A(n_614), .Y(n_773) );
BUFx3_ASAP7_75t_L g1073 ( .A(n_614), .Y(n_1073) );
INVx2_ASAP7_75t_L g1127 ( .A(n_614), .Y(n_1127) );
BUFx2_ASAP7_75t_L g1136 ( .A(n_614), .Y(n_1136) );
OAI22xp33_ASAP7_75t_L g1065 ( .A1(n_615), .A2(n_1066), .B1(n_1067), .B2(n_1068), .Y(n_1065) );
INVx2_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
INVx2_ASAP7_75t_L g692 ( .A(n_618), .Y(n_692) );
INVx2_ASAP7_75t_SL g938 ( .A(n_618), .Y(n_938) );
INVx1_ASAP7_75t_L g948 ( .A(n_618), .Y(n_948) );
INVx2_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
AOI22xp5_ASAP7_75t_L g1793 ( .A1(n_621), .A2(n_1786), .B1(n_1794), .B2(n_1795), .Y(n_1793) );
INVx1_ASAP7_75t_SL g1794 ( .A(n_622), .Y(n_1794) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
AND2x4_ASAP7_75t_L g638 ( .A(n_626), .B(n_639), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g1144 ( .A(n_626), .B(n_1145), .Y(n_1144) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
AOI22xp5_ASAP7_75t_L g632 ( .A1(n_633), .A2(n_634), .B1(n_725), .B2(n_726), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
NAND3xp33_ASAP7_75t_SL g635 ( .A(n_636), .B(n_649), .C(n_682), .Y(n_635) );
AOI21xp33_ASAP7_75t_L g636 ( .A1(n_637), .A2(n_643), .B(n_644), .Y(n_636) );
AOI221xp5_ASAP7_75t_L g857 ( .A1(n_637), .A2(n_825), .B1(n_858), .B2(n_860), .C(n_861), .Y(n_857) );
AOI21xp5_ASAP7_75t_L g973 ( .A1(n_637), .A2(n_974), .B(n_975), .Y(n_973) );
AOI221xp5_ASAP7_75t_L g983 ( .A1(n_637), .A2(n_858), .B1(n_984), .B2(n_985), .C(n_986), .Y(n_983) );
NAND2xp5_ASAP7_75t_L g1177 ( .A(n_637), .B(n_1178), .Y(n_1177) );
AOI221xp5_ASAP7_75t_L g1196 ( .A1(n_637), .A2(n_858), .B1(n_1197), .B2(n_1198), .C(n_1199), .Y(n_1196) );
AOI21xp5_ASAP7_75t_L g1441 ( .A1(n_637), .A2(n_1442), .B(n_1443), .Y(n_1441) );
INVx8_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
OR2x2_ASAP7_75t_L g639 ( .A(n_640), .B(n_642), .Y(n_639) );
INVx1_ASAP7_75t_L g741 ( .A(n_640), .Y(n_741) );
BUFx3_ASAP7_75t_L g834 ( .A(n_640), .Y(n_834) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
BUFx6f_ASAP7_75t_L g962 ( .A(n_641), .Y(n_962) );
INVx1_ASAP7_75t_L g676 ( .A(n_642), .Y(n_676) );
INVx1_ASAP7_75t_L g679 ( .A(n_642), .Y(n_679) );
INVx2_ASAP7_75t_L g1494 ( .A(n_646), .Y(n_1494) );
NAND2xp5_ASAP7_75t_L g1088 ( .A(n_647), .B(n_1089), .Y(n_1088) );
NOR3xp33_ASAP7_75t_L g649 ( .A(n_650), .B(n_672), .C(n_680), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_651), .B(n_658), .Y(n_650) );
AOI22xp33_ASAP7_75t_L g651 ( .A1(n_652), .A2(n_653), .B1(n_655), .B2(n_656), .Y(n_651) );
AOI22xp33_ASAP7_75t_L g1207 ( .A1(n_653), .A2(n_656), .B1(n_1208), .B2(n_1209), .Y(n_1207) );
INVx1_ASAP7_75t_L g1420 ( .A(n_653), .Y(n_1420) );
AND2x4_ASAP7_75t_L g656 ( .A(n_654), .B(n_657), .Y(n_656) );
AND2x4_ASAP7_75t_L g680 ( .A(n_654), .B(n_681), .Y(n_680) );
AND2x4_ASAP7_75t_SL g972 ( .A(n_654), .B(n_657), .Y(n_972) );
A2O1A1Ixp33_ASAP7_75t_L g1497 ( .A1(n_654), .A2(n_660), .B(n_1473), .C(n_1498), .Y(n_1497) );
AOI22xp33_ASAP7_75t_L g863 ( .A1(n_656), .A2(n_808), .B1(n_814), .B2(n_864), .Y(n_863) );
AOI22xp33_ASAP7_75t_L g987 ( .A1(n_656), .A2(n_864), .B1(n_988), .B2(n_989), .Y(n_987) );
INVx1_ASAP7_75t_L g1421 ( .A(n_656), .Y(n_1421) );
AOI33xp33_ASAP7_75t_L g658 ( .A1(n_659), .A2(n_662), .A3(n_663), .B1(n_667), .B2(n_669), .B3(n_671), .Y(n_658) );
AOI22xp33_ASAP7_75t_L g1095 ( .A1(n_660), .A2(n_850), .B1(n_1090), .B2(n_1096), .Y(n_1095) );
AOI22xp33_ASAP7_75t_L g1051 ( .A1(n_661), .A2(n_874), .B1(n_1052), .B2(n_1053), .Y(n_1051) );
BUFx3_ASAP7_75t_L g991 ( .A(n_662), .Y(n_991) );
AOI33xp33_ASAP7_75t_L g1185 ( .A1(n_662), .A2(n_1186), .A3(n_1187), .B1(n_1189), .B2(n_1191), .B3(n_1192), .Y(n_1185) );
AOI33xp33_ASAP7_75t_L g1200 ( .A1(n_662), .A2(n_669), .A3(n_1201), .B1(n_1204), .B2(n_1205), .B3(n_1206), .Y(n_1200) );
INVx8_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
OAI22xp5_ASAP7_75t_L g1503 ( .A1(n_665), .A2(n_1504), .B1(n_1505), .B2(n_1506), .Y(n_1503) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
OR2x2_ASAP7_75t_L g673 ( .A(n_674), .B(n_675), .Y(n_673) );
OR2x6_ASAP7_75t_L g862 ( .A(n_674), .B(n_675), .Y(n_862) );
INVxp67_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
AND2x2_ASAP7_75t_L g1174 ( .A(n_676), .B(n_1175), .Y(n_1174) );
INVx2_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
INVx2_ASAP7_75t_L g856 ( .A(n_678), .Y(n_856) );
AOI22xp33_ASAP7_75t_L g976 ( .A1(n_678), .A2(n_930), .B1(n_931), .B2(n_977), .Y(n_976) );
AOI22xp33_ASAP7_75t_L g1023 ( .A1(n_678), .A2(n_1005), .B1(n_1006), .B2(n_1024), .Y(n_1023) );
AND2x4_ASAP7_75t_L g977 ( .A(n_679), .B(n_978), .Y(n_977) );
AND2x4_ASAP7_75t_L g1024 ( .A(n_679), .B(n_978), .Y(n_1024) );
INVx3_ASAP7_75t_L g866 ( .A(n_680), .Y(n_866) );
NOR3xp33_ASAP7_75t_L g951 ( .A(n_680), .B(n_952), .C(n_968), .Y(n_951) );
INVx3_ASAP7_75t_L g1193 ( .A(n_680), .Y(n_1193) );
OAI21xp5_ASAP7_75t_L g682 ( .A1(n_683), .A2(n_700), .B(n_721), .Y(n_682) );
INVx2_ASAP7_75t_SL g684 ( .A(n_685), .Y(n_684) );
AOI22xp33_ASAP7_75t_SL g822 ( .A1(n_685), .A2(n_823), .B1(n_824), .B2(n_825), .Y(n_822) );
AOI221xp5_ASAP7_75t_L g1007 ( .A1(n_685), .A2(n_694), .B1(n_984), .B2(n_1008), .C(n_1013), .Y(n_1007) );
INVx3_ASAP7_75t_L g1165 ( .A(n_685), .Y(n_1165) );
AOI221xp5_ASAP7_75t_L g1215 ( .A1(n_685), .A2(n_694), .B1(n_1197), .B2(n_1216), .C(n_1217), .Y(n_1215) );
HB1xp67_ASAP7_75t_L g693 ( .A(n_686), .Y(n_693) );
BUFx2_ASAP7_75t_L g1131 ( .A(n_686), .Y(n_1131) );
INVx1_ASAP7_75t_L g1836 ( .A(n_686), .Y(n_1836) );
AOI21xp5_ASAP7_75t_L g687 ( .A1(n_688), .A2(n_691), .B(n_694), .Y(n_687) );
AOI221xp5_ASAP7_75t_L g812 ( .A1(n_694), .A2(n_813), .B1(n_814), .B2(n_815), .C(n_820), .Y(n_812) );
AOI21xp5_ASAP7_75t_L g932 ( .A1(n_694), .A2(n_933), .B(n_937), .Y(n_932) );
AOI21xp5_ASAP7_75t_L g1166 ( .A1(n_694), .A2(n_1167), .B(n_1168), .Y(n_1166) );
INVx1_ASAP7_75t_L g1449 ( .A(n_694), .Y(n_1449) );
AOI22xp33_ASAP7_75t_L g695 ( .A1(n_696), .A2(n_697), .B1(n_698), .B2(n_699), .Y(n_695) );
AOI22xp33_ASAP7_75t_L g929 ( .A1(n_697), .A2(n_699), .B1(n_930), .B2(n_931), .Y(n_929) );
AOI22xp33_ASAP7_75t_L g1004 ( .A1(n_697), .A2(n_823), .B1(n_1005), .B2(n_1006), .Y(n_1004) );
AOI22xp33_ASAP7_75t_L g1169 ( .A1(n_697), .A2(n_699), .B1(n_1170), .B2(n_1171), .Y(n_1169) );
AOI22xp33_ASAP7_75t_L g1219 ( .A1(n_697), .A2(n_699), .B1(n_1220), .B2(n_1221), .Y(n_1219) );
INVx1_ASAP7_75t_L g1460 ( .A(n_697), .Y(n_1460) );
BUFx6f_ASAP7_75t_L g823 ( .A(n_699), .Y(n_823) );
HB1xp67_ASAP7_75t_L g1452 ( .A(n_699), .Y(n_1452) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
INVx2_ASAP7_75t_L g941 ( .A(n_702), .Y(n_941) );
INVx4_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
INVx2_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
BUFx3_ASAP7_75t_L g813 ( .A(n_704), .Y(n_813) );
BUFx2_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVx2_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
INVx2_ASAP7_75t_L g1453 ( .A(n_707), .Y(n_1453) );
NOR2x1_ASAP7_75t_L g707 ( .A(n_708), .B(n_709), .Y(n_707) );
INVx1_ASAP7_75t_L g1479 ( .A(n_709), .Y(n_1479) );
OAI211xp5_ASAP7_75t_SL g710 ( .A1(n_711), .A2(n_712), .B(n_714), .C(n_718), .Y(n_710) );
OAI22xp5_ASAP7_75t_L g1234 ( .A1(n_712), .A2(n_1235), .B1(n_1236), .B2(n_1237), .Y(n_1234) );
HB1xp67_ASAP7_75t_L g1341 ( .A(n_712), .Y(n_1341) );
INVx2_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
INVx2_ASAP7_75t_L g1075 ( .A(n_713), .Y(n_1075) );
INVx3_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
INVx2_ASAP7_75t_L g802 ( .A(n_716), .Y(n_802) );
INVx2_ASAP7_75t_L g946 ( .A(n_716), .Y(n_946) );
INVx1_ASAP7_75t_L g1017 ( .A(n_716), .Y(n_1017) );
OAI221xp5_ASAP7_75t_L g1154 ( .A1(n_716), .A2(n_944), .B1(n_1071), .B2(n_1155), .C(n_1156), .Y(n_1154) );
INVx1_ASAP7_75t_L g1352 ( .A(n_717), .Y(n_1352) );
INVxp67_ASAP7_75t_L g1372 ( .A(n_717), .Y(n_1372) );
BUFx6f_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx3_ASAP7_75t_L g1140 ( .A(n_720), .Y(n_1140) );
AOI21xp5_ASAP7_75t_L g1210 ( .A1(n_721), .A2(n_1211), .B(n_1222), .Y(n_1210) );
INVx1_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
OAI21xp33_ASAP7_75t_L g1092 ( .A1(n_722), .A2(n_1093), .B(n_1109), .Y(n_1092) );
INVx1_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
A2O1A1Ixp33_ASAP7_75t_SL g728 ( .A1(n_723), .A2(n_729), .B(n_752), .C(n_757), .Y(n_728) );
INVx1_ASAP7_75t_L g827 ( .A(n_723), .Y(n_827) );
BUFx2_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
HB1xp67_ASAP7_75t_L g950 ( .A(n_724), .Y(n_950) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
OR2x2_ASAP7_75t_L g727 ( .A(n_728), .B(n_761), .Y(n_727) );
OAI21xp33_ASAP7_75t_L g732 ( .A1(n_733), .A2(n_737), .B(n_743), .Y(n_732) );
OAI22xp5_ASAP7_75t_L g772 ( .A1(n_734), .A2(n_744), .B1(n_773), .B2(n_774), .Y(n_772) );
OAI22xp5_ASAP7_75t_L g737 ( .A1(n_738), .A2(n_739), .B1(n_740), .B2(n_742), .Y(n_737) );
INVx1_ASAP7_75t_L g880 ( .A(n_738), .Y(n_880) );
INVx1_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
OAI22xp5_ASAP7_75t_L g775 ( .A1(n_742), .A2(n_769), .B1(n_776), .B2(n_778), .Y(n_775) );
OAI211xp5_ASAP7_75t_L g743 ( .A1(n_744), .A2(n_745), .B(n_747), .C(n_750), .Y(n_743) );
OAI21xp5_ASAP7_75t_SL g1781 ( .A1(n_745), .A2(n_1782), .B(n_1783), .Y(n_1781) );
INVx3_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
INVx2_ASAP7_75t_L g843 ( .A(n_746), .Y(n_843) );
INVx2_ASAP7_75t_L g1103 ( .A(n_746), .Y(n_1103) );
BUFx2_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
BUFx2_ASAP7_75t_L g1041 ( .A(n_751), .Y(n_1041) );
INVx1_ASAP7_75t_L g1263 ( .A(n_751), .Y(n_1263) );
NAND2xp5_ASAP7_75t_L g757 ( .A(n_758), .B(n_759), .Y(n_757) );
INVx1_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
NAND3xp33_ASAP7_75t_L g761 ( .A(n_762), .B(n_782), .C(n_786), .Y(n_761) );
NOR2xp33_ASAP7_75t_SL g762 ( .A(n_763), .B(n_781), .Y(n_762) );
OAI33xp33_ASAP7_75t_L g763 ( .A1(n_764), .A2(n_765), .A3(n_770), .B1(n_772), .B2(n_775), .B3(n_779), .Y(n_763) );
OAI33xp33_ASAP7_75t_L g1230 ( .A1(n_764), .A2(n_1231), .A3(n_1234), .B1(n_1238), .B2(n_1243), .B3(n_1248), .Y(n_1230) );
OAI22xp5_ASAP7_75t_SL g1304 ( .A1(n_764), .A2(n_1305), .B1(n_1307), .B2(n_1308), .Y(n_1304) );
OAI22xp5_ASAP7_75t_L g765 ( .A1(n_766), .A2(n_767), .B1(n_768), .B2(n_769), .Y(n_765) );
OAI221xp5_ASAP7_75t_L g1308 ( .A1(n_774), .A2(n_1280), .B1(n_1285), .B2(n_1309), .C(n_1310), .Y(n_1308) );
OAI221xp5_ASAP7_75t_L g1446 ( .A1(n_776), .A2(n_1346), .B1(n_1426), .B2(n_1438), .C(n_1447), .Y(n_1446) );
INVx2_ASAP7_75t_L g776 ( .A(n_777), .Y(n_776) );
INVx2_ASAP7_75t_L g779 ( .A(n_780), .Y(n_779) );
INVx2_ASAP7_75t_L g1248 ( .A(n_780), .Y(n_1248) );
AOI21xp5_ASAP7_75t_L g920 ( .A1(n_783), .A2(n_921), .B(n_922), .Y(n_920) );
INVx2_ASAP7_75t_L g783 ( .A(n_784), .Y(n_783) );
XOR2xp5_ASAP7_75t_L g788 ( .A(n_789), .B(n_867), .Y(n_788) );
XNOR2x1_ASAP7_75t_L g789 ( .A(n_790), .B(n_791), .Y(n_789) );
AND2x2_ASAP7_75t_L g791 ( .A(n_792), .B(n_857), .Y(n_791) );
AOI221xp5_ASAP7_75t_L g792 ( .A1(n_793), .A2(n_795), .B1(n_796), .B2(n_826), .C(n_828), .Y(n_792) );
INVx2_ASAP7_75t_L g793 ( .A(n_794), .Y(n_793) );
NAND3xp33_ASAP7_75t_L g796 ( .A(n_797), .B(n_812), .C(n_822), .Y(n_796) );
AOI222xp33_ASAP7_75t_L g797 ( .A1(n_798), .A2(n_803), .B1(n_806), .B2(n_808), .C1(n_809), .C2(n_811), .Y(n_797) );
BUFx2_ASAP7_75t_L g799 ( .A(n_800), .Y(n_799) );
INVx2_ASAP7_75t_L g800 ( .A(n_801), .Y(n_800) );
INVx2_ASAP7_75t_L g935 ( .A(n_801), .Y(n_935) );
HB1xp67_ASAP7_75t_L g804 ( .A(n_805), .Y(n_804) );
HB1xp67_ASAP7_75t_L g821 ( .A(n_805), .Y(n_821) );
INVx1_ASAP7_75t_L g1020 ( .A(n_806), .Y(n_1020) );
AOI222xp33_ASAP7_75t_L g1212 ( .A1(n_806), .A2(n_813), .B1(n_1208), .B2(n_1209), .C1(n_1213), .C2(n_1214), .Y(n_1212) );
AOI22xp33_ASAP7_75t_SL g1480 ( .A1(n_806), .A2(n_1481), .B1(n_1482), .B2(n_1483), .Y(n_1480) );
INVx2_ASAP7_75t_L g809 ( .A(n_810), .Y(n_809) );
AOI222xp33_ASAP7_75t_L g1014 ( .A1(n_813), .A2(n_988), .B1(n_989), .B2(n_1015), .C1(n_1018), .C2(n_1019), .Y(n_1014) );
INVx1_ASAP7_75t_L g816 ( .A(n_817), .Y(n_816) );
HB1xp67_ASAP7_75t_SL g818 ( .A(n_819), .Y(n_818) );
INVx2_ASAP7_75t_L g826 ( .A(n_827), .Y(n_826) );
OAI22xp5_ASAP7_75t_L g829 ( .A1(n_830), .A2(n_831), .B1(n_833), .B2(n_834), .Y(n_829) );
INVx1_ASAP7_75t_L g831 ( .A(n_832), .Y(n_831) );
INVx1_ASAP7_75t_L g1425 ( .A(n_832), .Y(n_1425) );
OAI22xp5_ASAP7_75t_L g1326 ( .A1(n_834), .A2(n_1327), .B1(n_1328), .B2(n_1329), .Y(n_1326) );
CKINVDCx20_ASAP7_75t_R g956 ( .A(n_835), .Y(n_956) );
BUFx8_ASAP7_75t_L g835 ( .A(n_836), .Y(n_835) );
BUFx2_ASAP7_75t_L g1318 ( .A(n_836), .Y(n_1318) );
BUFx4f_ASAP7_75t_L g1428 ( .A(n_836), .Y(n_1428) );
OAI22xp33_ASAP7_75t_L g837 ( .A1(n_838), .A2(n_839), .B1(n_842), .B2(n_843), .Y(n_837) );
OAI22xp33_ASAP7_75t_L g1331 ( .A1(n_839), .A2(n_1332), .B1(n_1333), .B2(n_1334), .Y(n_1331) );
INVx2_ASAP7_75t_L g839 ( .A(n_840), .Y(n_839) );
INVx1_ASAP7_75t_L g840 ( .A(n_841), .Y(n_840) );
OAI22xp33_ASAP7_75t_L g1510 ( .A1(n_841), .A2(n_876), .B1(n_1511), .B2(n_1512), .Y(n_1510) );
OAI22xp5_ASAP7_75t_L g1771 ( .A1(n_841), .A2(n_1772), .B1(n_1773), .B2(n_1774), .Y(n_1771) );
INVx1_ASAP7_75t_L g845 ( .A(n_846), .Y(n_845) );
INVx1_ASAP7_75t_L g851 ( .A(n_852), .Y(n_851) );
BUFx2_ASAP7_75t_L g852 ( .A(n_853), .Y(n_852) );
BUFx2_ASAP7_75t_L g1000 ( .A(n_853), .Y(n_1000) );
BUFx2_ASAP7_75t_L g1192 ( .A(n_853), .Y(n_1192) );
INVx3_ASAP7_75t_L g853 ( .A(n_854), .Y(n_853) );
INVx3_ASAP7_75t_L g967 ( .A(n_854), .Y(n_967) );
INVxp67_ASAP7_75t_L g1418 ( .A(n_856), .Y(n_1418) );
NAND2xp5_ASAP7_75t_L g1183 ( .A(n_858), .B(n_1184), .Y(n_1183) );
INVx3_ASAP7_75t_L g858 ( .A(n_859), .Y(n_858) );
AOI22xp5_ASAP7_75t_L g1180 ( .A1(n_864), .A2(n_972), .B1(n_1181), .B2(n_1182), .Y(n_1180) );
INVx2_ASAP7_75t_L g864 ( .A(n_865), .Y(n_864) );
NAND3xp33_ASAP7_75t_SL g986 ( .A(n_866), .B(n_987), .C(n_990), .Y(n_986) );
XNOR2xp5_ASAP7_75t_L g867 ( .A(n_868), .B(n_923), .Y(n_867) );
OR2x2_ASAP7_75t_L g869 ( .A(n_870), .B(n_894), .Y(n_869) );
A2O1A1Ixp33_ASAP7_75t_L g870 ( .A1(n_871), .A2(n_884), .B(n_888), .C(n_890), .Y(n_870) );
NOR3xp33_ASAP7_75t_L g871 ( .A(n_872), .B(n_873), .C(n_879), .Y(n_871) );
INVx2_ASAP7_75t_L g1112 ( .A(n_876), .Y(n_1112) );
BUFx6f_ASAP7_75t_L g1333 ( .A(n_876), .Y(n_1333) );
OAI22xp5_ASAP7_75t_L g905 ( .A1(n_883), .A2(n_906), .B1(n_907), .B2(n_909), .Y(n_905) );
A2O1A1Ixp33_ASAP7_75t_L g1256 ( .A1(n_888), .A2(n_1257), .B(n_1260), .C(n_1270), .Y(n_1256) );
INVx2_ASAP7_75t_L g888 ( .A(n_889), .Y(n_888) );
INVx1_ASAP7_75t_L g1021 ( .A(n_889), .Y(n_1021) );
AOI21xp5_ASAP7_75t_L g1029 ( .A1(n_889), .A2(n_1030), .B(n_1055), .Y(n_1029) );
NAND2xp5_ASAP7_75t_L g890 ( .A(n_891), .B(n_892), .Y(n_890) );
INVx1_ASAP7_75t_L g892 ( .A(n_893), .Y(n_892) );
NAND4xp25_ASAP7_75t_L g894 ( .A(n_895), .B(n_898), .C(n_918), .D(n_920), .Y(n_894) );
INVx1_ASAP7_75t_L g901 ( .A(n_902), .Y(n_901) );
INVx1_ASAP7_75t_L g1448 ( .A(n_902), .Y(n_1448) );
INVx1_ASAP7_75t_L g903 ( .A(n_904), .Y(n_903) );
INVx4_ASAP7_75t_L g907 ( .A(n_908), .Y(n_907) );
INVx3_ASAP7_75t_L g1067 ( .A(n_908), .Y(n_1067) );
BUFx6f_ASAP7_75t_L g1160 ( .A(n_908), .Y(n_1160) );
HB1xp67_ASAP7_75t_L g1339 ( .A(n_909), .Y(n_1339) );
INVx2_ASAP7_75t_L g1347 ( .A(n_909), .Y(n_1347) );
OAI22xp5_ASAP7_75t_L g912 ( .A1(n_913), .A2(n_914), .B1(n_916), .B2(n_917), .Y(n_912) );
INVx1_ASAP7_75t_L g914 ( .A(n_915), .Y(n_914) );
OAI22xp5_ASAP7_75t_L g1243 ( .A1(n_917), .A2(n_1244), .B1(n_1246), .B2(n_1247), .Y(n_1243) );
NOR3xp33_ASAP7_75t_L g1303 ( .A(n_922), .B(n_1304), .C(n_1311), .Y(n_1303) );
AND4x1_ASAP7_75t_L g924 ( .A(n_925), .B(n_951), .C(n_973), .D(n_976), .Y(n_924) );
OAI21xp33_ASAP7_75t_L g925 ( .A1(n_926), .A2(n_940), .B(n_950), .Y(n_925) );
INVx2_ASAP7_75t_L g927 ( .A(n_928), .Y(n_927) );
OAI211xp5_ASAP7_75t_L g942 ( .A1(n_943), .A2(n_944), .B(n_945), .C(n_947), .Y(n_942) );
A2O1A1Ixp33_ASAP7_75t_L g1276 ( .A1(n_950), .A2(n_1277), .B(n_1291), .C(n_1298), .Y(n_1276) );
OAI22xp5_ASAP7_75t_L g952 ( .A1(n_953), .A2(n_957), .B1(n_960), .B2(n_966), .Y(n_952) );
OAI21xp5_ASAP7_75t_L g953 ( .A1(n_954), .A2(n_955), .B(n_956), .Y(n_953) );
INVx1_ASAP7_75t_L g1190 ( .A(n_954), .Y(n_1190) );
OAI22xp5_ASAP7_75t_L g1115 ( .A1(n_961), .A2(n_1116), .B1(n_1117), .B2(n_1118), .Y(n_1115) );
CKINVDCx8_ASAP7_75t_R g961 ( .A(n_962), .Y(n_961) );
INVx3_ASAP7_75t_L g1269 ( .A(n_962), .Y(n_1269) );
INVx3_ASAP7_75t_L g1289 ( .A(n_962), .Y(n_1289) );
INVx3_ASAP7_75t_L g1773 ( .A(n_962), .Y(n_1773) );
AOI22xp5_ASAP7_75t_L g1785 ( .A1(n_965), .A2(n_978), .B1(n_1766), .B2(n_1786), .Y(n_1785) );
CKINVDCx5p33_ASAP7_75t_R g966 ( .A(n_967), .Y(n_966) );
INVx1_ASAP7_75t_L g969 ( .A(n_970), .Y(n_969) );
INVx1_ASAP7_75t_L g971 ( .A(n_972), .Y(n_971) );
AOI22xp33_ASAP7_75t_L g1173 ( .A1(n_977), .A2(n_1170), .B1(n_1171), .B2(n_1174), .Y(n_1173) );
AOI22xp33_ASAP7_75t_L g1223 ( .A1(n_977), .A2(n_1174), .B1(n_1220), .B2(n_1221), .Y(n_1223) );
XNOR2xp5_ASAP7_75t_L g979 ( .A(n_980), .B(n_1025), .Y(n_979) );
XNOR2x1_ASAP7_75t_L g1313 ( .A(n_980), .B(n_1025), .Y(n_1313) );
BUFx3_ASAP7_75t_L g980 ( .A(n_981), .Y(n_980) );
NAND2xp5_ASAP7_75t_L g982 ( .A(n_983), .B(n_1002), .Y(n_982) );
AOI33xp33_ASAP7_75t_L g990 ( .A1(n_991), .A2(n_992), .A3(n_996), .B1(n_998), .B2(n_1000), .B3(n_1001), .Y(n_990) );
INVx1_ASAP7_75t_L g993 ( .A(n_994), .Y(n_993) );
INVx1_ASAP7_75t_L g1330 ( .A(n_1000), .Y(n_1330) );
AOI21xp5_ASAP7_75t_SL g1002 ( .A1(n_1003), .A2(n_1021), .B(n_1022), .Y(n_1002) );
NAND3xp33_ASAP7_75t_SL g1003 ( .A(n_1004), .B(n_1007), .C(n_1014), .Y(n_1003) );
INVx2_ASAP7_75t_L g1009 ( .A(n_1010), .Y(n_1009) );
INVx1_ASAP7_75t_L g1010 ( .A(n_1011), .Y(n_1010) );
INVx1_ASAP7_75t_L g1011 ( .A(n_1012), .Y(n_1011) );
BUFx2_ASAP7_75t_L g1839 ( .A(n_1012), .Y(n_1839) );
INVx1_ASAP7_75t_L g1019 ( .A(n_1020), .Y(n_1019) );
O2A1O1Ixp33_ASAP7_75t_SL g1152 ( .A1(n_1021), .A2(n_1153), .B(n_1164), .C(n_1172), .Y(n_1152) );
OAI31xp33_ASAP7_75t_L g1444 ( .A1(n_1021), .A2(n_1445), .A3(n_1450), .B(n_1459), .Y(n_1444) );
NAND2xp5_ASAP7_75t_L g1490 ( .A(n_1024), .B(n_1491), .Y(n_1490) );
XNOR2x1_ASAP7_75t_L g1025 ( .A(n_1026), .B(n_1147), .Y(n_1025) );
XNOR2x2_ASAP7_75t_L g1026 ( .A(n_1027), .B(n_1083), .Y(n_1026) );
AOI21xp5_ASAP7_75t_L g1027 ( .A1(n_1028), .A2(n_1081), .B(n_1082), .Y(n_1027) );
AND3x1_ASAP7_75t_L g1028 ( .A(n_1029), .B(n_1056), .C(n_1062), .Y(n_1028) );
AOI31xp33_ASAP7_75t_L g1082 ( .A1(n_1029), .A2(n_1056), .A3(n_1062), .B(n_1081), .Y(n_1082) );
NAND3xp33_ASAP7_75t_SL g1030 ( .A(n_1031), .B(n_1042), .C(n_1046), .Y(n_1030) );
AOI22xp5_ASAP7_75t_L g1031 ( .A1(n_1032), .A2(n_1035), .B1(n_1036), .B2(n_1039), .Y(n_1031) );
INVx2_ASAP7_75t_L g1037 ( .A(n_1038), .Y(n_1037) );
OAI22xp5_ASAP7_75t_L g1778 ( .A1(n_1038), .A2(n_1289), .B1(n_1779), .B2(n_1780), .Y(n_1778) );
NOR3xp33_ASAP7_75t_L g1260 ( .A(n_1045), .B(n_1261), .C(n_1266), .Y(n_1260) );
NOR3xp33_ASAP7_75t_L g1277 ( .A(n_1045), .B(n_1278), .C(n_1283), .Y(n_1277) );
NOR2xp33_ASAP7_75t_L g1842 ( .A(n_1045), .B(n_1843), .Y(n_1842) );
INVxp67_ASAP7_75t_L g1094 ( .A(n_1047), .Y(n_1094) );
INVx1_ASAP7_75t_L g1047 ( .A(n_1048), .Y(n_1047) );
OAI22xp5_ASAP7_75t_L g1287 ( .A1(n_1050), .A2(n_1288), .B1(n_1289), .B2(n_1290), .Y(n_1287) );
INVx2_ASAP7_75t_L g1437 ( .A(n_1050), .Y(n_1437) );
AND2x2_ASAP7_75t_L g1056 ( .A(n_1057), .B(n_1059), .Y(n_1056) );
NAND2xp5_ASAP7_75t_L g1059 ( .A(n_1060), .B(n_1061), .Y(n_1059) );
INVx2_ASAP7_75t_SL g1456 ( .A(n_1067), .Y(n_1456) );
OAI221xp5_ASAP7_75t_L g1070 ( .A1(n_1071), .A2(n_1074), .B1(n_1075), .B2(n_1076), .C(n_1077), .Y(n_1070) );
OAI22xp5_ASAP7_75t_L g1342 ( .A1(n_1071), .A2(n_1137), .B1(n_1321), .B2(n_1334), .Y(n_1342) );
INVx3_ASAP7_75t_L g1071 ( .A(n_1072), .Y(n_1071) );
INVx2_ASAP7_75t_L g1072 ( .A(n_1073), .Y(n_1072) );
OAI221xp5_ASAP7_75t_L g1305 ( .A1(n_1073), .A2(n_1129), .B1(n_1281), .B2(n_1288), .C(n_1306), .Y(n_1305) );
BUFx6f_ASAP7_75t_L g1078 ( .A(n_1079), .Y(n_1078) );
INVx1_ASAP7_75t_L g1084 ( .A(n_1085), .Y(n_1084) );
NAND3xp33_ASAP7_75t_L g1085 ( .A(n_1086), .B(n_1092), .C(n_1119), .Y(n_1085) );
NAND2xp5_ASAP7_75t_L g1802 ( .A(n_1088), .B(n_1803), .Y(n_1802) );
OAI211xp5_ASAP7_75t_L g1093 ( .A1(n_1094), .A2(n_1095), .B(n_1097), .C(n_1100), .Y(n_1093) );
OAI211xp5_ASAP7_75t_L g1100 ( .A1(n_1101), .A2(n_1102), .B(n_1104), .C(n_1107), .Y(n_1100) );
OAI221xp5_ASAP7_75t_L g1133 ( .A1(n_1101), .A2(n_1113), .B1(n_1134), .B2(n_1137), .C(n_1138), .Y(n_1133) );
HB1xp67_ASAP7_75t_L g1102 ( .A(n_1103), .Y(n_1102) );
INVx1_ASAP7_75t_L g1105 ( .A(n_1106), .Y(n_1105) );
OAI22xp5_ASAP7_75t_L g1268 ( .A1(n_1106), .A2(n_1235), .B1(n_1247), .B2(n_1269), .Y(n_1268) );
INVx1_ASAP7_75t_L g1111 ( .A(n_1112), .Y(n_1111) );
OAI221xp5_ASAP7_75t_L g1125 ( .A1(n_1117), .A2(n_1126), .B1(n_1128), .B2(n_1129), .C(n_1130), .Y(n_1125) );
NOR3xp33_ASAP7_75t_L g1119 ( .A(n_1120), .B(n_1132), .C(n_1142), .Y(n_1119) );
INVxp67_ASAP7_75t_L g1121 ( .A(n_1122), .Y(n_1121) );
HB1xp67_ASAP7_75t_L g1122 ( .A(n_1123), .Y(n_1122) );
INVx2_ASAP7_75t_SL g1123 ( .A(n_1124), .Y(n_1123) );
OAI22xp5_ASAP7_75t_L g1340 ( .A1(n_1126), .A2(n_1323), .B1(n_1328), .B2(n_1341), .Y(n_1340) );
INVx2_ASAP7_75t_L g1126 ( .A(n_1127), .Y(n_1126) );
BUFx2_ASAP7_75t_L g1240 ( .A(n_1127), .Y(n_1240) );
INVx2_ASAP7_75t_L g1309 ( .A(n_1127), .Y(n_1309) );
INVx2_ASAP7_75t_L g1134 ( .A(n_1135), .Y(n_1134) );
INVx4_ASAP7_75t_L g1236 ( .A(n_1135), .Y(n_1236) );
INVx2_ASAP7_75t_L g1471 ( .A(n_1135), .Y(n_1471) );
INVx4_ASAP7_75t_L g1135 ( .A(n_1136), .Y(n_1135) );
INVx2_ASAP7_75t_L g1139 ( .A(n_1140), .Y(n_1139) );
INVx1_ASAP7_75t_L g1218 ( .A(n_1140), .Y(n_1218) );
INVx1_ASAP7_75t_L g1143 ( .A(n_1144), .Y(n_1143) );
NAND2xp5_ASAP7_75t_L g1804 ( .A(n_1144), .B(n_1805), .Y(n_1804) );
XNOR2xp5_ASAP7_75t_L g1147 ( .A(n_1148), .B(n_1224), .Y(n_1147) );
XNOR2xp5_ASAP7_75t_L g1148 ( .A(n_1149), .B(n_1194), .Y(n_1148) );
NOR2x1p5_ASAP7_75t_L g1150 ( .A(n_1151), .B(n_1176), .Y(n_1150) );
INVx1_ASAP7_75t_L g1151 ( .A(n_1152), .Y(n_1151) );
OAI22xp5_ASAP7_75t_L g1157 ( .A1(n_1158), .A2(n_1159), .B1(n_1161), .B2(n_1162), .Y(n_1157) );
INVx2_ASAP7_75t_L g1159 ( .A(n_1160), .Y(n_1159) );
BUFx3_ASAP7_75t_L g1162 ( .A(n_1163), .Y(n_1162) );
AOI22xp33_ASAP7_75t_L g1492 ( .A1(n_1174), .A2(n_1483), .B1(n_1493), .B2(n_1494), .Y(n_1492) );
INVx2_ASAP7_75t_L g1265 ( .A(n_1175), .Y(n_1265) );
INVx2_ASAP7_75t_L g1294 ( .A(n_1175), .Y(n_1294) );
NAND2xp5_ASAP7_75t_L g1176 ( .A(n_1177), .B(n_1179), .Y(n_1176) );
AND4x1_ASAP7_75t_L g1179 ( .A(n_1180), .B(n_1183), .C(n_1185), .D(n_1193), .Y(n_1179) );
NAND3xp33_ASAP7_75t_L g1199 ( .A(n_1193), .B(n_1200), .C(n_1207), .Y(n_1199) );
AND2x2_ASAP7_75t_L g1195 ( .A(n_1196), .B(n_1210), .Y(n_1195) );
NAND3xp33_ASAP7_75t_L g1211 ( .A(n_1212), .B(n_1215), .C(n_1219), .Y(n_1211) );
XNOR2x1_ASAP7_75t_L g1224 ( .A(n_1225), .B(n_1272), .Y(n_1224) );
XNOR2x1_ASAP7_75t_L g1225 ( .A(n_1226), .B(n_1227), .Y(n_1225) );
NOR2x1_ASAP7_75t_L g1227 ( .A(n_1228), .B(n_1256), .Y(n_1227) );
NAND3xp33_ASAP7_75t_L g1228 ( .A(n_1229), .B(n_1250), .C(n_1254), .Y(n_1228) );
NOR2xp33_ASAP7_75t_L g1229 ( .A(n_1230), .B(n_1249), .Y(n_1229) );
INVx4_ASAP7_75t_L g1239 ( .A(n_1240), .Y(n_1239) );
INVx1_ASAP7_75t_L g1244 ( .A(n_1245), .Y(n_1244) );
INVx1_ASAP7_75t_L g1262 ( .A(n_1263), .Y(n_1262) );
OAI22xp5_ASAP7_75t_L g1507 ( .A1(n_1265), .A2(n_1505), .B1(n_1508), .B2(n_1509), .Y(n_1507) );
INVx2_ASAP7_75t_L g1272 ( .A(n_1273), .Y(n_1272) );
XNOR2x1_ASAP7_75t_L g1273 ( .A(n_1274), .B(n_1275), .Y(n_1273) );
OR2x2_ASAP7_75t_L g1275 ( .A(n_1276), .B(n_1299), .Y(n_1275) );
OAI22xp5_ASAP7_75t_L g1322 ( .A1(n_1289), .A2(n_1323), .B1(n_1324), .B2(n_1325), .Y(n_1322) );
INVx1_ASAP7_75t_L g1344 ( .A(n_1307), .Y(n_1344) );
INVx2_ASAP7_75t_L g1312 ( .A(n_1313), .Y(n_1312) );
INVx1_ASAP7_75t_L g1409 ( .A(n_1314), .Y(n_1409) );
NAND3xp33_ASAP7_75t_L g1315 ( .A(n_1316), .B(n_1348), .C(n_1379), .Y(n_1315) );
NOR2xp33_ASAP7_75t_L g1316 ( .A(n_1317), .B(n_1335), .Y(n_1316) );
OAI33xp33_ASAP7_75t_L g1317 ( .A1(n_1318), .A2(n_1319), .A3(n_1322), .B1(n_1326), .B2(n_1330), .B3(n_1331), .Y(n_1317) );
OAI22xp5_ASAP7_75t_SL g1336 ( .A1(n_1320), .A2(n_1332), .B1(n_1337), .B2(n_1339), .Y(n_1336) );
OAI22xp5_ASAP7_75t_L g1345 ( .A1(n_1325), .A2(n_1329), .B1(n_1337), .B2(n_1346), .Y(n_1345) );
OAI22xp5_ASAP7_75t_L g1429 ( .A1(n_1333), .A2(n_1430), .B1(n_1432), .B2(n_1433), .Y(n_1429) );
INVx2_ASAP7_75t_L g1337 ( .A(n_1338), .Y(n_1337) );
INVx2_ASAP7_75t_L g1343 ( .A(n_1344), .Y(n_1343) );
OAI221xp5_ASAP7_75t_L g1454 ( .A1(n_1346), .A2(n_1432), .B1(n_1455), .B2(n_1457), .C(n_1458), .Y(n_1454) );
INVx2_ASAP7_75t_L g1346 ( .A(n_1347), .Y(n_1346) );
OAI31xp33_ASAP7_75t_L g1348 ( .A1(n_1349), .A2(n_1361), .A3(n_1368), .B(n_1375), .Y(n_1348) );
INVx3_ASAP7_75t_L g1350 ( .A(n_1351), .Y(n_1350) );
AOI22xp33_ASAP7_75t_L g1353 ( .A1(n_1354), .A2(n_1355), .B1(n_1357), .B2(n_1358), .Y(n_1353) );
AOI22xp33_ASAP7_75t_L g1388 ( .A1(n_1354), .A2(n_1389), .B1(n_1393), .B2(n_1396), .Y(n_1388) );
INVx2_ASAP7_75t_L g1358 ( .A(n_1359), .Y(n_1358) );
INVx2_ASAP7_75t_L g1359 ( .A(n_1360), .Y(n_1359) );
HB1xp67_ASAP7_75t_L g1362 ( .A(n_1363), .Y(n_1362) );
INVx2_ASAP7_75t_L g1365 ( .A(n_1366), .Y(n_1365) );
INVx2_ASAP7_75t_L g1366 ( .A(n_1367), .Y(n_1366) );
INVx1_ASAP7_75t_L g1369 ( .A(n_1370), .Y(n_1369) );
NAND2xp5_ASAP7_75t_L g1525 ( .A(n_1370), .B(n_1526), .Y(n_1525) );
AND2x4_ASAP7_75t_SL g1807 ( .A(n_1370), .B(n_1808), .Y(n_1807) );
INVx3_ASAP7_75t_L g1370 ( .A(n_1371), .Y(n_1370) );
INVx3_ASAP7_75t_SL g1373 ( .A(n_1374), .Y(n_1373) );
BUFx3_ASAP7_75t_L g1375 ( .A(n_1376), .Y(n_1375) );
AND2x4_ASAP7_75t_L g1376 ( .A(n_1377), .B(n_1378), .Y(n_1376) );
INVx1_ASAP7_75t_L g1526 ( .A(n_1377), .Y(n_1526) );
NOR2xp33_ASAP7_75t_L g1808 ( .A(n_1377), .B(n_1518), .Y(n_1808) );
OAI31xp33_ASAP7_75t_L g1379 ( .A1(n_1380), .A2(n_1385), .A3(n_1397), .B(n_1403), .Y(n_1379) );
INVx2_ASAP7_75t_L g1382 ( .A(n_1383), .Y(n_1382) );
CKINVDCx8_ASAP7_75t_R g1386 ( .A(n_1387), .Y(n_1386) );
BUFx3_ASAP7_75t_L g1389 ( .A(n_1390), .Y(n_1389) );
AND2x2_ASAP7_75t_L g1390 ( .A(n_1391), .B(n_1392), .Y(n_1390) );
AND2x4_ASAP7_75t_L g1394 ( .A(n_1391), .B(n_1395), .Y(n_1394) );
BUFx6f_ASAP7_75t_L g1393 ( .A(n_1394), .Y(n_1393) );
INVx1_ASAP7_75t_L g1398 ( .A(n_1399), .Y(n_1398) );
INVx2_ASAP7_75t_SL g1399 ( .A(n_1400), .Y(n_1399) );
BUFx3_ASAP7_75t_L g1401 ( .A(n_1402), .Y(n_1401) );
BUFx2_ASAP7_75t_L g1403 ( .A(n_1404), .Y(n_1403) );
AND2x2_ASAP7_75t_SL g1404 ( .A(n_1405), .B(n_1407), .Y(n_1404) );
INVx1_ASAP7_75t_SL g1405 ( .A(n_1406), .Y(n_1405) );
INVx1_ASAP7_75t_L g1407 ( .A(n_1408), .Y(n_1407) );
CKINVDCx5p33_ASAP7_75t_R g1410 ( .A(n_1411), .Y(n_1410) );
HB1xp67_ASAP7_75t_L g1411 ( .A(n_1412), .Y(n_1411) );
OAI22xp33_ASAP7_75t_L g1412 ( .A1(n_1413), .A2(n_1462), .B1(n_1463), .B2(n_1514), .Y(n_1412) );
INVx2_ASAP7_75t_L g1414 ( .A(n_1415), .Y(n_1414) );
AND3x2_ASAP7_75t_L g1415 ( .A(n_1416), .B(n_1441), .C(n_1444), .Y(n_1415) );
AOI211xp5_ASAP7_75t_SL g1416 ( .A1(n_1417), .A2(n_1418), .B(n_1419), .C(n_1422), .Y(n_1416) );
BUFx3_ASAP7_75t_L g1427 ( .A(n_1428), .Y(n_1427) );
OAI33xp33_ASAP7_75t_L g1499 ( .A1(n_1428), .A2(n_1500), .A3(n_1503), .B1(n_1507), .B2(n_1510), .B3(n_1513), .Y(n_1499) );
INVx2_ASAP7_75t_L g1430 ( .A(n_1431), .Y(n_1430) );
INVx2_ASAP7_75t_L g1436 ( .A(n_1437), .Y(n_1436) );
INVxp67_ASAP7_75t_L g1451 ( .A(n_1452), .Y(n_1451) );
INVx2_ASAP7_75t_L g1455 ( .A(n_1456), .Y(n_1455) );
INVx1_ASAP7_75t_L g1462 ( .A(n_1463), .Y(n_1462) );
HB1xp67_ASAP7_75t_L g1463 ( .A(n_1464), .Y(n_1463) );
INVx2_ASAP7_75t_L g1466 ( .A(n_1467), .Y(n_1466) );
OR2x2_ASAP7_75t_L g1467 ( .A(n_1468), .B(n_1489), .Y(n_1467) );
AOI21xp5_ASAP7_75t_L g1469 ( .A1(n_1470), .A2(n_1475), .B(n_1476), .Y(n_1469) );
NAND2xp5_ASAP7_75t_L g1476 ( .A(n_1477), .B(n_1480), .Y(n_1476) );
AOI22xp5_ASAP7_75t_L g1484 ( .A1(n_1485), .A2(n_1486), .B1(n_1487), .B2(n_1488), .Y(n_1484) );
NAND3xp33_ASAP7_75t_SL g1489 ( .A(n_1490), .B(n_1492), .C(n_1495), .Y(n_1489) );
NOR2xp33_ASAP7_75t_SL g1495 ( .A(n_1496), .B(n_1499), .Y(n_1495) );
BUFx3_ASAP7_75t_L g1515 ( .A(n_1516), .Y(n_1515) );
INVx3_ASAP7_75t_L g1516 ( .A(n_1517), .Y(n_1516) );
OR2x2_ASAP7_75t_L g1517 ( .A(n_1518), .B(n_1524), .Y(n_1517) );
INVx1_ASAP7_75t_L g1518 ( .A(n_1519), .Y(n_1518) );
NOR2xp33_ASAP7_75t_L g1519 ( .A(n_1520), .B(n_1522), .Y(n_1519) );
NOR2xp33_ASAP7_75t_L g1813 ( .A(n_1520), .B(n_1523), .Y(n_1813) );
INVx1_ASAP7_75t_L g1860 ( .A(n_1520), .Y(n_1860) );
HB1xp67_ASAP7_75t_L g1520 ( .A(n_1521), .Y(n_1520) );
INVx1_ASAP7_75t_L g1522 ( .A(n_1523), .Y(n_1522) );
NOR2xp33_ASAP7_75t_L g1862 ( .A(n_1523), .B(n_1860), .Y(n_1862) );
INVx1_ASAP7_75t_L g1524 ( .A(n_1525), .Y(n_1524) );
OAI221xp5_ASAP7_75t_L g1527 ( .A1(n_1528), .A2(n_1756), .B1(n_1759), .B2(n_1806), .C(n_1809), .Y(n_1527) );
AND5x1_ASAP7_75t_L g1528 ( .A(n_1529), .B(n_1670), .C(n_1717), .D(n_1739), .E(n_1752), .Y(n_1528) );
OAI31xp33_ASAP7_75t_L g1529 ( .A1(n_1530), .A2(n_1608), .A3(n_1647), .B(n_1661), .Y(n_1529) );
OAI221xp5_ASAP7_75t_L g1530 ( .A1(n_1531), .A2(n_1559), .B1(n_1570), .B2(n_1577), .C(n_1578), .Y(n_1530) );
NAND2x1_ASAP7_75t_L g1531 ( .A(n_1532), .B(n_1547), .Y(n_1531) );
NAND2xp5_ASAP7_75t_SL g1623 ( .A(n_1532), .B(n_1624), .Y(n_1623) );
CKINVDCx5p33_ASAP7_75t_R g1644 ( .A(n_1532), .Y(n_1644) );
OAI21xp33_ASAP7_75t_L g1684 ( .A1(n_1532), .A2(n_1597), .B(n_1685), .Y(n_1684) );
NOR2xp33_ASAP7_75t_L g1690 ( .A(n_1532), .B(n_1691), .Y(n_1690) );
AND2x2_ASAP7_75t_L g1694 ( .A(n_1532), .B(n_1600), .Y(n_1694) );
NOR2x1_ASAP7_75t_L g1699 ( .A(n_1532), .B(n_1700), .Y(n_1699) );
OAI22xp5_ASAP7_75t_SL g1722 ( .A1(n_1532), .A2(n_1678), .B1(n_1723), .B2(n_1727), .Y(n_1722) );
AND2x2_ASAP7_75t_L g1750 ( .A(n_1532), .B(n_1751), .Y(n_1750) );
INVx4_ASAP7_75t_L g1532 ( .A(n_1533), .Y(n_1532) );
INVx4_ASAP7_75t_L g1571 ( .A(n_1533), .Y(n_1571) );
OR2x2_ASAP7_75t_L g1604 ( .A(n_1533), .B(n_1548), .Y(n_1604) );
NAND2xp5_ASAP7_75t_SL g1606 ( .A(n_1533), .B(n_1548), .Y(n_1606) );
NOR2xp33_ASAP7_75t_L g1637 ( .A(n_1533), .B(n_1638), .Y(n_1637) );
NOR3xp33_ASAP7_75t_L g1658 ( .A(n_1533), .B(n_1659), .C(n_1660), .Y(n_1658) );
NOR2xp33_ASAP7_75t_L g1677 ( .A(n_1533), .B(n_1581), .Y(n_1677) );
NOR2xp33_ASAP7_75t_L g1702 ( .A(n_1533), .B(n_1703), .Y(n_1702) );
AND2x4_ASAP7_75t_SL g1533 ( .A(n_1534), .B(n_1542), .Y(n_1533) );
AND2x4_ASAP7_75t_L g1535 ( .A(n_1536), .B(n_1537), .Y(n_1535) );
AND2x6_ASAP7_75t_L g1540 ( .A(n_1536), .B(n_1541), .Y(n_1540) );
AND2x6_ASAP7_75t_L g1543 ( .A(n_1536), .B(n_1544), .Y(n_1543) );
AND2x2_ASAP7_75t_L g1545 ( .A(n_1536), .B(n_1546), .Y(n_1545) );
AND2x2_ASAP7_75t_L g1551 ( .A(n_1536), .B(n_1546), .Y(n_1551) );
AND2x2_ASAP7_75t_L g1564 ( .A(n_1536), .B(n_1546), .Y(n_1564) );
NAND2xp5_ASAP7_75t_L g1665 ( .A(n_1536), .B(n_1537), .Y(n_1665) );
AND2x2_ASAP7_75t_L g1537 ( .A(n_1538), .B(n_1539), .Y(n_1537) );
INVx2_ASAP7_75t_L g1667 ( .A(n_1540), .Y(n_1667) );
INVx2_ASAP7_75t_L g1758 ( .A(n_1543), .Y(n_1758) );
OAI21xp5_ASAP7_75t_L g1859 ( .A1(n_1544), .A2(n_1860), .B(n_1861), .Y(n_1859) );
AND2x2_ASAP7_75t_L g1547 ( .A(n_1548), .B(n_1552), .Y(n_1547) );
INVx1_ASAP7_75t_L g1574 ( .A(n_1548), .Y(n_1574) );
OR2x2_ASAP7_75t_L g1625 ( .A(n_1548), .B(n_1626), .Y(n_1625) );
OR2x2_ASAP7_75t_L g1682 ( .A(n_1548), .B(n_1553), .Y(n_1682) );
NAND2xp5_ASAP7_75t_L g1695 ( .A(n_1548), .B(n_1556), .Y(n_1695) );
OR2x2_ASAP7_75t_L g1703 ( .A(n_1548), .B(n_1593), .Y(n_1703) );
AND2x2_ASAP7_75t_L g1726 ( .A(n_1548), .B(n_1593), .Y(n_1726) );
AND2x2_ASAP7_75t_L g1548 ( .A(n_1549), .B(n_1550), .Y(n_1548) );
AND2x2_ASAP7_75t_L g1591 ( .A(n_1549), .B(n_1550), .Y(n_1591) );
INVx1_ASAP7_75t_L g1700 ( .A(n_1552), .Y(n_1700) );
AND2x2_ASAP7_75t_L g1716 ( .A(n_1552), .B(n_1653), .Y(n_1716) );
AND2x2_ASAP7_75t_L g1552 ( .A(n_1553), .B(n_1556), .Y(n_1552) );
NAND2xp5_ASAP7_75t_L g1575 ( .A(n_1553), .B(n_1576), .Y(n_1575) );
OR2x2_ASAP7_75t_L g1581 ( .A(n_1553), .B(n_1556), .Y(n_1581) );
INVx2_ASAP7_75t_L g1593 ( .A(n_1553), .Y(n_1593) );
AOI332xp33_ASAP7_75t_L g1636 ( .A1(n_1553), .A2(n_1591), .A3(n_1629), .B1(n_1637), .B2(n_1639), .B3(n_1642), .C1(n_1645), .C2(n_1646), .Y(n_1636) );
NAND2x1p5_ASAP7_75t_L g1553 ( .A(n_1554), .B(n_1555), .Y(n_1553) );
INVx1_ASAP7_75t_L g1576 ( .A(n_1556), .Y(n_1576) );
AND2x2_ASAP7_75t_L g1592 ( .A(n_1556), .B(n_1593), .Y(n_1592) );
INVx1_ASAP7_75t_L g1626 ( .A(n_1556), .Y(n_1626) );
OR2x2_ASAP7_75t_L g1691 ( .A(n_1556), .B(n_1591), .Y(n_1691) );
NAND3xp33_ASAP7_75t_L g1735 ( .A(n_1556), .B(n_1561), .C(n_1662), .Y(n_1735) );
AND2x2_ASAP7_75t_L g1556 ( .A(n_1557), .B(n_1558), .Y(n_1556) );
OAI21xp33_ASAP7_75t_L g1697 ( .A1(n_1559), .A2(n_1698), .B(n_1701), .Y(n_1697) );
INVx1_ASAP7_75t_L g1559 ( .A(n_1560), .Y(n_1559) );
AND2x2_ASAP7_75t_L g1560 ( .A(n_1561), .B(n_1565), .Y(n_1560) );
INVx3_ASAP7_75t_L g1584 ( .A(n_1561), .Y(n_1584) );
INVx1_ASAP7_75t_L g1643 ( .A(n_1561), .Y(n_1643) );
AND2x2_ASAP7_75t_L g1649 ( .A(n_1561), .B(n_1566), .Y(n_1649) );
OR2x2_ASAP7_75t_L g1660 ( .A(n_1561), .B(n_1566), .Y(n_1660) );
NOR2xp33_ASAP7_75t_SL g1711 ( .A(n_1561), .B(n_1663), .Y(n_1711) );
OAI322xp33_ASAP7_75t_L g1753 ( .A1(n_1561), .A2(n_1599), .A3(n_1602), .B1(n_1648), .B2(n_1682), .C1(n_1754), .C2(n_1755), .Y(n_1753) );
AND2x2_ASAP7_75t_L g1561 ( .A(n_1562), .B(n_1563), .Y(n_1561) );
INVx1_ASAP7_75t_L g1565 ( .A(n_1566), .Y(n_1565) );
INVx2_ASAP7_75t_L g1577 ( .A(n_1566), .Y(n_1577) );
OR2x2_ASAP7_75t_L g1585 ( .A(n_1566), .B(n_1586), .Y(n_1585) );
AND2x2_ASAP7_75t_L g1621 ( .A(n_1566), .B(n_1584), .Y(n_1621) );
AND2x2_ASAP7_75t_L g1629 ( .A(n_1566), .B(n_1600), .Y(n_1629) );
OR2x2_ASAP7_75t_L g1638 ( .A(n_1566), .B(n_1587), .Y(n_1638) );
INVx2_ASAP7_75t_L g1566 ( .A(n_1567), .Y(n_1566) );
OR2x2_ASAP7_75t_L g1598 ( .A(n_1567), .B(n_1586), .Y(n_1598) );
NAND2xp5_ASAP7_75t_L g1567 ( .A(n_1568), .B(n_1569), .Y(n_1567) );
NAND2xp5_ASAP7_75t_L g1570 ( .A(n_1571), .B(n_1572), .Y(n_1570) );
CKINVDCx5p33_ASAP7_75t_R g1596 ( .A(n_1571), .Y(n_1596) );
NOR2xp33_ASAP7_75t_L g1610 ( .A(n_1571), .B(n_1611), .Y(n_1610) );
AND2x2_ASAP7_75t_L g1707 ( .A(n_1571), .B(n_1616), .Y(n_1707) );
OR2x2_ASAP7_75t_L g1721 ( .A(n_1571), .B(n_1686), .Y(n_1721) );
INVx1_ASAP7_75t_L g1572 ( .A(n_1573), .Y(n_1572) );
OAI211xp5_ASAP7_75t_L g1718 ( .A1(n_1573), .A2(n_1655), .B(n_1676), .C(n_1719), .Y(n_1718) );
OR2x2_ASAP7_75t_L g1573 ( .A(n_1574), .B(n_1575), .Y(n_1573) );
AND2x2_ASAP7_75t_L g1579 ( .A(n_1574), .B(n_1580), .Y(n_1579) );
NOR2xp33_ASAP7_75t_L g1613 ( .A(n_1574), .B(n_1593), .Y(n_1613) );
AND2x2_ASAP7_75t_L g1645 ( .A(n_1574), .B(n_1592), .Y(n_1645) );
AND2x2_ASAP7_75t_L g1714 ( .A(n_1574), .B(n_1699), .Y(n_1714) );
OR2x2_ASAP7_75t_L g1746 ( .A(n_1574), .B(n_1581), .Y(n_1746) );
OR2x2_ASAP7_75t_L g1605 ( .A(n_1575), .B(n_1606), .Y(n_1605) );
NAND2xp5_ASAP7_75t_L g1640 ( .A(n_1575), .B(n_1641), .Y(n_1640) );
OR2x2_ASAP7_75t_L g1686 ( .A(n_1575), .B(n_1591), .Y(n_1686) );
INVx1_ASAP7_75t_L g1751 ( .A(n_1575), .Y(n_1751) );
INVx1_ASAP7_75t_L g1678 ( .A(n_1577), .Y(n_1678) );
NAND2xp5_ASAP7_75t_L g1725 ( .A(n_1577), .B(n_1662), .Y(n_1725) );
AOI221xp5_ASAP7_75t_L g1578 ( .A1(n_1579), .A2(n_1582), .B1(n_1590), .B2(n_1594), .C(n_1601), .Y(n_1578) );
AND2x2_ASAP7_75t_L g1656 ( .A(n_1579), .B(n_1596), .Y(n_1656) );
AND2x2_ASAP7_75t_L g1652 ( .A(n_1580), .B(n_1653), .Y(n_1652) );
INVx1_ASAP7_75t_L g1580 ( .A(n_1581), .Y(n_1580) );
OR2x2_ASAP7_75t_L g1631 ( .A(n_1581), .B(n_1604), .Y(n_1631) );
INVx1_ASAP7_75t_L g1582 ( .A(n_1583), .Y(n_1582) );
OR2x2_ASAP7_75t_L g1583 ( .A(n_1584), .B(n_1585), .Y(n_1583) );
NAND2xp5_ASAP7_75t_L g1599 ( .A(n_1584), .B(n_1600), .Y(n_1599) );
OR2x2_ASAP7_75t_L g1607 ( .A(n_1584), .B(n_1600), .Y(n_1607) );
AND2x2_ASAP7_75t_L g1615 ( .A(n_1584), .B(n_1616), .Y(n_1615) );
OR2x2_ASAP7_75t_L g1635 ( .A(n_1584), .B(n_1598), .Y(n_1635) );
CKINVDCx14_ASAP7_75t_R g1696 ( .A(n_1584), .Y(n_1696) );
OR2x2_ASAP7_75t_L g1738 ( .A(n_1584), .B(n_1620), .Y(n_1738) );
CKINVDCx5p33_ASAP7_75t_R g1616 ( .A(n_1585), .Y(n_1616) );
INVx1_ASAP7_75t_L g1620 ( .A(n_1586), .Y(n_1620) );
NOR2xp33_ASAP7_75t_L g1728 ( .A(n_1586), .B(n_1729), .Y(n_1728) );
INVx1_ASAP7_75t_L g1586 ( .A(n_1587), .Y(n_1586) );
INVx1_ASAP7_75t_L g1600 ( .A(n_1587), .Y(n_1600) );
NAND2xp5_ASAP7_75t_L g1587 ( .A(n_1588), .B(n_1589), .Y(n_1587) );
INVx1_ASAP7_75t_L g1659 ( .A(n_1590), .Y(n_1659) );
AOI22xp5_ASAP7_75t_L g1723 ( .A1(n_1590), .A2(n_1646), .B1(n_1724), .B2(n_1726), .Y(n_1723) );
AND2x2_ASAP7_75t_L g1590 ( .A(n_1591), .B(n_1592), .Y(n_1590) );
NAND2xp5_ASAP7_75t_L g1676 ( .A(n_1591), .B(n_1677), .Y(n_1676) );
NAND2xp5_ASAP7_75t_L g1602 ( .A(n_1592), .B(n_1603), .Y(n_1602) );
NAND2xp5_ASAP7_75t_L g1633 ( .A(n_1592), .B(n_1634), .Y(n_1633) );
INVx1_ASAP7_75t_L g1641 ( .A(n_1592), .Y(n_1641) );
OAI311xp33_ASAP7_75t_L g1672 ( .A1(n_1593), .A2(n_1596), .A3(n_1673), .B1(n_1674), .C1(n_1688), .Y(n_1672) );
NAND2xp5_ASAP7_75t_L g1594 ( .A(n_1595), .B(n_1599), .Y(n_1594) );
NAND2xp5_ASAP7_75t_L g1595 ( .A(n_1596), .B(n_1597), .Y(n_1595) );
AND2x2_ASAP7_75t_L g1734 ( .A(n_1596), .B(n_1616), .Y(n_1734) );
O2A1O1Ixp33_ASAP7_75t_L g1752 ( .A1(n_1597), .A2(n_1675), .B(n_1740), .C(n_1753), .Y(n_1752) );
CKINVDCx5p33_ASAP7_75t_R g1597 ( .A(n_1598), .Y(n_1597) );
INVx2_ASAP7_75t_L g1655 ( .A(n_1600), .Y(n_1655) );
AND2x2_ASAP7_75t_L g1683 ( .A(n_1600), .B(n_1644), .Y(n_1683) );
AOI21xp33_ASAP7_75t_L g1601 ( .A1(n_1602), .A2(n_1605), .B(n_1607), .Y(n_1601) );
INVx1_ASAP7_75t_L g1603 ( .A(n_1604), .Y(n_1603) );
NOR2xp33_ASAP7_75t_L g1709 ( .A(n_1605), .B(n_1655), .Y(n_1709) );
INVx1_ASAP7_75t_L g1653 ( .A(n_1606), .Y(n_1653) );
O2A1O1Ixp33_ASAP7_75t_L g1712 ( .A1(n_1607), .A2(n_1646), .B(n_1713), .C(n_1715), .Y(n_1712) );
INVx1_ASAP7_75t_L g1744 ( .A(n_1607), .Y(n_1744) );
OAI211xp5_ASAP7_75t_SL g1608 ( .A1(n_1609), .A2(n_1614), .B(n_1617), .C(n_1636), .Y(n_1608) );
INVx1_ASAP7_75t_L g1609 ( .A(n_1610), .Y(n_1609) );
INVx1_ASAP7_75t_L g1611 ( .A(n_1612), .Y(n_1611) );
HB1xp67_ASAP7_75t_L g1612 ( .A(n_1613), .Y(n_1612) );
INVx1_ASAP7_75t_L g1614 ( .A(n_1615), .Y(n_1614) );
AOI211xp5_ASAP7_75t_L g1617 ( .A1(n_1618), .A2(n_1622), .B(n_1627), .C(n_1632), .Y(n_1617) );
INVx1_ASAP7_75t_L g1618 ( .A(n_1619), .Y(n_1618) );
NAND2xp5_ASAP7_75t_L g1619 ( .A(n_1620), .B(n_1621), .Y(n_1619) );
INVx1_ASAP7_75t_L g1651 ( .A(n_1620), .Y(n_1651) );
O2A1O1Ixp33_ASAP7_75t_L g1708 ( .A1(n_1620), .A2(n_1677), .B(n_1685), .C(n_1709), .Y(n_1708) );
AOI211xp5_ASAP7_75t_L g1717 ( .A1(n_1621), .A2(n_1718), .B(n_1722), .C(n_1730), .Y(n_1717) );
INVxp67_ASAP7_75t_SL g1622 ( .A(n_1623), .Y(n_1622) );
INVx1_ASAP7_75t_L g1624 ( .A(n_1625), .Y(n_1624) );
INVxp67_ASAP7_75t_SL g1627 ( .A(n_1628), .Y(n_1627) );
NAND2xp5_ASAP7_75t_L g1628 ( .A(n_1629), .B(n_1630), .Y(n_1628) );
NAND2xp5_ASAP7_75t_L g1687 ( .A(n_1629), .B(n_1645), .Y(n_1687) );
INVx1_ASAP7_75t_L g1630 ( .A(n_1631), .Y(n_1630) );
INVx1_ASAP7_75t_L g1632 ( .A(n_1633), .Y(n_1632) );
INVx1_ASAP7_75t_L g1634 ( .A(n_1635), .Y(n_1634) );
AOI21xp33_ASAP7_75t_L g1747 ( .A1(n_1635), .A2(n_1748), .B(n_1749), .Y(n_1747) );
INVx1_ASAP7_75t_L g1754 ( .A(n_1637), .Y(n_1754) );
INVx1_ASAP7_75t_L g1646 ( .A(n_1638), .Y(n_1646) );
OR2x2_ASAP7_75t_L g1673 ( .A(n_1638), .B(n_1643), .Y(n_1673) );
INVx1_ASAP7_75t_L g1639 ( .A(n_1640), .Y(n_1639) );
AND2x2_ASAP7_75t_L g1642 ( .A(n_1643), .B(n_1644), .Y(n_1642) );
OAI21xp33_ASAP7_75t_SL g1741 ( .A1(n_1643), .A2(n_1742), .B(n_1743), .Y(n_1741) );
INVx1_ASAP7_75t_L g1731 ( .A(n_1645), .Y(n_1731) );
OAI21xp33_ASAP7_75t_L g1736 ( .A1(n_1646), .A2(n_1720), .B(n_1737), .Y(n_1736) );
OAI211xp5_ASAP7_75t_L g1647 ( .A1(n_1648), .A2(n_1650), .B(n_1654), .C(n_1657), .Y(n_1647) );
INVx1_ASAP7_75t_L g1648 ( .A(n_1649), .Y(n_1648) );
NAND2xp5_ASAP7_75t_L g1701 ( .A(n_1649), .B(n_1702), .Y(n_1701) );
NAND2xp5_ASAP7_75t_L g1650 ( .A(n_1651), .B(n_1652), .Y(n_1650) );
AND2x2_ASAP7_75t_L g1689 ( .A(n_1651), .B(n_1690), .Y(n_1689) );
NAND2xp5_ASAP7_75t_L g1715 ( .A(n_1651), .B(n_1716), .Y(n_1715) );
INVx1_ASAP7_75t_L g1729 ( .A(n_1652), .Y(n_1729) );
NAND2xp5_ASAP7_75t_L g1654 ( .A(n_1655), .B(n_1656), .Y(n_1654) );
NAND2xp5_ASAP7_75t_SL g1719 ( .A(n_1655), .B(n_1720), .Y(n_1719) );
OR2x2_ASAP7_75t_L g1732 ( .A(n_1655), .B(n_1660), .Y(n_1732) );
INVx1_ASAP7_75t_L g1748 ( .A(n_1656), .Y(n_1748) );
INVx1_ASAP7_75t_L g1657 ( .A(n_1658), .Y(n_1657) );
INVx1_ASAP7_75t_L g1671 ( .A(n_1661), .Y(n_1671) );
INVx2_ASAP7_75t_L g1661 ( .A(n_1662), .Y(n_1661) );
INVx1_ASAP7_75t_L g1662 ( .A(n_1663), .Y(n_1662) );
INVx1_ASAP7_75t_L g1663 ( .A(n_1664), .Y(n_1663) );
OAI221xp5_ASAP7_75t_L g1664 ( .A1(n_1665), .A2(n_1666), .B1(n_1667), .B2(n_1668), .C(n_1669), .Y(n_1664) );
AOI211xp5_ASAP7_75t_L g1670 ( .A1(n_1671), .A2(n_1672), .B(n_1704), .C(n_1712), .Y(n_1670) );
AOI221xp5_ASAP7_75t_L g1739 ( .A1(n_1671), .A2(n_1685), .B1(n_1740), .B2(n_1741), .C(n_1747), .Y(n_1739) );
INVx1_ASAP7_75t_L g1740 ( .A(n_1673), .Y(n_1740) );
AOI21xp5_ASAP7_75t_SL g1674 ( .A1(n_1675), .A2(n_1678), .B(n_1679), .Y(n_1674) );
INVx1_ASAP7_75t_L g1675 ( .A(n_1676), .Y(n_1675) );
NAND3xp33_ASAP7_75t_L g1680 ( .A(n_1678), .B(n_1681), .C(n_1683), .Y(n_1680) );
NAND3xp33_ASAP7_75t_SL g1679 ( .A(n_1680), .B(n_1684), .C(n_1687), .Y(n_1679) );
INVx1_ASAP7_75t_L g1681 ( .A(n_1682), .Y(n_1681) );
INVx1_ASAP7_75t_L g1685 ( .A(n_1686), .Y(n_1685) );
O2A1O1Ixp33_ASAP7_75t_L g1688 ( .A1(n_1689), .A2(n_1692), .B(n_1696), .C(n_1697), .Y(n_1688) );
INVxp67_ASAP7_75t_SL g1755 ( .A(n_1692), .Y(n_1755) );
NOR2xp33_ASAP7_75t_L g1692 ( .A(n_1693), .B(n_1695), .Y(n_1692) );
INVx1_ASAP7_75t_L g1693 ( .A(n_1694), .Y(n_1693) );
INVx1_ASAP7_75t_L g1705 ( .A(n_1695), .Y(n_1705) );
INVx1_ASAP7_75t_L g1698 ( .A(n_1699), .Y(n_1698) );
O2A1O1Ixp33_ASAP7_75t_SL g1704 ( .A1(n_1705), .A2(n_1706), .B(n_1708), .C(n_1710), .Y(n_1704) );
INVx1_ASAP7_75t_L g1706 ( .A(n_1707), .Y(n_1706) );
INVx1_ASAP7_75t_L g1710 ( .A(n_1711), .Y(n_1710) );
INVx1_ASAP7_75t_L g1713 ( .A(n_1714), .Y(n_1713) );
INVx1_ASAP7_75t_L g1742 ( .A(n_1716), .Y(n_1742) );
INVx1_ASAP7_75t_L g1720 ( .A(n_1721), .Y(n_1720) );
INVx1_ASAP7_75t_L g1724 ( .A(n_1725), .Y(n_1724) );
INVx1_ASAP7_75t_L g1727 ( .A(n_1728), .Y(n_1727) );
OAI221xp5_ASAP7_75t_L g1730 ( .A1(n_1731), .A2(n_1732), .B1(n_1733), .B2(n_1735), .C(n_1736), .Y(n_1730) );
INVx1_ASAP7_75t_L g1733 ( .A(n_1734), .Y(n_1733) );
INVx1_ASAP7_75t_L g1737 ( .A(n_1738), .Y(n_1737) );
NAND2xp5_ASAP7_75t_L g1743 ( .A(n_1744), .B(n_1745), .Y(n_1743) );
INVx1_ASAP7_75t_L g1745 ( .A(n_1746), .Y(n_1745) );
INVx1_ASAP7_75t_L g1749 ( .A(n_1750), .Y(n_1749) );
CKINVDCx20_ASAP7_75t_R g1756 ( .A(n_1757), .Y(n_1756) );
CKINVDCx20_ASAP7_75t_R g1757 ( .A(n_1758), .Y(n_1757) );
INVx1_ASAP7_75t_L g1759 ( .A(n_1760), .Y(n_1759) );
HB1xp67_ASAP7_75t_L g1760 ( .A(n_1761), .Y(n_1760) );
XNOR2xp5_ASAP7_75t_L g1761 ( .A(n_1762), .B(n_1763), .Y(n_1761) );
NOR2x1_ASAP7_75t_L g1763 ( .A(n_1764), .B(n_1787), .Y(n_1763) );
NAND2xp5_ASAP7_75t_L g1764 ( .A(n_1765), .B(n_1768), .Y(n_1764) );
OAI211xp5_ASAP7_75t_L g1798 ( .A1(n_1776), .A2(n_1799), .B(n_1800), .C(n_1801), .Y(n_1798) );
NAND3xp33_ASAP7_75t_L g1787 ( .A(n_1788), .B(n_1802), .C(n_1804), .Y(n_1787) );
NOR3xp33_ASAP7_75t_SL g1788 ( .A(n_1789), .B(n_1796), .C(n_1797), .Y(n_1788) );
OAI21xp5_ASAP7_75t_SL g1789 ( .A1(n_1790), .A2(n_1792), .B(n_1793), .Y(n_1789) );
INVx3_ASAP7_75t_L g1806 ( .A(n_1807), .Y(n_1806) );
HB1xp67_ASAP7_75t_L g1810 ( .A(n_1811), .Y(n_1810) );
BUFx3_ASAP7_75t_L g1811 ( .A(n_1812), .Y(n_1811) );
BUFx3_ASAP7_75t_L g1812 ( .A(n_1813), .Y(n_1812) );
INVxp33_ASAP7_75t_SL g1814 ( .A(n_1815), .Y(n_1814) );
HB1xp67_ASAP7_75t_L g1816 ( .A(n_1817), .Y(n_1816) );
INVx1_ASAP7_75t_L g1817 ( .A(n_1818), .Y(n_1817) );
NAND3xp33_ASAP7_75t_L g1818 ( .A(n_1819), .B(n_1821), .C(n_1840), .Y(n_1818) );
NOR2xp33_ASAP7_75t_L g1821 ( .A(n_1822), .B(n_1826), .Y(n_1821) );
NAND3xp33_ASAP7_75t_SL g1826 ( .A(n_1827), .B(n_1830), .C(n_1833), .Y(n_1826) );
INVx1_ASAP7_75t_L g1835 ( .A(n_1836), .Y(n_1835) );
INVx1_ASAP7_75t_L g1838 ( .A(n_1839), .Y(n_1838) );
NAND3xp33_ASAP7_75t_L g1841 ( .A(n_1842), .B(n_1846), .C(n_1851), .Y(n_1841) );
INVx1_ASAP7_75t_L g1844 ( .A(n_1845), .Y(n_1844) );
AOI22xp33_ASAP7_75t_L g1846 ( .A1(n_1847), .A2(n_1848), .B1(n_1849), .B2(n_1850), .Y(n_1846) );
INVx1_ASAP7_75t_L g1855 ( .A(n_1856), .Y(n_1855) );
HB1xp67_ASAP7_75t_L g1858 ( .A(n_1859), .Y(n_1858) );
INVx1_ASAP7_75t_L g1861 ( .A(n_1862), .Y(n_1861) );
endmodule