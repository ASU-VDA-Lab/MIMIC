module real_aes_4100_n_8 (n_4, n_0, n_3, n_5, n_2, n_7, n_6, n_1, n_8);
input n_4;
input n_0;
input n_3;
input n_5;
input n_2;
input n_7;
input n_6;
input n_1;
output n_8;
wire n_17;
wire n_28;
wire n_22;
wire n_13;
wire n_24;
wire n_12;
wire n_19;
wire n_25;
wire n_14;
wire n_11;
wire n_16;
wire n_15;
wire n_27;
wire n_9;
wire n_23;
wire n_29;
wire n_20;
wire n_18;
wire n_26;
wire n_21;
wire n_10;
INVx1_ASAP7_75t_L g13 ( .A(n_0), .Y(n_13) );
NAND2xp5_ASAP7_75t_L g24 ( .A(n_0), .B(n_4), .Y(n_24) );
INVxp67_ASAP7_75t_L g18 ( .A(n_1), .Y(n_18) );
NAND3xp33_ASAP7_75t_L g15 ( .A(n_2), .B(n_16), .C(n_18), .Y(n_15) );
HB1xp67_ASAP7_75t_L g29 ( .A(n_3), .Y(n_29) );
NOR2xp33_ASAP7_75t_L g12 ( .A(n_4), .B(n_13), .Y(n_12) );
AND2x2_ASAP7_75t_L g16 ( .A(n_5), .B(n_17), .Y(n_16) );
INVx1_ASAP7_75t_L g28 ( .A(n_5), .Y(n_28) );
BUFx3_ASAP7_75t_L g20 ( .A(n_6), .Y(n_20) );
BUFx8_ASAP7_75t_SL g25 ( .A(n_6), .Y(n_25) );
INVx1_ASAP7_75t_L g17 ( .A(n_7), .Y(n_17) );
AOI221xp5_ASAP7_75t_L g8 ( .A1(n_9), .A2(n_19), .B1(n_21), .B2(n_25), .C(n_26), .Y(n_8) );
CKINVDCx5p33_ASAP7_75t_R g9 ( .A(n_10), .Y(n_9) );
INVx8_ASAP7_75t_L g10 ( .A(n_11), .Y(n_10) );
AND2x6_ASAP7_75t_SL g11 ( .A(n_12), .B(n_14), .Y(n_11) );
INVx1_ASAP7_75t_L g14 ( .A(n_15), .Y(n_14) );
OR2x2_ASAP7_75t_SL g23 ( .A(n_15), .B(n_24), .Y(n_23) );
NAND3xp33_ASAP7_75t_L g27 ( .A(n_17), .B(n_28), .C(n_29), .Y(n_27) );
CKINVDCx20_ASAP7_75t_R g19 ( .A(n_20), .Y(n_19) );
CKINVDCx11_ASAP7_75t_R g21 ( .A(n_22), .Y(n_21) );
BUFx12f_ASAP7_75t_L g22 ( .A(n_23), .Y(n_22) );
CKINVDCx5p33_ASAP7_75t_R g26 ( .A(n_27), .Y(n_26) );
endmodule