module fake_jpeg_29344_n_128 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_128);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_128;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_8),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_3),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_27),
.B(n_0),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_28),
.B(n_36),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_19),
.B(n_8),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_17),
.B(n_7),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_41),
.Y(n_45)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

INVx13_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

INVx13_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_19),
.B(n_9),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_42),
.B(n_22),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_30),
.A2(n_26),
.B1(n_22),
.B2(n_21),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_43),
.A2(n_29),
.B1(n_16),
.B2(n_23),
.Y(n_63)
);

AOI21xp33_ASAP7_75t_L g44 ( 
.A1(n_36),
.A2(n_23),
.B(n_18),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_44),
.B(n_50),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_33),
.B(n_21),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_52),
.B(n_54),
.Y(n_66)
);

AND2x4_ASAP7_75t_L g54 ( 
.A(n_28),
.B(n_0),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_42),
.B(n_20),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_56),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_32),
.B(n_20),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_61),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_63),
.Y(n_87)
);

INVx1_ASAP7_75t_SL g64 ( 
.A(n_55),
.Y(n_64)
);

INVx1_ASAP7_75t_SL g82 ( 
.A(n_64),
.Y(n_82)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_57),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_65),
.Y(n_77)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_67),
.B(n_69),
.Y(n_80)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_54),
.A2(n_39),
.B1(n_38),
.B2(n_18),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_70),
.A2(n_71),
.B1(n_74),
.B2(n_60),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_47),
.A2(n_29),
.B1(n_31),
.B2(n_34),
.Y(n_71)
);

OAI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_48),
.A2(n_31),
.B1(n_35),
.B2(n_40),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_72),
.A2(n_59),
.B1(n_51),
.B2(n_60),
.Y(n_86)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_73),
.Y(n_83)
);

OA22x2_ASAP7_75t_L g74 ( 
.A1(n_54),
.A2(n_48),
.B1(n_55),
.B2(n_49),
.Y(n_74)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_57),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_76),
.B(n_65),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_78),
.A2(n_84),
.B1(n_74),
.B2(n_64),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_68),
.B(n_45),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_79),
.B(n_81),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_68),
.B(n_75),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_70),
.A2(n_47),
.B1(n_49),
.B2(n_59),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_85),
.Y(n_93)
);

OR2x2_ASAP7_75t_L g90 ( 
.A(n_86),
.B(n_60),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_89),
.A2(n_90),
.B1(n_86),
.B2(n_93),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_80),
.B(n_75),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_91),
.B(n_92),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_SL g92 ( 
.A(n_78),
.B(n_66),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_87),
.B(n_66),
.C(n_62),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_94),
.A2(n_96),
.B(n_84),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_82),
.B(n_58),
.Y(n_95)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_95),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_87),
.B(n_74),
.C(n_67),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_97),
.B(n_77),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g98 ( 
.A1(n_96),
.A2(n_82),
.B(n_69),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_98),
.A2(n_102),
.B(n_94),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_SL g108 ( 
.A(n_100),
.B(n_58),
.Y(n_108)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_88),
.Y(n_101)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_101),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_SL g102 ( 
.A1(n_92),
.A2(n_74),
.B(n_54),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_104),
.B(n_83),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_103),
.B(n_83),
.C(n_90),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_106),
.B(n_108),
.C(n_73),
.Y(n_113)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_99),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_107),
.B(n_76),
.Y(n_114)
);

OAI322xp33_ASAP7_75t_L g109 ( 
.A1(n_102),
.A2(n_53),
.A3(n_13),
.B1(n_14),
.B2(n_12),
.C1(n_4),
.C2(n_11),
.Y(n_109)
);

NOR3xp33_ASAP7_75t_SL g115 ( 
.A(n_109),
.B(n_4),
.C(n_14),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_110),
.A2(n_97),
.B1(n_77),
.B2(n_98),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_111),
.B(n_113),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_112),
.B(n_106),
.C(n_104),
.Y(n_119)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_114),
.Y(n_117)
);

NAND4xp25_ASAP7_75t_L g116 ( 
.A(n_115),
.B(n_13),
.C(n_105),
.D(n_108),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_116),
.A2(n_1),
.B(n_2),
.Y(n_122)
);

MAJx2_ASAP7_75t_L g120 ( 
.A(n_119),
.B(n_112),
.C(n_115),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_120),
.B(n_121),
.C(n_122),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_118),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_120),
.A2(n_119),
.B(n_117),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_124),
.B(n_2),
.Y(n_125)
);

BUFx24_ASAP7_75t_SL g126 ( 
.A(n_125),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_126),
.B(n_123),
.C(n_3),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_127),
.B(n_3),
.Y(n_128)
);


endmodule