module fake_jpeg_26264_n_298 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_298);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_298;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_288;
wire n_272;
wire n_284;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_14),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

INVx2_ASAP7_75t_SL g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

INVx11_ASAP7_75t_SL g23 ( 
.A(n_11),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVx13_ASAP7_75t_L g31 ( 
.A(n_21),
.Y(n_31)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

AND2x2_ASAP7_75t_SL g41 ( 
.A(n_33),
.B(n_36),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_18),
.B(n_0),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_35),
.B(n_18),
.Y(n_52)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_38),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_35),
.B(n_20),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_43),
.B(n_44),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_35),
.B(n_15),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_32),
.A2(n_18),
.B1(n_20),
.B2(n_24),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_45),
.A2(n_31),
.B1(n_36),
.B2(n_33),
.Y(n_65)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_47),
.Y(n_55)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_50),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_35),
.A2(n_20),
.B1(n_18),
.B2(n_28),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_51),
.A2(n_36),
.B1(n_33),
.B2(n_26),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_52),
.B(n_31),
.Y(n_63)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_31),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_53),
.B(n_31),
.Y(n_70)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_32),
.Y(n_54)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

INVx1_ASAP7_75t_SL g107 ( 
.A(n_56),
.Y(n_107)
);

A2O1A1Ixp33_ASAP7_75t_L g58 ( 
.A1(n_43),
.A2(n_35),
.B(n_19),
.C(n_25),
.Y(n_58)
);

XNOR2xp5_ASAP7_75t_L g82 ( 
.A(n_58),
.B(n_72),
.Y(n_82)
);

OAI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_51),
.A2(n_32),
.B1(n_25),
.B2(n_19),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_59),
.A2(n_75),
.B1(n_33),
.B2(n_36),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_44),
.B(n_24),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_61),
.B(n_64),
.Y(n_89)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_62),
.B(n_71),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_63),
.A2(n_42),
.B1(n_33),
.B2(n_36),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_52),
.B(n_28),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_65),
.A2(n_48),
.B1(n_40),
.B2(n_31),
.Y(n_88)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_66),
.Y(n_83)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_67),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_68),
.A2(n_48),
.B1(n_39),
.B2(n_36),
.Y(n_94)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_70),
.Y(n_99)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_L g72 ( 
.A(n_45),
.B(n_15),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_41),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_73),
.Y(n_102)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_74),
.B(n_46),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_40),
.A2(n_22),
.B1(n_31),
.B2(n_29),
.Y(n_75)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_41),
.Y(n_77)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_77),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_50),
.B(n_19),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_78),
.B(n_79),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_41),
.B(n_21),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_41),
.B(n_37),
.C(n_34),
.Y(n_80)
);

XOR2xp5_ASAP7_75t_L g84 ( 
.A(n_80),
.B(n_31),
.Y(n_84)
);

NOR2x1_ASAP7_75t_R g81 ( 
.A(n_58),
.B(n_41),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_81),
.B(n_57),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_84),
.B(n_37),
.C(n_38),
.Y(n_111)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_76),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_85),
.B(n_87),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_88),
.A2(n_90),
.B1(n_104),
.B2(n_67),
.Y(n_113)
);

OA22x2_ASAP7_75t_L g90 ( 
.A1(n_73),
.A2(n_53),
.B1(n_42),
.B2(n_40),
.Y(n_90)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_76),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_92),
.B(n_95),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_77),
.A2(n_53),
.B1(n_42),
.B2(n_15),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_93),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_94),
.A2(n_98),
.B1(n_64),
.B2(n_61),
.Y(n_110)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_76),
.Y(n_95)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_55),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_96),
.B(n_103),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_97),
.B(n_38),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_68),
.A2(n_72),
.B1(n_63),
.B2(n_57),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_62),
.A2(n_28),
.B1(n_48),
.B2(n_39),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_100),
.A2(n_56),
.B1(n_66),
.B2(n_69),
.Y(n_116)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_101),
.Y(n_114)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_55),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_80),
.A2(n_33),
.B1(n_38),
.B2(n_37),
.Y(n_104)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_63),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_108),
.B(n_38),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_109),
.A2(n_113),
.B(n_121),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_110),
.B(n_129),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_111),
.B(n_122),
.C(n_34),
.Y(n_159)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_107),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_112),
.B(n_118),
.Y(n_144)
);

A2O1A1Ixp33_ASAP7_75t_SL g139 ( 
.A1(n_116),
.A2(n_88),
.B(n_90),
.C(n_97),
.Y(n_139)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_107),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_81),
.A2(n_74),
.B1(n_71),
.B2(n_69),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_120),
.A2(n_126),
.B1(n_128),
.B2(n_92),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_84),
.B(n_38),
.C(n_37),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_91),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_123),
.Y(n_156)
);

BUFx2_ASAP7_75t_L g124 ( 
.A(n_103),
.Y(n_124)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_124),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_82),
.B(n_27),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_125),
.B(n_135),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_104),
.A2(n_60),
.B1(n_22),
.B2(n_29),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_98),
.B(n_60),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_127),
.B(n_132),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_89),
.A2(n_22),
.B1(n_29),
.B2(n_24),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_96),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_94),
.A2(n_38),
.B1(n_37),
.B2(n_34),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_131),
.A2(n_95),
.B1(n_85),
.B2(n_83),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_106),
.B(n_26),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_99),
.B(n_22),
.Y(n_133)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_133),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_134),
.A2(n_105),
.B(n_86),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_82),
.B(n_38),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_135),
.B(n_90),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_119),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_137),
.B(n_141),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_139),
.A2(n_147),
.B1(n_130),
.B2(n_131),
.Y(n_171)
);

OAI32xp33_ASAP7_75t_L g140 ( 
.A1(n_109),
.A2(n_102),
.A3(n_108),
.B1(n_105),
.B2(n_89),
.Y(n_140)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_140),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_117),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_143),
.A2(n_153),
.B(n_16),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_145),
.B(n_152),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_116),
.Y(n_146)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_146),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_130),
.A2(n_99),
.B1(n_90),
.B2(n_86),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_148),
.A2(n_160),
.B1(n_153),
.B2(n_141),
.Y(n_188)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_124),
.Y(n_149)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_149),
.Y(n_169)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_124),
.Y(n_150)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_150),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_110),
.B(n_89),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_134),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_127),
.B(n_83),
.Y(n_154)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_154),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_SL g186 ( 
.A(n_157),
.B(n_166),
.Y(n_186)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_126),
.Y(n_158)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_158),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_159),
.B(n_164),
.C(n_34),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_160),
.A2(n_37),
.B1(n_34),
.B2(n_30),
.Y(n_181)
);

NAND4xp25_ASAP7_75t_SL g161 ( 
.A(n_115),
.B(n_46),
.C(n_27),
.D(n_30),
.Y(n_161)
);

HB1xp67_ASAP7_75t_L g183 ( 
.A(n_161),
.Y(n_183)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_120),
.Y(n_162)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_162),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_111),
.B(n_38),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_163),
.B(n_165),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_125),
.B(n_37),
.C(n_34),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_122),
.B(n_37),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_121),
.B(n_27),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_156),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_168),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_144),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_170),
.B(n_195),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_171),
.A2(n_176),
.B1(n_178),
.B2(n_182),
.Y(n_212)
);

OA21x2_ASAP7_75t_L g173 ( 
.A1(n_145),
.A2(n_113),
.B(n_114),
.Y(n_173)
);

INVx1_ASAP7_75t_SL g211 ( 
.A(n_173),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_138),
.A2(n_123),
.B(n_132),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_175),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_162),
.A2(n_114),
.B1(n_118),
.B2(n_129),
.Y(n_176)
);

OAI21xp33_ASAP7_75t_L g177 ( 
.A1(n_136),
.A2(n_128),
.B(n_112),
.Y(n_177)
);

XOR2x1_ASAP7_75t_L g204 ( 
.A(n_177),
.B(n_191),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_151),
.A2(n_26),
.B1(n_30),
.B2(n_17),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_143),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_179),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_181),
.A2(n_184),
.B1(n_188),
.B2(n_190),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_158),
.A2(n_30),
.B1(n_17),
.B2(n_16),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_139),
.A2(n_17),
.B1(n_16),
.B2(n_34),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_187),
.B(n_159),
.C(n_165),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_154),
.A2(n_17),
.B1(n_16),
.B2(n_34),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_139),
.A2(n_14),
.B1(n_13),
.B2(n_12),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_194),
.A2(n_155),
.B1(n_150),
.B2(n_149),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_138),
.A2(n_0),
.B(n_1),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_186),
.B(n_157),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_197),
.B(n_203),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_199),
.B(n_201),
.C(n_207),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_187),
.B(n_163),
.C(n_164),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_186),
.B(n_166),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_185),
.B(n_136),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_206),
.B(n_192),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_172),
.B(n_152),
.C(n_139),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g208 ( 
.A(n_176),
.B(n_194),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_208),
.B(n_214),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_175),
.B(n_139),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_209),
.B(n_215),
.C(n_216),
.Y(n_227)
);

OR2x2_ASAP7_75t_L g219 ( 
.A(n_210),
.B(n_171),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_174),
.A2(n_140),
.B1(n_142),
.B2(n_161),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_172),
.B(n_142),
.C(n_13),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_167),
.B(n_13),
.C(n_11),
.Y(n_216)
);

FAx1_ASAP7_75t_SL g217 ( 
.A(n_192),
.B(n_11),
.CI(n_10),
.CON(n_217),
.SN(n_217)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_217),
.B(n_216),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_167),
.B(n_10),
.C(n_1),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_218),
.B(n_195),
.C(n_191),
.Y(n_228)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_219),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_220),
.B(n_226),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_200),
.B(n_173),
.Y(n_221)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_221),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_213),
.A2(n_181),
.B1(n_170),
.B2(n_193),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_223),
.B(n_228),
.Y(n_246)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_225),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_208),
.A2(n_180),
.B1(n_196),
.B2(n_190),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_199),
.B(n_196),
.C(n_173),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_229),
.B(n_232),
.C(n_235),
.Y(n_251)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_217),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_230),
.B(n_231),
.Y(n_242)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_215),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_201),
.B(n_184),
.C(n_178),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_205),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_233),
.B(n_234),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_211),
.B(n_189),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_207),
.B(n_189),
.C(n_169),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_224),
.B(n_202),
.C(n_197),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_237),
.B(n_243),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_222),
.A2(n_213),
.B1(n_204),
.B2(n_211),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_239),
.B(n_244),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_SL g241 ( 
.A(n_236),
.B(n_203),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_241),
.B(n_250),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_224),
.B(n_235),
.C(n_229),
.Y(n_243)
);

BUFx24_ASAP7_75t_SL g244 ( 
.A(n_236),
.Y(n_244)
);

BUFx24_ASAP7_75t_SL g247 ( 
.A(n_219),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_247),
.B(n_169),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_227),
.B(n_209),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_245),
.B(n_227),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_252),
.B(n_253),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_251),
.B(n_232),
.C(n_228),
.Y(n_253)
);

INVx1_ASAP7_75t_SL g254 ( 
.A(n_248),
.Y(n_254)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_254),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_241),
.B(n_204),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_255),
.B(n_256),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_250),
.B(n_218),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_251),
.B(n_198),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_258),
.B(n_261),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_249),
.A2(n_212),
.B(n_182),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_260),
.B(n_262),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_246),
.B(n_183),
.Y(n_261)
);

INVxp67_ASAP7_75t_SL g262 ( 
.A(n_242),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_263),
.B(n_262),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_254),
.A2(n_240),
.B1(n_238),
.B2(n_2),
.Y(n_267)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_267),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_256),
.B(n_0),
.C(n_1),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_269),
.B(n_272),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_257),
.B(n_0),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_270),
.B(n_274),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_264),
.B(n_255),
.C(n_259),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_273),
.B(n_2),
.Y(n_276)
);

OAI21x1_ASAP7_75t_L g274 ( 
.A1(n_262),
.A2(n_2),
.B(n_3),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_276),
.B(n_277),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_271),
.B(n_4),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_275),
.B(n_4),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_279),
.B(n_280),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_268),
.B(n_5),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_SL g283 ( 
.A(n_272),
.B(n_5),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_283),
.B(n_6),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_278),
.B(n_266),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_285),
.A2(n_287),
.B(n_265),
.Y(n_292)
);

OAI21x1_ASAP7_75t_L g287 ( 
.A1(n_282),
.A2(n_269),
.B(n_270),
.Y(n_287)
);

A2O1A1Ixp33_ASAP7_75t_SL g290 ( 
.A1(n_288),
.A2(n_280),
.B(n_7),
.C(n_8),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_281),
.A2(n_265),
.B1(n_7),
.B2(n_8),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_289),
.A2(n_6),
.B(n_7),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_290),
.B(n_291),
.Y(n_293)
);

AOI321xp33_ASAP7_75t_L g294 ( 
.A1(n_293),
.A2(n_292),
.A3(n_286),
.B1(n_284),
.B2(n_9),
.C(n_8),
.Y(n_294)
);

HB1xp67_ASAP7_75t_L g295 ( 
.A(n_294),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_295),
.B(n_6),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_296),
.B(n_6),
.C(n_7),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_297),
.A2(n_9),
.B(n_286),
.Y(n_298)
);


endmodule