module real_jpeg_3888_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_0),
.Y(n_61)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_0),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_0),
.Y(n_82)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_0),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_0),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_0),
.Y(n_93)
);

BUFx5_ASAP7_75t_L g101 ( 
.A(n_0),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_0),
.Y(n_150)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_1),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_2),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_3),
.A2(n_46),
.B1(n_49),
.B2(n_50),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_3),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_3),
.A2(n_49),
.B1(n_82),
.B2(n_83),
.Y(n_81)
);

OAI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_3),
.A2(n_49),
.B1(n_141),
.B2(n_143),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_3),
.A2(n_49),
.B1(n_189),
.B2(n_191),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_4),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_4),
.A2(n_66),
.B1(n_119),
.B2(n_120),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_4),
.A2(n_66),
.B1(n_174),
.B2(n_178),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_4),
.A2(n_31),
.B1(n_66),
.B2(n_203),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_4),
.B(n_73),
.Y(n_238)
);

O2A1O1Ixp33_ASAP7_75t_L g254 ( 
.A1(n_4),
.A2(n_255),
.B(n_257),
.C(n_263),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_4),
.B(n_28),
.C(n_160),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_4),
.B(n_146),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_4),
.B(n_319),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_4),
.B(n_164),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_5),
.A2(n_88),
.B1(n_89),
.B2(n_90),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_5),
.Y(n_89)
);

OAI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_5),
.A2(n_89),
.B1(n_133),
.B2(n_134),
.Y(n_132)
);

OAI22xp33_ASAP7_75t_SL g272 ( 
.A1(n_5),
.A2(n_89),
.B1(n_273),
.B2(n_274),
.Y(n_272)
);

AOI22xp33_ASAP7_75t_L g293 ( 
.A1(n_5),
.A2(n_89),
.B1(n_294),
.B2(n_296),
.Y(n_293)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_6),
.Y(n_108)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g311 ( 
.A(n_7),
.Y(n_311)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_8),
.Y(n_60)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_8),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_8),
.Y(n_80)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_8),
.Y(n_97)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_10),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g14 ( 
.A1(n_11),
.A2(n_15),
.B1(n_18),
.B2(n_19),
.Y(n_14)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_12),
.A2(n_27),
.B1(n_28),
.B2(n_30),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_12),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_12),
.A2(n_27),
.B1(n_209),
.B2(n_211),
.Y(n_208)
);

BUFx5_ASAP7_75t_L g160 ( 
.A(n_13),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_13),
.Y(n_161)
);

BUFx3_ASAP7_75t_L g166 ( 
.A(n_13),
.Y(n_166)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_13),
.Y(n_170)
);

INVx13_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

INVx8_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

INVx13_ASAP7_75t_L g18 ( 
.A(n_17),
.Y(n_18)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_225),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_223),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_194),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_22),
.B(n_194),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_135),
.C(n_179),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_23),
.B(n_242),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_70),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_24),
.B(n_71),
.C(n_102),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g24 ( 
.A(n_25),
.B(n_52),
.Y(n_24)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_25),
.B(n_52),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_36),
.B(n_39),
.Y(n_25)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_26),
.A2(n_181),
.B(n_182),
.Y(n_180)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_29),
.Y(n_168)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_29),
.Y(n_297)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx4_ASAP7_75t_SL g31 ( 
.A(n_32),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_35),
.Y(n_205)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_38),
.Y(n_184)
);

INVx4_ASAP7_75t_L g319 ( 
.A(n_38),
.Y(n_319)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_39),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_45),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_40),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_40),
.B(n_202),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_40),
.A2(n_202),
.B(n_266),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_40),
.B(n_293),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_43),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx4_ASAP7_75t_L g200 ( 
.A(n_43),
.Y(n_200)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_45),
.B(n_183),
.Y(n_182)
);

INVx1_ASAP7_75t_SL g46 ( 
.A(n_47),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_48),
.Y(n_167)
);

BUFx8_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g317 ( 
.A(n_51),
.Y(n_317)
);

AOI32xp33_ASAP7_75t_L g52 ( 
.A1(n_53),
.A2(n_58),
.A3(n_61),
.B1(n_62),
.B2(n_67),
.Y(n_52)
);

HB1xp67_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_54),
.Y(n_133)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx5_ASAP7_75t_L g119 ( 
.A(n_56),
.Y(n_119)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_57),
.Y(n_68)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_57),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_57),
.Y(n_77)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_57),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_57),
.Y(n_144)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVxp33_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_63),
.A2(n_66),
.B(n_150),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_64),
.B(n_66),
.Y(n_63)
);

INVx1_ASAP7_75t_SL g90 ( 
.A(n_64),
.Y(n_90)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

OAI21xp33_ASAP7_75t_L g257 ( 
.A1(n_66),
.A2(n_258),
.B(n_260),
.Y(n_257)
);

NAND2xp33_ASAP7_75t_SL g67 ( 
.A(n_68),
.B(n_69),
.Y(n_67)
);

HB1xp67_ASAP7_75t_L g131 ( 
.A(n_68),
.Y(n_131)
);

AO22x1_ASAP7_75t_SL g73 ( 
.A1(n_69),
.A2(n_74),
.B1(n_76),
.B2(n_78),
.Y(n_73)
);

XOR2xp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_102),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_86),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_81),
.Y(n_72)
);

NOR2x1_ASAP7_75t_L g91 ( 
.A(n_73),
.B(n_92),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_73),
.B(n_87),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_74),
.A2(n_128),
.B1(n_130),
.B2(n_131),
.Y(n_127)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx6_ASAP7_75t_SL g76 ( 
.A(n_77),
.Y(n_76)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_80),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_81),
.B(n_91),
.Y(n_220)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_91),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_91),
.B(n_149),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_93),
.A2(n_94),
.B1(n_98),
.B2(n_100),
.Y(n_92)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_124),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_117),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_105),
.B(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_105),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_109),
.B1(n_111),
.B2(n_114),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_107),
.Y(n_116)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_108),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g130 ( 
.A(n_108),
.Y(n_130)
);

INVx3_ASAP7_75t_L g259 ( 
.A(n_108),
.Y(n_259)
);

BUFx5_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx11_ASAP7_75t_L g113 ( 
.A(n_110),
.Y(n_113)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_110),
.Y(n_158)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_110),
.Y(n_163)
);

BUFx3_ASAP7_75t_L g177 ( 
.A(n_110),
.Y(n_177)
);

BUFx3_ASAP7_75t_L g193 ( 
.A(n_110),
.Y(n_193)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_110),
.Y(n_262)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_111),
.Y(n_190)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx6_ASAP7_75t_L g276 ( 
.A(n_113),
.Y(n_276)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVxp67_ASAP7_75t_SL g117 ( 
.A(n_118),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_118),
.A2(n_125),
.B(n_146),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_118),
.B(n_125),
.Y(n_334)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_119),
.Y(n_134)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

BUFx12f_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_122),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_124),
.B(n_236),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_125),
.B(n_132),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_126),
.B(n_139),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx4_ASAP7_75t_L g256 ( 
.A(n_129),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_132),
.B(n_146),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_135),
.B(n_179),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_147),
.C(n_152),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_136),
.A2(n_152),
.B1(n_230),
.B2(n_231),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_136),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_137),
.B(n_145),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_140),
.B(n_146),
.Y(n_236)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx3_ASAP7_75t_L g264 ( 
.A(n_144),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_145),
.B(n_334),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_SL g228 ( 
.A(n_147),
.B(n_229),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_148),
.B(n_151),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_151),
.B(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_152),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_153),
.A2(n_171),
.B(n_172),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_154),
.B(n_173),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_154),
.B(n_188),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_154),
.B(n_272),
.Y(n_271)
);

NOR2x1_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_164),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_159),
.B1(n_161),
.B2(n_162),
.Y(n_155)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_158),
.Y(n_273)
);

INVx4_ASAP7_75t_SL g159 ( 
.A(n_160),
.Y(n_159)
);

INVx5_ASAP7_75t_L g210 ( 
.A(n_162),
.Y(n_210)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_163),
.Y(n_178)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_164),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_164),
.B(n_188),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_164),
.B(n_272),
.Y(n_288)
);

AO22x1_ASAP7_75t_SL g164 ( 
.A1(n_165),
.A2(n_167),
.B1(n_168),
.B2(n_169),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx4_ASAP7_75t_L g295 ( 
.A(n_167),
.Y(n_295)
);

BUFx5_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_171),
.A2(n_208),
.B(n_214),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_171),
.B(n_172),
.Y(n_270)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx4_ASAP7_75t_SL g213 ( 
.A(n_178),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_185),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_180),
.B(n_185),
.Y(n_216)
);

OR2x2_ASAP7_75t_L g239 ( 
.A(n_182),
.B(n_240),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g322 ( 
.A(n_182),
.B(n_292),
.Y(n_322)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

AND2x2_ASAP7_75t_SL g185 ( 
.A(n_186),
.B(n_187),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_186),
.B(n_288),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_187),
.B(n_271),
.Y(n_299)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_196),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_215),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_207),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_206),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_199),
.B(n_291),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_201),
.Y(n_199)
);

INVx1_ASAP7_75t_SL g266 ( 
.A(n_200),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx4_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx8_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_206),
.B(n_308),
.Y(n_307)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_214),
.B(n_288),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_217),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_218),
.A2(n_219),
.B1(n_221),
.B2(n_222),
.Y(n_217)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_218),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_219),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_226),
.A2(n_243),
.B(n_346),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_241),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_227),
.B(n_241),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_232),
.C(n_234),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_228),
.B(n_247),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_232),
.A2(n_233),
.B1(n_234),
.B2(n_248),
.Y(n_247)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_234),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_237),
.C(n_239),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_235),
.B(n_251),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_237),
.A2(n_238),
.B1(n_239),
.B2(n_252),
.Y(n_251)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g252 ( 
.A(n_239),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_240),
.B(n_309),
.Y(n_320)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g244 ( 
.A1(n_245),
.A2(n_277),
.B(n_345),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_246),
.B(n_249),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_246),
.B(n_249),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_253),
.C(n_267),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g340 ( 
.A(n_250),
.B(n_341),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_253),
.A2(n_267),
.B1(n_268),
.B2(n_342),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_253),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_265),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g335 ( 
.A1(n_254),
.A2(n_265),
.B1(n_336),
.B2(n_337),
.Y(n_335)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_254),
.Y(n_337)
);

INVx8_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx6_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

BUFx3_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx4_ASAP7_75t_L g285 ( 
.A(n_262),
.Y(n_285)
);

INVx4_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_265),
.Y(n_336)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_271),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx3_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx6_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_278),
.A2(n_339),
.B(n_344),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_279),
.A2(n_327),
.B(n_338),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_280),
.A2(n_303),
.B(n_326),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_289),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_281),
.B(n_289),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_287),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_282),
.A2(n_283),
.B1(n_287),
.B2(n_306),
.Y(n_305)
);

CKINVDCx16_ASAP7_75t_R g282 ( 
.A(n_283),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_286),
.Y(n_283)
);

INVx4_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_287),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_298),
.Y(n_289)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_290),
.Y(n_329)
);

INVxp67_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_293),
.B(n_310),
.Y(n_309)
);

INVx6_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx6_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_299),
.A2(n_300),
.B1(n_301),
.B2(n_302),
.Y(n_298)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_299),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_300),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_300),
.B(n_301),
.C(n_329),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_304),
.A2(n_312),
.B(n_325),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_305),
.B(n_307),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_305),
.B(n_307),
.Y(n_325)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_313),
.A2(n_321),
.B(n_324),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_320),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_318),
.Y(n_314)
);

INVx1_ASAP7_75t_SL g315 ( 
.A(n_316),
.Y(n_315)
);

INVx3_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_322),
.B(n_323),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_322),
.B(n_323),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_330),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_328),
.B(n_330),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_331),
.B(n_335),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_332),
.B(n_333),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_332),
.B(n_333),
.C(n_335),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_340),
.B(n_343),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_340),
.B(n_343),
.Y(n_344)
);


endmodule