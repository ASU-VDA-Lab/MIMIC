module fake_jpeg_21640_n_168 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_168);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_168;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_57;
wire n_21;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_140;
wire n_96;

BUFx3_ASAP7_75t_L g11 ( 
.A(n_9),
.Y(n_11)
);

BUFx12f_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

BUFx5_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

BUFx24_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

INVx11_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_10),
.Y(n_17)
);

BUFx6f_ASAP7_75t_SL g18 ( 
.A(n_3),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_15),
.Y(n_22)
);

INVx4_ASAP7_75t_SL g38 ( 
.A(n_22),
.Y(n_38)
);

INVx5_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

BUFx4f_ASAP7_75t_SL g32 ( 
.A(n_24),
.Y(n_32)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_25),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_18),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_26),
.B(n_29),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

INVx4_ASAP7_75t_SL g39 ( 
.A(n_28),
.Y(n_39)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_18),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_30),
.B(n_12),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_26),
.A2(n_14),
.B1(n_19),
.B2(n_17),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_40),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g34 ( 
.A(n_29),
.B(n_12),
.C(n_20),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_42),
.Y(n_43)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_26),
.A2(n_14),
.B1(n_19),
.B2(n_17),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_29),
.B(n_12),
.C(n_20),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_36),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_44),
.B(n_49),
.Y(n_59)
);

MAJx2_ASAP7_75t_L g46 ( 
.A(n_37),
.B(n_18),
.C(n_29),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_46),
.B(n_50),
.C(n_56),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_38),
.A2(n_16),
.B1(n_29),
.B2(n_23),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_38),
.A2(n_16),
.B1(n_23),
.B2(n_30),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_33),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_31),
.B(n_28),
.Y(n_50)
);

INVx2_ASAP7_75t_R g52 ( 
.A(n_38),
.Y(n_52)
);

OAI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_52),
.A2(n_53),
.B1(n_39),
.B2(n_35),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_35),
.A2(n_16),
.B1(n_23),
.B2(n_30),
.Y(n_53)
);

BUFx2_ASAP7_75t_L g54 ( 
.A(n_32),
.Y(n_54)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_54),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_31),
.Y(n_55)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_55),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_34),
.B(n_28),
.Y(n_56)
);

XOR2xp5_ASAP7_75t_L g57 ( 
.A(n_56),
.B(n_42),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_57),
.B(n_70),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_44),
.B(n_21),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_58),
.B(n_69),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_61),
.A2(n_67),
.B1(n_43),
.B2(n_51),
.Y(n_77)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_54),
.Y(n_65)
);

INVx3_ASAP7_75t_SL g75 ( 
.A(n_65),
.Y(n_75)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_66),
.Y(n_79)
);

OAI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_49),
.A2(n_55),
.B1(n_51),
.B2(n_45),
.Y(n_67)
);

AND2x6_ASAP7_75t_L g69 ( 
.A(n_43),
.B(n_13),
.Y(n_69)
);

AND2x6_ASAP7_75t_L g70 ( 
.A(n_43),
.B(n_13),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_59),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_72),
.B(n_82),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_69),
.A2(n_70),
.B1(n_63),
.B2(n_68),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_73),
.A2(n_83),
.B1(n_60),
.B2(n_24),
.Y(n_93)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_62),
.Y(n_74)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_74),
.Y(n_94)
);

OR2x2_ASAP7_75t_L g76 ( 
.A(n_68),
.B(n_52),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_76),
.B(n_77),
.Y(n_97)
);

OA21x2_ASAP7_75t_L g78 ( 
.A1(n_64),
.A2(n_45),
.B(n_52),
.Y(n_78)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_78),
.Y(n_96)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_62),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_80),
.Y(n_88)
);

INVx1_ASAP7_75t_SL g82 ( 
.A(n_65),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_64),
.A2(n_46),
.B1(n_39),
.B2(n_41),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_83),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_84),
.B(n_89),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_76),
.B(n_57),
.C(n_46),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_86),
.B(n_87),
.C(n_73),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g87 ( 
.A(n_71),
.B(n_60),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_72),
.B(n_21),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_74),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_90),
.B(n_91),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_81),
.B(n_14),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_79),
.B(n_54),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_92),
.B(n_95),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_93),
.A2(n_22),
.B(n_25),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_76),
.Y(n_95)
);

HB1xp67_ASAP7_75t_L g98 ( 
.A(n_97),
.Y(n_98)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_98),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_SL g118 ( 
.A(n_101),
.B(n_88),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_96),
.A2(n_78),
.B1(n_77),
.B2(n_80),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_102),
.A2(n_106),
.B1(n_110),
.B2(n_84),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_96),
.A2(n_71),
.B(n_78),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_103),
.A2(n_109),
.B1(n_75),
.B2(n_41),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_86),
.B(n_78),
.C(n_81),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_104),
.B(n_105),
.Y(n_112)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_94),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_90),
.A2(n_79),
.B1(n_75),
.B2(n_82),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_97),
.B(n_75),
.C(n_28),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_107),
.B(n_108),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_93),
.A2(n_87),
.B(n_95),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_94),
.Y(n_109)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_113),
.Y(n_127)
);

HB1xp67_ASAP7_75t_L g114 ( 
.A(n_106),
.Y(n_114)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_114),
.Y(n_130)
);

HB1xp67_ASAP7_75t_L g115 ( 
.A(n_107),
.Y(n_115)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_115),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_101),
.B(n_85),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_117),
.B(n_118),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_119),
.B(n_120),
.Y(n_128)
);

NOR3xp33_ASAP7_75t_SL g120 ( 
.A(n_100),
.B(n_13),
.C(n_11),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_99),
.A2(n_39),
.B1(n_35),
.B2(n_24),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_121),
.A2(n_25),
.B(n_22),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_104),
.A2(n_103),
.B1(n_111),
.B2(n_110),
.Y(n_123)
);

AO221x1_ASAP7_75t_L g125 ( 
.A1(n_123),
.A2(n_11),
.B1(n_12),
.B2(n_32),
.C(n_20),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_101),
.B(n_11),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_124),
.B(n_28),
.C(n_27),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_125),
.A2(n_24),
.B1(n_112),
.B2(n_120),
.Y(n_140)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_131),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_132),
.B(n_24),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_117),
.B(n_27),
.C(n_32),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_133),
.B(n_124),
.C(n_118),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_122),
.A2(n_32),
.B(n_1),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_134),
.B(n_121),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_135),
.A2(n_140),
.B1(n_131),
.B2(n_127),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_126),
.B(n_116),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_137),
.B(n_138),
.Y(n_147)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_134),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_139),
.B(n_129),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_130),
.A2(n_7),
.B(n_2),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_141),
.A2(n_132),
.B(n_133),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_142),
.B(n_143),
.Y(n_148)
);

NOR3xp33_ASAP7_75t_SL g143 ( 
.A(n_128),
.B(n_6),
.C(n_2),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_144),
.B(n_145),
.Y(n_153)
);

MAJx2_ASAP7_75t_L g146 ( 
.A(n_139),
.B(n_129),
.C(n_126),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_146),
.A2(n_143),
.B(n_3),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_136),
.B(n_142),
.Y(n_149)
);

OR2x2_ASAP7_75t_L g152 ( 
.A(n_149),
.B(n_148),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_150),
.B(n_27),
.C(n_3),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_151),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_152),
.B(n_154),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_147),
.B(n_27),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_147),
.B(n_7),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_155),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_160)
);

NOR2xp67_ASAP7_75t_L g157 ( 
.A(n_156),
.B(n_7),
.Y(n_157)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_157),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_160),
.B(n_153),
.C(n_5),
.Y(n_162)
);

AO21x1_ASAP7_75t_L g165 ( 
.A1(n_162),
.A2(n_8),
.B(n_9),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_159),
.B(n_5),
.C(n_6),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_163),
.A2(n_158),
.B(n_8),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_164),
.A2(n_165),
.B(n_161),
.Y(n_166)
);

O2A1O1Ixp33_ASAP7_75t_SL g167 ( 
.A1(n_166),
.A2(n_0),
.B(n_10),
.C(n_157),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_167),
.B(n_0),
.Y(n_168)
);


endmodule