module fake_jpeg_13279_n_111 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_111);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_111;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_106;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

BUFx12_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_2),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

BUFx10_ASAP7_75t_L g45 ( 
.A(n_4),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_12),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_48),
.Y(n_60)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_40),
.A2(n_15),
.B1(n_34),
.B2(n_33),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_50),
.B(n_4),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_43),
.B(n_0),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_51),
.B(n_52),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_0),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_39),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_53),
.B(n_54),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_44),
.B(n_1),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_44),
.B(n_2),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_55),
.B(n_5),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_53),
.B(n_3),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_57),
.B(n_61),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_59),
.B(n_6),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_49),
.B(n_5),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_62),
.B(n_67),
.Y(n_79)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_63),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_64),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_65),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_52),
.B(n_6),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_58),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_68),
.B(n_69),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_66),
.B(n_37),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_73),
.B(n_7),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_63),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_74),
.B(n_36),
.Y(n_83)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_60),
.Y(n_76)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_76),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_56),
.B(n_36),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_77),
.B(n_14),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_64),
.A2(n_47),
.B1(n_46),
.B2(n_45),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_78),
.A2(n_65),
.B1(n_60),
.B2(n_64),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_L g80 ( 
.A1(n_59),
.A2(n_45),
.B(n_37),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_80),
.A2(n_42),
.B(n_8),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_81),
.B(n_83),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_72),
.A2(n_42),
.B1(n_39),
.B2(n_9),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_84),
.B(n_87),
.Y(n_98)
);

NAND3xp33_ASAP7_75t_L g94 ( 
.A(n_85),
.B(n_88),
.C(n_90),
.Y(n_94)
);

OAI22xp33_ASAP7_75t_L g87 ( 
.A1(n_72),
.A2(n_20),
.B1(n_28),
.B2(n_27),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_80),
.B(n_18),
.C(n_26),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_89),
.B(n_70),
.C(n_79),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_79),
.B(n_7),
.Y(n_90)
);

NAND2xp67_ASAP7_75t_SL g91 ( 
.A(n_69),
.B(n_19),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_91),
.B(n_92),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_93),
.B(n_95),
.C(n_100),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_82),
.B(n_73),
.C(n_78),
.Y(n_95)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_86),
.Y(n_97)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_97),
.B(n_8),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_89),
.B(n_87),
.C(n_91),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_96),
.A2(n_84),
.B1(n_75),
.B2(n_71),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_101),
.A2(n_98),
.B1(n_94),
.B2(n_99),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_99),
.B(n_21),
.Y(n_102)
);

OAI221xp5_ASAP7_75t_L g106 ( 
.A1(n_102),
.A2(n_104),
.B1(n_9),
.B2(n_10),
.C(n_11),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_105),
.B(n_106),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_107),
.Y(n_108)
);

OR2x2_ASAP7_75t_L g109 ( 
.A(n_108),
.B(n_102),
.Y(n_109)
);

AOI321xp33_ASAP7_75t_L g110 ( 
.A1(n_109),
.A2(n_103),
.A3(n_23),
.B1(n_13),
.B2(n_22),
.C(n_25),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_110),
.B(n_35),
.Y(n_111)
);


endmodule