module fake_jpeg_10694_n_260 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_260);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_260;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_219;
wire n_70;
wire n_121;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_96;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx2_ASAP7_75t_SL g19 ( 
.A(n_13),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_12),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_5),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_12),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

INVx13_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_34),
.Y(n_36)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_26),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_37),
.B(n_43),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

INVx13_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_20),
.B(n_0),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_15),
.Y(n_44)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_19),
.Y(n_46)
);

HB1xp67_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

INVx2_ASAP7_75t_SL g47 ( 
.A(n_22),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_47),
.B(n_22),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_36),
.A2(n_41),
.B1(n_40),
.B2(n_21),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_50),
.A2(n_54),
.B1(n_56),
.B2(n_64),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_47),
.A2(n_19),
.B1(n_17),
.B2(n_21),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_51),
.A2(n_29),
.B1(n_17),
.B2(n_44),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_42),
.A2(n_21),
.B1(n_15),
.B2(n_23),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_37),
.B(n_30),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_55),
.B(n_61),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_42),
.A2(n_15),
.B1(n_18),
.B2(n_23),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_43),
.B(n_30),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_57),
.B(n_31),
.Y(n_101)
);

NAND2xp33_ASAP7_75t_SL g92 ( 
.A(n_59),
.B(n_47),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_45),
.B(n_33),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_44),
.A2(n_23),
.B1(n_18),
.B2(n_25),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_48),
.B(n_32),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_68),
.B(n_78),
.Y(n_114)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_60),
.Y(n_69)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_69),
.Y(n_124)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_60),
.Y(n_71)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_71),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_61),
.B(n_33),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_72),
.B(n_82),
.Y(n_112)
);

CKINVDCx12_ASAP7_75t_R g73 ( 
.A(n_49),
.Y(n_73)
);

INVx13_ASAP7_75t_L g116 ( 
.A(n_73),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_SL g74 ( 
.A1(n_55),
.A2(n_46),
.B(n_47),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_74),
.A2(n_109),
.B(n_26),
.Y(n_140)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_66),
.Y(n_75)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_75),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_59),
.B(n_38),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_76),
.B(n_87),
.Y(n_122)
);

OR2x2_ASAP7_75t_L g77 ( 
.A(n_53),
.B(n_24),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_77),
.B(n_79),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_48),
.B(n_20),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_65),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_57),
.B(n_27),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_80),
.Y(n_130)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_62),
.Y(n_81)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_81),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_53),
.B(n_16),
.Y(n_82)
);

OR2x2_ASAP7_75t_L g83 ( 
.A(n_58),
.B(n_16),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_83),
.B(n_84),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_58),
.B(n_32),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_59),
.Y(n_85)
);

INVx13_ASAP7_75t_L g128 ( 
.A(n_85),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_49),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_86),
.B(n_89),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_66),
.B(n_38),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_52),
.B(n_27),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_88),
.A2(n_97),
.B1(n_103),
.B2(n_104),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_52),
.B(n_25),
.Y(n_89)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_62),
.Y(n_90)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_90),
.Y(n_119)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_63),
.Y(n_91)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_91),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_92),
.B(n_93),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_52),
.B(n_25),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_50),
.B(n_31),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_94),
.Y(n_117)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_63),
.Y(n_95)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_95),
.Y(n_136)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_67),
.Y(n_96)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_96),
.Y(n_111)
);

NOR3xp33_ASAP7_75t_L g97 ( 
.A(n_67),
.B(n_16),
.C(n_24),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_64),
.B(n_22),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_98),
.A2(n_107),
.B(n_28),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_67),
.B(n_24),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_99),
.A2(n_101),
.B1(n_102),
.B2(n_106),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_54),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_100),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_56),
.B(n_33),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_60),
.Y(n_103)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_49),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_57),
.B(n_28),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_48),
.B(n_28),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_108),
.A2(n_86),
.B1(n_104),
.B2(n_77),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_59),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_70),
.A2(n_23),
.B1(n_18),
.B2(n_17),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_113),
.A2(n_129),
.B1(n_87),
.B2(n_96),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_115),
.B(n_93),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_105),
.A2(n_18),
.B1(n_35),
.B2(n_39),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_118),
.A2(n_123),
.B1(n_125),
.B2(n_89),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_98),
.A2(n_109),
.B1(n_85),
.B2(n_79),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_98),
.A2(n_39),
.B1(n_35),
.B2(n_26),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_70),
.A2(n_26),
.B1(n_1),
.B2(n_2),
.Y(n_129)
);

AND2x6_ASAP7_75t_L g134 ( 
.A(n_74),
.B(n_0),
.Y(n_134)
);

NOR3xp33_ASAP7_75t_SL g156 ( 
.A(n_134),
.B(n_1),
.C(n_4),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_138),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_140),
.B(n_76),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_132),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_141),
.B(n_145),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_142),
.A2(n_144),
.B1(n_150),
.B2(n_154),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_143),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_120),
.A2(n_72),
.B1(n_83),
.B2(n_99),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_132),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_114),
.B(n_82),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_146),
.B(n_157),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_147),
.B(n_151),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_140),
.A2(n_103),
.B(n_76),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_148),
.A2(n_164),
.B(n_124),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_118),
.A2(n_95),
.B1(n_69),
.B2(n_71),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_122),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_112),
.B(n_87),
.C(n_75),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_152),
.B(n_131),
.C(n_136),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_153),
.B(n_156),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_112),
.A2(n_91),
.B1(n_90),
.B2(n_81),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_113),
.A2(n_26),
.B1(n_3),
.B2(n_4),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_155),
.A2(n_125),
.B1(n_115),
.B2(n_111),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_117),
.B(n_1),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_122),
.Y(n_158)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_158),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_139),
.B(n_4),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_159),
.B(n_160),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_133),
.B(n_6),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_137),
.B(n_6),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_161),
.B(n_129),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_130),
.B(n_6),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_162),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_134),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_163),
.A2(n_130),
.B1(n_119),
.B2(n_135),
.Y(n_172)
);

AND2x4_ASAP7_75t_L g164 ( 
.A(n_128),
.B(n_14),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_122),
.Y(n_165)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_165),
.Y(n_178)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_126),
.Y(n_166)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_166),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_143),
.A2(n_110),
.B(n_137),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_167),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_SL g197 ( 
.A(n_170),
.B(n_152),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_143),
.A2(n_137),
.B(n_127),
.Y(n_171)
);

HB1xp67_ASAP7_75t_L g190 ( 
.A(n_171),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_172),
.B(n_164),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_175),
.A2(n_179),
.B1(n_164),
.B2(n_150),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_149),
.A2(n_128),
.B1(n_124),
.B2(n_136),
.Y(n_179)
);

NOR3xp33_ASAP7_75t_L g198 ( 
.A(n_180),
.B(n_185),
.C(n_164),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_184),
.B(n_151),
.C(n_158),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_148),
.A2(n_119),
.B(n_131),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_166),
.Y(n_186)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_186),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_149),
.A2(n_135),
.B(n_116),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_188),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_192),
.A2(n_187),
.B1(n_180),
.B2(n_185),
.Y(n_219)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_183),
.Y(n_193)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_193),
.Y(n_210)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_183),
.Y(n_194)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_194),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_195),
.A2(n_198),
.B(n_188),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_196),
.B(n_200),
.C(n_202),
.Y(n_208)
);

XNOR2x1_ASAP7_75t_L g221 ( 
.A(n_197),
.B(n_190),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_168),
.B(n_145),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_199),
.B(n_203),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_168),
.B(n_161),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_171),
.B(n_165),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_187),
.A2(n_141),
.B1(n_153),
.B2(n_155),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_186),
.Y(n_204)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_204),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_184),
.B(n_154),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_205),
.B(n_167),
.C(n_182),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_177),
.B(n_147),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_206),
.B(n_173),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_207),
.B(n_213),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_209),
.B(n_214),
.C(n_216),
.Y(n_231)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_191),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_197),
.B(n_196),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_200),
.B(n_181),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_215),
.B(n_220),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_202),
.B(n_169),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_205),
.B(n_169),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_217),
.B(n_221),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_219),
.A2(n_203),
.B1(n_175),
.B2(n_179),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_218),
.A2(n_192),
.B1(n_201),
.B2(n_189),
.Y(n_222)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_222),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_219),
.A2(n_201),
.B1(n_176),
.B2(n_172),
.Y(n_224)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_224),
.Y(n_240)
);

OA21x2_ASAP7_75t_SL g226 ( 
.A1(n_221),
.A2(n_178),
.B(n_182),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_226),
.A2(n_228),
.B1(n_208),
.B2(n_212),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_220),
.A2(n_178),
.B(n_156),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_227),
.B(n_232),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_210),
.B(n_163),
.Y(n_230)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_230),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_209),
.A2(n_174),
.B(n_164),
.Y(n_232)
);

BUFx12_ASAP7_75t_L g233 ( 
.A(n_216),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_233),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_231),
.B(n_214),
.C(n_208),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_234),
.B(n_238),
.C(n_231),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_225),
.B(n_174),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_236),
.B(n_217),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_235),
.A2(n_229),
.B(n_237),
.Y(n_242)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_242),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_241),
.A2(n_230),
.B1(n_227),
.B2(n_211),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_243),
.B(n_239),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_244),
.B(n_246),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_245),
.B(n_247),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_240),
.B(n_241),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_234),
.B(n_223),
.C(n_232),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_251),
.B(n_239),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_250),
.B(n_244),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_252),
.B(n_253),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_248),
.B(n_240),
.C(n_223),
.Y(n_254)
);

AOI322xp5_ASAP7_75t_L g256 ( 
.A1(n_254),
.A2(n_249),
.A3(n_233),
.B1(n_224),
.B2(n_222),
.C1(n_116),
.C2(n_111),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_256),
.B(n_170),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_257),
.B(n_255),
.C(n_233),
.Y(n_258)
);

AOI321xp33_ASAP7_75t_SL g259 ( 
.A1(n_258),
.A2(n_121),
.A3(n_10),
.B1(n_12),
.B2(n_13),
.C(n_14),
.Y(n_259)
);

BUFx24_ASAP7_75t_SL g260 ( 
.A(n_259),
.Y(n_260)
);


endmodule