module real_jpeg_26388_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_148;
wire n_373;
wire n_375;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_0),
.B(n_39),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_0),
.B(n_28),
.Y(n_52)
);

CKINVDCx14_ASAP7_75t_R g237 ( 
.A(n_0),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_0),
.B(n_87),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_0),
.B(n_94),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_0),
.B(n_61),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_0),
.B(n_50),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_0),
.B(n_35),
.Y(n_369)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_2),
.B(n_58),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_2),
.B(n_159),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_2),
.B(n_87),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_2),
.B(n_94),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_2),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_2),
.B(n_50),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_2),
.B(n_35),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_3),
.B(n_119),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_3),
.B(n_87),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_3),
.B(n_94),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_3),
.B(n_61),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_3),
.B(n_50),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_3),
.B(n_35),
.Y(n_271)
);

CKINVDCx14_ASAP7_75t_R g283 ( 
.A(n_3),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_3),
.B(n_39),
.Y(n_328)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_4),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g95 ( 
.A(n_5),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_6),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_7),
.B(n_150),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_7),
.B(n_87),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_7),
.B(n_94),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_7),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_7),
.B(n_35),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_7),
.B(n_28),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_7),
.B(n_39),
.Y(n_355)
);

INVx8_ASAP7_75t_SL g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_9),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_10),
.B(n_87),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_10),
.B(n_17),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_10),
.B(n_94),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_10),
.B(n_61),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_10),
.B(n_50),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_10),
.B(n_35),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_10),
.B(n_28),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_10),
.B(n_58),
.Y(n_256)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_12),
.B(n_83),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_12),
.B(n_87),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_12),
.B(n_94),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_12),
.B(n_61),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_12),
.B(n_50),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_12),
.B(n_35),
.Y(n_223)
);

CKINVDCx14_ASAP7_75t_R g252 ( 
.A(n_12),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_12),
.B(n_58),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_13),
.B(n_24),
.Y(n_23)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_13),
.B(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_13),
.B(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_13),
.B(n_94),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_14),
.B(n_39),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_14),
.B(n_159),
.Y(n_194)
);

CKINVDCx14_ASAP7_75t_R g234 ( 
.A(n_14),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_14),
.B(n_94),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_14),
.B(n_61),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_14),
.B(n_50),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_14),
.B(n_35),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_14),
.B(n_28),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_15),
.B(n_61),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_15),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_15),
.B(n_87),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_15),
.B(n_50),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_15),
.B(n_35),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_15),
.B(n_28),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_16),
.B(n_94),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_16),
.B(n_87),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_16),
.B(n_109),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_16),
.B(n_61),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_16),
.B(n_50),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_16),
.B(n_35),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_16),
.B(n_28),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_16),
.B(n_39),
.Y(n_238)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_17),
.Y(n_84)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_17),
.Y(n_110)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_17),
.Y(n_120)
);

INVx6_ASAP7_75t_L g151 ( 
.A(n_17),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_66),
.Y(n_18)
);

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_21),
.B1(n_42),
.B2(n_43),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_21),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_33),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_26),
.B1(n_31),
.B2(n_32),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_23),
.Y(n_31)
);

INVx11_ASAP7_75t_L g199 ( 
.A(n_24),
.Y(n_199)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_25),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_26),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_SL g33 ( 
.A(n_26),
.B(n_34),
.C(n_38),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_26),
.A2(n_32),
.B1(n_34),
.B2(n_51),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_27),
.B(n_30),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_27),
.B(n_252),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_27),
.B(n_283),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_27),
.B(n_247),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g27 ( 
.A(n_28),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_30),
.B(n_60),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_30),
.B(n_110),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_30),
.B(n_235),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_34),
.A2(n_48),
.B1(n_49),
.B2(n_51),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_34),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

XNOR2xp5_ASAP7_75t_L g64 ( 
.A(n_38),
.B(n_65),
.Y(n_64)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_43),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_63),
.C(n_64),
.Y(n_43)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_44),
.B(n_386),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_54),
.C(n_55),
.Y(n_44)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_45),
.B(n_384),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_46),
.A2(n_47),
.B1(n_52),
.B2(n_53),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_47),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_L g374 ( 
.A1(n_48),
.A2(n_49),
.B1(n_59),
.B2(n_342),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_49),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_49),
.B(n_56),
.C(n_59),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_49),
.B(n_51),
.C(n_53),
.Y(n_63)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_50),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_52),
.Y(n_53)
);

XNOR2xp5_ASAP7_75t_L g384 ( 
.A(n_54),
.B(n_55),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_56),
.A2(n_57),
.B1(n_374),
.B2(n_375),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_57),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g341 ( 
.A1(n_59),
.A2(n_314),
.B1(n_315),
.B2(n_342),
.Y(n_341)
);

CKINVDCx16_ASAP7_75t_R g342 ( 
.A(n_59),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_SL g372 ( 
.A(n_59),
.B(n_315),
.C(n_340),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_60),
.B(n_213),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_60),
.B(n_247),
.Y(n_246)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

XNOR2xp5_ASAP7_75t_L g386 ( 
.A(n_63),
.B(n_64),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_385),
.C(n_387),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_379),
.C(n_380),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_361),
.C(n_362),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_332),
.C(n_333),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_307),
.C(n_308),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_275),
.C(n_276),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_240),
.C(n_241),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_205),
.C(n_206),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_174),
.C(n_175),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_153),
.C(n_154),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_133),
.C(n_134),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_111),
.C(n_112),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_96),
.C(n_101),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_80),
.A2(n_81),
.B1(n_90),
.B2(n_91),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_80),
.B(n_92),
.C(n_93),
.Y(n_111)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_82),
.A2(n_85),
.B1(n_86),
.B2(n_89),
.Y(n_81)
);

CKINVDCx14_ASAP7_75t_R g89 ( 
.A(n_82),
.Y(n_89)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx8_ASAP7_75t_L g159 ( 
.A(n_84),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_85),
.B(n_89),
.Y(n_115)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx4_ASAP7_75t_L g235 ( 
.A(n_87),
.Y(n_235)
);

BUFx12f_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_SL g91 ( 
.A(n_92),
.B(n_93),
.Y(n_91)
);

INVx13_ASAP7_75t_L g105 ( 
.A(n_94),
.Y(n_105)
);

BUFx24_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_97),
.B(n_99),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_97),
.A2(n_98),
.B1(n_99),
.B2(n_100),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_98),
.Y(n_97)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_103),
.C(n_106),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_105),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_104),
.B(n_199),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_108),
.Y(n_106)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_110),
.B(n_237),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_124),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_114),
.A2(n_115),
.B1(n_116),
.B2(n_117),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_114),
.B(n_117),
.C(n_124),
.Y(n_133)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_118),
.A2(n_121),
.B1(n_122),
.B2(n_123),
.Y(n_117)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_118),
.Y(n_123)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_121),
.B(n_123),
.Y(n_143)
);

CKINVDCx14_ASAP7_75t_R g121 ( 
.A(n_122),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_125),
.A2(n_126),
.B1(n_127),
.B2(n_132),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_125),
.Y(n_132)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_128),
.A2(n_129),
.B1(n_130),
.B2(n_131),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_128),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_129),
.B(n_131),
.C(n_132),
.Y(n_136)
);

CKINVDCx14_ASAP7_75t_R g129 ( 
.A(n_130),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_SL g134 ( 
.A(n_135),
.B(n_142),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_137),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_136),
.B(n_137),
.C(n_142),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_139),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_138),
.B(n_140),
.C(n_141),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_141),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_SL g142 ( 
.A(n_143),
.B(n_144),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_143),
.B(n_145),
.C(n_146),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_146),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_147),
.A2(n_148),
.B1(n_149),
.B2(n_152),
.Y(n_146)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_147),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_148),
.B(n_152),
.Y(n_172)
);

CKINVDCx14_ASAP7_75t_R g148 ( 
.A(n_149),
.Y(n_148)
);

INVx5_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_168),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_155),
.B(n_169),
.C(n_173),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_SL g155 ( 
.A(n_156),
.B(n_164),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_163),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_157),
.B(n_163),
.C(n_164),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_158),
.A2(n_160),
.B1(n_161),
.B2(n_162),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_158),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_160),
.B(n_162),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_161),
.Y(n_160)
);

BUFx24_ASAP7_75t_SL g392 ( 
.A(n_164),
.Y(n_392)
);

FAx1_ASAP7_75t_SL g164 ( 
.A(n_165),
.B(n_166),
.CI(n_167),
.CON(n_164),
.SN(n_164)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_165),
.B(n_166),
.C(n_167),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_173),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_169),
.Y(n_191)
);

FAx1_ASAP7_75t_SL g169 ( 
.A(n_170),
.B(n_171),
.CI(n_172),
.CON(n_169),
.SN(n_169)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_190),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_178),
.B1(n_179),
.B2(n_180),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_178),
.B(n_179),
.C(n_190),
.Y(n_205)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_SL g180 ( 
.A(n_181),
.B(n_185),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_181),
.B(n_186),
.C(n_189),
.Y(n_209)
);

BUFx24_ASAP7_75t_SL g389 ( 
.A(n_181),
.Y(n_389)
);

FAx1_ASAP7_75t_SL g181 ( 
.A(n_182),
.B(n_183),
.CI(n_184),
.CON(n_181),
.SN(n_181)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_182),
.B(n_183),
.C(n_184),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_186),
.A2(n_187),
.B1(n_188),
.B2(n_189),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_189),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_SL g190 ( 
.A(n_191),
.B(n_192),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_191),
.B(n_197),
.C(n_203),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_193),
.A2(n_197),
.B1(n_203),
.B2(n_204),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_193),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_194),
.A2(n_195),
.B(n_196),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_194),
.B(n_195),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_196),
.B(n_230),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_196),
.B(n_230),
.C(n_231),
.Y(n_265)
);

CKINVDCx16_ASAP7_75t_R g204 ( 
.A(n_197),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_200),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_198),
.B(n_201),
.C(n_202),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_202),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_207),
.A2(n_208),
.B1(n_226),
.B2(n_239),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_207),
.B(n_227),
.C(n_228),
.Y(n_240)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_SL g208 ( 
.A(n_209),
.B(n_210),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_209),
.B(n_211),
.C(n_219),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_219),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_214),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_212),
.B(n_215),
.C(n_218),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_213),
.B(n_250),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_215),
.A2(n_216),
.B1(n_217),
.B2(n_218),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_216),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_217),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_225),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_221),
.A2(n_222),
.B1(n_223),
.B2(n_224),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_221),
.B(n_224),
.C(n_225),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_222),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_223),
.Y(n_224)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_226),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_SL g226 ( 
.A(n_227),
.B(n_228),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_231),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_SL g231 ( 
.A(n_232),
.B(n_238),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_236),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_233),
.B(n_236),
.C(n_238),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_235),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_242),
.A2(n_243),
.B1(n_273),
.B2(n_274),
.Y(n_241)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_242),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_243),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_SL g243 ( 
.A(n_244),
.B(n_264),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_244),
.B(n_264),
.C(n_273),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_253),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_245),
.B(n_254),
.C(n_255),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_248),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_246),
.B(n_249),
.C(n_251),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_251),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_255),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_256),
.A2(n_257),
.B1(n_258),
.B2(n_263),
.Y(n_255)
);

CKINVDCx16_ASAP7_75t_R g263 ( 
.A(n_256),
.Y(n_263)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_259),
.A2(n_260),
.B1(n_261),
.B2(n_262),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_259),
.A2(n_260),
.B1(n_285),
.B2(n_286),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_259),
.B(n_262),
.C(n_263),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_259),
.B(n_282),
.C(n_285),
.Y(n_330)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_262),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_266),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_265),
.B(n_267),
.C(n_268),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_268),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_272),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_271),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_270),
.B(n_271),
.C(n_272),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_278),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_277),
.B(n_279),
.C(n_306),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_279),
.A2(n_280),
.B1(n_293),
.B2(n_306),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_287),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_281),
.B(n_288),
.C(n_289),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_SL g281 ( 
.A(n_282),
.B(n_284),
.Y(n_281)
);

CKINVDCx14_ASAP7_75t_R g286 ( 
.A(n_285),
.Y(n_286)
);

AOI22xp33_ASAP7_75t_L g313 ( 
.A1(n_285),
.A2(n_286),
.B1(n_314),
.B2(n_315),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_SL g346 ( 
.A(n_285),
.B(n_312),
.C(n_315),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_289),
.Y(n_287)
);

BUFx24_ASAP7_75t_SL g388 ( 
.A(n_289),
.Y(n_388)
);

FAx1_ASAP7_75t_SL g289 ( 
.A(n_290),
.B(n_291),
.CI(n_292),
.CON(n_289),
.SN(n_289)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_290),
.B(n_291),
.C(n_292),
.Y(n_317)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_293),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_295),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_294),
.B(n_296),
.C(n_297),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_297),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_298),
.A2(n_299),
.B1(n_300),
.B2(n_305),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_298),
.B(n_301),
.C(n_303),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_299),
.Y(n_298)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_300),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_301),
.A2(n_302),
.B1(n_303),
.B2(n_304),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_301),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_302),
.A2(n_303),
.B1(n_328),
.B2(n_329),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_303),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_303),
.B(n_329),
.C(n_330),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_331),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_322),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_310),
.B(n_322),
.C(n_331),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_316),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_311),
.B(n_317),
.C(n_318),
.Y(n_349)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_313),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_315),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_318),
.Y(n_316)
);

BUFx24_ASAP7_75t_SL g391 ( 
.A(n_318),
.Y(n_391)
);

FAx1_ASAP7_75t_SL g318 ( 
.A(n_319),
.B(n_320),
.CI(n_321),
.CON(n_318),
.SN(n_318)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_319),
.B(n_320),
.C(n_321),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_SL g322 ( 
.A(n_323),
.B(n_324),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_323),
.B(n_325),
.C(n_326),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_326),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_330),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_328),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_334),
.B(n_335),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_334),
.B(n_336),
.C(n_348),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_336),
.A2(n_337),
.B1(n_347),
.B2(n_348),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_338),
.A2(n_339),
.B1(n_343),
.B2(n_344),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_338),
.B(n_345),
.C(n_346),
.Y(n_364)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_340),
.B(n_341),
.Y(n_339)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

XOR2xp5_ASAP7_75t_L g344 ( 
.A(n_345),
.B(n_346),
.Y(n_344)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_349),
.B(n_350),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_349),
.B(n_351),
.C(n_354),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_351),
.A2(n_352),
.B1(n_353),
.B2(n_354),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

CKINVDCx16_ASAP7_75t_R g353 ( 
.A(n_354),
.Y(n_353)
);

XOR2xp5_ASAP7_75t_L g354 ( 
.A(n_355),
.B(n_356),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_355),
.B(n_357),
.C(n_360),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_357),
.A2(n_358),
.B1(n_359),
.B2(n_360),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_358),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_359),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_363),
.A2(n_376),
.B1(n_377),
.B2(n_378),
.Y(n_362)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_363),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_SL g363 ( 
.A(n_364),
.B(n_365),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_364),
.B(n_365),
.C(n_378),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_366),
.B(n_371),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_366),
.B(n_372),
.C(n_373),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_367),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_367),
.B(n_383),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_367),
.B(n_381),
.C(n_383),
.Y(n_387)
);

FAx1_ASAP7_75t_SL g367 ( 
.A(n_368),
.B(n_369),
.CI(n_370),
.CON(n_367),
.SN(n_367)
);

XNOR2xp5_ASAP7_75t_L g371 ( 
.A(n_372),
.B(n_373),
.Y(n_371)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_374),
.Y(n_375)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_376),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_381),
.B(n_382),
.Y(n_380)
);


endmodule