module fake_jpeg_29159_n_9 (n_3, n_2, n_1, n_0, n_4, n_9);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;

output n_9;

wire n_8;
wire n_6;
wire n_5;
wire n_7;

NAND2xp5_ASAP7_75t_SL g5 ( 
.A(n_4),
.B(n_1),
.Y(n_5)
);

INVx1_ASAP7_75t_L g6 ( 
.A(n_2),
.Y(n_6)
);

MAJIxp5_ASAP7_75t_L g7 ( 
.A(n_5),
.B(n_0),
.C(n_1),
.Y(n_7)
);

FAx1_ASAP7_75t_SL g8 ( 
.A(n_7),
.B(n_0),
.CI(n_2),
.CON(n_8),
.SN(n_8)
);

AOI332xp33_ASAP7_75t_L g9 ( 
.A1(n_8),
.A2(n_3),
.A3(n_6),
.B1(n_5),
.B2(n_7),
.B3(n_2),
.C1(n_0),
.C2(n_1),
.Y(n_9)
);


endmodule