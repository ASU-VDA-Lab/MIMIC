module real_jpeg_22437_n_18 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_329, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_329;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_215;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_0),
.A2(n_31),
.B1(n_32),
.B2(n_98),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_0),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_0),
.A2(n_25),
.B1(n_26),
.B2(n_98),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_0),
.A2(n_47),
.B1(n_48),
.B2(n_98),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_0),
.A2(n_42),
.B1(n_43),
.B2(n_98),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_1),
.A2(n_42),
.B1(n_43),
.B2(n_88),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_1),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_1),
.A2(n_47),
.B1(n_48),
.B2(n_88),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_1),
.A2(n_31),
.B1(n_32),
.B2(n_88),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_1),
.A2(n_25),
.B1(n_26),
.B2(n_88),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_2),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_2),
.B(n_30),
.Y(n_132)
);

AOI21xp33_ASAP7_75t_L g153 ( 
.A1(n_2),
.A2(n_44),
.B(n_47),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_2),
.A2(n_42),
.B1(n_43),
.B2(n_103),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_2),
.A2(n_82),
.B1(n_83),
.B2(n_161),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_2),
.B(n_58),
.Y(n_175)
);

AOI21xp33_ASAP7_75t_L g192 ( 
.A1(n_2),
.A2(n_32),
.B(n_193),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g23 ( 
.A1(n_3),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_3),
.A2(n_24),
.B1(n_31),
.B2(n_32),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_3),
.A2(n_24),
.B1(n_47),
.B2(n_48),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_3),
.A2(n_24),
.B1(n_42),
.B2(n_43),
.Y(n_265)
);

OAI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_4),
.A2(n_25),
.B1(n_26),
.B2(n_105),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_4),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_4),
.A2(n_31),
.B1(n_32),
.B2(n_105),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_4),
.A2(n_42),
.B1(n_43),
.B2(n_105),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_4),
.A2(n_47),
.B1(n_48),
.B2(n_105),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_5),
.A2(n_25),
.B1(n_26),
.B2(n_66),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_5),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_5),
.A2(n_47),
.B1(n_48),
.B2(n_66),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g232 ( 
.A1(n_5),
.A2(n_42),
.B1(n_43),
.B2(n_66),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_SL g278 ( 
.A1(n_5),
.A2(n_31),
.B1(n_32),
.B2(n_66),
.Y(n_278)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_6),
.A2(n_31),
.B1(n_32),
.B2(n_100),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_6),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_6),
.A2(n_47),
.B1(n_48),
.B2(n_100),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_6),
.A2(n_42),
.B1(n_43),
.B2(n_100),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g239 ( 
.A1(n_6),
.A2(n_25),
.B1(n_26),
.B2(n_100),
.Y(n_239)
);

BUFx16f_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_8),
.A2(n_25),
.B1(n_26),
.B2(n_63),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_8),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_8),
.A2(n_42),
.B1(n_43),
.B2(n_63),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_8),
.A2(n_47),
.B1(n_48),
.B2(n_63),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_8),
.A2(n_31),
.B1(n_32),
.B2(n_63),
.Y(n_259)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_9),
.Y(n_83)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_9),
.Y(n_120)
);

BUFx12_ASAP7_75t_L g47 ( 
.A(n_10),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_11),
.A2(n_25),
.B1(n_26),
.B2(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_11),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_11),
.A2(n_35),
.B1(n_42),
.B2(n_43),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_11),
.A2(n_31),
.B1(n_32),
.B2(n_35),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_11),
.A2(n_35),
.B1(n_47),
.B2(n_48),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_12),
.A2(n_42),
.B1(n_43),
.B2(n_94),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_12),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_12),
.A2(n_31),
.B1(n_32),
.B2(n_94),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g180 ( 
.A1(n_12),
.A2(n_47),
.B1(n_48),
.B2(n_94),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_12),
.A2(n_25),
.B1(n_26),
.B2(n_94),
.Y(n_255)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx13_ASAP7_75t_L g54 ( 
.A(n_14),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_14),
.A2(n_42),
.B1(n_43),
.B2(n_54),
.Y(n_56)
);

OAI32xp33_ASAP7_75t_L g187 ( 
.A1(n_14),
.A2(n_32),
.A3(n_43),
.B1(n_188),
.B2(n_189),
.Y(n_187)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

BUFx3_ASAP7_75t_SL g43 ( 
.A(n_17),
.Y(n_43)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_72),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_71),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_36),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_22),
.B(n_36),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_27),
.B1(n_30),
.B2(n_34),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_23),
.A2(n_27),
.B1(n_30),
.B2(n_70),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_25),
.Y(n_26)
);

O2A1O1Ixp33_ASAP7_75t_L g27 ( 
.A1(n_25),
.A2(n_28),
.B(n_29),
.C(n_30),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_25),
.B(n_28),
.Y(n_29)
);

HAxp5_ASAP7_75t_SL g102 ( 
.A(n_25),
.B(n_103),
.CON(n_102),
.SN(n_102)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_27),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_27),
.A2(n_30),
.B1(n_102),
.B2(n_104),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_27),
.A2(n_30),
.B1(n_285),
.B2(n_286),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_28),
.A2(n_31),
.B1(n_32),
.B2(n_33),
.Y(n_30)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_28),
.B(n_32),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_29),
.A2(n_31),
.B1(n_102),
.B2(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_30),
.Y(n_64)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_31),
.Y(n_32)
);

A2O1A1Ixp33_ASAP7_75t_L g53 ( 
.A1(n_31),
.A2(n_54),
.B(n_55),
.C(n_56),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_31),
.B(n_54),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_31),
.B(n_103),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_67),
.C(n_69),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_37),
.A2(n_38),
.B1(n_324),
.B2(n_326),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_38),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_50),
.C(n_59),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g294 ( 
.A1(n_39),
.A2(n_295),
.B1(n_296),
.B2(n_298),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_39),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_39),
.A2(n_50),
.B1(n_298),
.B2(n_311),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_SL g39 ( 
.A1(n_40),
.A2(n_46),
.B(n_49),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_40),
.A2(n_46),
.B1(n_87),
.B2(n_89),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_40),
.A2(n_46),
.B1(n_87),
.B2(n_93),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_40),
.A2(n_46),
.B1(n_156),
.B2(n_157),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_40),
.A2(n_46),
.B1(n_157),
.B2(n_178),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_40),
.A2(n_46),
.B1(n_178),
.B2(n_196),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_40),
.A2(n_46),
.B1(n_93),
.B2(n_196),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_40),
.A2(n_46),
.B1(n_89),
.B2(n_232),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_40),
.A2(n_46),
.B1(n_232),
.B2(n_265),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_40),
.A2(n_46),
.B1(n_49),
.B2(n_265),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_46),
.Y(n_40)
);

OAI22xp33_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_43),
.B1(n_44),
.B2(n_45),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_42),
.B(n_54),
.Y(n_188)
);

INVx2_ASAP7_75t_SL g42 ( 
.A(n_43),
.Y(n_42)
);

A2O1A1Ixp33_ASAP7_75t_L g152 ( 
.A1(n_43),
.A2(n_45),
.B(n_103),
.C(n_153),
.Y(n_152)
);

OA22x2_ASAP7_75t_L g46 ( 
.A1(n_44),
.A2(n_45),
.B1(n_47),
.B2(n_48),
.Y(n_46)
);

CKINVDCx9p33_ASAP7_75t_R g44 ( 
.A(n_45),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_46),
.B(n_103),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g48 ( 
.A(n_47),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_47),
.B(n_83),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_48),
.B(n_166),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_50),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_51),
.A2(n_52),
.B1(n_57),
.B2(n_58),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_51),
.A2(n_52),
.B1(n_58),
.B2(n_297),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_SL g68 ( 
.A1(n_52),
.A2(n_57),
.B(n_58),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_52),
.A2(n_58),
.B1(n_129),
.B2(n_131),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_52),
.A2(n_58),
.B1(n_258),
.B2(n_259),
.Y(n_257)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_53),
.A2(n_56),
.B1(n_97),
.B2(n_99),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_53),
.A2(n_56),
.B1(n_99),
.B2(n_113),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_53),
.A2(n_56),
.B1(n_130),
.B2(n_192),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_53),
.A2(n_56),
.B1(n_113),
.B2(n_241),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_53),
.A2(n_56),
.B1(n_277),
.B2(n_278),
.Y(n_276)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_56),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_59),
.A2(n_60),
.B1(n_309),
.B2(n_310),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_60),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_61),
.A2(n_62),
.B1(n_64),
.B2(n_65),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_61),
.A2(n_64),
.B1(n_110),
.B2(n_111),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_61),
.A2(n_64),
.B1(n_111),
.B2(n_239),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_61),
.A2(n_64),
.B1(n_239),
.B2(n_255),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_61),
.A2(n_62),
.B1(n_64),
.B2(n_300),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_65),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_67),
.A2(n_68),
.B1(n_69),
.B2(n_325),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_68),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_69),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_321),
.B(n_327),
.Y(n_72)
);

OAI321xp33_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_290),
.A3(n_313),
.B1(n_319),
.B2(n_320),
.C(n_329),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_269),
.B(n_289),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_SL g75 ( 
.A1(n_76),
.A2(n_245),
.B(n_268),
.Y(n_75)
);

O2A1O1Ixp33_ASAP7_75t_SL g76 ( 
.A1(n_77),
.A2(n_136),
.B(n_221),
.C(n_244),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_121),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_78),
.B(n_121),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_106),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_90),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_80),
.B(n_90),
.C(n_106),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_86),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_81),
.B(n_86),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_83),
.B1(n_84),
.B2(n_85),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_82),
.A2(n_84),
.B1(n_119),
.B2(n_120),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_82),
.A2(n_119),
.B1(n_120),
.B2(n_135),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_82),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_82),
.A2(n_146),
.B1(n_161),
.B2(n_162),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_82),
.A2(n_83),
.B1(n_149),
.B2(n_180),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_82),
.A2(n_135),
.B1(n_162),
.B2(n_180),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_82),
.A2(n_85),
.B1(n_162),
.B2(n_230),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_82),
.A2(n_162),
.B(n_230),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_83),
.B(n_103),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_95),
.C(n_101),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_91),
.A2(n_92),
.B1(n_95),
.B2(n_96),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_96),
.Y(n_95)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_97),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_SL g122 ( 
.A(n_101),
.B(n_123),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_104),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_SL g106 ( 
.A(n_107),
.B(n_115),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_108),
.A2(n_109),
.B1(n_112),
.B2(n_114),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_108),
.B(n_114),
.C(n_115),
.Y(n_224)
);

CKINVDCx14_ASAP7_75t_R g108 ( 
.A(n_109),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_112),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_118),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_116),
.B(n_118),
.Y(n_125)
);

INVx5_ASAP7_75t_L g147 ( 
.A(n_120),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_124),
.C(n_126),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_122),
.B(n_218),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_124),
.A2(n_125),
.B1(n_126),
.B2(n_127),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_125),
.Y(n_124)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_132),
.C(n_133),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_128),
.B(n_206),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_132),
.A2(n_133),
.B1(n_134),
.B2(n_207),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_132),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_134),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_137),
.B(n_220),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_138),
.A2(n_215),
.B(n_219),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_139),
.A2(n_201),
.B(n_214),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_140),
.A2(n_182),
.B(n_200),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_141),
.A2(n_170),
.B(n_181),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_142),
.A2(n_158),
.B(n_169),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_150),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_143),
.B(n_150),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_145),
.B1(n_147),
.B2(n_148),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_147),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_149),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_152),
.B1(n_154),
.B2(n_155),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_152),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_152),
.B(n_154),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_155),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_159),
.A2(n_164),
.B(n_168),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_163),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_160),
.B(n_163),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_167),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_172),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_171),
.B(n_172),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_179),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_174),
.A2(n_175),
.B1(n_176),
.B2(n_177),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_174),
.B(n_177),
.C(n_179),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_175),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_177),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_184),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_183),
.B(n_184),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_185),
.A2(n_190),
.B1(n_198),
.B2(n_199),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_185),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_187),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_186),
.B(n_187),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_189),
.Y(n_193)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_190),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_191),
.A2(n_194),
.B1(n_195),
.B2(n_197),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_191),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_194),
.B(n_197),
.C(n_198),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_195),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_203),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_202),
.B(n_203),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_204),
.A2(n_205),
.B1(n_208),
.B2(n_209),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_204),
.B(n_211),
.C(n_212),
.Y(n_216)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_210),
.A2(n_211),
.B1(n_212),
.B2(n_213),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_210),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_211),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_217),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_216),
.B(n_217),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_223),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_222),
.B(n_223),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_224),
.A2(n_225),
.B1(n_226),
.B2(n_243),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g243 ( 
.A(n_224),
.Y(n_243)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_227),
.A2(n_228),
.B1(n_233),
.B2(n_234),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_227),
.B(n_234),
.C(n_243),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_228),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_231),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_229),
.B(n_231),
.Y(n_251)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_236),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_235),
.B(n_237),
.C(n_242),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_237),
.A2(n_238),
.B1(n_240),
.B2(n_242),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_238),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_240),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_241),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_247),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_246),
.B(n_247),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_267),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_249),
.A2(n_250),
.B1(n_260),
.B2(n_261),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_249),
.B(n_261),
.C(n_267),
.Y(n_270)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_252),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_251),
.B(n_253),
.C(n_257),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_253),
.A2(n_254),
.B1(n_256),
.B2(n_257),
.Y(n_252)
);

CKINVDCx16_ASAP7_75t_R g253 ( 
.A(n_254),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_255),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_257),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_259),
.Y(n_277)
);

CKINVDCx16_ASAP7_75t_R g260 ( 
.A(n_261),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_262),
.A2(n_263),
.B1(n_264),
.B2(n_266),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_262),
.A2(n_263),
.B1(n_283),
.B2(n_284),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_263),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_263),
.B(n_264),
.Y(n_281)
);

AOI21xp33_ASAP7_75t_L g304 ( 
.A1(n_263),
.A2(n_281),
.B(n_284),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_264),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_271),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_270),
.B(n_271),
.Y(n_289)
);

AOI22xp33_ASAP7_75t_SL g271 ( 
.A1(n_272),
.A2(n_273),
.B1(n_287),
.B2(n_288),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_280),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_274),
.B(n_280),
.C(n_288),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_275),
.A2(n_276),
.B(n_279),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_275),
.B(n_276),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_278),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_279),
.B(n_292),
.C(n_303),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_279),
.A2(n_292),
.B1(n_293),
.B2(n_318),
.Y(n_317)
);

CKINVDCx14_ASAP7_75t_R g318 ( 
.A(n_279),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_282),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_284),
.Y(n_283)
);

CKINVDCx16_ASAP7_75t_R g300 ( 
.A(n_286),
.Y(n_300)
);

CKINVDCx16_ASAP7_75t_R g288 ( 
.A(n_287),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_305),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_291),
.B(n_305),
.Y(n_320)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_294),
.A2(n_299),
.B1(n_301),
.B2(n_302),
.Y(n_293)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_294),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_296),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_296),
.B(n_298),
.C(n_299),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_299),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_299),
.A2(n_302),
.B1(n_307),
.B2(n_308),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_299),
.B(n_307),
.C(n_312),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_303),
.A2(n_304),
.B1(n_316),
.B2(n_317),
.Y(n_315)
);

CKINVDCx14_ASAP7_75t_R g303 ( 
.A(n_304),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_312),
.Y(n_305)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

CKINVDCx16_ASAP7_75t_R g309 ( 
.A(n_310),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_315),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_314),
.B(n_315),
.Y(n_319)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_322),
.B(n_323),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_322),
.B(n_323),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_324),
.Y(n_326)
);


endmodule