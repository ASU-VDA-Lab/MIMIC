module fake_aes_2489_n_652 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_71, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_652);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_71;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_652;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_73;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_72;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_260;
wire n_78;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_363;
wire n_409;
wire n_315;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_75;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_74;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g72 ( .A(n_0), .Y(n_72) );
INVx1_ASAP7_75t_L g73 ( .A(n_36), .Y(n_73) );
INVxp67_ASAP7_75t_L g74 ( .A(n_15), .Y(n_74) );
INVx1_ASAP7_75t_L g75 ( .A(n_21), .Y(n_75) );
INVxp67_ASAP7_75t_L g76 ( .A(n_66), .Y(n_76) );
HB1xp67_ASAP7_75t_L g77 ( .A(n_20), .Y(n_77) );
INVx4_ASAP7_75t_R g78 ( .A(n_31), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_58), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_60), .Y(n_80) );
INVxp67_ASAP7_75t_L g81 ( .A(n_24), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_25), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_15), .Y(n_83) );
CKINVDCx20_ASAP7_75t_R g84 ( .A(n_64), .Y(n_84) );
INVx2_ASAP7_75t_L g85 ( .A(n_4), .Y(n_85) );
INVx2_ASAP7_75t_L g86 ( .A(n_71), .Y(n_86) );
CKINVDCx5p33_ASAP7_75t_R g87 ( .A(n_8), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_5), .Y(n_88) );
INVxp33_ASAP7_75t_SL g89 ( .A(n_42), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_1), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_44), .Y(n_91) );
CKINVDCx20_ASAP7_75t_R g92 ( .A(n_21), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_54), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_48), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_19), .Y(n_95) );
CKINVDCx5p33_ASAP7_75t_R g96 ( .A(n_49), .Y(n_96) );
INVx1_ASAP7_75t_SL g97 ( .A(n_50), .Y(n_97) );
INVxp33_ASAP7_75t_SL g98 ( .A(n_55), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_39), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_41), .Y(n_100) );
BUFx3_ASAP7_75t_L g101 ( .A(n_35), .Y(n_101) );
CKINVDCx20_ASAP7_75t_R g102 ( .A(n_16), .Y(n_102) );
CKINVDCx5p33_ASAP7_75t_R g103 ( .A(n_11), .Y(n_103) );
NOR2xp67_ASAP7_75t_L g104 ( .A(n_30), .B(n_7), .Y(n_104) );
CKINVDCx20_ASAP7_75t_R g105 ( .A(n_68), .Y(n_105) );
INVxp67_ASAP7_75t_SL g106 ( .A(n_16), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_1), .Y(n_107) );
CKINVDCx5p33_ASAP7_75t_R g108 ( .A(n_8), .Y(n_108) );
INVxp67_ASAP7_75t_SL g109 ( .A(n_40), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_37), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_59), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_47), .Y(n_112) );
CKINVDCx16_ASAP7_75t_R g113 ( .A(n_51), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_9), .Y(n_114) );
CKINVDCx5p33_ASAP7_75t_R g115 ( .A(n_14), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_12), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_57), .Y(n_117) );
CKINVDCx16_ASAP7_75t_R g118 ( .A(n_13), .Y(n_118) );
INVxp33_ASAP7_75t_SL g119 ( .A(n_38), .Y(n_119) );
NOR2xp33_ASAP7_75t_R g120 ( .A(n_113), .B(n_29), .Y(n_120) );
CKINVDCx5p33_ASAP7_75t_R g121 ( .A(n_84), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_73), .Y(n_122) );
CKINVDCx20_ASAP7_75t_R g123 ( .A(n_118), .Y(n_123) );
BUFx3_ASAP7_75t_L g124 ( .A(n_101), .Y(n_124) );
AND2x6_ASAP7_75t_L g125 ( .A(n_101), .B(n_28), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_73), .Y(n_126) );
CKINVDCx5p33_ASAP7_75t_R g127 ( .A(n_105), .Y(n_127) );
CKINVDCx5p33_ASAP7_75t_R g128 ( .A(n_87), .Y(n_128) );
BUFx6f_ASAP7_75t_L g129 ( .A(n_86), .Y(n_129) );
INVx3_ASAP7_75t_L g130 ( .A(n_85), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_79), .Y(n_131) );
NAND2xp33_ASAP7_75t_R g132 ( .A(n_119), .B(n_32), .Y(n_132) );
CKINVDCx5p33_ASAP7_75t_R g133 ( .A(n_103), .Y(n_133) );
CKINVDCx5p33_ASAP7_75t_R g134 ( .A(n_108), .Y(n_134) );
CKINVDCx5p33_ASAP7_75t_R g135 ( .A(n_115), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_79), .Y(n_136) );
CKINVDCx5p33_ASAP7_75t_R g137 ( .A(n_89), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_80), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_80), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_77), .B(n_0), .Y(n_140) );
CKINVDCx20_ASAP7_75t_R g141 ( .A(n_92), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_74), .B(n_86), .Y(n_142) );
INVx3_ASAP7_75t_L g143 ( .A(n_85), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g144 ( .A(n_82), .B(n_2), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_82), .Y(n_145) );
HB1xp67_ASAP7_75t_L g146 ( .A(n_72), .Y(n_146) );
BUFx6f_ASAP7_75t_L g147 ( .A(n_91), .Y(n_147) );
CKINVDCx5p33_ASAP7_75t_R g148 ( .A(n_98), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_91), .Y(n_149) );
INVx3_ASAP7_75t_L g150 ( .A(n_93), .Y(n_150) );
INVx3_ASAP7_75t_L g151 ( .A(n_93), .Y(n_151) );
CKINVDCx5p33_ASAP7_75t_R g152 ( .A(n_96), .Y(n_152) );
HB1xp67_ASAP7_75t_L g153 ( .A(n_72), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_94), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_94), .Y(n_155) );
BUFx6f_ASAP7_75t_L g156 ( .A(n_99), .Y(n_156) );
CKINVDCx5p33_ASAP7_75t_R g157 ( .A(n_102), .Y(n_157) );
AND2x2_ASAP7_75t_L g158 ( .A(n_75), .B(n_2), .Y(n_158) );
BUFx6f_ASAP7_75t_L g159 ( .A(n_117), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_99), .Y(n_160) );
CKINVDCx5p33_ASAP7_75t_R g161 ( .A(n_97), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_147), .Y(n_162) );
NOR2xp33_ASAP7_75t_L g163 ( .A(n_142), .B(n_81), .Y(n_163) );
NOR2xp33_ASAP7_75t_L g164 ( .A(n_137), .B(n_76), .Y(n_164) );
BUFx3_ASAP7_75t_L g165 ( .A(n_124), .Y(n_165) );
AND2x6_ASAP7_75t_L g166 ( .A(n_158), .B(n_117), .Y(n_166) );
BUFx2_ASAP7_75t_L g167 ( .A(n_128), .Y(n_167) );
NOR2xp33_ASAP7_75t_L g168 ( .A(n_148), .B(n_100), .Y(n_168) );
AND2x4_ASAP7_75t_L g169 ( .A(n_146), .B(n_116), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_147), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_147), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_147), .Y(n_172) );
INVx2_ASAP7_75t_L g173 ( .A(n_129), .Y(n_173) );
INVxp67_ASAP7_75t_L g174 ( .A(n_133), .Y(n_174) );
BUFx6f_ASAP7_75t_L g175 ( .A(n_129), .Y(n_175) );
INVx2_ASAP7_75t_L g176 ( .A(n_129), .Y(n_176) );
BUFx6f_ASAP7_75t_L g177 ( .A(n_129), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_147), .Y(n_178) );
BUFx6f_ASAP7_75t_L g179 ( .A(n_129), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_122), .B(n_100), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_147), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_156), .Y(n_182) );
INVx1_ASAP7_75t_L g183 ( .A(n_156), .Y(n_183) );
OAI22xp5_ASAP7_75t_L g184 ( .A1(n_134), .A2(n_116), .B1(n_114), .B2(n_83), .Y(n_184) );
INVx4_ASAP7_75t_L g185 ( .A(n_125), .Y(n_185) );
BUFx3_ASAP7_75t_L g186 ( .A(n_124), .Y(n_186) );
INVx1_ASAP7_75t_L g187 ( .A(n_156), .Y(n_187) );
NAND3xp33_ASAP7_75t_L g188 ( .A(n_153), .B(n_114), .C(n_83), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_156), .Y(n_189) );
NOR2xp33_ASAP7_75t_L g190 ( .A(n_152), .B(n_112), .Y(n_190) );
AND2x2_ASAP7_75t_L g191 ( .A(n_122), .B(n_75), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_156), .Y(n_192) );
NOR2xp33_ASAP7_75t_L g193 ( .A(n_135), .B(n_112), .Y(n_193) );
INVx2_ASAP7_75t_L g194 ( .A(n_129), .Y(n_194) );
INVx1_ASAP7_75t_L g195 ( .A(n_156), .Y(n_195) );
INVx1_ASAP7_75t_L g196 ( .A(n_159), .Y(n_196) );
INVxp67_ASAP7_75t_L g197 ( .A(n_161), .Y(n_197) );
INVx1_ASAP7_75t_L g198 ( .A(n_159), .Y(n_198) );
BUFx2_ASAP7_75t_L g199 ( .A(n_120), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_159), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_126), .B(n_111), .Y(n_201) );
INVx2_ASAP7_75t_L g202 ( .A(n_159), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_126), .B(n_111), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_159), .Y(n_204) );
HB1xp67_ASAP7_75t_L g205 ( .A(n_157), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_131), .B(n_110), .Y(n_206) );
AND2x2_ASAP7_75t_L g207 ( .A(n_131), .B(n_88), .Y(n_207) );
A2O1A1Ixp33_ASAP7_75t_L g208 ( .A1(n_136), .A2(n_110), .B(n_107), .C(n_88), .Y(n_208) );
NOR2xp33_ASAP7_75t_L g209 ( .A(n_136), .B(n_109), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_159), .Y(n_210) );
CKINVDCx16_ASAP7_75t_R g211 ( .A(n_123), .Y(n_211) );
INVx2_ASAP7_75t_L g212 ( .A(n_124), .Y(n_212) );
INVx2_ASAP7_75t_L g213 ( .A(n_150), .Y(n_213) );
INVx2_ASAP7_75t_L g214 ( .A(n_150), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_138), .B(n_107), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_138), .B(n_95), .Y(n_216) );
OAI221xp5_ASAP7_75t_L g217 ( .A1(n_140), .A2(n_95), .B1(n_90), .B2(n_106), .C(n_104), .Y(n_217) );
INVx2_ASAP7_75t_L g218 ( .A(n_150), .Y(n_218) );
AND2x4_ASAP7_75t_L g219 ( .A(n_150), .B(n_90), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_151), .Y(n_220) );
OAI22xp5_ASAP7_75t_L g221 ( .A1(n_139), .A2(n_78), .B1(n_4), .B2(n_5), .Y(n_221) );
AND2x2_ASAP7_75t_L g222 ( .A(n_139), .B(n_3), .Y(n_222) );
NOR2xp33_ASAP7_75t_L g223 ( .A(n_145), .B(n_34), .Y(n_223) );
AND2x2_ASAP7_75t_L g224 ( .A(n_169), .B(n_121), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_163), .B(n_160), .Y(n_225) );
NAND2xp33_ASAP7_75t_SL g226 ( .A(n_185), .B(n_127), .Y(n_226) );
BUFx12f_ASAP7_75t_L g227 ( .A(n_167), .Y(n_227) );
AND2x2_ASAP7_75t_L g228 ( .A(n_169), .B(n_158), .Y(n_228) );
NAND2xp5_ASAP7_75t_SL g229 ( .A(n_185), .B(n_169), .Y(n_229) );
HB1xp67_ASAP7_75t_L g230 ( .A(n_221), .Y(n_230) );
BUFx6f_ASAP7_75t_L g231 ( .A(n_185), .Y(n_231) );
HB1xp67_ASAP7_75t_L g232 ( .A(n_166), .Y(n_232) );
NOR2xp33_ASAP7_75t_L g233 ( .A(n_190), .B(n_160), .Y(n_233) );
INVx2_ASAP7_75t_L g234 ( .A(n_213), .Y(n_234) );
INVx3_ASAP7_75t_L g235 ( .A(n_219), .Y(n_235) );
NOR3xp33_ASAP7_75t_SL g236 ( .A(n_211), .B(n_132), .C(n_144), .Y(n_236) );
CKINVDCx8_ASAP7_75t_R g237 ( .A(n_211), .Y(n_237) );
OAI21xp33_ASAP7_75t_SL g238 ( .A1(n_180), .A2(n_155), .B(n_154), .Y(n_238) );
INVx6_ASAP7_75t_L g239 ( .A(n_219), .Y(n_239) );
AND2x2_ASAP7_75t_L g240 ( .A(n_197), .B(n_155), .Y(n_240) );
AND2x4_ASAP7_75t_L g241 ( .A(n_191), .B(n_154), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_166), .B(n_149), .Y(n_242) );
HB1xp67_ASAP7_75t_L g243 ( .A(n_166), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_166), .B(n_149), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_222), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_222), .Y(n_246) );
NAND2xp5_ASAP7_75t_SL g247 ( .A(n_220), .B(n_151), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_166), .B(n_145), .Y(n_248) );
AND2x4_ASAP7_75t_L g249 ( .A(n_191), .B(n_151), .Y(n_249) );
BUFx6f_ASAP7_75t_L g250 ( .A(n_175), .Y(n_250) );
INVx2_ASAP7_75t_SL g251 ( .A(n_166), .Y(n_251) );
BUFx2_ASAP7_75t_L g252 ( .A(n_167), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_166), .B(n_151), .Y(n_253) );
AND2x4_ASAP7_75t_SL g254 ( .A(n_205), .B(n_141), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_219), .Y(n_255) );
INVx6_ASAP7_75t_L g256 ( .A(n_219), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_207), .B(n_125), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_207), .B(n_125), .Y(n_258) );
AND2x4_ASAP7_75t_L g259 ( .A(n_188), .B(n_130), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_209), .B(n_125), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_220), .Y(n_261) );
AOI21xp5_ASAP7_75t_L g262 ( .A1(n_212), .A2(n_143), .B(n_130), .Y(n_262) );
AND2x2_ASAP7_75t_L g263 ( .A(n_174), .B(n_130), .Y(n_263) );
INVx2_ASAP7_75t_L g264 ( .A(n_213), .Y(n_264) );
NOR2xp33_ASAP7_75t_R g265 ( .A(n_199), .B(n_125), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_214), .Y(n_266) );
INVx2_ASAP7_75t_SL g267 ( .A(n_199), .Y(n_267) );
OR2x6_ASAP7_75t_L g268 ( .A(n_184), .B(n_143), .Y(n_268) );
AND2x4_ASAP7_75t_L g269 ( .A(n_208), .B(n_130), .Y(n_269) );
NOR2xp33_ASAP7_75t_R g270 ( .A(n_164), .B(n_125), .Y(n_270) );
BUFx12f_ASAP7_75t_L g271 ( .A(n_175), .Y(n_271) );
NOR2x1_ASAP7_75t_L g272 ( .A(n_217), .B(n_143), .Y(n_272) );
AND2x4_ASAP7_75t_L g273 ( .A(n_193), .B(n_143), .Y(n_273) );
NAND2xp5_ASAP7_75t_SL g274 ( .A(n_214), .B(n_125), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_218), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_201), .B(n_3), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_203), .B(n_6), .Y(n_277) );
BUFx2_ASAP7_75t_L g278 ( .A(n_206), .Y(n_278) );
AND2x4_ASAP7_75t_L g279 ( .A(n_168), .B(n_6), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_215), .B(n_7), .Y(n_280) );
INVx2_ASAP7_75t_SL g281 ( .A(n_216), .Y(n_281) );
AOI22xp33_ASAP7_75t_L g282 ( .A1(n_218), .A2(n_9), .B1(n_10), .B2(n_11), .Y(n_282) );
OR2x6_ASAP7_75t_L g283 ( .A(n_165), .B(n_10), .Y(n_283) );
BUFx3_ASAP7_75t_L g284 ( .A(n_165), .Y(n_284) );
OR2x2_ASAP7_75t_L g285 ( .A(n_212), .B(n_12), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_186), .Y(n_286) );
NAND2xp5_ASAP7_75t_SL g287 ( .A(n_186), .B(n_45), .Y(n_287) );
NAND2xp5_ASAP7_75t_SL g288 ( .A(n_223), .B(n_46), .Y(n_288) );
OR2x2_ASAP7_75t_L g289 ( .A(n_162), .B(n_13), .Y(n_289) );
OAI22xp5_ASAP7_75t_L g290 ( .A1(n_230), .A2(n_210), .B1(n_204), .B2(n_162), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_261), .Y(n_291) );
OAI22xp5_ASAP7_75t_L g292 ( .A1(n_230), .A2(n_210), .B1(n_204), .B2(n_170), .Y(n_292) );
INVxp67_ASAP7_75t_L g293 ( .A(n_278), .Y(n_293) );
INVx2_ASAP7_75t_L g294 ( .A(n_234), .Y(n_294) );
BUFx3_ASAP7_75t_L g295 ( .A(n_271), .Y(n_295) );
AND2x4_ASAP7_75t_L g296 ( .A(n_229), .B(n_14), .Y(n_296) );
BUFx2_ASAP7_75t_L g297 ( .A(n_252), .Y(n_297) );
HB1xp67_ASAP7_75t_L g298 ( .A(n_283), .Y(n_298) );
BUFx2_ASAP7_75t_L g299 ( .A(n_283), .Y(n_299) );
INVx2_ASAP7_75t_L g300 ( .A(n_234), .Y(n_300) );
INVx2_ASAP7_75t_L g301 ( .A(n_264), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_281), .B(n_182), .Y(n_302) );
INVxp67_ASAP7_75t_SL g303 ( .A(n_232), .Y(n_303) );
O2A1O1Ixp33_ASAP7_75t_SL g304 ( .A1(n_288), .A2(n_183), .B(n_200), .C(n_198), .Y(n_304) );
AOI22xp33_ASAP7_75t_L g305 ( .A1(n_279), .A2(n_182), .B1(n_200), .B2(n_198), .Y(n_305) );
OAI221xp5_ASAP7_75t_L g306 ( .A1(n_245), .A2(n_170), .B1(n_196), .B2(n_195), .C(n_171), .Y(n_306) );
BUFx4f_ASAP7_75t_L g307 ( .A(n_251), .Y(n_307) );
OAI21xp5_ASAP7_75t_L g308 ( .A1(n_257), .A2(n_181), .B(n_196), .Y(n_308) );
OA21x2_ASAP7_75t_L g309 ( .A1(n_274), .A2(n_171), .B(n_195), .Y(n_309) );
HB1xp67_ASAP7_75t_L g310 ( .A(n_283), .Y(n_310) );
AND2x4_ASAP7_75t_L g311 ( .A(n_229), .B(n_17), .Y(n_311) );
AND2x2_ASAP7_75t_L g312 ( .A(n_241), .B(n_17), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_255), .Y(n_313) );
AOI21xp5_ASAP7_75t_L g314 ( .A1(n_274), .A2(n_172), .B(n_178), .Y(n_314) );
NAND2x1p5_ASAP7_75t_L g315 ( .A(n_231), .B(n_172), .Y(n_315) );
HB1xp67_ASAP7_75t_L g316 ( .A(n_232), .Y(n_316) );
HB1xp67_ASAP7_75t_L g317 ( .A(n_243), .Y(n_317) );
INVx2_ASAP7_75t_L g318 ( .A(n_264), .Y(n_318) );
BUFx6f_ASAP7_75t_L g319 ( .A(n_231), .Y(n_319) );
INVx6_ASAP7_75t_L g320 ( .A(n_271), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_266), .Y(n_321) );
NAND2x1p5_ASAP7_75t_L g322 ( .A(n_231), .B(n_181), .Y(n_322) );
NOR2xp33_ASAP7_75t_L g323 ( .A(n_267), .B(n_18), .Y(n_323) );
NOR2xp33_ASAP7_75t_L g324 ( .A(n_224), .B(n_18), .Y(n_324) );
NAND2xp5_ASAP7_75t_SL g325 ( .A(n_265), .B(n_178), .Y(n_325) );
BUFx2_ASAP7_75t_L g326 ( .A(n_227), .Y(n_326) );
INVx3_ASAP7_75t_L g327 ( .A(n_231), .Y(n_327) );
INVx2_ASAP7_75t_L g328 ( .A(n_275), .Y(n_328) );
BUFx3_ASAP7_75t_L g329 ( .A(n_284), .Y(n_329) );
INVx2_ASAP7_75t_SL g330 ( .A(n_239), .Y(n_330) );
INVx3_ASAP7_75t_L g331 ( .A(n_284), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_233), .B(n_183), .Y(n_332) );
AOI22xp33_ASAP7_75t_SL g333 ( .A1(n_279), .A2(n_19), .B1(n_20), .B2(n_22), .Y(n_333) );
BUFx3_ASAP7_75t_L g334 ( .A(n_239), .Y(n_334) );
AOI22xp33_ASAP7_75t_L g335 ( .A1(n_246), .A2(n_187), .B1(n_192), .B2(n_189), .Y(n_335) );
INVx3_ASAP7_75t_L g336 ( .A(n_235), .Y(n_336) );
AOI21xp5_ASAP7_75t_L g337 ( .A1(n_258), .A2(n_187), .B(n_192), .Y(n_337) );
CKINVDCx5p33_ASAP7_75t_R g338 ( .A(n_227), .Y(n_338) );
INVx2_ASAP7_75t_L g339 ( .A(n_235), .Y(n_339) );
CKINVDCx20_ASAP7_75t_R g340 ( .A(n_338), .Y(n_340) );
AND2x4_ASAP7_75t_L g341 ( .A(n_295), .B(n_241), .Y(n_341) );
OR2x2_ASAP7_75t_L g342 ( .A(n_293), .B(n_254), .Y(n_342) );
OAI22xp5_ASAP7_75t_L g343 ( .A1(n_299), .A2(n_233), .B1(n_241), .B2(n_243), .Y(n_343) );
AOI22xp33_ASAP7_75t_L g344 ( .A1(n_296), .A2(n_279), .B1(n_256), .B2(n_239), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_312), .Y(n_345) );
CKINVDCx14_ASAP7_75t_R g346 ( .A(n_326), .Y(n_346) );
AOI21xp5_ASAP7_75t_L g347 ( .A1(n_337), .A2(n_260), .B(n_225), .Y(n_347) );
INVx4_ASAP7_75t_L g348 ( .A(n_320), .Y(n_348) );
INVx2_ASAP7_75t_L g349 ( .A(n_294), .Y(n_349) );
AO31x2_ASAP7_75t_L g350 ( .A1(n_290), .A2(n_276), .A3(n_277), .B(n_280), .Y(n_350) );
CKINVDCx20_ASAP7_75t_R g351 ( .A(n_326), .Y(n_351) );
NAND2xp33_ASAP7_75t_R g352 ( .A(n_299), .B(n_265), .Y(n_352) );
AOI221xp5_ASAP7_75t_L g353 ( .A1(n_293), .A2(n_228), .B1(n_240), .B2(n_263), .C(n_249), .Y(n_353) );
BUFx2_ASAP7_75t_L g354 ( .A(n_295), .Y(n_354) );
AOI22xp33_ASAP7_75t_L g355 ( .A1(n_296), .A2(n_256), .B1(n_268), .B2(n_259), .Y(n_355) );
BUFx3_ASAP7_75t_L g356 ( .A(n_295), .Y(n_356) );
AOI21xp5_ASAP7_75t_L g357 ( .A1(n_337), .A2(n_253), .B(n_247), .Y(n_357) );
OAI221xp5_ASAP7_75t_L g358 ( .A1(n_324), .A2(n_237), .B1(n_268), .B2(n_236), .C(n_238), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_312), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_312), .B(n_249), .Y(n_360) );
INVx4_ASAP7_75t_L g361 ( .A(n_320), .Y(n_361) );
AOI221xp5_ASAP7_75t_L g362 ( .A1(n_297), .A2(n_269), .B1(n_273), .B2(n_254), .C(n_259), .Y(n_362) );
NOR2xp33_ASAP7_75t_L g363 ( .A(n_297), .B(n_256), .Y(n_363) );
OA21x2_ASAP7_75t_L g364 ( .A1(n_314), .A2(n_288), .B(n_287), .Y(n_364) );
AOI21xp33_ASAP7_75t_L g365 ( .A1(n_298), .A2(n_310), .B(n_323), .Y(n_365) );
OR2x2_ASAP7_75t_L g366 ( .A(n_298), .B(n_268), .Y(n_366) );
CKINVDCx5p33_ASAP7_75t_R g367 ( .A(n_320), .Y(n_367) );
OAI221xp5_ASAP7_75t_L g368 ( .A1(n_310), .A2(n_272), .B1(n_242), .B2(n_244), .C(n_248), .Y(n_368) );
OAI21xp33_ASAP7_75t_SL g369 ( .A1(n_291), .A2(n_282), .B(n_285), .Y(n_369) );
OAI22xp5_ASAP7_75t_L g370 ( .A1(n_303), .A2(n_282), .B1(n_273), .B2(n_289), .Y(n_370) );
AOI22xp33_ASAP7_75t_L g371 ( .A1(n_362), .A2(n_296), .B1(n_311), .B2(n_333), .Y(n_371) );
INVx2_ASAP7_75t_L g372 ( .A(n_349), .Y(n_372) );
HB1xp67_ASAP7_75t_L g373 ( .A(n_349), .Y(n_373) );
NAND2xp5_ASAP7_75t_SL g374 ( .A(n_356), .B(n_226), .Y(n_374) );
AOI21xp5_ASAP7_75t_L g375 ( .A1(n_347), .A2(n_304), .B(n_314), .Y(n_375) );
AND2x4_ASAP7_75t_L g376 ( .A(n_356), .B(n_291), .Y(n_376) );
AOI22xp33_ASAP7_75t_L g377 ( .A1(n_355), .A2(n_296), .B1(n_311), .B2(n_333), .Y(n_377) );
INVx1_ASAP7_75t_SL g378 ( .A(n_341), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_345), .Y(n_379) );
AND2x4_ASAP7_75t_L g380 ( .A(n_348), .B(n_328), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_359), .Y(n_381) );
AOI22xp33_ASAP7_75t_SL g382 ( .A1(n_346), .A2(n_311), .B1(n_296), .B2(n_320), .Y(n_382) );
AOI22xp33_ASAP7_75t_L g383 ( .A1(n_353), .A2(n_311), .B1(n_273), .B2(n_269), .Y(n_383) );
OR2x2_ASAP7_75t_L g384 ( .A(n_360), .B(n_328), .Y(n_384) );
AOI22xp33_ASAP7_75t_L g385 ( .A1(n_358), .A2(n_311), .B1(n_269), .B2(n_334), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_350), .Y(n_386) );
AND2x2_ASAP7_75t_L g387 ( .A(n_341), .B(n_328), .Y(n_387) );
AND2x2_ASAP7_75t_L g388 ( .A(n_341), .B(n_344), .Y(n_388) );
OAI22xp33_ASAP7_75t_L g389 ( .A1(n_370), .A2(n_321), .B1(n_303), .B2(n_332), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_350), .Y(n_390) );
AOI222xp33_ASAP7_75t_L g391 ( .A1(n_343), .A2(n_313), .B1(n_321), .B2(n_226), .C1(n_332), .C2(n_334), .Y(n_391) );
OAI21xp5_ASAP7_75t_L g392 ( .A1(n_369), .A2(n_292), .B(n_290), .Y(n_392) );
AOI22xp33_ASAP7_75t_L g393 ( .A1(n_366), .A2(n_334), .B1(n_320), .B2(n_330), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_350), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_350), .B(n_313), .Y(n_395) );
AOI22xp33_ASAP7_75t_L g396 ( .A1(n_365), .A2(n_330), .B1(n_336), .B2(n_316), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_357), .Y(n_397) );
AND2x2_ASAP7_75t_L g398 ( .A(n_387), .B(n_294), .Y(n_398) );
INVx2_ASAP7_75t_L g399 ( .A(n_372), .Y(n_399) );
BUFx10_ASAP7_75t_L g400 ( .A(n_380), .Y(n_400) );
OAI211xp5_ASAP7_75t_L g401 ( .A1(n_382), .A2(n_346), .B(n_342), .C(n_354), .Y(n_401) );
AND2x2_ASAP7_75t_L g402 ( .A(n_387), .B(n_294), .Y(n_402) );
BUFx2_ASAP7_75t_L g403 ( .A(n_373), .Y(n_403) );
OAI211xp5_ASAP7_75t_L g404 ( .A1(n_382), .A2(n_363), .B(n_351), .C(n_367), .Y(n_404) );
AOI21xp5_ASAP7_75t_L g405 ( .A1(n_389), .A2(n_364), .B(n_287), .Y(n_405) );
INVx2_ASAP7_75t_L g406 ( .A(n_372), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_373), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_379), .B(n_351), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_372), .Y(n_409) );
AOI21xp5_ASAP7_75t_L g410 ( .A1(n_389), .A2(n_364), .B(n_318), .Y(n_410) );
AOI22xp5_ASAP7_75t_L g411 ( .A1(n_371), .A2(n_377), .B1(n_383), .B2(n_388), .Y(n_411) );
AOI22xp33_ASAP7_75t_L g412 ( .A1(n_388), .A2(n_368), .B1(n_361), .B2(n_348), .Y(n_412) );
AOI22xp33_ASAP7_75t_SL g413 ( .A1(n_392), .A2(n_361), .B1(n_348), .B2(n_340), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_379), .B(n_361), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_386), .Y(n_415) );
OR2x2_ASAP7_75t_L g416 ( .A(n_395), .B(n_318), .Y(n_416) );
AOI22xp33_ASAP7_75t_L g417 ( .A1(n_391), .A2(n_316), .B1(n_317), .B2(n_330), .Y(n_417) );
HB1xp67_ASAP7_75t_L g418 ( .A(n_380), .Y(n_418) );
AOI221xp5_ASAP7_75t_L g419 ( .A1(n_381), .A2(n_292), .B1(n_306), .B2(n_262), .C(n_305), .Y(n_419) );
AOI21xp5_ASAP7_75t_L g420 ( .A1(n_395), .A2(n_364), .B(n_300), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_386), .Y(n_421) );
OAI221xp5_ASAP7_75t_L g422 ( .A1(n_385), .A2(n_352), .B1(n_306), .B2(n_336), .C(n_335), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_390), .Y(n_423) );
INVxp67_ASAP7_75t_L g424 ( .A(n_376), .Y(n_424) );
AOI22xp33_ASAP7_75t_SL g425 ( .A1(n_392), .A2(n_340), .B1(n_352), .B2(n_329), .Y(n_425) );
CKINVDCx8_ASAP7_75t_R g426 ( .A(n_380), .Y(n_426) );
HB1xp67_ASAP7_75t_L g427 ( .A(n_380), .Y(n_427) );
INVx2_ASAP7_75t_L g428 ( .A(n_397), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_390), .Y(n_429) );
AND2x2_ASAP7_75t_L g430 ( .A(n_381), .B(n_300), .Y(n_430) );
OAI221xp5_ASAP7_75t_L g431 ( .A1(n_396), .A2(n_336), .B1(n_335), .B2(n_339), .C(n_302), .Y(n_431) );
AOI22xp33_ASAP7_75t_L g432 ( .A1(n_391), .A2(n_317), .B1(n_339), .B2(n_329), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_384), .B(n_336), .Y(n_433) );
BUFx3_ASAP7_75t_L g434 ( .A(n_426), .Y(n_434) );
INVx1_ASAP7_75t_SL g435 ( .A(n_403), .Y(n_435) );
AOI22xp33_ASAP7_75t_L g436 ( .A1(n_411), .A2(n_376), .B1(n_378), .B2(n_394), .Y(n_436) );
HB1xp67_ASAP7_75t_L g437 ( .A(n_403), .Y(n_437) );
BUFx3_ASAP7_75t_L g438 ( .A(n_426), .Y(n_438) );
AND2x2_ASAP7_75t_L g439 ( .A(n_409), .B(n_394), .Y(n_439) );
OAI22xp5_ASAP7_75t_L g440 ( .A1(n_411), .A2(n_384), .B1(n_378), .B2(n_376), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_415), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_415), .B(n_421), .Y(n_442) );
AND2x2_ASAP7_75t_L g443 ( .A(n_409), .B(n_397), .Y(n_443) );
INVx2_ASAP7_75t_L g444 ( .A(n_428), .Y(n_444) );
CKINVDCx5p33_ASAP7_75t_R g445 ( .A(n_408), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_421), .Y(n_446) );
AND2x2_ASAP7_75t_L g447 ( .A(n_399), .B(n_406), .Y(n_447) );
AND2x2_ASAP7_75t_L g448 ( .A(n_399), .B(n_376), .Y(n_448) );
OR2x2_ASAP7_75t_L g449 ( .A(n_407), .B(n_318), .Y(n_449) );
OR2x2_ASAP7_75t_L g450 ( .A(n_407), .B(n_301), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_423), .Y(n_451) );
OR2x2_ASAP7_75t_L g452 ( .A(n_416), .B(n_301), .Y(n_452) );
NAND2xp5_ASAP7_75t_SL g453 ( .A(n_413), .B(n_374), .Y(n_453) );
BUFx2_ASAP7_75t_SL g454 ( .A(n_400), .Y(n_454) );
AND2x2_ASAP7_75t_L g455 ( .A(n_399), .B(n_301), .Y(n_455) );
AOI22xp33_ASAP7_75t_L g456 ( .A1(n_425), .A2(n_393), .B1(n_329), .B2(n_331), .Y(n_456) );
INVx2_ASAP7_75t_L g457 ( .A(n_428), .Y(n_457) );
OAI33xp33_ASAP7_75t_L g458 ( .A1(n_423), .A2(n_189), .A3(n_22), .B1(n_23), .B2(n_176), .B3(n_173), .Y(n_458) );
NAND3xp33_ASAP7_75t_L g459 ( .A(n_428), .B(n_375), .C(n_179), .Y(n_459) );
AND2x2_ASAP7_75t_L g460 ( .A(n_406), .B(n_300), .Y(n_460) );
AND2x2_ASAP7_75t_L g461 ( .A(n_406), .B(n_23), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_429), .Y(n_462) );
NOR2x1_ASAP7_75t_L g463 ( .A(n_401), .B(n_375), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_429), .B(n_331), .Y(n_464) );
AND2x2_ASAP7_75t_L g465 ( .A(n_416), .B(n_309), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_420), .Y(n_466) );
NAND3xp33_ASAP7_75t_L g467 ( .A(n_412), .B(n_175), .C(n_177), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_430), .B(n_331), .Y(n_468) );
INVx2_ASAP7_75t_L g469 ( .A(n_430), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_418), .B(n_331), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_427), .Y(n_471) );
INVx2_ASAP7_75t_L g472 ( .A(n_400), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_410), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_400), .Y(n_474) );
AND2x2_ASAP7_75t_L g475 ( .A(n_398), .B(n_309), .Y(n_475) );
AOI221xp5_ASAP7_75t_L g476 ( .A1(n_417), .A2(n_302), .B1(n_339), .B2(n_247), .C(n_308), .Y(n_476) );
INVx2_ASAP7_75t_L g477 ( .A(n_400), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_398), .B(n_309), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_402), .Y(n_479) );
OR2x2_ASAP7_75t_L g480 ( .A(n_424), .B(n_309), .Y(n_480) );
INVx2_ASAP7_75t_SL g481 ( .A(n_414), .Y(n_481) );
INVxp67_ASAP7_75t_L g482 ( .A(n_402), .Y(n_482) );
HB1xp67_ASAP7_75t_L g483 ( .A(n_433), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_405), .Y(n_484) );
AND2x2_ASAP7_75t_L g485 ( .A(n_439), .B(n_432), .Y(n_485) );
OR2x2_ASAP7_75t_L g486 ( .A(n_482), .B(n_404), .Y(n_486) );
INVxp67_ASAP7_75t_L g487 ( .A(n_454), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_441), .Y(n_488) );
AND2x4_ASAP7_75t_SL g489 ( .A(n_472), .B(n_327), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_441), .Y(n_490) );
INVx2_ASAP7_75t_L g491 ( .A(n_444), .Y(n_491) );
OR2x2_ASAP7_75t_L g492 ( .A(n_435), .B(n_422), .Y(n_492) );
INVx2_ASAP7_75t_L g493 ( .A(n_444), .Y(n_493) );
AND2x2_ASAP7_75t_L g494 ( .A(n_439), .B(n_419), .Y(n_494) );
AND4x1_ASAP7_75t_L g495 ( .A(n_467), .B(n_26), .C(n_27), .D(n_33), .Y(n_495) );
NOR2xp33_ASAP7_75t_L g496 ( .A(n_445), .B(n_431), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_482), .B(n_309), .Y(n_497) );
INVx2_ASAP7_75t_SL g498 ( .A(n_472), .Y(n_498) );
OAI22xp5_ASAP7_75t_SL g499 ( .A1(n_434), .A2(n_319), .B1(n_327), .B2(n_322), .Y(n_499) );
OAI21xp33_ASAP7_75t_SL g500 ( .A1(n_453), .A2(n_325), .B(n_308), .Y(n_500) );
OR2x2_ASAP7_75t_L g501 ( .A(n_435), .B(n_173), .Y(n_501) );
INVx2_ASAP7_75t_L g502 ( .A(n_444), .Y(n_502) );
OR2x2_ASAP7_75t_L g503 ( .A(n_437), .B(n_471), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_479), .B(n_286), .Y(n_504) );
AND2x2_ASAP7_75t_L g505 ( .A(n_446), .B(n_194), .Y(n_505) );
INVx2_ASAP7_75t_L g506 ( .A(n_457), .Y(n_506) );
INVx3_ASAP7_75t_L g507 ( .A(n_477), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_479), .B(n_176), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_451), .Y(n_509) );
AOI21xp33_ASAP7_75t_L g510 ( .A1(n_463), .A2(n_179), .B(n_177), .Y(n_510) );
AND2x2_ASAP7_75t_L g511 ( .A(n_451), .B(n_179), .Y(n_511) );
INVx2_ASAP7_75t_L g512 ( .A(n_457), .Y(n_512) );
OR2x2_ASAP7_75t_L g513 ( .A(n_471), .B(n_175), .Y(n_513) );
NOR2xp33_ASAP7_75t_R g514 ( .A(n_434), .B(n_327), .Y(n_514) );
NAND2xp5_ASAP7_75t_SL g515 ( .A(n_467), .B(n_319), .Y(n_515) );
AND2x2_ASAP7_75t_L g516 ( .A(n_462), .B(n_175), .Y(n_516) );
NOR3xp33_ASAP7_75t_L g517 ( .A(n_458), .B(n_202), .C(n_327), .Y(n_517) );
AND2x2_ASAP7_75t_L g518 ( .A(n_443), .B(n_469), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_442), .Y(n_519) );
NOR4xp25_ASAP7_75t_SL g520 ( .A(n_476), .B(n_43), .C(n_52), .D(n_53), .Y(n_520) );
NOR4xp25_ASAP7_75t_L g521 ( .A(n_440), .B(n_56), .C(n_61), .D(n_62), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_442), .Y(n_522) );
OR2x2_ASAP7_75t_L g523 ( .A(n_469), .B(n_179), .Y(n_523) );
AND2x2_ASAP7_75t_L g524 ( .A(n_443), .B(n_179), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_483), .B(n_177), .Y(n_525) );
NOR2xp33_ASAP7_75t_R g526 ( .A(n_434), .B(n_63), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_461), .Y(n_527) );
AND2x2_ASAP7_75t_L g528 ( .A(n_448), .B(n_177), .Y(n_528) );
OR2x2_ASAP7_75t_L g529 ( .A(n_481), .B(n_65), .Y(n_529) );
INVx2_ASAP7_75t_L g530 ( .A(n_457), .Y(n_530) );
OR2x2_ASAP7_75t_L g531 ( .A(n_481), .B(n_67), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_461), .Y(n_532) );
NAND2xp33_ASAP7_75t_SL g533 ( .A(n_477), .B(n_270), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_449), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_449), .Y(n_535) );
AND2x2_ASAP7_75t_L g536 ( .A(n_448), .B(n_177), .Y(n_536) );
AND2x2_ASAP7_75t_L g537 ( .A(n_447), .B(n_69), .Y(n_537) );
AOI21xp33_ASAP7_75t_L g538 ( .A1(n_496), .A2(n_463), .B(n_474), .Y(n_538) );
OR2x2_ASAP7_75t_L g539 ( .A(n_518), .B(n_452), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_503), .Y(n_540) );
XNOR2xp5_ASAP7_75t_L g541 ( .A(n_518), .B(n_454), .Y(n_541) );
INVx3_ASAP7_75t_L g542 ( .A(n_507), .Y(n_542) );
OAI21xp33_ASAP7_75t_SL g543 ( .A1(n_487), .A2(n_450), .B(n_452), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_519), .B(n_436), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_522), .B(n_465), .Y(n_545) );
NAND3xp33_ASAP7_75t_SL g546 ( .A(n_526), .B(n_476), .C(n_456), .Y(n_546) );
INVx2_ASAP7_75t_L g547 ( .A(n_491), .Y(n_547) );
OAI211xp5_ASAP7_75t_SL g548 ( .A1(n_500), .A2(n_470), .B(n_466), .C(n_468), .Y(n_548) );
AOI21xp33_ASAP7_75t_L g549 ( .A1(n_486), .A2(n_466), .B(n_473), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_488), .Y(n_550) );
OAI21xp5_ASAP7_75t_L g551 ( .A1(n_521), .A2(n_450), .B(n_459), .Y(n_551) );
AOI21xp5_ASAP7_75t_L g552 ( .A1(n_515), .A2(n_458), .B(n_459), .Y(n_552) );
AOI211x1_ASAP7_75t_L g553 ( .A1(n_495), .A2(n_464), .B(n_470), .C(n_468), .Y(n_553) );
NOR2x1_ASAP7_75t_L g554 ( .A(n_515), .B(n_438), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_494), .B(n_465), .Y(n_555) );
NAND3xp33_ASAP7_75t_L g556 ( .A(n_492), .B(n_484), .C(n_473), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_494), .B(n_464), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_490), .Y(n_558) );
O2A1O1Ixp33_ASAP7_75t_L g559 ( .A1(n_504), .A2(n_484), .B(n_438), .C(n_480), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_509), .Y(n_560) );
AOI322xp5_ASAP7_75t_L g561 ( .A1(n_485), .A2(n_475), .A3(n_478), .B1(n_460), .B2(n_455), .C1(n_480), .C2(n_70), .Y(n_561) );
HB1xp67_ASAP7_75t_L g562 ( .A(n_498), .Y(n_562) );
AOI21xp5_ASAP7_75t_L g563 ( .A1(n_533), .A2(n_478), .B(n_460), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_534), .B(n_475), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_535), .B(n_319), .Y(n_565) );
INVx3_ASAP7_75t_SL g566 ( .A(n_489), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_513), .Y(n_567) );
AOI22xp33_ASAP7_75t_L g568 ( .A1(n_485), .A2(n_319), .B1(n_270), .B2(n_315), .Y(n_568) );
AND2x2_ASAP7_75t_L g569 ( .A(n_507), .B(n_512), .Y(n_569) );
INVxp67_ASAP7_75t_SL g570 ( .A(n_513), .Y(n_570) );
OAI21xp5_ASAP7_75t_SL g571 ( .A1(n_492), .A2(n_315), .B(n_322), .Y(n_571) );
OAI22xp5_ASAP7_75t_L g572 ( .A1(n_529), .A2(n_319), .B1(n_307), .B2(n_322), .Y(n_572) );
NAND2x1_ASAP7_75t_L g573 ( .A(n_507), .B(n_319), .Y(n_573) );
INVxp33_ASAP7_75t_L g574 ( .A(n_526), .Y(n_574) );
INVx2_ASAP7_75t_L g575 ( .A(n_493), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_493), .Y(n_576) );
O2A1O1Ixp33_ASAP7_75t_L g577 ( .A1(n_531), .A2(n_315), .B(n_322), .C(n_307), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_502), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_527), .B(n_319), .Y(n_579) );
AOI21xp5_ASAP7_75t_L g580 ( .A1(n_533), .A2(n_307), .B(n_315), .Y(n_580) );
INVxp67_ASAP7_75t_L g581 ( .A(n_562), .Y(n_581) );
AOI321xp33_ASAP7_75t_L g582 ( .A1(n_559), .A2(n_532), .A3(n_537), .B1(n_525), .B2(n_517), .C(n_528), .Y(n_582) );
INVx2_ASAP7_75t_L g583 ( .A(n_547), .Y(n_583) );
AND2x2_ASAP7_75t_L g584 ( .A(n_540), .B(n_498), .Y(n_584) );
NOR3xp33_ASAP7_75t_SL g585 ( .A(n_546), .B(n_499), .C(n_497), .Y(n_585) );
NOR3xp33_ASAP7_75t_SL g586 ( .A(n_543), .B(n_508), .C(n_510), .Y(n_586) );
NOR2xp33_ASAP7_75t_L g587 ( .A(n_538), .B(n_574), .Y(n_587) );
AOI22xp5_ASAP7_75t_L g588 ( .A1(n_574), .A2(n_544), .B1(n_571), .B2(n_557), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_550), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_558), .Y(n_590) );
NOR3xp33_ASAP7_75t_SL g591 ( .A(n_551), .B(n_514), .C(n_520), .Y(n_591) );
NAND3xp33_ASAP7_75t_L g592 ( .A(n_556), .B(n_511), .C(n_516), .Y(n_592) );
AOI321xp33_ASAP7_75t_R g593 ( .A1(n_555), .A2(n_512), .A3(n_530), .B1(n_506), .B2(n_505), .C(n_511), .Y(n_593) );
NOR3xp33_ASAP7_75t_SL g594 ( .A(n_548), .B(n_489), .C(n_536), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_560), .Y(n_595) );
INVxp33_ASAP7_75t_L g596 ( .A(n_554), .Y(n_596) );
NAND2xp33_ASAP7_75t_SL g597 ( .A(n_566), .B(n_530), .Y(n_597) );
NOR2xp33_ASAP7_75t_L g598 ( .A(n_549), .B(n_506), .Y(n_598) );
AND2x2_ASAP7_75t_L g599 ( .A(n_541), .B(n_536), .Y(n_599) );
OAI22xp33_ASAP7_75t_L g600 ( .A1(n_566), .A2(n_501), .B1(n_523), .B2(n_524), .Y(n_600) );
XOR2x2_ASAP7_75t_L g601 ( .A(n_553), .B(n_524), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_570), .Y(n_602) );
NAND2xp33_ASAP7_75t_R g603 ( .A(n_542), .B(n_528), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_570), .B(n_505), .Y(n_604) );
AND2x2_ASAP7_75t_L g605 ( .A(n_569), .B(n_523), .Y(n_605) );
AND2x2_ASAP7_75t_L g606 ( .A(n_539), .B(n_501), .Y(n_606) );
NOR2x1_ASAP7_75t_L g607 ( .A(n_573), .B(n_250), .Y(n_607) );
INVxp67_ASAP7_75t_L g608 ( .A(n_562), .Y(n_608) );
NOR4xp75_ASAP7_75t_L g609 ( .A(n_564), .B(n_250), .C(n_545), .D(n_572), .Y(n_609) );
O2A1O1Ixp33_ASAP7_75t_SL g610 ( .A1(n_561), .A2(n_250), .B(n_577), .C(n_552), .Y(n_610) );
OAI22xp5_ASAP7_75t_L g611 ( .A1(n_588), .A2(n_567), .B1(n_542), .B2(n_563), .Y(n_611) );
XNOR2xp5_ASAP7_75t_L g612 ( .A(n_601), .B(n_568), .Y(n_612) );
NAND4xp75_ASAP7_75t_L g613 ( .A(n_591), .B(n_580), .C(n_565), .D(n_569), .Y(n_613) );
HB1xp67_ASAP7_75t_L g614 ( .A(n_581), .Y(n_614) );
OAI22xp5_ASAP7_75t_L g615 ( .A1(n_593), .A2(n_568), .B1(n_576), .B2(n_578), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_602), .Y(n_616) );
BUFx2_ASAP7_75t_L g617 ( .A(n_597), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_589), .Y(n_618) );
XNOR2xp5_ASAP7_75t_L g619 ( .A(n_601), .B(n_579), .Y(n_619) );
AND2x4_ASAP7_75t_L g620 ( .A(n_608), .B(n_547), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_590), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_595), .Y(n_622) );
INVx2_ASAP7_75t_L g623 ( .A(n_583), .Y(n_623) );
OAI21xp5_ASAP7_75t_SL g624 ( .A1(n_596), .A2(n_587), .B(n_592), .Y(n_624) );
INVx1_ASAP7_75t_SL g625 ( .A(n_597), .Y(n_625) );
XNOR2x1_ASAP7_75t_L g626 ( .A(n_609), .B(n_575), .Y(n_626) );
NOR3xp33_ASAP7_75t_L g627 ( .A(n_613), .B(n_610), .C(n_600), .Y(n_627) );
AOI211xp5_ASAP7_75t_L g628 ( .A1(n_624), .A2(n_610), .B(n_598), .C(n_599), .Y(n_628) );
AOI211xp5_ASAP7_75t_L g629 ( .A1(n_612), .A2(n_598), .B(n_604), .C(n_584), .Y(n_629) );
OAI211xp5_ASAP7_75t_SL g630 ( .A1(n_625), .A2(n_585), .B(n_586), .C(n_582), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_616), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_614), .Y(n_632) );
XNOR2x1_ASAP7_75t_L g633 ( .A(n_612), .B(n_606), .Y(n_633) );
AOI221x1_ASAP7_75t_L g634 ( .A1(n_611), .A2(n_605), .B1(n_603), .B2(n_594), .C(n_607), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_615), .B(n_603), .Y(n_635) );
NOR2xp33_ASAP7_75t_L g636 ( .A(n_619), .B(n_622), .Y(n_636) );
AO22x2_ASAP7_75t_L g637 ( .A1(n_613), .A2(n_626), .B1(n_618), .B2(n_621), .Y(n_637) );
OAI211xp5_ASAP7_75t_L g638 ( .A1(n_623), .A2(n_624), .B(n_617), .C(n_587), .Y(n_638) );
OAI21xp33_ASAP7_75t_L g639 ( .A1(n_626), .A2(n_624), .B(n_612), .Y(n_639) );
NAND3xp33_ASAP7_75t_L g640 ( .A(n_620), .B(n_624), .C(n_612), .Y(n_640) );
INVx2_ASAP7_75t_SL g641 ( .A(n_632), .Y(n_641) );
HB1xp67_ASAP7_75t_L g642 ( .A(n_631), .Y(n_642) );
AND2x4_ASAP7_75t_L g643 ( .A(n_634), .B(n_640), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_639), .B(n_633), .Y(n_644) );
OAI22xp5_ASAP7_75t_L g645 ( .A1(n_643), .A2(n_637), .B1(n_635), .B2(n_629), .Y(n_645) );
XNOR2xp5_ASAP7_75t_L g646 ( .A(n_644), .B(n_628), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_642), .Y(n_647) );
INVx2_ASAP7_75t_L g648 ( .A(n_647), .Y(n_648) );
HB1xp67_ASAP7_75t_L g649 ( .A(n_646), .Y(n_649) );
OAI32xp33_ASAP7_75t_L g650 ( .A1(n_649), .A2(n_645), .A3(n_627), .B1(n_643), .B2(n_641), .Y(n_650) );
AOI22xp5_ASAP7_75t_L g651 ( .A1(n_650), .A2(n_648), .B1(n_638), .B2(n_630), .Y(n_651) );
AOI21xp5_ASAP7_75t_L g652 ( .A1(n_651), .A2(n_630), .B(n_636), .Y(n_652) );
endmodule