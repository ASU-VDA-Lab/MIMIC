module real_aes_9312_n_282 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_281, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_274, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_269, n_152, n_198, n_201, n_122, n_7, n_228, n_272, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_275, n_69, n_279, n_46, n_109, n_59, n_25, n_203, n_236, n_278, n_73, n_77, n_218, n_81, n_133, n_48, n_267, n_270, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_273, n_138, n_50, n_114, n_276, n_89, n_170, n_277, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_271, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_258, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_280, n_38, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_268, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_282);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_281;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_274;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_269;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_272;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_275;
input n_69;
input n_279;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_278;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_267;
input n_270;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_273;
input n_138;
input n_50;
input n_114;
input n_276;
input n_89;
input n_170;
input n_277;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_271;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_280;
input n_38;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_268;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_282;
wire n_476;
wire n_599;
wire n_887;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_1591;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_1423;
wire n_571;
wire n_549;
wire n_1034;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1468;
wire n_870;
wire n_1248;
wire n_1602;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_1520;
wire n_1453;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_292;
wire n_1379;
wire n_400;
wire n_1597;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_553;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1225;
wire n_1441;
wire n_875;
wire n_1199;
wire n_951;
wire n_1382;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_1599;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_1537;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_1607;
wire n_455;
wire n_682;
wire n_812;
wire n_817;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_1588;
wire n_363;
wire n_1317;
wire n_417;
wire n_323;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1589;
wire n_947;
wire n_970;
wire n_1149;
wire n_368;
wire n_527;
wire n_1342;
wire n_1440;
wire n_1346;
wire n_552;
wire n_1383;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_805;
wire n_1600;
wire n_619;
wire n_1250;
wire n_1095;
wire n_1284;
wire n_360;
wire n_1583;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_488;
wire n_501;
wire n_1380;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1502;
wire n_404;
wire n_1073;
wire n_728;
wire n_1301;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_306;
wire n_1003;
wire n_346;
wire n_293;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1587;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_290;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1510;
wire n_1495;
wire n_712;
wire n_422;
wire n_861;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_1445;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_652;
wire n_1538;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_1488;
wire n_337;
wire n_1572;
wire n_1514;
wire n_480;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_635;
wire n_792;
wire n_1392;
wire n_1542;
wire n_665;
wire n_667;
wire n_991;
wire n_1556;
wire n_580;
wire n_1004;
wire n_1370;
wire n_1417;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_328;
wire n_1260;
wire n_355;
wire n_1606;
wire n_1129;
wire n_1285;
wire n_1014;
wire n_742;
wire n_1385;
wire n_461;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_1594;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1613;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_948;
wire n_1499;
wire n_399;
wire n_700;
wire n_1269;
wire n_677;
wire n_378;
wire n_591;
wire n_1518;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1577;
wire n_1406;
wire n_550;
wire n_966;
wire n_333;
wire n_1568;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1612;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_1611;
wire n_992;
wire n_813;
wire n_1338;
wire n_981;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1189;
wire n_1070;
wire n_535;
wire n_882;
wire n_1210;
wire n_1456;
wire n_746;
wire n_656;
wire n_1614;
wire n_1148;
wire n_860;
wire n_748;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_311;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_617;
wire n_602;
wire n_402;
wire n_733;
wire n_1404;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_286;
wire n_1011;
wire n_416;
wire n_1567;
wire n_1569;
wire n_895;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_645;
wire n_1145;
wire n_1529;
wire n_557;
wire n_777;
wire n_985;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_296;
wire n_1347;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_735;
wire n_1179;
wire n_334;
wire n_1171;
wire n_569;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_1580;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1551;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_354;
wire n_720;
wire n_1026;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_643;
wire n_1403;
wire n_486;
wire n_291;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_1513;
wire n_1194;
wire n_389;
wire n_1609;
wire n_1462;
wire n_701;
wire n_809;
wire n_1532;
wire n_679;
wire n_520;
wire n_926;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_300;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1474;
wire n_721;
wire n_1431;
wire n_1133;
wire n_1593;
wire n_313;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1162;
wire n_1463;
wire n_762;
wire n_1524;
wire n_325;
wire n_1298;
wire n_442;
wire n_740;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_459;
wire n_1172;
wire n_998;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_1578;
wire n_473;
wire n_967;
wire n_1159;
wire n_474;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_307;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_285;
wire n_1377;
wire n_800;
wire n_778;
wire n_1175;
wire n_1170;
wire n_522;
wire n_1475;
wire n_943;
wire n_977;
wire n_287;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1333;
wire n_577;
wire n_1610;
wire n_759;
wire n_1235;
wire n_299;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_766;
wire n_852;
wire n_1268;
wire n_1113;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_865;
wire n_594;
wire n_856;
wire n_1146;
wire n_1435;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_1540;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_1470;
wire n_816;
wire n_625;
wire n_953;
wire n_289;
wire n_1565;
wire n_1373;
wire n_1558;
wire n_716;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_370;
wire n_352;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_284;
wire n_316;
wire n_1168;
wire n_1598;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1263;
wire n_1411;
wire n_1115;
wire n_310;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_1555;
wire n_324;
wire n_664;
wire n_367;
wire n_1017;
wire n_936;
wire n_581;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1608;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_1560;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1414;
wire n_502;
wire n_434;
wire n_769;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_1450;
wire n_1603;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_288;
wire n_303;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_366;
wire n_1083;
wire n_727;
wire n_397;
wire n_1056;
wire n_1592;
wire n_1605;
wire n_663;
wire n_588;
wire n_1448;
wire n_707;
wire n_915;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1038;
wire n_1085;
wire n_295;
wire n_845;
wire n_1127;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_1581;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1355;
wire n_309;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_1496;
wire n_524;
wire n_1378;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_525;
wire n_1226;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_929;
wire n_1143;
wire n_1190;
wire n_543;
wire n_305;
wire n_585;
wire n_465;
wire n_719;
wire n_1457;
wire n_1343;
wire n_1604;
wire n_1156;
wire n_988;
wire n_1466;
wire n_921;
wire n_1396;
wire n_1176;
wire n_640;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_1211;
wire n_650;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_1480;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1407;
wire n_1104;
wire n_1061;
wire n_849;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1590;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_1596;
wire n_987;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_319;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_376;
wire n_308;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_460;
wire n_317;
wire n_1595;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1381;
wire n_1582;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1541;
wire n_1272;
wire n_408;
wire n_578;
wire n_372;
wire n_892;
wire n_938;
wire n_327;
wire n_774;
wire n_466;
wire n_1584;
wire n_559;
wire n_1277;
wire n_1049;
wire n_984;
wire n_301;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_532;
wire n_1025;
wire n_298;
wire n_924;
wire n_1264;
wire n_1527;
wire n_297;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_304;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1318;
wire n_1290;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_1100;
wire n_398;
wire n_1519;
wire n_425;
wire n_879;
wire n_331;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1547;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1356;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1249;
wire n_1416;
wire n_387;
wire n_1239;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_302;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_1252;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1430;
wire n_1481;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1536;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1601;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1573;
wire n_1130;
wire n_794;
wire n_283;
wire n_314;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1253;
wire n_312;
wire n_1183;
wire n_335;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_338;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1412;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_340;
wire n_483;
wire n_394;
wire n_729;
wire n_1280;
wire n_1323;
wire n_1352;
wire n_1097;
wire n_703;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_342;
wire n_348;
wire n_1528;
wire n_603;
wire n_1288;
wire n_868;
wire n_1024;
wire n_1144;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_429;
AO221x1_ASAP7_75t_L g1345 ( .A1(n_0), .A2(n_177), .B1(n_1263), .B2(n_1336), .C(n_1346), .Y(n_1345) );
CKINVDCx5p33_ASAP7_75t_R g1558 ( .A(n_1), .Y(n_1558) );
OAI221xp5_ASAP7_75t_L g496 ( .A1(n_2), .A2(n_497), .B1(n_500), .B2(n_509), .C(n_512), .Y(n_496) );
AOI21xp33_ASAP7_75t_L g567 ( .A1(n_2), .A2(n_568), .B(n_570), .Y(n_567) );
INVx1_ASAP7_75t_L g1105 ( .A(n_3), .Y(n_1105) );
OAI221xp5_ASAP7_75t_L g1129 ( .A1(n_3), .A2(n_86), .B1(n_1130), .B2(n_1131), .C(n_1132), .Y(n_1129) );
AOI22xp33_ASAP7_75t_L g1112 ( .A1(n_4), .A2(n_279), .B1(n_335), .B2(n_562), .Y(n_1112) );
INVx1_ASAP7_75t_L g1141 ( .A(n_4), .Y(n_1141) );
INVx1_ASAP7_75t_L g1207 ( .A(n_5), .Y(n_1207) );
OAI221xp5_ASAP7_75t_L g1234 ( .A1(n_5), .A2(n_37), .B1(n_1062), .B2(n_1235), .C(n_1236), .Y(n_1234) );
AOI22xp33_ASAP7_75t_SL g687 ( .A1(n_6), .A2(n_89), .B1(n_679), .B2(n_680), .Y(n_687) );
INVxp67_ASAP7_75t_SL g716 ( .A(n_6), .Y(n_716) );
HB1xp67_ASAP7_75t_L g296 ( .A(n_7), .Y(n_296) );
AND2x2_ASAP7_75t_L g387 ( .A(n_7), .B(n_388), .Y(n_387) );
INVx1_ASAP7_75t_L g442 ( .A(n_7), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_7), .B(n_218), .Y(n_449) );
AOI22xp33_ASAP7_75t_L g757 ( .A1(n_8), .A2(n_26), .B1(n_679), .B2(n_758), .Y(n_757) );
AOI22xp33_ASAP7_75t_L g784 ( .A1(n_8), .A2(n_219), .B1(n_708), .B2(n_785), .Y(n_784) );
CKINVDCx5p33_ASAP7_75t_R g828 ( .A(n_9), .Y(n_828) );
INVx1_ASAP7_75t_L g424 ( .A(n_10), .Y(n_424) );
INVxp67_ASAP7_75t_L g1052 ( .A(n_11), .Y(n_1052) );
OAI222xp33_ASAP7_75t_L g1066 ( .A1(n_11), .A2(n_52), .B1(n_270), .B2(n_349), .C1(n_622), .C2(n_1067), .Y(n_1066) );
AOI22xp5_ASAP7_75t_L g1288 ( .A1(n_12), .A2(n_133), .B1(n_1263), .B2(n_1269), .Y(n_1288) );
OAI221xp5_ASAP7_75t_L g884 ( .A1(n_13), .A2(n_463), .B1(n_817), .B2(n_885), .C(n_891), .Y(n_884) );
INVx1_ASAP7_75t_L g907 ( .A(n_13), .Y(n_907) );
INVx1_ASAP7_75t_L g433 ( .A(n_14), .Y(n_433) );
XNOR2x2_ASAP7_75t_L g1153 ( .A(n_15), .B(n_1154), .Y(n_1153) );
OAI211xp5_ASAP7_75t_L g1549 ( .A1(n_16), .A2(n_1550), .B(n_1551), .C(n_1582), .Y(n_1549) );
CKINVDCx5p33_ASAP7_75t_R g1568 ( .A(n_17), .Y(n_1568) );
OAI221xp5_ASAP7_75t_L g517 ( .A1(n_18), .A2(n_30), .B1(n_518), .B2(n_521), .C(n_522), .Y(n_517) );
CKINVDCx5p33_ASAP7_75t_R g578 ( .A(n_18), .Y(n_578) );
AOI221xp5_ASAP7_75t_L g879 ( .A1(n_19), .A2(n_65), .B1(n_438), .B2(n_523), .C(n_880), .Y(n_879) );
INVx1_ASAP7_75t_L g912 ( .A(n_19), .Y(n_912) );
INVx1_ASAP7_75t_L g874 ( .A(n_20), .Y(n_874) );
AOI22xp33_ASAP7_75t_L g909 ( .A1(n_20), .A2(n_68), .B1(n_699), .B2(n_709), .Y(n_909) );
INVx1_ASAP7_75t_L g1486 ( .A(n_21), .Y(n_1486) );
AO22x2_ASAP7_75t_L g916 ( .A1(n_22), .A2(n_917), .B1(n_972), .B2(n_973), .Y(n_916) );
CKINVDCx14_ASAP7_75t_R g972 ( .A(n_22), .Y(n_972) );
AOI22xp33_ASAP7_75t_SL g1210 ( .A1(n_23), .A2(n_249), .B1(n_765), .B2(n_1211), .Y(n_1210) );
AOI221xp5_ASAP7_75t_L g1242 ( .A1(n_23), .A2(n_78), .B1(n_555), .B2(n_634), .C(n_1243), .Y(n_1242) );
CKINVDCx5p33_ASAP7_75t_R g829 ( .A(n_24), .Y(n_829) );
AOI221xp5_ASAP7_75t_L g1109 ( .A1(n_25), .A2(n_47), .B1(n_555), .B2(n_948), .C(n_1110), .Y(n_1109) );
INVx1_ASAP7_75t_L g1142 ( .A(n_25), .Y(n_1142) );
AOI221xp5_ASAP7_75t_L g780 ( .A1(n_26), .A2(n_101), .B1(n_631), .B2(n_781), .C(n_783), .Y(n_780) );
AOI22xp33_ASAP7_75t_L g1212 ( .A1(n_27), .A2(n_78), .B1(n_1213), .B2(n_1215), .Y(n_1212) );
AOI22xp33_ASAP7_75t_L g1244 ( .A1(n_27), .A2(n_249), .B1(n_1077), .B2(n_1245), .Y(n_1244) );
AO221x2_ASAP7_75t_L g1333 ( .A1(n_28), .A2(n_195), .B1(n_1334), .B2(n_1336), .C(n_1338), .Y(n_1333) );
AOI22xp5_ASAP7_75t_L g1502 ( .A1(n_29), .A2(n_247), .B1(n_708), .B2(n_1503), .Y(n_1502) );
OAI22xp5_ASAP7_75t_L g1533 ( .A1(n_29), .A2(n_247), .B1(n_383), .B2(n_466), .Y(n_1533) );
CKINVDCx5p33_ASAP7_75t_R g577 ( .A(n_30), .Y(n_577) );
CKINVDCx5p33_ASAP7_75t_R g892 ( .A(n_31), .Y(n_892) );
INVx1_ASAP7_75t_L g806 ( .A(n_32), .Y(n_806) );
AOI22xp33_ASAP7_75t_L g849 ( .A1(n_32), .A2(n_246), .B1(n_322), .B2(n_850), .Y(n_849) );
INVx2_ASAP7_75t_L g318 ( .A(n_33), .Y(n_318) );
OR2x2_ASAP7_75t_L g477 ( .A(n_33), .B(n_366), .Y(n_477) );
AOI221xp5_ASAP7_75t_L g612 ( .A1(n_34), .A2(n_208), .B1(n_613), .B2(n_614), .C(n_616), .Y(n_612) );
INVx1_ASAP7_75t_L g626 ( .A(n_34), .Y(n_626) );
AO22x1_ASAP7_75t_L g869 ( .A1(n_35), .A2(n_870), .B1(n_914), .B2(n_915), .Y(n_869) );
INVx1_ASAP7_75t_L g915 ( .A(n_35), .Y(n_915) );
INVx1_ASAP7_75t_L g1053 ( .A(n_36), .Y(n_1053) );
INVx1_ASAP7_75t_L g1206 ( .A(n_37), .Y(n_1206) );
OAI221xp5_ASAP7_75t_L g1559 ( .A1(n_38), .A2(n_232), .B1(n_1036), .B2(n_1560), .C(n_1562), .Y(n_1559) );
INVx1_ASAP7_75t_L g1595 ( .A(n_38), .Y(n_1595) );
BUFx2_ASAP7_75t_L g320 ( .A(n_39), .Y(n_320) );
BUFx2_ASAP7_75t_L g354 ( .A(n_39), .Y(n_354) );
INVx1_ASAP7_75t_L g368 ( .A(n_39), .Y(n_368) );
OR2x2_ASAP7_75t_L g520 ( .A(n_39), .B(n_449), .Y(n_520) );
AOI22xp33_ASAP7_75t_SL g763 ( .A1(n_40), .A2(n_170), .B1(n_683), .B2(n_684), .Y(n_763) );
INVxp33_ASAP7_75t_SL g790 ( .A(n_40), .Y(n_790) );
INVx1_ASAP7_75t_L g920 ( .A(n_41), .Y(n_920) );
AOI21xp33_ASAP7_75t_L g962 ( .A1(n_41), .A2(n_699), .B(n_783), .Y(n_962) );
INVx1_ASAP7_75t_L g592 ( .A(n_42), .Y(n_592) );
INVxp33_ASAP7_75t_SL g754 ( .A(n_43), .Y(n_754) );
AOI221xp5_ASAP7_75t_L g773 ( .A1(n_43), .A2(n_230), .B1(n_327), .B2(n_347), .C(n_774), .Y(n_773) );
AOI22xp33_ASAP7_75t_SL g507 ( .A1(n_44), .A2(n_182), .B1(n_450), .B2(n_508), .Y(n_507) );
INVx1_ASAP7_75t_L g558 ( .A(n_44), .Y(n_558) );
CKINVDCx5p33_ASAP7_75t_R g824 ( .A(n_45), .Y(n_824) );
CKINVDCx5p33_ASAP7_75t_R g933 ( .A(n_46), .Y(n_933) );
INVx1_ASAP7_75t_L g1136 ( .A(n_47), .Y(n_1136) );
CKINVDCx5p33_ASAP7_75t_R g1114 ( .A(n_48), .Y(n_1114) );
AOI22xp33_ASAP7_75t_SL g678 ( .A1(n_49), .A2(n_203), .B1(n_679), .B2(n_680), .Y(n_678) );
AOI221xp5_ASAP7_75t_L g717 ( .A1(n_49), .A2(n_261), .B1(n_347), .B2(n_718), .C(n_721), .Y(n_717) );
AOI22xp33_ASAP7_75t_L g513 ( .A1(n_50), .A2(n_98), .B1(n_468), .B2(n_514), .Y(n_513) );
OAI22xp5_ASAP7_75t_L g538 ( .A1(n_50), .A2(n_98), .B1(n_539), .B2(n_543), .Y(n_538) );
INVx1_ASAP7_75t_L g1041 ( .A(n_51), .Y(n_1041) );
INVxp67_ASAP7_75t_L g1050 ( .A(n_52), .Y(n_1050) );
OAI221xp5_ASAP7_75t_L g963 ( .A1(n_53), .A2(n_236), .B1(n_964), .B2(n_965), .C(n_967), .Y(n_963) );
INVx1_ASAP7_75t_L g970 ( .A(n_53), .Y(n_970) );
INVx1_ASAP7_75t_L g890 ( .A(n_54), .Y(n_890) );
AOI22xp33_ASAP7_75t_L g905 ( .A1(n_54), .A2(n_165), .B1(n_323), .B2(n_709), .Y(n_905) );
AOI22xp33_ASAP7_75t_L g1218 ( .A1(n_55), .A2(n_64), .B1(n_1219), .B2(n_1221), .Y(n_1218) );
INVx1_ASAP7_75t_L g1247 ( .A(n_55), .Y(n_1247) );
INVx1_ASAP7_75t_L g602 ( .A(n_56), .Y(n_602) );
OAI22xp5_ASAP7_75t_L g881 ( .A1(n_57), .A2(n_178), .B1(n_835), .B2(n_882), .Y(n_881) );
OAI22xp5_ASAP7_75t_SL g898 ( .A1(n_57), .A2(n_178), .B1(n_359), .B2(n_371), .Y(n_898) );
AOI22xp33_ASAP7_75t_L g1158 ( .A1(n_58), .A2(n_61), .B1(n_614), .B2(n_1159), .Y(n_1158) );
OAI22xp5_ASAP7_75t_L g1200 ( .A1(n_58), .A2(n_77), .B1(n_487), .B2(n_1201), .Y(n_1200) );
CKINVDCx5p33_ASAP7_75t_R g369 ( .A(n_59), .Y(n_369) );
INVx1_ASAP7_75t_L g1347 ( .A(n_60), .Y(n_1347) );
INVxp67_ASAP7_75t_SL g1198 ( .A(n_61), .Y(n_1198) );
INVx1_ASAP7_75t_L g503 ( .A(n_62), .Y(n_503) );
AOI21xp33_ASAP7_75t_L g554 ( .A1(n_62), .A2(n_555), .B(n_556), .Y(n_554) );
AOI22xp33_ASAP7_75t_SL g686 ( .A1(n_63), .A2(n_105), .B1(n_683), .B2(n_684), .Y(n_686) );
INVxp33_ASAP7_75t_SL g730 ( .A(n_63), .Y(n_730) );
INVx1_ASAP7_75t_L g1241 ( .A(n_64), .Y(n_1241) );
OAI22xp5_ASAP7_75t_L g913 ( .A1(n_65), .A2(n_124), .B1(n_479), .B2(n_487), .Y(n_913) );
INVx1_ASAP7_75t_L g1175 ( .A(n_66), .Y(n_1175) );
AOI22xp33_ASAP7_75t_L g1496 ( .A1(n_67), .A2(n_81), .B1(n_328), .B2(n_1497), .Y(n_1496) );
INVxp67_ASAP7_75t_L g1523 ( .A(n_67), .Y(n_1523) );
INVx1_ASAP7_75t_L g875 ( .A(n_68), .Y(n_875) );
AOI22xp33_ASAP7_75t_SL g991 ( .A1(n_69), .A2(n_126), .B1(n_992), .B2(n_993), .Y(n_991) );
AOI221xp5_ASAP7_75t_L g1017 ( .A1(n_69), .A2(n_156), .B1(n_556), .B2(n_1018), .C(n_1020), .Y(n_1017) );
AOI22xp33_ASAP7_75t_L g346 ( .A1(n_70), .A2(n_217), .B1(n_347), .B2(n_348), .Y(n_346) );
OAI22xp33_ASAP7_75t_L g382 ( .A1(n_70), .A2(n_277), .B1(n_383), .B2(n_393), .Y(n_382) );
XNOR2xp5_ASAP7_75t_L g1546 ( .A(n_71), .B(n_1547), .Y(n_1546) );
AO22x2_ASAP7_75t_L g795 ( .A1(n_72), .A2(n_796), .B1(n_797), .B2(n_866), .Y(n_795) );
INVx1_ASAP7_75t_L g866 ( .A(n_72), .Y(n_866) );
CKINVDCx5p33_ASAP7_75t_R g831 ( .A(n_73), .Y(n_831) );
INVx1_ASAP7_75t_L g1557 ( .A(n_74), .Y(n_1557) );
AOI221xp5_ASAP7_75t_L g1601 ( .A1(n_74), .A2(n_151), .B1(n_855), .B2(n_1602), .C(n_1604), .Y(n_1601) );
CKINVDCx5p33_ASAP7_75t_R g376 ( .A(n_75), .Y(n_376) );
INVx1_ASAP7_75t_L g1348 ( .A(n_76), .Y(n_1348) );
AOI221xp5_ASAP7_75t_L g1161 ( .A1(n_77), .A2(n_206), .B1(n_438), .B2(n_1162), .C(n_1164), .Y(n_1161) );
INVxp33_ASAP7_75t_SL g984 ( .A(n_79), .Y(n_984) );
AOI22xp33_ASAP7_75t_SL g1012 ( .A1(n_79), .A2(n_220), .B1(n_323), .B2(n_709), .Y(n_1012) );
OAI22xp5_ASAP7_75t_L g799 ( .A1(n_80), .A2(n_211), .B1(n_800), .B2(n_801), .Y(n_799) );
AOI22xp33_ASAP7_75t_SL g858 ( .A1(n_80), .A2(n_211), .B1(n_859), .B2(n_860), .Y(n_858) );
INVxp67_ASAP7_75t_L g1521 ( .A(n_81), .Y(n_1521) );
AOI221xp5_ASAP7_75t_L g597 ( .A1(n_82), .A2(n_155), .B1(n_426), .B2(n_598), .C(n_599), .Y(n_597) );
AOI22xp33_ASAP7_75t_L g636 ( .A1(n_82), .A2(n_99), .B1(n_637), .B2(n_638), .Y(n_636) );
CKINVDCx5p33_ASAP7_75t_R g822 ( .A(n_83), .Y(n_822) );
INVx1_ASAP7_75t_L g1576 ( .A(n_84), .Y(n_1576) );
OAI22xp5_ASAP7_75t_L g1605 ( .A1(n_84), .A2(n_254), .B1(n_543), .B2(n_546), .Y(n_1605) );
INVxp67_ASAP7_75t_SL g982 ( .A(n_85), .Y(n_982) );
OAI221xp5_ASAP7_75t_L g1008 ( .A1(n_85), .A2(n_228), .B1(n_965), .B2(n_1009), .C(n_1010), .Y(n_1008) );
INVx1_ASAP7_75t_L g1106 ( .A(n_86), .Y(n_1106) );
CKINVDCx5p33_ASAP7_75t_R g506 ( .A(n_87), .Y(n_506) );
AO221x1_ASAP7_75t_L g1298 ( .A1(n_88), .A2(n_144), .B1(n_1263), .B2(n_1269), .C(n_1299), .Y(n_1298) );
INVxp33_ASAP7_75t_L g728 ( .A(n_89), .Y(n_728) );
INVx1_ASAP7_75t_L g601 ( .A(n_90), .Y(n_601) );
AOI221xp5_ASAP7_75t_L g630 ( .A1(n_90), .A2(n_155), .B1(n_631), .B2(n_632), .C(n_634), .Y(n_630) );
INVx1_ASAP7_75t_L g1340 ( .A(n_91), .Y(n_1340) );
AOI221xp5_ASAP7_75t_L g1081 ( .A1(n_92), .A2(n_167), .B1(n_1082), .B2(n_1083), .C(n_1084), .Y(n_1081) );
OAI221xp5_ASAP7_75t_L g1086 ( .A1(n_92), .A2(n_191), .B1(n_1087), .B2(n_1088), .C(n_1090), .Y(n_1086) );
CKINVDCx5p33_ASAP7_75t_R g833 ( .A(n_93), .Y(n_833) );
AO221x1_ASAP7_75t_L g1290 ( .A1(n_94), .A2(n_192), .B1(n_1263), .B2(n_1269), .C(n_1291), .Y(n_1290) );
INVx1_ASAP7_75t_L g1295 ( .A(n_95), .Y(n_1295) );
INVx1_ASAP7_75t_L g317 ( .A(n_96), .Y(n_317) );
INVx1_ASAP7_75t_L g366 ( .A(n_96), .Y(n_366) );
INVx1_ASAP7_75t_L g617 ( .A(n_97), .Y(n_617) );
OAI221xp5_ASAP7_75t_L g621 ( .A1(n_97), .A2(n_208), .B1(n_622), .B2(n_624), .C(n_625), .Y(n_621) );
INVxp67_ASAP7_75t_SL g600 ( .A(n_99), .Y(n_600) );
INVxp67_ASAP7_75t_SL g659 ( .A(n_100), .Y(n_659) );
OAI22xp33_ASAP7_75t_L g700 ( .A1(n_100), .A2(n_235), .B1(n_701), .B2(n_703), .Y(n_700) );
AOI22xp33_ASAP7_75t_SL g760 ( .A1(n_101), .A2(n_219), .B1(n_683), .B2(n_761), .Y(n_760) );
NAND2xp33_ASAP7_75t_SL g1101 ( .A(n_102), .B(n_1102), .Y(n_1101) );
INVx1_ASAP7_75t_L g1125 ( .A(n_102), .Y(n_1125) );
OAI221xp5_ASAP7_75t_L g819 ( .A1(n_103), .A2(n_393), .B1(n_820), .B2(n_825), .C(n_830), .Y(n_819) );
AOI22xp33_ASAP7_75t_SL g854 ( .A1(n_103), .A2(n_142), .B1(n_855), .B2(n_857), .Y(n_854) );
INVx1_ASAP7_75t_L g1493 ( .A(n_104), .Y(n_1493) );
INVxp67_ASAP7_75t_SL g697 ( .A(n_105), .Y(n_697) );
OAI22xp33_ASAP7_75t_L g532 ( .A1(n_106), .A2(n_171), .B1(n_533), .B2(n_536), .Y(n_532) );
AOI22xp33_ASAP7_75t_L g566 ( .A1(n_106), .A2(n_231), .B1(n_324), .B2(n_562), .Y(n_566) );
INVx1_ASAP7_75t_L g609 ( .A(n_107), .Y(n_609) );
AOI221xp5_ASAP7_75t_L g641 ( .A1(n_107), .A2(n_164), .B1(n_570), .B2(n_642), .C(n_643), .Y(n_641) );
OAI22xp5_ASAP7_75t_L g525 ( .A1(n_108), .A2(n_231), .B1(n_526), .B2(n_529), .Y(n_525) );
INVx1_ASAP7_75t_L g564 ( .A(n_108), .Y(n_564) );
XNOR2xp5_ASAP7_75t_L g1031 ( .A(n_109), .B(n_1032), .Y(n_1031) );
INVx1_ASAP7_75t_L g1177 ( .A(n_110), .Y(n_1177) );
AOI221xp5_ASAP7_75t_L g1183 ( .A1(n_110), .A2(n_273), .B1(n_852), .B2(n_1184), .C(n_1186), .Y(n_1183) );
INVxp33_ASAP7_75t_SL g988 ( .A(n_111), .Y(n_988) );
AOI21xp33_ASAP7_75t_L g1013 ( .A1(n_111), .A2(n_778), .B(n_1014), .Y(n_1013) );
OAI22xp5_ASAP7_75t_L g738 ( .A1(n_112), .A2(n_739), .B1(n_740), .B2(n_794), .Y(n_738) );
INVx1_ASAP7_75t_L g794 ( .A(n_112), .Y(n_794) );
INVxp67_ASAP7_75t_L g1039 ( .A(n_113), .Y(n_1039) );
AOI221xp5_ASAP7_75t_L g1070 ( .A1(n_113), .A2(n_187), .B1(n_555), .B2(n_948), .C(n_1071), .Y(n_1070) );
OAI21xp33_ASAP7_75t_L g583 ( .A1(n_114), .A2(n_584), .B(n_619), .Y(n_583) );
INVx1_ASAP7_75t_L g653 ( .A(n_114), .Y(n_653) );
CKINVDCx20_ASAP7_75t_R g1094 ( .A(n_115), .Y(n_1094) );
INVx1_ASAP7_75t_L g618 ( .A(n_116), .Y(n_618) );
CKINVDCx5p33_ASAP7_75t_R g768 ( .A(n_117), .Y(n_768) );
AOI22xp33_ASAP7_75t_L g1262 ( .A1(n_118), .A2(n_242), .B1(n_1263), .B2(n_1269), .Y(n_1262) );
INVx1_ASAP7_75t_L g1581 ( .A(n_119), .Y(n_1581) );
OAI211xp5_ASAP7_75t_SL g1583 ( .A1(n_119), .A2(n_1584), .B(n_1585), .C(n_1591), .Y(n_1583) );
INVx1_ASAP7_75t_L g753 ( .A(n_120), .Y(n_753) );
AOI22xp33_ASAP7_75t_SL g1500 ( .A1(n_121), .A2(n_176), .B1(n_1499), .B2(n_1501), .Y(n_1500) );
OAI221xp5_ASAP7_75t_L g1519 ( .A1(n_121), .A2(n_463), .B1(n_1179), .B2(n_1520), .C(n_1527), .Y(n_1519) );
AOI22xp33_ASAP7_75t_L g1000 ( .A1(n_122), .A2(n_185), .B1(n_680), .B2(n_1001), .Y(n_1000) );
INVxp33_ASAP7_75t_SL g1024 ( .A(n_122), .Y(n_1024) );
CKINVDCx5p33_ASAP7_75t_R g1117 ( .A(n_123), .Y(n_1117) );
AOI22xp33_ASAP7_75t_L g877 ( .A1(n_124), .A2(n_143), .B1(n_613), .B2(n_878), .Y(n_877) );
AOI22xp33_ASAP7_75t_SL g764 ( .A1(n_125), .A2(n_147), .B1(n_679), .B2(n_765), .Y(n_764) );
INVxp33_ASAP7_75t_L g789 ( .A(n_125), .Y(n_789) );
AOI22xp33_ASAP7_75t_L g1021 ( .A1(n_126), .A2(n_129), .B1(n_327), .B2(n_1022), .Y(n_1021) );
INVxp33_ASAP7_75t_SL g1489 ( .A(n_127), .Y(n_1489) );
AOI221xp5_ASAP7_75t_L g1514 ( .A1(n_127), .A2(n_172), .B1(n_438), .B2(n_765), .C(n_1515), .Y(n_1514) );
INVx1_ASAP7_75t_L g1301 ( .A(n_128), .Y(n_1301) );
AOI22xp33_ASAP7_75t_L g995 ( .A1(n_129), .A2(n_156), .B1(n_996), .B2(n_997), .Y(n_995) );
INVx1_ASAP7_75t_L g815 ( .A(n_130), .Y(n_815) );
AOI22xp33_ASAP7_75t_L g851 ( .A1(n_130), .A2(n_154), .B1(n_852), .B2(n_853), .Y(n_851) );
INVx1_ASAP7_75t_L g288 ( .A(n_131), .Y(n_288) );
INVx1_ASAP7_75t_L g1026 ( .A(n_132), .Y(n_1026) );
INVx1_ASAP7_75t_L g1118 ( .A(n_134), .Y(n_1118) );
AOI22xp33_ASAP7_75t_L g1498 ( .A1(n_135), .A2(n_200), .B1(n_785), .B2(n_1499), .Y(n_1498) );
INVxp67_ASAP7_75t_SL g1532 ( .A(n_135), .Y(n_1532) );
CKINVDCx5p33_ASAP7_75t_R g930 ( .A(n_136), .Y(n_930) );
AOI22xp33_ASAP7_75t_L g999 ( .A1(n_137), .A2(n_196), .B1(n_996), .B2(n_997), .Y(n_999) );
INVxp67_ASAP7_75t_SL g1007 ( .A(n_137), .Y(n_1007) );
AOI22xp33_ASAP7_75t_L g1216 ( .A1(n_138), .A2(n_209), .B1(n_1159), .B2(n_1217), .Y(n_1216) );
INVx1_ASAP7_75t_L g1248 ( .A(n_138), .Y(n_1248) );
AOI22xp5_ASAP7_75t_L g1283 ( .A1(n_139), .A2(n_222), .B1(n_1271), .B2(n_1277), .Y(n_1283) );
INVxp67_ASAP7_75t_SL g745 ( .A(n_140), .Y(n_745) );
OAI22xp5_ASAP7_75t_L g772 ( .A1(n_140), .A2(n_281), .B1(n_701), .B2(n_703), .Y(n_772) );
OAI221xp5_ASAP7_75t_SL g605 ( .A1(n_141), .A2(n_253), .B1(n_606), .B2(n_607), .C(n_608), .Y(n_605) );
AOI22xp33_ASAP7_75t_L g644 ( .A1(n_141), .A2(n_253), .B1(n_323), .B2(n_645), .Y(n_644) );
OAI221xp5_ASAP7_75t_L g802 ( .A1(n_142), .A2(n_463), .B1(n_803), .B2(n_809), .C(n_817), .Y(n_802) );
INVx1_ASAP7_75t_L g911 ( .A(n_143), .Y(n_911) );
INVx1_ASAP7_75t_L g1300 ( .A(n_145), .Y(n_1300) );
AOI22xp33_ASAP7_75t_SL g1099 ( .A1(n_146), .A2(n_238), .B1(n_328), .B2(n_1100), .Y(n_1099) );
INVx1_ASAP7_75t_L g1128 ( .A(n_146), .Y(n_1128) );
INVxp67_ASAP7_75t_SL g787 ( .A(n_147), .Y(n_787) );
XOR2xp5_ASAP7_75t_L g493 ( .A(n_148), .B(n_494), .Y(n_493) );
AOI22xp5_ASAP7_75t_L g1270 ( .A1(n_149), .A2(n_280), .B1(n_1271), .B2(n_1277), .Y(n_1270) );
AOI22xp5_ASAP7_75t_L g1284 ( .A1(n_150), .A2(n_199), .B1(n_1263), .B2(n_1269), .Y(n_1284) );
INVx1_ASAP7_75t_L g1555 ( .A(n_151), .Y(n_1555) );
INVx1_ASAP7_75t_L g986 ( .A(n_152), .Y(n_986) );
INVx1_ASAP7_75t_L g1181 ( .A(n_153), .Y(n_1181) );
INVx1_ASAP7_75t_L g812 ( .A(n_154), .Y(n_812) );
INVx1_ASAP7_75t_L g751 ( .A(n_157), .Y(n_751) );
OAI222xp33_ASAP7_75t_L g1034 ( .A1(n_158), .A2(n_186), .B1(n_272), .B2(n_536), .C1(n_1035), .C2(n_1036), .Y(n_1034) );
INVx1_ASAP7_75t_L g1060 ( .A(n_158), .Y(n_1060) );
CKINVDCx5p33_ASAP7_75t_R g1224 ( .A(n_159), .Y(n_1224) );
CKINVDCx5p33_ASAP7_75t_R g936 ( .A(n_160), .Y(n_936) );
INVx1_ASAP7_75t_L g1251 ( .A(n_161), .Y(n_1251) );
CKINVDCx5p33_ASAP7_75t_R g1108 ( .A(n_162), .Y(n_1108) );
AOI22xp33_ASAP7_75t_L g321 ( .A1(n_163), .A2(n_263), .B1(n_322), .B2(n_327), .Y(n_321) );
INVx1_ASAP7_75t_L g406 ( .A(n_163), .Y(n_406) );
INVx1_ASAP7_75t_L g611 ( .A(n_164), .Y(n_611) );
INVx1_ASAP7_75t_L g888 ( .A(n_165), .Y(n_888) );
INVx1_ASAP7_75t_L g1223 ( .A(n_166), .Y(n_1223) );
AOI22xp33_ASAP7_75t_L g1237 ( .A1(n_166), .A2(n_245), .B1(n_324), .B2(n_350), .Y(n_1237) );
OAI332xp33_ASAP7_75t_L g1037 ( .A1(n_167), .A2(n_509), .A3(n_941), .B1(n_1038), .B2(n_1042), .B3(n_1045), .C1(n_1051), .C2(n_1056), .Y(n_1037) );
INVx1_ASAP7_75t_L g921 ( .A(n_168), .Y(n_921) );
AOI22xp33_ASAP7_75t_SL g961 ( .A1(n_168), .A2(n_214), .B1(n_709), .B2(n_786), .Y(n_961) );
OAI22xp5_ASAP7_75t_L g1166 ( .A1(n_169), .A2(n_193), .B1(n_835), .B2(n_882), .Y(n_1166) );
OAI221xp5_ASAP7_75t_L g1194 ( .A1(n_169), .A2(n_193), .B1(n_865), .B2(n_1195), .C(n_1196), .Y(n_1194) );
INVxp67_ASAP7_75t_SL g771 ( .A(n_170), .Y(n_771) );
INVx1_ASAP7_75t_L g572 ( .A(n_171), .Y(n_572) );
INVxp33_ASAP7_75t_SL g1487 ( .A(n_172), .Y(n_1487) );
CKINVDCx5p33_ASAP7_75t_R g694 ( .A(n_173), .Y(n_694) );
CKINVDCx5p33_ASAP7_75t_R g436 ( .A(n_174), .Y(n_436) );
CKINVDCx5p33_ASAP7_75t_R g837 ( .A(n_175), .Y(n_837) );
OAI211xp5_ASAP7_75t_SL g1509 ( .A1(n_176), .A2(n_393), .B(n_1510), .C(n_1516), .Y(n_1509) );
XNOR2xp5_ASAP7_75t_L g1481 ( .A(n_177), .B(n_1482), .Y(n_1481) );
AOI22xp33_ASAP7_75t_L g1540 ( .A1(n_177), .A2(n_1541), .B1(n_1545), .B2(n_1607), .Y(n_1540) );
INVxp67_ASAP7_75t_SL g1571 ( .A(n_179), .Y(n_1571) );
AOI221xp5_ASAP7_75t_L g1589 ( .A1(n_179), .A2(n_212), .B1(n_631), .B2(n_781), .C(n_1590), .Y(n_1589) );
XOR2x2_ASAP7_75t_L g654 ( .A(n_180), .B(n_655), .Y(n_654) );
AOI22xp33_ASAP7_75t_L g345 ( .A1(n_181), .A2(n_277), .B1(n_334), .B2(n_340), .Y(n_345) );
OAI22xp33_ASAP7_75t_L g462 ( .A1(n_181), .A2(n_217), .B1(n_463), .B2(n_466), .Y(n_462) );
INVx1_ASAP7_75t_L g553 ( .A(n_182), .Y(n_553) );
OAI22xp5_ASAP7_75t_L g939 ( .A1(n_183), .A2(n_205), .B1(n_940), .B2(n_941), .Y(n_939) );
INVx1_ASAP7_75t_L g952 ( .A(n_183), .Y(n_952) );
OAI22xp5_ASAP7_75t_L g942 ( .A1(n_184), .A2(n_233), .B1(n_533), .B2(n_536), .Y(n_942) );
AOI22xp33_ASAP7_75t_SL g955 ( .A1(n_184), .A2(n_205), .B1(n_699), .B2(n_709), .Y(n_955) );
INVxp67_ASAP7_75t_SL g1016 ( .A(n_185), .Y(n_1016) );
INVx1_ASAP7_75t_L g1075 ( .A(n_186), .Y(n_1075) );
INVx1_ASAP7_75t_L g1043 ( .A(n_187), .Y(n_1043) );
CKINVDCx5p33_ASAP7_75t_R g931 ( .A(n_188), .Y(n_931) );
HB1xp67_ASAP7_75t_L g290 ( .A(n_189), .Y(n_290) );
AND3x2_ASAP7_75t_L g1267 ( .A(n_189), .B(n_288), .C(n_1268), .Y(n_1267) );
NAND2xp5_ASAP7_75t_L g1276 ( .A(n_189), .B(n_288), .Y(n_1276) );
OA332x1_ASAP7_75t_L g918 ( .A1(n_190), .A2(n_497), .A3(n_509), .B1(n_919), .B2(n_924), .B3(n_928), .C1(n_932), .C2(n_937), .Y(n_918) );
AOI21xp5_ASAP7_75t_L g956 ( .A1(n_190), .A2(n_957), .B(n_958), .Y(n_956) );
INVx1_ASAP7_75t_L g1080 ( .A(n_191), .Y(n_1080) );
INVx2_ASAP7_75t_L g301 ( .A(n_194), .Y(n_301) );
INVxp33_ASAP7_75t_SL g1025 ( .A(n_196), .Y(n_1025) );
CKINVDCx5p33_ASAP7_75t_R g670 ( .A(n_197), .Y(n_670) );
OAI211xp5_ASAP7_75t_L g872 ( .A1(n_198), .A2(n_393), .B(n_873), .C(n_876), .Y(n_872) );
INVx1_ASAP7_75t_L g908 ( .A(n_198), .Y(n_908) );
INVxp67_ASAP7_75t_SL g1529 ( .A(n_200), .Y(n_1529) );
INVx1_ASAP7_75t_L g588 ( .A(n_201), .Y(n_588) );
INVxp33_ASAP7_75t_SL g672 ( .A(n_202), .Y(n_672) );
AOI221xp5_ASAP7_75t_L g705 ( .A1(n_202), .A2(n_248), .B1(n_706), .B2(n_708), .C(n_710), .Y(n_705) );
AOI22xp33_ASAP7_75t_L g723 ( .A1(n_203), .A2(n_229), .B1(n_645), .B2(n_724), .Y(n_723) );
INVx1_ASAP7_75t_L g1174 ( .A(n_204), .Y(n_1174) );
INVxp67_ASAP7_75t_SL g1199 ( .A(n_206), .Y(n_1199) );
INVx1_ASAP7_75t_L g1268 ( .A(n_207), .Y(n_1268) );
INVx1_ASAP7_75t_L g1233 ( .A(n_209), .Y(n_1233) );
AOI22xp33_ASAP7_75t_L g515 ( .A1(n_210), .A2(n_271), .B1(n_450), .B2(n_508), .Y(n_515) );
OAI22xp5_ASAP7_75t_L g545 ( .A1(n_210), .A2(n_271), .B1(n_546), .B2(n_548), .Y(n_545) );
INVxp67_ASAP7_75t_SL g1565 ( .A(n_212), .Y(n_1565) );
AOI22xp33_ASAP7_75t_L g333 ( .A1(n_213), .A2(n_257), .B1(n_334), .B2(n_340), .Y(n_333) );
INVx1_ASAP7_75t_L g418 ( .A(n_213), .Y(n_418) );
INVx1_ASAP7_75t_L g925 ( .A(n_214), .Y(n_925) );
CKINVDCx5p33_ASAP7_75t_R g1249 ( .A(n_215), .Y(n_1249) );
OAI211xp5_ASAP7_75t_L g1156 ( .A1(n_216), .A2(n_393), .B(n_1157), .C(n_1167), .Y(n_1156) );
AOI221xp5_ASAP7_75t_L g1188 ( .A1(n_216), .A2(n_224), .B1(n_334), .B2(n_718), .C(n_1189), .Y(n_1188) );
INVx1_ASAP7_75t_L g303 ( .A(n_218), .Y(n_303) );
INVx2_ASAP7_75t_L g388 ( .A(n_218), .Y(n_388) );
INVxp33_ASAP7_75t_SL g989 ( .A(n_220), .Y(n_989) );
INVx1_ASAP7_75t_L g1168 ( .A(n_221), .Y(n_1168) );
AOI22xp5_ASAP7_75t_L g1287 ( .A1(n_223), .A2(n_237), .B1(n_1271), .B2(n_1277), .Y(n_1287) );
OAI221xp5_ASAP7_75t_L g1170 ( .A1(n_224), .A2(n_463), .B1(n_1171), .B2(n_1176), .C(n_1179), .Y(n_1170) );
INVx1_ASAP7_75t_L g896 ( .A(n_225), .Y(n_896) );
INVx1_ASAP7_75t_L g1292 ( .A(n_226), .Y(n_1292) );
INVx1_ASAP7_75t_L g1226 ( .A(n_227), .Y(n_1226) );
AOI21xp33_ASAP7_75t_L g1238 ( .A1(n_227), .A2(n_570), .B(n_1014), .Y(n_1238) );
INVxp67_ASAP7_75t_SL g981 ( .A(n_228), .Y(n_981) );
AOI22xp33_ASAP7_75t_SL g682 ( .A1(n_229), .A2(n_261), .B1(n_683), .B2(n_684), .Y(n_682) );
INVxp33_ASAP7_75t_SL g749 ( .A(n_230), .Y(n_749) );
INVx1_ASAP7_75t_L g1597 ( .A(n_232), .Y(n_1597) );
INVx1_ASAP7_75t_L g968 ( .A(n_233), .Y(n_968) );
INVx1_ASAP7_75t_L g453 ( .A(n_234), .Y(n_453) );
INVxp67_ASAP7_75t_SL g662 ( .A(n_235), .Y(n_662) );
INVx1_ASAP7_75t_L g971 ( .A(n_236), .Y(n_971) );
XOR2xp5_ASAP7_75t_L g309 ( .A(n_237), .B(n_310), .Y(n_309) );
INVx1_ASAP7_75t_L g1123 ( .A(n_238), .Y(n_1123) );
CKINVDCx5p33_ASAP7_75t_R g1115 ( .A(n_239), .Y(n_1115) );
INVx1_ASAP7_75t_L g667 ( .A(n_240), .Y(n_667) );
INVx1_ASAP7_75t_L g429 ( .A(n_241), .Y(n_429) );
INVx1_ASAP7_75t_L g1490 ( .A(n_243), .Y(n_1490) );
INVx1_ASAP7_75t_L g1570 ( .A(n_244), .Y(n_1570) );
INVx1_ASAP7_75t_L g1227 ( .A(n_245), .Y(n_1227) );
INVx1_ASAP7_75t_L g808 ( .A(n_246), .Y(n_808) );
INVxp33_ASAP7_75t_SL g664 ( .A(n_248), .Y(n_664) );
INVx1_ASAP7_75t_L g1266 ( .A(n_250), .Y(n_1266) );
NAND2xp5_ASAP7_75t_L g1279 ( .A(n_250), .B(n_1274), .Y(n_1279) );
INVx1_ASAP7_75t_L g1063 ( .A(n_251), .Y(n_1063) );
INVx1_ASAP7_75t_L g1573 ( .A(n_252), .Y(n_1573) );
OAI211xp5_ASAP7_75t_L g1592 ( .A1(n_252), .A2(n_1593), .B(n_1594), .C(n_1598), .Y(n_1592) );
INVx1_ASAP7_75t_L g1578 ( .A(n_254), .Y(n_1578) );
INVx1_ASAP7_75t_L g1044 ( .A(n_255), .Y(n_1044) );
INVx1_ASAP7_75t_L g1494 ( .A(n_256), .Y(n_1494) );
INVx1_ASAP7_75t_L g414 ( .A(n_257), .Y(n_414) );
AO22x1_ASAP7_75t_L g1319 ( .A1(n_258), .A2(n_267), .B1(n_1269), .B2(n_1320), .Y(n_1319) );
CKINVDCx5p33_ASAP7_75t_R g893 ( .A(n_259), .Y(n_893) );
INVx2_ASAP7_75t_L g300 ( .A(n_260), .Y(n_300) );
AO22x1_ASAP7_75t_L g1321 ( .A1(n_262), .A2(n_274), .B1(n_1271), .B2(n_1277), .Y(n_1321) );
INVx1_ASAP7_75t_L g400 ( .A(n_263), .Y(n_400) );
AOI21xp33_ASAP7_75t_L g1104 ( .A1(n_264), .A2(n_335), .B(n_570), .Y(n_1104) );
INVx1_ASAP7_75t_L g1127 ( .A(n_264), .Y(n_1127) );
CKINVDCx5p33_ASAP7_75t_R g926 ( .A(n_265), .Y(n_926) );
CKINVDCx5p33_ASAP7_75t_R g1507 ( .A(n_266), .Y(n_1507) );
CKINVDCx5p33_ASAP7_75t_R g1554 ( .A(n_268), .Y(n_1554) );
INVx1_ASAP7_75t_L g1169 ( .A(n_269), .Y(n_1169) );
INVxp67_ASAP7_75t_L g1046 ( .A(n_270), .Y(n_1046) );
INVx1_ASAP7_75t_L g1064 ( .A(n_272), .Y(n_1064) );
AOI21xp33_ASAP7_75t_L g1178 ( .A1(n_273), .A2(n_510), .B(n_1162), .Y(n_1178) );
BUFx3_ASAP7_75t_L g326 ( .A(n_275), .Y(n_326) );
INVx1_ASAP7_75t_L g332 ( .A(n_275), .Y(n_332) );
INVx1_ASAP7_75t_L g325 ( .A(n_276), .Y(n_325) );
BUFx3_ASAP7_75t_L g331 ( .A(n_276), .Y(n_331) );
INVx1_ASAP7_75t_L g1004 ( .A(n_278), .Y(n_1004) );
INVx1_ASAP7_75t_L g1138 ( .A(n_279), .Y(n_1138) );
INVxp67_ASAP7_75t_SL g746 ( .A(n_281), .Y(n_746) );
AOI21xp5_ASAP7_75t_L g282 ( .A1(n_283), .A2(n_304), .B(n_1254), .Y(n_282) );
BUFx12f_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
BUFx3_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
AND2x4_ASAP7_75t_L g285 ( .A(n_286), .B(n_291), .Y(n_285) );
AND2x4_ASAP7_75t_L g1539 ( .A(n_286), .B(n_292), .Y(n_1539) );
NOR2xp33_ASAP7_75t_SL g286 ( .A(n_287), .B(n_289), .Y(n_286) );
INVx1_ASAP7_75t_SL g1544 ( .A(n_287), .Y(n_1544) );
NAND2xp5_ASAP7_75t_L g1614 ( .A(n_287), .B(n_289), .Y(n_1614) );
HB1xp67_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
AND2x2_ASAP7_75t_L g1543 ( .A(n_289), .B(n_1544), .Y(n_1543) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
NOR2xp33_ASAP7_75t_L g292 ( .A(n_293), .B(n_297), .Y(n_292) );
INVxp67_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
HB1xp67_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
AND2x2_ASAP7_75t_L g421 ( .A(n_295), .B(n_303), .Y(n_421) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
OR2x2_ASAP7_75t_L g510 ( .A(n_296), .B(n_511), .Y(n_510) );
OR2x6_ASAP7_75t_L g297 ( .A(n_298), .B(n_302), .Y(n_297) );
BUFx2_ASAP7_75t_L g417 ( .A(n_298), .Y(n_417) );
INVx1_ASAP7_75t_L g435 ( .A(n_298), .Y(n_435) );
OR2x2_ASAP7_75t_L g536 ( .A(n_298), .B(n_520), .Y(n_536) );
OAI22xp33_ASAP7_75t_L g599 ( .A1(n_298), .A2(n_431), .B1(n_600), .B2(n_601), .Y(n_599) );
OAI22xp33_ASAP7_75t_L g616 ( .A1(n_298), .A2(n_431), .B1(n_617), .B2(n_618), .Y(n_616) );
INVx2_ASAP7_75t_SL g814 ( .A(n_298), .Y(n_814) );
BUFx6f_ASAP7_75t_L g929 ( .A(n_298), .Y(n_929) );
INVx2_ASAP7_75t_SL g1531 ( .A(n_298), .Y(n_1531) );
BUFx6f_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_300), .B(n_301), .Y(n_299) );
AND2x4_ASAP7_75t_L g391 ( .A(n_300), .B(n_392), .Y(n_391) );
INVx1_ASAP7_75t_L g397 ( .A(n_300), .Y(n_397) );
INVx2_ASAP7_75t_L g405 ( .A(n_300), .Y(n_405) );
INVx1_ASAP7_75t_L g413 ( .A(n_300), .Y(n_413) );
AND2x2_ASAP7_75t_L g452 ( .A(n_300), .B(n_301), .Y(n_452) );
INVx2_ASAP7_75t_L g392 ( .A(n_301), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_301), .B(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g412 ( .A(n_301), .Y(n_412) );
INVx1_ASAP7_75t_L g459 ( .A(n_301), .Y(n_459) );
INVx1_ASAP7_75t_L g470 ( .A(n_301), .Y(n_470) );
INVx2_ASAP7_75t_SL g302 ( .A(n_303), .Y(n_302) );
XNOR2xp5_ASAP7_75t_L g304 ( .A(n_305), .B(n_1027), .Y(n_304) );
XOR2xp5_ASAP7_75t_L g305 ( .A(n_306), .B(n_976), .Y(n_305) );
XNOR2x2_ASAP7_75t_L g306 ( .A(n_307), .B(n_736), .Y(n_306) );
AO22x2_ASAP7_75t_L g307 ( .A1(n_308), .A2(n_654), .B1(n_734), .B2(n_735), .Y(n_307) );
INVx1_ASAP7_75t_L g734 ( .A(n_308), .Y(n_734) );
XNOR2xp5_ASAP7_75t_L g308 ( .A(n_309), .B(n_492), .Y(n_308) );
NAND4xp75_ASAP7_75t_L g310 ( .A(n_311), .B(n_381), .C(n_473), .D(n_482), .Y(n_310) );
AND2x2_ASAP7_75t_SL g311 ( .A(n_312), .B(n_357), .Y(n_311) );
AOI33xp33_ASAP7_75t_L g312 ( .A1(n_313), .A2(n_321), .A3(n_333), .B1(n_345), .B2(n_346), .B3(n_351), .Y(n_312) );
AOI33xp33_ASAP7_75t_L g1495 ( .A1(n_313), .A2(n_1496), .A3(n_1498), .B1(n_1500), .B2(n_1502), .B3(n_1505), .Y(n_1495) );
CKINVDCx5p33_ASAP7_75t_R g313 ( .A(n_314), .Y(n_313) );
CKINVDCx5p33_ASAP7_75t_R g848 ( .A(n_314), .Y(n_848) );
INVx2_ASAP7_75t_L g1187 ( .A(n_314), .Y(n_1187) );
OR2x6_ASAP7_75t_L g314 ( .A(n_315), .B(n_319), .Y(n_314) );
INVx1_ASAP7_75t_L g1111 ( .A(n_315), .Y(n_1111) );
INVx2_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
INVx2_ASAP7_75t_SL g556 ( .A(n_316), .Y(n_556) );
BUFx3_ASAP7_75t_L g635 ( .A(n_316), .Y(n_635) );
INVx1_ASAP7_75t_L g783 ( .A(n_316), .Y(n_783) );
INVx1_ASAP7_75t_L g901 ( .A(n_316), .Y(n_901) );
AND2x2_ASAP7_75t_L g316 ( .A(n_317), .B(n_318), .Y(n_316) );
AND2x4_ASAP7_75t_L g355 ( .A(n_317), .B(n_356), .Y(n_355) );
INVx2_ASAP7_75t_L g356 ( .A(n_318), .Y(n_356) );
AND2x2_ASAP7_75t_L g516 ( .A(n_319), .B(n_439), .Y(n_516) );
AND2x4_ASAP7_75t_L g596 ( .A(n_319), .B(n_421), .Y(n_596) );
INVx2_ASAP7_75t_L g649 ( .A(n_319), .Y(n_649) );
AND2x4_ASAP7_75t_L g677 ( .A(n_319), .B(n_421), .Y(n_677) );
BUFx2_ASAP7_75t_L g793 ( .A(n_319), .Y(n_793) );
OR2x2_ASAP7_75t_L g900 ( .A(n_319), .B(n_901), .Y(n_900) );
INVx2_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
BUFx2_ASAP7_75t_L g472 ( .A(n_320), .Y(n_472) );
OR2x6_ASAP7_75t_L g509 ( .A(n_320), .B(n_510), .Y(n_509) );
BUFx2_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
BUFx3_ASAP7_75t_L g347 ( .A(n_323), .Y(n_347) );
INVx1_ASAP7_75t_L g707 ( .A(n_323), .Y(n_707) );
BUFx6f_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
INVx2_ASAP7_75t_SL g485 ( .A(n_324), .Y(n_485) );
BUFx6f_ASAP7_75t_L g541 ( .A(n_324), .Y(n_541) );
BUFx6f_ASAP7_75t_L g555 ( .A(n_324), .Y(n_555) );
BUFx6f_ASAP7_75t_L g699 ( .A(n_324), .Y(n_699) );
BUFx3_ASAP7_75t_L g1100 ( .A(n_324), .Y(n_1100) );
HB1xp67_ASAP7_75t_L g1600 ( .A(n_324), .Y(n_1600) );
AND2x4_ASAP7_75t_L g324 ( .A(n_325), .B(n_326), .Y(n_324) );
INVx1_ASAP7_75t_L g491 ( .A(n_325), .Y(n_491) );
INVx2_ASAP7_75t_L g338 ( .A(n_326), .Y(n_338) );
AND2x2_ASAP7_75t_L g344 ( .A(n_326), .B(n_331), .Y(n_344) );
BUFx2_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
INVx2_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
OR2x6_ASAP7_75t_L g479 ( .A(n_329), .B(n_476), .Y(n_479) );
OR2x2_ASAP7_75t_L g1201 ( .A(n_329), .B(n_476), .Y(n_1201) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
BUFx6f_ASAP7_75t_L g350 ( .A(n_330), .Y(n_350) );
INVx2_ASAP7_75t_L g544 ( .A(n_330), .Y(n_544) );
BUFx6f_ASAP7_75t_L g709 ( .A(n_330), .Y(n_709) );
AND2x4_ASAP7_75t_L g330 ( .A(n_331), .B(n_332), .Y(n_330) );
INVx2_ASAP7_75t_L g339 ( .A(n_331), .Y(n_339) );
INVx1_ASAP7_75t_L g490 ( .A(n_332), .Y(n_490) );
BUFx2_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
AND2x2_ASAP7_75t_L g474 ( .A(n_335), .B(n_475), .Y(n_474) );
A2O1A1Ixp33_ASAP7_75t_L g571 ( .A1(n_335), .A2(n_572), .B(n_573), .C(n_579), .Y(n_571) );
INVx2_ASAP7_75t_SL g335 ( .A(n_336), .Y(n_335) );
INVx1_ASAP7_75t_L g724 ( .A(n_336), .Y(n_724) );
INVx1_ASAP7_75t_L g957 ( .A(n_336), .Y(n_957) );
INVx2_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
AND2x2_ASAP7_75t_L g481 ( .A(n_337), .B(n_364), .Y(n_481) );
INVx6_ASAP7_75t_L g569 ( .A(n_337), .Y(n_569) );
BUFx2_ASAP7_75t_L g1245 ( .A(n_337), .Y(n_1245) );
AND2x4_ASAP7_75t_L g337 ( .A(n_338), .B(n_339), .Y(n_337) );
INVx1_ASAP7_75t_L g362 ( .A(n_338), .Y(n_362) );
INVx1_ASAP7_75t_L g374 ( .A(n_339), .Y(n_374) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
AND2x4_ASAP7_75t_L g725 ( .A(n_342), .B(n_726), .Y(n_725) );
INVx1_ASAP7_75t_L g1185 ( .A(n_342), .Y(n_1185) );
BUFx6f_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
INVx1_ASAP7_75t_L g379 ( .A(n_343), .Y(n_379) );
BUFx6f_ASAP7_75t_L g643 ( .A(n_343), .Y(n_643) );
INVx2_ASAP7_75t_L g1103 ( .A(n_343), .Y(n_1103) );
BUFx6f_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
BUFx6f_ASAP7_75t_L g550 ( .A(n_344), .Y(n_550) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
INVx2_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx1_ASAP7_75t_L g624 ( .A(n_350), .Y(n_624) );
BUFx6f_ASAP7_75t_L g645 ( .A(n_350), .Y(n_645) );
BUFx6f_ASAP7_75t_L g946 ( .A(n_350), .Y(n_946) );
INVx1_ASAP7_75t_L g1069 ( .A(n_350), .Y(n_1069) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
OAI22xp5_ASAP7_75t_SL g899 ( .A1(n_352), .A2(n_900), .B1(n_902), .B2(n_906), .Y(n_899) );
INVx4_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
BUFx4f_ASAP7_75t_L g862 ( .A(n_353), .Y(n_862) );
AOI221xp5_ASAP7_75t_L g1182 ( .A1(n_353), .A2(n_1183), .B1(n_1187), .B2(n_1188), .C(n_1194), .Y(n_1182) );
BUFx4f_ASAP7_75t_L g1505 ( .A(n_353), .Y(n_1505) );
AND2x4_ASAP7_75t_L g353 ( .A(n_354), .B(n_355), .Y(n_353) );
AND2x4_ASAP7_75t_L g480 ( .A(n_354), .B(n_481), .Y(n_480) );
CKINVDCx5p33_ASAP7_75t_R g570 ( .A(n_355), .Y(n_570) );
HB1xp67_ASAP7_75t_L g713 ( .A(n_355), .Y(n_713) );
INVx2_ASAP7_75t_L g778 ( .A(n_355), .Y(n_778) );
INVx2_ASAP7_75t_SL g958 ( .A(n_355), .Y(n_958) );
INVx1_ASAP7_75t_L g1084 ( .A(n_355), .Y(n_1084) );
AND2x4_ASAP7_75t_L g364 ( .A(n_356), .B(n_365), .Y(n_364) );
AOI221xp5_ASAP7_75t_L g357 ( .A1(n_358), .A2(n_369), .B1(n_370), .B2(n_376), .C(n_377), .Y(n_357) );
AOI22xp5_ASAP7_75t_L g845 ( .A1(n_358), .A2(n_831), .B1(n_833), .B2(n_846), .Y(n_845) );
AOI22xp33_ASAP7_75t_L g1492 ( .A1(n_358), .A2(n_846), .B1(n_1493), .B2(n_1494), .Y(n_1492) );
INVx2_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
OR2x6_ASAP7_75t_L g359 ( .A(n_360), .B(n_363), .Y(n_359) );
OR2x2_ASAP7_75t_L g703 ( .A(n_360), .B(n_704), .Y(n_703) );
OR2x2_ASAP7_75t_L g1196 ( .A(n_360), .B(n_363), .Y(n_1196) );
INVx2_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
AOI22xp5_ASAP7_75t_L g575 ( .A1(n_361), .A2(n_576), .B1(n_577), .B2(n_578), .Y(n_575) );
AND2x4_ASAP7_75t_L g628 ( .A(n_361), .B(n_364), .Y(n_628) );
AND2x2_ASAP7_75t_L g966 ( .A(n_361), .B(n_364), .Y(n_966) );
BUFx3_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx2_ASAP7_75t_SL g375 ( .A(n_363), .Y(n_375) );
INVx1_ASAP7_75t_L g380 ( .A(n_363), .Y(n_380) );
NAND2x1p5_ASAP7_75t_L g363 ( .A(n_364), .B(n_367), .Y(n_363) );
BUFx2_ASAP7_75t_L g580 ( .A(n_364), .Y(n_580) );
AND2x4_ASAP7_75t_L g627 ( .A(n_364), .B(n_576), .Y(n_627) );
AND2x4_ASAP7_75t_L g702 ( .A(n_364), .B(n_576), .Y(n_702) );
INVx1_ASAP7_75t_L g704 ( .A(n_364), .Y(n_704) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
OR2x6_ASAP7_75t_L g689 ( .A(n_367), .B(n_440), .Y(n_689) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
OR2x2_ASAP7_75t_L g476 ( .A(n_368), .B(n_477), .Y(n_476) );
AND2x4_ASAP7_75t_L g499 ( .A(n_368), .B(n_387), .Y(n_499) );
AOI22xp33_ASAP7_75t_L g456 ( .A1(n_369), .A2(n_376), .B1(n_457), .B2(n_460), .Y(n_456) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVx2_ASAP7_75t_L g846 ( .A(n_371), .Y(n_846) );
NAND2x1p5_ASAP7_75t_L g371 ( .A(n_372), .B(n_375), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
INVx2_ASAP7_75t_L g576 ( .A(n_373), .Y(n_576) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
NOR3xp33_ASAP7_75t_L g897 ( .A(n_377), .B(n_898), .C(n_899), .Y(n_897) );
AND2x2_ASAP7_75t_L g377 ( .A(n_378), .B(n_380), .Y(n_377) );
HB1xp67_ASAP7_75t_L g1020 ( .A(n_378), .Y(n_1020) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g865 ( .A(n_380), .B(n_720), .Y(n_865) );
OAI31xp33_ASAP7_75t_L g381 ( .A1(n_382), .A2(n_398), .A3(n_462), .B(n_471), .Y(n_381) );
INVx3_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
INVx3_ASAP7_75t_L g801 ( .A(n_384), .Y(n_801) );
AOI22xp33_ASAP7_75t_L g873 ( .A1(n_384), .A2(n_467), .B1(n_874), .B2(n_875), .Y(n_873) );
AOI22xp33_ASAP7_75t_L g1167 ( .A1(n_384), .A2(n_467), .B1(n_1168), .B2(n_1169), .Y(n_1167) );
AND2x4_ASAP7_75t_L g384 ( .A(n_385), .B(n_389), .Y(n_384) );
AND2x4_ASAP7_75t_L g394 ( .A(n_385), .B(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx2_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
AND2x4_ASAP7_75t_L g464 ( .A(n_387), .B(n_465), .Y(n_464) );
AND2x2_ASAP7_75t_L g467 ( .A(n_387), .B(n_468), .Y(n_467) );
INVx1_ASAP7_75t_L g441 ( .A(n_388), .Y(n_441) );
INVx1_ASAP7_75t_L g511 ( .A(n_388), .Y(n_511) );
INVx1_ASAP7_75t_L g1526 ( .A(n_389), .Y(n_1526) );
INVx2_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g514 ( .A(n_390), .Y(n_514) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
BUFx6f_ASAP7_75t_L g408 ( .A(n_391), .Y(n_408) );
INVx3_ASAP7_75t_L g428 ( .A(n_391), .Y(n_428) );
AND2x4_ASAP7_75t_L g396 ( .A(n_392), .B(n_397), .Y(n_396) );
INVx8_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
BUFx6f_ASAP7_75t_L g759 ( .A(n_395), .Y(n_759) );
BUFx3_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
BUFx6f_ASAP7_75t_L g508 ( .A(n_396), .Y(n_508) );
BUFx3_ASAP7_75t_L g523 ( .A(n_396), .Y(n_523) );
BUFx6f_ASAP7_75t_L g531 ( .A(n_396), .Y(n_531) );
BUFx2_ASAP7_75t_L g594 ( .A(n_396), .Y(n_594) );
OAI221xp5_ASAP7_75t_L g398 ( .A1(n_399), .A2(n_409), .B1(n_422), .B2(n_430), .C(n_443), .Y(n_398) );
OAI22xp5_ASAP7_75t_L g399 ( .A1(n_400), .A2(n_401), .B1(n_406), .B2(n_407), .Y(n_399) );
INVx2_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx2_ASAP7_75t_SL g423 ( .A(n_402), .Y(n_423) );
INVx2_ASAP7_75t_L g1040 ( .A(n_402), .Y(n_1040) );
INVx2_ASAP7_75t_L g1513 ( .A(n_402), .Y(n_1513) );
BUFx3_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g606 ( .A(n_403), .Y(n_606) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g502 ( .A(n_404), .Y(n_502) );
BUFx2_ASAP7_75t_L g887 ( .A(n_404), .Y(n_887) );
INVx1_ASAP7_75t_L g461 ( .A(n_405), .Y(n_461) );
AND2x4_ASAP7_75t_L g468 ( .A(n_405), .B(n_469), .Y(n_468) );
OAI22xp5_ASAP7_75t_L g932 ( .A1(n_407), .A2(n_933), .B1(n_934), .B2(n_936), .Y(n_932) );
INVx2_ASAP7_75t_SL g407 ( .A(n_408), .Y(n_407) );
INVx2_ASAP7_75t_SL g685 ( .A(n_408), .Y(n_685) );
INVx4_ASAP7_75t_L g762 ( .A(n_408), .Y(n_762) );
INVx2_ASAP7_75t_SL g807 ( .A(n_408), .Y(n_807) );
INVx2_ASAP7_75t_SL g998 ( .A(n_408), .Y(n_998) );
OAI221xp5_ASAP7_75t_L g409 ( .A1(n_410), .A2(n_414), .B1(n_415), .B2(n_418), .C(n_419), .Y(n_409) );
OAI21xp5_ASAP7_75t_SL g1176 ( .A1(n_410), .A2(n_1177), .B(n_1178), .Y(n_1176) );
INVx2_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx3_ASAP7_75t_L g455 ( .A(n_411), .Y(n_455) );
BUFx2_ASAP7_75t_L g811 ( .A(n_411), .Y(n_811) );
INVx2_ASAP7_75t_L g818 ( .A(n_411), .Y(n_818) );
AND2x2_ASAP7_75t_L g411 ( .A(n_412), .B(n_413), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_412), .B(n_413), .Y(n_432) );
INVx1_ASAP7_75t_L g591 ( .A(n_413), .Y(n_591) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g1140 ( .A(n_416), .Y(n_1140) );
INVx2_ASAP7_75t_SL g1146 ( .A(n_416), .Y(n_1146) );
INVx2_ASAP7_75t_SL g416 ( .A(n_417), .Y(n_416) );
OAI221xp5_ASAP7_75t_L g1527 ( .A1(n_419), .A2(n_1528), .B1(n_1529), .B2(n_1530), .C(n_1532), .Y(n_1527) );
INVx2_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
BUFx2_ASAP7_75t_SL g816 ( .A(n_421), .Y(n_816) );
OAI22xp5_ASAP7_75t_L g422 ( .A1(n_423), .A2(n_424), .B1(n_425), .B2(n_429), .Y(n_422) );
BUFx2_ASAP7_75t_L g1522 ( .A(n_423), .Y(n_1522) );
AOI22xp5_ASAP7_75t_L g482 ( .A1(n_424), .A2(n_433), .B1(n_483), .B2(n_486), .Y(n_482) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx2_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx2_ASAP7_75t_L g878 ( .A(n_427), .Y(n_878) );
INVx3_ASAP7_75t_L g1575 ( .A(n_427), .Y(n_1575) );
BUFx6f_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx3_ASAP7_75t_L g505 ( .A(n_428), .Y(n_505) );
INVx3_ASAP7_75t_L g535 ( .A(n_428), .Y(n_535) );
AOI222xp33_ASAP7_75t_L g473 ( .A1(n_429), .A2(n_436), .B1(n_453), .B2(n_474), .C1(n_478), .C2(n_480), .Y(n_473) );
OAI221xp5_ASAP7_75t_L g430 ( .A1(n_431), .A2(n_433), .B1(n_434), .B2(n_436), .C(n_437), .Y(n_430) );
BUFx3_ASAP7_75t_L g927 ( .A(n_431), .Y(n_927) );
OAI22xp33_ASAP7_75t_L g928 ( .A1(n_431), .A2(n_929), .B1(n_930), .B2(n_931), .Y(n_928) );
INVx2_ASAP7_75t_L g1055 ( .A(n_431), .Y(n_1055) );
BUFx6f_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
OAI22xp5_ASAP7_75t_SL g1051 ( .A1(n_434), .A2(n_1052), .B1(n_1053), .B2(n_1054), .Y(n_1051) );
INVx2_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx1_ASAP7_75t_L g823 ( .A(n_435), .Y(n_823) );
OAI221xp5_ASAP7_75t_L g820 ( .A1(n_437), .A2(n_821), .B1(n_822), .B2(n_823), .C(n_824), .Y(n_820) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx2_ASAP7_75t_SL g438 ( .A(n_439), .Y(n_438) );
INVx2_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
NAND2x1p5_ASAP7_75t_L g440 ( .A(n_441), .B(n_442), .Y(n_440) );
AOI21xp5_ASAP7_75t_L g443 ( .A1(n_444), .A2(n_453), .B(n_454), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
NOR2xp67_ASAP7_75t_L g839 ( .A(n_445), .B(n_649), .Y(n_839) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_446), .B(n_450), .Y(n_445) );
AND2x2_ASAP7_75t_L g832 ( .A(n_446), .B(n_587), .Y(n_832) );
AND2x2_ASAP7_75t_L g1518 ( .A(n_446), .B(n_587), .Y(n_1518) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
AOI21xp33_ASAP7_75t_L g454 ( .A1(n_447), .A2(n_455), .B(n_456), .Y(n_454) );
OR2x6_ASAP7_75t_L g817 ( .A(n_447), .B(n_818), .Y(n_817) );
OR2x6_ASAP7_75t_L g835 ( .A(n_447), .B(n_461), .Y(n_835) );
INVx1_ASAP7_75t_L g883 ( .A(n_447), .Y(n_883) );
OR2x2_ASAP7_75t_L g1179 ( .A(n_447), .B(n_818), .Y(n_1179) );
INVx2_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
AND2x2_ASAP7_75t_L g498 ( .A(n_450), .B(n_499), .Y(n_498) );
INVx2_ASAP7_75t_SL g450 ( .A(n_451), .Y(n_450) );
INVx2_ASAP7_75t_SL g610 ( .A(n_451), .Y(n_610) );
INVx2_ASAP7_75t_L g1211 ( .A(n_451), .Y(n_1211) );
INVx3_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
BUFx6f_ASAP7_75t_L g465 ( .A(n_452), .Y(n_465) );
OAI221xp5_ASAP7_75t_L g891 ( .A1(n_455), .A2(n_813), .B1(n_816), .B2(n_892), .C(n_893), .Y(n_891) );
INVx1_ASAP7_75t_L g1580 ( .A(n_455), .Y(n_1580) );
NAND2x1_ASAP7_75t_SL g518 ( .A(n_457), .B(n_519), .Y(n_518) );
NAND2x1p5_ASAP7_75t_L g882 ( .A(n_457), .B(n_883), .Y(n_882) );
INVx2_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
HB1xp67_ASAP7_75t_L g587 ( .A(n_459), .Y(n_587) );
NAND2x1p5_ASAP7_75t_L g521 ( .A(n_460), .B(n_519), .Y(n_521) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
CKINVDCx6p67_ASAP7_75t_R g463 ( .A(n_464), .Y(n_463) );
BUFx6f_ASAP7_75t_L g880 ( .A(n_465), .Y(n_880) );
INVx3_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVx3_ASAP7_75t_L g800 ( .A(n_467), .Y(n_800) );
BUFx6f_ASAP7_75t_L g528 ( .A(n_468), .Y(n_528) );
BUFx6f_ASAP7_75t_L g598 ( .A(n_468), .Y(n_598) );
BUFx6f_ASAP7_75t_L g613 ( .A(n_468), .Y(n_613) );
BUFx2_ASAP7_75t_L g996 ( .A(n_468), .Y(n_996) );
INVx1_ASAP7_75t_L g1160 ( .A(n_468), .Y(n_1160) );
INVx1_ASAP7_75t_L g1214 ( .A(n_468), .Y(n_1214) );
INVx1_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
INVx2_ASAP7_75t_L g581 ( .A(n_471), .Y(n_581) );
BUFx8_ASAP7_75t_SL g894 ( .A(n_471), .Y(n_894) );
OAI31xp33_ASAP7_75t_L g1508 ( .A1(n_471), .A2(n_1509), .A3(n_1519), .B(n_1533), .Y(n_1508) );
INVx2_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
BUFx2_ASAP7_75t_L g733 ( .A(n_472), .Y(n_733) );
AOI22xp33_ASAP7_75t_L g843 ( .A1(n_474), .A2(n_483), .B1(n_824), .B2(n_828), .Y(n_843) );
AOI221xp5_ASAP7_75t_L g910 ( .A1(n_474), .A2(n_483), .B1(n_911), .B2(n_912), .C(n_913), .Y(n_910) );
AOI221xp5_ASAP7_75t_L g1197 ( .A1(n_474), .A2(n_483), .B1(n_1198), .B2(n_1199), .C(n_1200), .Y(n_1197) );
AOI22xp33_ASAP7_75t_L g1488 ( .A1(n_474), .A2(n_483), .B1(n_1489), .B2(n_1490), .Y(n_1488) );
AND2x2_ASAP7_75t_L g483 ( .A(n_475), .B(n_484), .Y(n_483) );
INVx1_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
OR2x6_ASAP7_75t_L g487 ( .A(n_476), .B(n_488), .Y(n_487) );
INVx2_ASAP7_75t_L g542 ( .A(n_477), .Y(n_542) );
OR2x2_ASAP7_75t_L g543 ( .A(n_477), .B(n_544), .Y(n_543) );
OR2x2_ASAP7_75t_L g546 ( .A(n_477), .B(n_547), .Y(n_546) );
A2O1A1Ixp33_ASAP7_75t_L g944 ( .A1(n_477), .A2(n_945), .B(n_947), .C(n_949), .Y(n_944) );
AOI22xp33_ASAP7_75t_L g842 ( .A1(n_478), .A2(n_486), .B1(n_822), .B2(n_829), .Y(n_842) );
AOI22xp33_ASAP7_75t_L g1485 ( .A1(n_478), .A2(n_486), .B1(n_1486), .B2(n_1487), .Y(n_1485) );
CKINVDCx6p67_ASAP7_75t_R g478 ( .A(n_479), .Y(n_478) );
INVx2_ASAP7_75t_L g693 ( .A(n_480), .Y(n_693) );
OR2x6_ASAP7_75t_L g838 ( .A(n_480), .B(n_839), .Y(n_838) );
INVx2_ASAP7_75t_L g647 ( .A(n_481), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g967 ( .A(n_481), .B(n_968), .Y(n_967) );
AOI22xp33_ASAP7_75t_L g947 ( .A1(n_484), .A2(n_931), .B1(n_933), .B2(n_948), .Y(n_947) );
INVx2_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
INVx1_ASAP7_75t_L g631 ( .A(n_485), .Y(n_631) );
OAI22xp5_ASAP7_75t_L g1186 ( .A1(n_485), .A2(n_624), .B1(n_1174), .B2(n_1175), .Y(n_1186) );
CKINVDCx6p67_ASAP7_75t_R g486 ( .A(n_487), .Y(n_486) );
OAI21xp33_ASAP7_75t_L g552 ( .A1(n_488), .A2(n_553), .B(n_554), .Y(n_552) );
OAI221xp5_ASAP7_75t_L g710 ( .A1(n_488), .A2(n_667), .B1(n_670), .B2(n_711), .C(n_713), .Y(n_710) );
INVx2_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
INVx1_ASAP7_75t_L g565 ( .A(n_489), .Y(n_565) );
INVx1_ASAP7_75t_L g574 ( .A(n_489), .Y(n_574) );
BUFx2_ASAP7_75t_L g776 ( .A(n_489), .Y(n_776) );
BUFx4f_ASAP7_75t_L g904 ( .A(n_489), .Y(n_904) );
AND2x2_ASAP7_75t_L g489 ( .A(n_490), .B(n_491), .Y(n_489) );
OR2x2_ASAP7_75t_L g547 ( .A(n_490), .B(n_491), .Y(n_547) );
XNOR2xp5_ASAP7_75t_L g492 ( .A(n_493), .B(n_582), .Y(n_492) );
NAND3xp33_ASAP7_75t_L g494 ( .A(n_495), .B(n_524), .C(n_537), .Y(n_494) );
NOR2xp33_ASAP7_75t_L g495 ( .A(n_496), .B(n_517), .Y(n_495) );
INVx1_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
AND2x2_ASAP7_75t_L g527 ( .A(n_499), .B(n_528), .Y(n_527) );
AND2x2_ASAP7_75t_L g530 ( .A(n_499), .B(n_531), .Y(n_530) );
AND2x2_ASAP7_75t_L g534 ( .A(n_499), .B(n_535), .Y(n_534) );
AOI22xp5_ASAP7_75t_L g604 ( .A1(n_499), .A2(n_516), .B1(n_605), .B2(n_612), .Y(n_604) );
AND2x4_ASAP7_75t_L g666 ( .A(n_499), .B(n_505), .Y(n_666) );
AND2x6_ASAP7_75t_L g668 ( .A(n_499), .B(n_523), .Y(n_668) );
AND2x4_ASAP7_75t_L g671 ( .A(n_499), .B(n_610), .Y(n_671) );
AND2x2_ASAP7_75t_L g673 ( .A(n_499), .B(n_528), .Y(n_673) );
AND2x2_ASAP7_75t_L g755 ( .A(n_499), .B(n_528), .Y(n_755) );
AND2x2_ASAP7_75t_L g1228 ( .A(n_499), .B(n_528), .Y(n_1228) );
OAI221xp5_ASAP7_75t_L g500 ( .A1(n_501), .A2(n_503), .B1(n_504), .B2(n_506), .C(n_507), .Y(n_500) );
INVx1_ASAP7_75t_L g827 ( .A(n_501), .Y(n_827) );
INVx1_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
INVx1_ASAP7_75t_L g935 ( .A(n_502), .Y(n_935) );
HB1xp67_ASAP7_75t_L g1173 ( .A(n_502), .Y(n_1173) );
INVx1_ASAP7_75t_SL g504 ( .A(n_505), .Y(n_504) );
INVx2_ASAP7_75t_L g607 ( .A(n_505), .Y(n_607) );
INVx1_ASAP7_75t_L g889 ( .A(n_505), .Y(n_889) );
BUFx3_ASAP7_75t_L g1149 ( .A(n_505), .Y(n_1149) );
OAI22xp5_ASAP7_75t_L g557 ( .A1(n_506), .A2(n_558), .B1(n_559), .B2(n_561), .Y(n_557) );
INVx2_ASAP7_75t_SL g1165 ( .A(n_508), .Y(n_1165) );
BUFx2_ASAP7_75t_L g1221 ( .A(n_508), .Y(n_1221) );
OAI33xp33_ASAP7_75t_L g1133 ( .A1(n_509), .A2(n_1134), .A3(n_1139), .B1(n_1143), .B2(n_1145), .B3(n_1147), .Y(n_1133) );
OAI33xp33_ASAP7_75t_L g1563 ( .A1(n_509), .A2(n_1143), .A3(n_1564), .B1(n_1569), .B2(n_1572), .B3(n_1577), .Y(n_1563) );
NAND3xp33_ASAP7_75t_L g512 ( .A(n_513), .B(n_515), .C(n_516), .Y(n_512) );
INVx1_ASAP7_75t_L g1137 ( .A(n_514), .Y(n_1137) );
HB1xp67_ASAP7_75t_L g1215 ( .A(n_514), .Y(n_1215) );
HB1xp67_ASAP7_75t_L g1130 ( .A(n_518), .Y(n_1130) );
INVx2_ASAP7_75t_L g1561 ( .A(n_518), .Y(n_1561) );
NAND2x1p5_ASAP7_75t_L g522 ( .A(n_519), .B(n_523), .Y(n_522) );
AND2x4_ASAP7_75t_L g586 ( .A(n_519), .B(n_587), .Y(n_586) );
AND2x4_ASAP7_75t_L g589 ( .A(n_519), .B(n_590), .Y(n_589) );
AND2x4_ASAP7_75t_L g593 ( .A(n_519), .B(n_594), .Y(n_593) );
INVx3_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
BUFx4f_ASAP7_75t_L g1036 ( .A(n_521), .Y(n_1036) );
BUFx4f_ASAP7_75t_L g1131 ( .A(n_521), .Y(n_1131) );
BUFx3_ASAP7_75t_L g1132 ( .A(n_522), .Y(n_1132) );
BUFx2_ASAP7_75t_L g1562 ( .A(n_522), .Y(n_1562) );
NOR2xp33_ASAP7_75t_SL g524 ( .A(n_525), .B(n_532), .Y(n_524) );
INVx1_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
INVx1_ASAP7_75t_L g940 ( .A(n_527), .Y(n_940) );
INVx1_ASAP7_75t_L g1035 ( .A(n_527), .Y(n_1035) );
AOI22xp33_ASAP7_75t_L g1126 ( .A1(n_527), .A2(n_671), .B1(n_1127), .B2(n_1128), .Y(n_1126) );
INVx1_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
INVxp67_ASAP7_75t_L g941 ( .A(n_530), .Y(n_941) );
INVx2_ASAP7_75t_SL g681 ( .A(n_531), .Y(n_681) );
BUFx6f_ASAP7_75t_L g765 ( .A(n_531), .Y(n_765) );
INVx2_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
INVx2_ASAP7_75t_L g615 ( .A(n_535), .Y(n_615) );
HB1xp67_ASAP7_75t_L g923 ( .A(n_535), .Y(n_923) );
INVx1_ASAP7_75t_L g1049 ( .A(n_535), .Y(n_1049) );
INVx2_ASAP7_75t_L g603 ( .A(n_536), .Y(n_603) );
AND2x4_ASAP7_75t_L g692 ( .A(n_536), .B(n_693), .Y(n_692) );
OAI31xp33_ASAP7_75t_SL g537 ( .A1(n_538), .A2(n_545), .A3(n_551), .B(n_581), .Y(n_537) );
INVx1_ASAP7_75t_L g1232 ( .A(n_539), .Y(n_1232) );
INVx1_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
AND2x2_ASAP7_75t_L g540 ( .A(n_541), .B(n_542), .Y(n_540) );
AOI22xp5_ASAP7_75t_L g625 ( .A1(n_541), .A2(n_550), .B1(n_618), .B2(n_626), .Y(n_625) );
INVx1_ASAP7_75t_L g1067 ( .A(n_541), .Y(n_1067) );
BUFx4f_ASAP7_75t_L g1191 ( .A(n_541), .Y(n_1191) );
AND2x4_ASAP7_75t_L g549 ( .A(n_542), .B(n_550), .Y(n_549) );
AOI222xp33_ASAP7_75t_L g620 ( .A1(n_542), .A2(n_588), .B1(n_592), .B2(n_621), .C1(n_627), .C2(n_628), .Y(n_620) );
AND2x4_ASAP7_75t_L g698 ( .A(n_542), .B(n_699), .Y(n_698) );
AOI221xp5_ASAP7_75t_L g1065 ( .A1(n_542), .A2(n_549), .B1(n_639), .B2(n_1053), .C(n_1066), .Y(n_1065) );
INVx4_ASAP7_75t_L g731 ( .A(n_543), .Y(n_731) );
INVx1_ASAP7_75t_L g562 ( .A(n_544), .Y(n_562) );
INVx2_ASAP7_75t_L g1079 ( .A(n_544), .Y(n_1079) );
INVx6_ASAP7_75t_L g729 ( .A(n_546), .Y(n_729) );
INVx1_ASAP7_75t_L g560 ( .A(n_547), .Y(n_560) );
INVx1_ASAP7_75t_L g623 ( .A(n_547), .Y(n_623) );
INVx2_ASAP7_75t_L g712 ( .A(n_547), .Y(n_712) );
INVx2_ASAP7_75t_SL g548 ( .A(n_549), .Y(n_548) );
BUFx6f_ASAP7_75t_L g715 ( .A(n_549), .Y(n_715) );
AOI221xp5_ASAP7_75t_L g1107 ( .A1(n_549), .A2(n_639), .B1(n_1108), .B2(n_1109), .C(n_1112), .Y(n_1107) );
HB1xp67_ASAP7_75t_L g1240 ( .A(n_549), .Y(n_1240) );
INVx2_ASAP7_75t_SL g633 ( .A(n_550), .Y(n_633) );
AND2x4_ASAP7_75t_L g639 ( .A(n_550), .B(n_580), .Y(n_639) );
BUFx6f_ASAP7_75t_L g720 ( .A(n_550), .Y(n_720) );
INVx1_ASAP7_75t_L g782 ( .A(n_550), .Y(n_782) );
BUFx3_ASAP7_75t_L g857 ( .A(n_550), .Y(n_857) );
BUFx4f_ASAP7_75t_L g948 ( .A(n_550), .Y(n_948) );
OAI211xp5_ASAP7_75t_SL g551 ( .A1(n_552), .A2(n_557), .B(n_563), .C(n_571), .Y(n_551) );
INVx2_ASAP7_75t_L g1019 ( .A(n_555), .Y(n_1019) );
BUFx3_ASAP7_75t_L g1074 ( .A(n_555), .Y(n_1074) );
INVx1_ASAP7_75t_L g722 ( .A(n_556), .Y(n_722) );
BUFx2_ASAP7_75t_L g1590 ( .A(n_556), .Y(n_1590) );
OAI221xp5_ASAP7_75t_L g774 ( .A1(n_559), .A2(n_751), .B1(n_753), .B2(n_775), .C(n_777), .Y(n_774) );
OAI221xp5_ASAP7_75t_L g906 ( .A1(n_559), .A2(n_903), .B1(n_907), .B2(n_908), .C(n_909), .Y(n_906) );
INVx2_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
INVx1_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
OAI211xp5_ASAP7_75t_L g563 ( .A1(n_564), .A2(n_565), .B(n_566), .C(n_567), .Y(n_563) );
OAI211xp5_ASAP7_75t_L g1236 ( .A1(n_565), .A2(n_1224), .B(n_1237), .C(n_1238), .Y(n_1236) );
BUFx6f_ASAP7_75t_L g637 ( .A(n_568), .Y(n_637) );
INVx1_ASAP7_75t_L g856 ( .A(n_568), .Y(n_856) );
INVx2_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
INVx2_ASAP7_75t_L g642 ( .A(n_569), .Y(n_642) );
INVx1_ASAP7_75t_L g786 ( .A(n_569), .Y(n_786) );
INVx2_ASAP7_75t_SL g1014 ( .A(n_569), .Y(n_1014) );
INVx1_ASAP7_75t_L g1083 ( .A(n_569), .Y(n_1083) );
NAND2xp33_ASAP7_75t_L g573 ( .A(n_574), .B(n_575), .Y(n_573) );
INVx1_ASAP7_75t_L g954 ( .A(n_574), .Y(n_954) );
BUFx3_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
NAND2xp5_ASAP7_75t_SL g582 ( .A(n_583), .B(n_650), .Y(n_582) );
INVx1_ASAP7_75t_L g652 ( .A(n_584), .Y(n_652) );
NAND3xp33_ASAP7_75t_SL g584 ( .A(n_585), .B(n_595), .C(n_604), .Y(n_584) );
AOI221xp5_ASAP7_75t_L g585 ( .A1(n_586), .A2(n_588), .B1(n_589), .B2(n_592), .C(n_593), .Y(n_585) );
INVx1_ASAP7_75t_L g661 ( .A(n_586), .Y(n_661) );
AOI221xp5_ASAP7_75t_L g742 ( .A1(n_586), .A2(n_743), .B1(n_745), .B2(n_746), .C(n_747), .Y(n_742) );
AOI221xp5_ASAP7_75t_L g969 ( .A1(n_586), .A2(n_589), .B1(n_593), .B2(n_970), .C(n_971), .Y(n_969) );
AOI221xp5_ASAP7_75t_L g980 ( .A1(n_586), .A2(n_589), .B1(n_593), .B2(n_981), .C(n_982), .Y(n_980) );
AOI21xp5_ASAP7_75t_L g1090 ( .A1(n_586), .A2(n_593), .B(n_1063), .Y(n_1090) );
AOI221xp5_ASAP7_75t_L g1205 ( .A1(n_586), .A2(n_589), .B1(n_593), .B2(n_1206), .C(n_1207), .Y(n_1205) );
HB1xp67_ASAP7_75t_L g658 ( .A(n_589), .Y(n_658) );
INVx1_ASAP7_75t_L g744 ( .A(n_589), .Y(n_744) );
INVx1_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
AOI221xp5_ASAP7_75t_L g657 ( .A1(n_593), .A2(n_658), .B1(n_659), .B2(n_660), .C(n_662), .Y(n_657) );
HB1xp67_ASAP7_75t_L g747 ( .A(n_593), .Y(n_747) );
AOI22xp33_ASAP7_75t_L g608 ( .A1(n_594), .A2(n_609), .B1(n_610), .B2(n_611), .Y(n_608) );
INVx1_ASAP7_75t_L g994 ( .A(n_594), .Y(n_994) );
AOI22xp5_ASAP7_75t_L g595 ( .A1(n_596), .A2(n_597), .B1(n_602), .B2(n_603), .Y(n_595) );
AOI33xp33_ASAP7_75t_L g990 ( .A1(n_596), .A2(n_688), .A3(n_991), .B1(n_995), .B2(n_999), .B3(n_1000), .Y(n_990) );
BUFx2_ASAP7_75t_L g1209 ( .A(n_596), .Y(n_1209) );
AOI22xp5_ASAP7_75t_L g640 ( .A1(n_602), .A2(n_641), .B1(n_644), .B2(n_646), .Y(n_640) );
INVx2_ASAP7_75t_L g805 ( .A(n_606), .Y(n_805) );
OAI22xp5_ASAP7_75t_L g1171 ( .A1(n_607), .A2(n_1172), .B1(n_1174), .B2(n_1175), .Y(n_1171) );
INVx1_ASAP7_75t_L g1217 ( .A(n_607), .Y(n_1217) );
BUFx3_ASAP7_75t_L g679 ( .A(n_610), .Y(n_679) );
INVx1_ASAP7_75t_L g1163 ( .A(n_610), .Y(n_1163) );
INVx1_ASAP7_75t_L g1220 ( .A(n_610), .Y(n_1220) );
BUFx3_ASAP7_75t_L g683 ( .A(n_613), .Y(n_683) );
INVx2_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
INVx1_ASAP7_75t_L g651 ( .A(n_619), .Y(n_651) );
AOI31xp33_ASAP7_75t_SL g619 ( .A1(n_620), .A2(n_629), .A3(n_640), .B(n_648), .Y(n_619) );
OAI221xp5_ASAP7_75t_SL g1068 ( .A1(n_622), .A2(n_1041), .B1(n_1044), .B2(n_1069), .C(n_1070), .Y(n_1068) );
INVx2_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
INVx1_ASAP7_75t_L g638 ( .A(n_624), .Y(n_638) );
INVx2_ASAP7_75t_L g1009 ( .A(n_627), .Y(n_1009) );
INVx4_ASAP7_75t_L g1062 ( .A(n_627), .Y(n_1062) );
AOI222xp33_ASAP7_75t_SL g1059 ( .A1(n_628), .A2(n_646), .B1(n_1060), .B2(n_1061), .C1(n_1063), .C2(n_1064), .Y(n_1059) );
AOI322xp5_ASAP7_75t_L g1098 ( .A1(n_628), .A2(n_702), .A3(n_1099), .B1(n_1101), .B2(n_1104), .C1(n_1105), .C2(n_1106), .Y(n_1098) );
INVx2_ASAP7_75t_SL g1235 ( .A(n_628), .Y(n_1235) );
AOI21xp5_ASAP7_75t_L g629 ( .A1(n_630), .A2(n_636), .B(n_639), .Y(n_629) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
INVx2_ASAP7_75t_L g853 ( .A(n_633), .Y(n_853) );
INVxp67_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
INVx3_ASAP7_75t_L g1071 ( .A(n_635), .Y(n_1071) );
INVx1_ASAP7_75t_L g949 ( .A(n_639), .Y(n_949) );
AOI221xp5_ASAP7_75t_L g1239 ( .A1(n_639), .A2(n_1240), .B1(n_1241), .B2(n_1242), .C(n_1244), .Y(n_1239) );
HB1xp67_ASAP7_75t_L g852 ( .A(n_642), .Y(n_852) );
AOI22xp33_ASAP7_75t_L g945 ( .A1(n_642), .A2(n_930), .B1(n_936), .B2(n_946), .Y(n_945) );
BUFx3_ASAP7_75t_L g1022 ( .A(n_642), .Y(n_1022) );
INVx2_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
INVx1_ASAP7_75t_L g1606 ( .A(n_648), .Y(n_1606) );
INVx2_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
NAND3xp33_ASAP7_75t_L g650 ( .A(n_651), .B(n_652), .C(n_653), .Y(n_650) );
INVx2_ASAP7_75t_L g735 ( .A(n_654), .Y(n_735) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_656), .B(n_690), .Y(n_655) );
AND4x1_ASAP7_75t_L g656 ( .A(n_657), .B(n_663), .C(n_669), .D(n_674), .Y(n_656) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
AOI22xp33_ASAP7_75t_L g663 ( .A1(n_664), .A2(n_665), .B1(n_667), .B2(n_668), .Y(n_663) );
BUFx2_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
BUFx2_ASAP7_75t_L g750 ( .A(n_666), .Y(n_750) );
BUFx2_ASAP7_75t_L g985 ( .A(n_666), .Y(n_985) );
BUFx2_ASAP7_75t_L g1089 ( .A(n_666), .Y(n_1089) );
BUFx2_ASAP7_75t_L g1124 ( .A(n_666), .Y(n_1124) );
AOI22xp33_ASAP7_75t_L g748 ( .A1(n_668), .A2(n_749), .B1(n_750), .B2(n_751), .Y(n_748) );
AOI22xp33_ASAP7_75t_L g983 ( .A1(n_668), .A2(n_984), .B1(n_985), .B2(n_986), .Y(n_983) );
AOI22xp33_ASAP7_75t_L g1122 ( .A1(n_668), .A2(n_1123), .B1(n_1124), .B2(n_1125), .Y(n_1122) );
AOI22xp33_ASAP7_75t_L g1222 ( .A1(n_668), .A2(n_1089), .B1(n_1223), .B2(n_1224), .Y(n_1222) );
AOI22xp33_ASAP7_75t_L g1553 ( .A1(n_668), .A2(n_1089), .B1(n_1554), .B2(n_1555), .Y(n_1553) );
AOI22xp33_ASAP7_75t_L g669 ( .A1(n_670), .A2(n_671), .B1(n_672), .B2(n_673), .Y(n_669) );
AOI22xp33_ASAP7_75t_L g752 ( .A1(n_671), .A2(n_753), .B1(n_754), .B2(n_755), .Y(n_752) );
AOI22xp33_ASAP7_75t_L g987 ( .A1(n_671), .A2(n_673), .B1(n_988), .B2(n_989), .Y(n_987) );
INVx1_ASAP7_75t_L g1087 ( .A(n_671), .Y(n_1087) );
AOI22xp33_ASAP7_75t_L g1225 ( .A1(n_671), .A2(n_1226), .B1(n_1227), .B2(n_1228), .Y(n_1225) );
AOI22xp33_ASAP7_75t_L g1556 ( .A1(n_671), .A2(n_673), .B1(n_1557), .B2(n_1558), .Y(n_1556) );
AOI33xp33_ASAP7_75t_L g674 ( .A1(n_675), .A2(n_678), .A3(n_682), .B1(n_686), .B2(n_687), .B3(n_688), .Y(n_674) );
AOI33xp33_ASAP7_75t_L g756 ( .A1(n_675), .A2(n_688), .A3(n_757), .B1(n_760), .B2(n_763), .B3(n_764), .Y(n_756) );
INVx2_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
INVx2_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
INVx2_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
OAI22xp5_ASAP7_75t_L g825 ( .A1(n_685), .A2(n_826), .B1(n_828), .B2(n_829), .Y(n_825) );
INVx1_ASAP7_75t_L g937 ( .A(n_688), .Y(n_937) );
INVx2_ASAP7_75t_L g1056 ( .A(n_688), .Y(n_1056) );
AOI33xp33_ASAP7_75t_L g1208 ( .A1(n_688), .A2(n_1209), .A3(n_1210), .B1(n_1212), .B2(n_1216), .B3(n_1218), .Y(n_1208) );
INVx6_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVx5_ASAP7_75t_L g1144 ( .A(n_689), .Y(n_1144) );
AOI21xp5_ASAP7_75t_L g690 ( .A1(n_691), .A2(n_694), .B(n_695), .Y(n_690) );
AOI21xp5_ASAP7_75t_L g1003 ( .A1(n_691), .A2(n_1004), .B(n_1005), .Y(n_1003) );
INVx1_ASAP7_75t_L g1550 ( .A(n_691), .Y(n_1550) );
INVx5_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
INVx1_ASAP7_75t_L g767 ( .A(n_692), .Y(n_767) );
INVx2_ASAP7_75t_SL g1119 ( .A(n_692), .Y(n_1119) );
INVx2_ASAP7_75t_L g1250 ( .A(n_692), .Y(n_1250) );
AOI31xp33_ASAP7_75t_L g695 ( .A1(n_696), .A2(n_714), .A3(n_727), .B(n_732), .Y(n_695) );
AOI211xp5_ASAP7_75t_L g696 ( .A1(n_697), .A2(n_698), .B(n_700), .C(n_705), .Y(n_696) );
AOI211xp5_ASAP7_75t_L g770 ( .A1(n_698), .A2(n_771), .B(n_772), .C(n_773), .Y(n_770) );
AOI21xp33_ASAP7_75t_SL g1006 ( .A1(n_698), .A2(n_1007), .B(n_1008), .Y(n_1006) );
NAND2xp5_ASAP7_75t_L g1116 ( .A(n_698), .B(n_1117), .Y(n_1116) );
INVx1_ASAP7_75t_L g1593 ( .A(n_698), .Y(n_1593) );
BUFx3_ASAP7_75t_L g859 ( .A(n_699), .Y(n_859) );
INVx2_ASAP7_75t_SL g1504 ( .A(n_699), .Y(n_1504) );
INVx2_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
INVx2_ASAP7_75t_SL g964 ( .A(n_702), .Y(n_964) );
AOI22xp33_ASAP7_75t_L g1594 ( .A1(n_702), .A2(n_1595), .B1(n_1596), .B2(n_1597), .Y(n_1594) );
INVx1_ASAP7_75t_L g1596 ( .A(n_703), .Y(n_1596) );
INVx1_ASAP7_75t_SL g726 ( .A(n_704), .Y(n_726) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
BUFx3_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
BUFx6f_ASAP7_75t_L g850 ( .A(n_709), .Y(n_850) );
INVx1_ASAP7_75t_L g861 ( .A(n_709), .Y(n_861) );
OAI221xp5_ASAP7_75t_L g902 ( .A1(n_711), .A2(n_892), .B1(n_893), .B2(n_903), .C(n_905), .Y(n_902) );
INVx2_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
HB1xp67_ASAP7_75t_L g1587 ( .A(n_712), .Y(n_1587) );
AOI221xp5_ASAP7_75t_L g714 ( .A1(n_715), .A2(n_716), .B1(n_717), .B2(n_723), .C(n_725), .Y(n_714) );
AOI221xp5_ASAP7_75t_L g779 ( .A1(n_715), .A2(n_725), .B1(n_780), .B2(n_784), .C(n_787), .Y(n_779) );
AOI221xp5_ASAP7_75t_L g1015 ( .A1(n_715), .A2(n_725), .B1(n_1016), .B2(n_1017), .C(n_1021), .Y(n_1015) );
INVx1_ASAP7_75t_L g1584 ( .A(n_715), .Y(n_1584) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
HB1xp67_ASAP7_75t_L g1499 ( .A(n_720), .Y(n_1499) );
INVx1_ASAP7_75t_L g1603 ( .A(n_720), .Y(n_1603) );
INVx1_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
INVx1_ASAP7_75t_L g1591 ( .A(n_725), .Y(n_1591) );
AOI22xp33_ASAP7_75t_L g727 ( .A1(n_728), .A2(n_729), .B1(n_730), .B2(n_731), .Y(n_727) );
AOI22xp33_ASAP7_75t_L g788 ( .A1(n_729), .A2(n_731), .B1(n_789), .B2(n_790), .Y(n_788) );
AOI22xp33_ASAP7_75t_L g1023 ( .A1(n_729), .A2(n_731), .B1(n_1024), .B2(n_1025), .Y(n_1023) );
AOI22xp33_ASAP7_75t_L g1113 ( .A1(n_729), .A2(n_731), .B1(n_1114), .B2(n_1115), .Y(n_1113) );
AOI22xp33_ASAP7_75t_L g1246 ( .A1(n_729), .A2(n_731), .B1(n_1247), .B2(n_1248), .Y(n_1246) );
INVx1_ASAP7_75t_L g1085 ( .A(n_732), .Y(n_1085) );
INVx2_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
OAI31xp33_ASAP7_75t_L g943 ( .A1(n_733), .A2(n_944), .A3(n_950), .B(n_963), .Y(n_943) );
AOI22xp5_ASAP7_75t_L g736 ( .A1(n_737), .A2(n_867), .B1(n_974), .B2(n_975), .Y(n_736) );
INVx1_ASAP7_75t_L g974 ( .A(n_737), .Y(n_974) );
XNOR2xp5_ASAP7_75t_L g737 ( .A(n_738), .B(n_795), .Y(n_737) );
INVx2_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
AND2x2_ASAP7_75t_L g740 ( .A(n_741), .B(n_766), .Y(n_740) );
AND4x1_ASAP7_75t_L g741 ( .A(n_742), .B(n_748), .C(n_752), .D(n_756), .Y(n_741) );
INVx1_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
HB1xp67_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
INVx2_ASAP7_75t_SL g761 ( .A(n_762), .Y(n_761) );
OAI22xp33_ASAP7_75t_L g1038 ( .A1(n_762), .A2(n_1039), .B1(n_1040), .B2(n_1041), .Y(n_1038) );
AOI21xp33_ASAP7_75t_SL g766 ( .A1(n_767), .A2(n_768), .B(n_769), .Y(n_766) );
AOI31xp33_ASAP7_75t_L g769 ( .A1(n_770), .A2(n_779), .A3(n_788), .B(n_791), .Y(n_769) );
INVx1_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
INVx1_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
BUFx2_ASAP7_75t_L g1604 ( .A(n_778), .Y(n_1604) );
INVx1_ASAP7_75t_L g781 ( .A(n_782), .Y(n_781) );
INVx1_ASAP7_75t_L g1082 ( .A(n_782), .Y(n_1082) );
HB1xp67_ASAP7_75t_L g785 ( .A(n_786), .Y(n_785) );
AOI31xp33_ASAP7_75t_L g1005 ( .A1(n_791), .A2(n_1006), .A3(n_1015), .B(n_1023), .Y(n_1005) );
INVx2_ASAP7_75t_L g791 ( .A(n_792), .Y(n_791) );
AOI22xp5_ASAP7_75t_L g1096 ( .A1(n_792), .A2(n_1097), .B1(n_1118), .B2(n_1119), .Y(n_1096) );
CKINVDCx8_ASAP7_75t_R g792 ( .A(n_793), .Y(n_792) );
OAI31xp33_ASAP7_75t_L g798 ( .A1(n_793), .A2(n_799), .A3(n_802), .B(n_819), .Y(n_798) );
OAI21xp5_ASAP7_75t_SL g1155 ( .A1(n_793), .A2(n_1156), .B(n_1170), .Y(n_1155) );
INVx1_ASAP7_75t_L g796 ( .A(n_797), .Y(n_796) );
NAND3xp33_ASAP7_75t_SL g797 ( .A(n_798), .B(n_836), .C(n_840), .Y(n_797) );
OAI22xp5_ASAP7_75t_L g803 ( .A1(n_804), .A2(n_806), .B1(n_807), .B2(n_808), .Y(n_803) );
INVx2_ASAP7_75t_L g804 ( .A(n_805), .Y(n_804) );
OAI221xp5_ASAP7_75t_L g809 ( .A1(n_810), .A2(n_812), .B1(n_813), .B2(n_815), .C(n_816), .Y(n_809) );
OAI22xp33_ASAP7_75t_L g1145 ( .A1(n_810), .A2(n_1108), .B1(n_1114), .B2(n_1146), .Y(n_1145) );
INVx1_ASAP7_75t_L g810 ( .A(n_811), .Y(n_810) );
INVx2_ASAP7_75t_L g821 ( .A(n_811), .Y(n_821) );
OAI22xp33_ASAP7_75t_L g924 ( .A1(n_813), .A2(n_925), .B1(n_926), .B2(n_927), .Y(n_924) );
OAI22xp33_ASAP7_75t_L g1042 ( .A1(n_813), .A2(n_818), .B1(n_1043), .B2(n_1044), .Y(n_1042) );
INVx3_ASAP7_75t_L g813 ( .A(n_814), .Y(n_813) );
INVx1_ASAP7_75t_L g826 ( .A(n_827), .Y(n_826) );
AOI22xp33_ASAP7_75t_L g830 ( .A1(n_831), .A2(n_832), .B1(n_833), .B2(n_834), .Y(n_830) );
AOI22xp33_ASAP7_75t_L g1516 ( .A1(n_834), .A2(n_1493), .B1(n_1494), .B2(n_1517), .Y(n_1516) );
CKINVDCx11_ASAP7_75t_R g834 ( .A(n_835), .Y(n_834) );
NAND2xp5_ASAP7_75t_L g836 ( .A(n_837), .B(n_838), .Y(n_836) );
NAND2xp5_ASAP7_75t_L g895 ( .A(n_838), .B(n_896), .Y(n_895) );
NAND2xp5_ASAP7_75t_L g1180 ( .A(n_838), .B(n_1181), .Y(n_1180) );
NAND2xp5_ASAP7_75t_L g1506 ( .A(n_838), .B(n_1507), .Y(n_1506) );
NOR2xp33_ASAP7_75t_L g840 ( .A(n_841), .B(n_844), .Y(n_840) );
NAND2xp5_ASAP7_75t_L g841 ( .A(n_842), .B(n_843), .Y(n_841) );
NAND3xp33_ASAP7_75t_SL g844 ( .A(n_845), .B(n_847), .C(n_863), .Y(n_844) );
INVx1_ASAP7_75t_L g1195 ( .A(n_846), .Y(n_1195) );
AOI33xp33_ASAP7_75t_L g847 ( .A1(n_848), .A2(n_849), .A3(n_851), .B1(n_854), .B2(n_858), .B3(n_862), .Y(n_847) );
INVx2_ASAP7_75t_L g855 ( .A(n_856), .Y(n_855) );
INVx1_ASAP7_75t_L g860 ( .A(n_861), .Y(n_860) );
NAND3xp33_ASAP7_75t_SL g1491 ( .A(n_863), .B(n_1492), .C(n_1495), .Y(n_1491) );
INVx1_ASAP7_75t_L g863 ( .A(n_864), .Y(n_863) );
INVx1_ASAP7_75t_L g864 ( .A(n_865), .Y(n_864) );
INVx1_ASAP7_75t_L g867 ( .A(n_868), .Y(n_867) );
HB1xp67_ASAP7_75t_L g975 ( .A(n_868), .Y(n_975) );
XNOR2x1_ASAP7_75t_L g868 ( .A(n_869), .B(n_916), .Y(n_868) );
INVx1_ASAP7_75t_L g914 ( .A(n_870), .Y(n_914) );
NAND4xp25_ASAP7_75t_L g870 ( .A(n_871), .B(n_895), .C(n_897), .D(n_910), .Y(n_870) );
OAI21xp5_ASAP7_75t_L g871 ( .A1(n_872), .A2(n_884), .B(n_894), .Y(n_871) );
AOI21xp5_ASAP7_75t_L g876 ( .A1(n_877), .A2(n_879), .B(n_881), .Y(n_876) );
HB1xp67_ASAP7_75t_L g992 ( .A(n_880), .Y(n_992) );
INVx1_ASAP7_75t_L g1002 ( .A(n_880), .Y(n_1002) );
OAI22xp5_ASAP7_75t_L g885 ( .A1(n_886), .A2(n_888), .B1(n_889), .B2(n_890), .Y(n_885) );
OAI22xp5_ASAP7_75t_L g919 ( .A1(n_886), .A2(n_920), .B1(n_921), .B2(n_922), .Y(n_919) );
BUFx2_ASAP7_75t_L g886 ( .A(n_887), .Y(n_886) );
INVx2_ASAP7_75t_L g1048 ( .A(n_887), .Y(n_1048) );
INVx2_ASAP7_75t_SL g903 ( .A(n_904), .Y(n_903) );
INVx1_ASAP7_75t_L g960 ( .A(n_904), .Y(n_960) );
INVx2_ASAP7_75t_L g1011 ( .A(n_904), .Y(n_1011) );
INVx1_ASAP7_75t_SL g973 ( .A(n_917), .Y(n_973) );
NAND4xp75_ASAP7_75t_L g917 ( .A(n_918), .B(n_938), .C(n_943), .D(n_969), .Y(n_917) );
INVx1_ASAP7_75t_L g922 ( .A(n_923), .Y(n_922) );
OAI211xp5_ASAP7_75t_L g959 ( .A1(n_926), .A2(n_960), .B(n_961), .C(n_962), .Y(n_959) );
OAI22xp33_ASAP7_75t_L g1139 ( .A1(n_927), .A2(n_1140), .B1(n_1141), .B2(n_1142), .Y(n_1139) );
BUFx3_ASAP7_75t_L g1528 ( .A(n_927), .Y(n_1528) );
OAI22xp33_ASAP7_75t_L g1569 ( .A1(n_929), .A2(n_1528), .B1(n_1570), .B2(n_1571), .Y(n_1569) );
OAI22xp33_ASAP7_75t_L g1577 ( .A1(n_929), .A2(n_1578), .B1(n_1579), .B2(n_1581), .Y(n_1577) );
BUFx2_ASAP7_75t_L g934 ( .A(n_935), .Y(n_934) );
BUFx2_ASAP7_75t_L g1135 ( .A(n_935), .Y(n_1135) );
NOR2x1_ASAP7_75t_L g938 ( .A(n_939), .B(n_942), .Y(n_938) );
INVx2_ASAP7_75t_SL g1588 ( .A(n_946), .Y(n_1588) );
NAND2xp5_ASAP7_75t_L g950 ( .A(n_951), .B(n_959), .Y(n_950) );
OAI211xp5_ASAP7_75t_L g951 ( .A1(n_952), .A2(n_953), .B(n_955), .C(n_956), .Y(n_951) );
INVx1_ASAP7_75t_L g953 ( .A(n_954), .Y(n_953) );
INVx3_ASAP7_75t_L g965 ( .A(n_966), .Y(n_965) );
HB1xp67_ASAP7_75t_L g976 ( .A(n_977), .Y(n_976) );
XNOR2x1_ASAP7_75t_L g977 ( .A(n_978), .B(n_1026), .Y(n_977) );
AND2x2_ASAP7_75t_L g978 ( .A(n_979), .B(n_1003), .Y(n_978) );
AND4x1_ASAP7_75t_L g979 ( .A(n_980), .B(n_983), .C(n_987), .D(n_990), .Y(n_979) );
OAI211xp5_ASAP7_75t_L g1010 ( .A1(n_986), .A2(n_1011), .B(n_1012), .C(n_1013), .Y(n_1010) );
INVx1_ASAP7_75t_L g993 ( .A(n_994), .Y(n_993) );
INVx1_ASAP7_75t_L g997 ( .A(n_998), .Y(n_997) );
OAI221xp5_ASAP7_75t_L g1510 ( .A1(n_998), .A2(n_1486), .B1(n_1490), .B2(n_1511), .C(n_1514), .Y(n_1510) );
INVx1_ASAP7_75t_L g1001 ( .A(n_1002), .Y(n_1001) );
INVx1_ASAP7_75t_L g1515 ( .A(n_1002), .Y(n_1515) );
INVx1_ASAP7_75t_L g1018 ( .A(n_1019), .Y(n_1018) );
XNOR2xp5_ASAP7_75t_L g1027 ( .A(n_1028), .B(n_1150), .Y(n_1027) );
XOR2xp5_ASAP7_75t_L g1028 ( .A(n_1029), .B(n_1091), .Y(n_1028) );
INVx1_ASAP7_75t_L g1029 ( .A(n_1030), .Y(n_1029) );
INVx1_ASAP7_75t_L g1030 ( .A(n_1031), .Y(n_1030) );
AND2x2_ASAP7_75t_L g1032 ( .A(n_1033), .B(n_1057), .Y(n_1032) );
NOR2xp33_ASAP7_75t_L g1033 ( .A(n_1034), .B(n_1037), .Y(n_1033) );
OAI22xp5_ASAP7_75t_L g1045 ( .A1(n_1046), .A2(n_1047), .B1(n_1049), .B2(n_1050), .Y(n_1045) );
OAI22xp5_ASAP7_75t_L g1564 ( .A1(n_1047), .A2(n_1565), .B1(n_1566), .B2(n_1568), .Y(n_1564) );
OAI22xp5_ASAP7_75t_L g1572 ( .A1(n_1047), .A2(n_1573), .B1(n_1574), .B2(n_1576), .Y(n_1572) );
INVx2_ASAP7_75t_L g1047 ( .A(n_1048), .Y(n_1047) );
INVx1_ASAP7_75t_L g1567 ( .A(n_1049), .Y(n_1567) );
INVx2_ASAP7_75t_L g1054 ( .A(n_1055), .Y(n_1054) );
AOI21xp5_ASAP7_75t_SL g1057 ( .A1(n_1058), .A2(n_1085), .B(n_1086), .Y(n_1057) );
NAND4xp25_ASAP7_75t_SL g1058 ( .A(n_1059), .B(n_1065), .C(n_1068), .D(n_1072), .Y(n_1058) );
INVx1_ASAP7_75t_L g1061 ( .A(n_1062), .Y(n_1061) );
INVx1_ASAP7_75t_L g1193 ( .A(n_1069), .Y(n_1193) );
OAI221xp5_ASAP7_75t_L g1072 ( .A1(n_1073), .A2(n_1075), .B1(n_1076), .B2(n_1080), .C(n_1081), .Y(n_1072) );
INVx1_ASAP7_75t_L g1073 ( .A(n_1074), .Y(n_1073) );
INVx1_ASAP7_75t_L g1076 ( .A(n_1077), .Y(n_1076) );
INVx1_ASAP7_75t_L g1077 ( .A(n_1078), .Y(n_1077) );
INVx2_ASAP7_75t_L g1078 ( .A(n_1079), .Y(n_1078) );
BUFx2_ASAP7_75t_L g1501 ( .A(n_1083), .Y(n_1501) );
AOI22xp5_ASAP7_75t_L g1229 ( .A1(n_1085), .A2(n_1230), .B1(n_1249), .B2(n_1250), .Y(n_1229) );
INVx1_ASAP7_75t_L g1088 ( .A(n_1089), .Y(n_1088) );
INVx1_ASAP7_75t_L g1091 ( .A(n_1092), .Y(n_1091) );
INVx1_ASAP7_75t_L g1092 ( .A(n_1093), .Y(n_1092) );
XNOR2xp5_ASAP7_75t_L g1093 ( .A(n_1094), .B(n_1095), .Y(n_1093) );
AND2x2_ASAP7_75t_L g1095 ( .A(n_1096), .B(n_1120), .Y(n_1095) );
NAND4xp25_ASAP7_75t_L g1097 ( .A(n_1098), .B(n_1107), .C(n_1113), .D(n_1116), .Y(n_1097) );
BUFx3_ASAP7_75t_L g1497 ( .A(n_1100), .Y(n_1497) );
INVx2_ASAP7_75t_L g1102 ( .A(n_1103), .Y(n_1102) );
INVx3_ASAP7_75t_L g1243 ( .A(n_1103), .Y(n_1243) );
INVx1_ASAP7_75t_L g1110 ( .A(n_1111), .Y(n_1110) );
OAI22xp5_ASAP7_75t_L g1147 ( .A1(n_1115), .A2(n_1117), .B1(n_1135), .B2(n_1148), .Y(n_1147) );
NOR3xp33_ASAP7_75t_SL g1120 ( .A(n_1121), .B(n_1129), .C(n_1133), .Y(n_1120) );
NAND2xp5_ASAP7_75t_L g1121 ( .A(n_1122), .B(n_1126), .Y(n_1121) );
OAI22xp5_ASAP7_75t_L g1134 ( .A1(n_1135), .A2(n_1136), .B1(n_1137), .B2(n_1138), .Y(n_1134) );
CKINVDCx8_ASAP7_75t_R g1143 ( .A(n_1144), .Y(n_1143) );
INVx1_ASAP7_75t_L g1148 ( .A(n_1149), .Y(n_1148) );
INVx1_ASAP7_75t_L g1150 ( .A(n_1151), .Y(n_1150) );
HB1xp67_ASAP7_75t_L g1151 ( .A(n_1152), .Y(n_1151) );
AO22x1_ASAP7_75t_SL g1152 ( .A1(n_1153), .A2(n_1202), .B1(n_1252), .B2(n_1253), .Y(n_1152) );
INVx1_ASAP7_75t_L g1252 ( .A(n_1153), .Y(n_1252) );
NAND4xp25_ASAP7_75t_L g1154 ( .A(n_1155), .B(n_1180), .C(n_1182), .D(n_1197), .Y(n_1154) );
AOI21xp5_ASAP7_75t_L g1157 ( .A1(n_1158), .A2(n_1161), .B(n_1166), .Y(n_1157) );
INVx2_ASAP7_75t_L g1159 ( .A(n_1160), .Y(n_1159) );
INVx1_ASAP7_75t_L g1162 ( .A(n_1163), .Y(n_1162) );
INVx2_ASAP7_75t_L g1164 ( .A(n_1165), .Y(n_1164) );
OAI22xp5_ASAP7_75t_L g1189 ( .A1(n_1168), .A2(n_1169), .B1(n_1190), .B2(n_1192), .Y(n_1189) );
INVx1_ASAP7_75t_L g1172 ( .A(n_1173), .Y(n_1172) );
INVx1_ASAP7_75t_L g1184 ( .A(n_1185), .Y(n_1184) );
INVx1_ASAP7_75t_L g1190 ( .A(n_1191), .Y(n_1190) );
INVx1_ASAP7_75t_L g1192 ( .A(n_1193), .Y(n_1192) );
INVx1_ASAP7_75t_L g1253 ( .A(n_1202), .Y(n_1253) );
XNOR2x1_ASAP7_75t_L g1202 ( .A(n_1203), .B(n_1251), .Y(n_1202) );
NAND2x1_ASAP7_75t_L g1203 ( .A(n_1204), .B(n_1229), .Y(n_1203) );
AND4x1_ASAP7_75t_L g1204 ( .A(n_1205), .B(n_1208), .C(n_1222), .D(n_1225), .Y(n_1204) );
INVx1_ASAP7_75t_L g1213 ( .A(n_1214), .Y(n_1213) );
INVx1_ASAP7_75t_L g1219 ( .A(n_1220), .Y(n_1219) );
NAND3xp33_ASAP7_75t_L g1230 ( .A(n_1231), .B(n_1239), .C(n_1246), .Y(n_1230) );
AOI21xp5_ASAP7_75t_SL g1231 ( .A1(n_1232), .A2(n_1233), .B(n_1234), .Y(n_1231) );
OAI22xp33_ASAP7_75t_L g1338 ( .A1(n_1251), .A2(n_1339), .B1(n_1340), .B2(n_1341), .Y(n_1338) );
OAI221xp5_ASAP7_75t_L g1254 ( .A1(n_1255), .A2(n_1477), .B1(n_1479), .B2(n_1534), .C(n_1540), .Y(n_1254) );
NOR4xp25_ASAP7_75t_L g1255 ( .A(n_1256), .B(n_1404), .C(n_1439), .D(n_1468), .Y(n_1255) );
NAND3xp33_ASAP7_75t_L g1256 ( .A(n_1257), .B(n_1350), .C(n_1376), .Y(n_1256) );
OAI21xp5_ASAP7_75t_L g1257 ( .A1(n_1258), .A2(n_1311), .B(n_1332), .Y(n_1257) );
AOI22xp5_ASAP7_75t_L g1258 ( .A1(n_1259), .A2(n_1302), .B1(n_1306), .B2(n_1310), .Y(n_1258) );
NOR2xp33_ASAP7_75t_L g1259 ( .A(n_1260), .B(n_1280), .Y(n_1259) );
AND2x2_ASAP7_75t_L g1331 ( .A(n_1260), .B(n_1324), .Y(n_1331) );
NOR2xp33_ASAP7_75t_L g1372 ( .A(n_1260), .B(n_1373), .Y(n_1372) );
INVx3_ASAP7_75t_L g1387 ( .A(n_1260), .Y(n_1387) );
NOR2xp33_ASAP7_75t_L g1406 ( .A(n_1260), .B(n_1312), .Y(n_1406) );
AOI21xp5_ASAP7_75t_L g1423 ( .A1(n_1260), .A2(n_1424), .B(n_1425), .Y(n_1423) );
AOI211xp5_ASAP7_75t_L g1440 ( .A1(n_1260), .A2(n_1416), .B(n_1441), .C(n_1446), .Y(n_1440) );
NAND2xp5_ASAP7_75t_L g1472 ( .A(n_1260), .B(n_1368), .Y(n_1472) );
CKINVDCx5p33_ASAP7_75t_R g1260 ( .A(n_1261), .Y(n_1260) );
INVx1_ASAP7_75t_L g1310 ( .A(n_1261), .Y(n_1310) );
INVx1_ASAP7_75t_SL g1317 ( .A(n_1261), .Y(n_1317) );
AND2x2_ASAP7_75t_L g1323 ( .A(n_1261), .B(n_1324), .Y(n_1323) );
AND2x2_ASAP7_75t_L g1354 ( .A(n_1261), .B(n_1318), .Y(n_1354) );
INVx1_ASAP7_75t_L g1367 ( .A(n_1261), .Y(n_1367) );
OR2x2_ASAP7_75t_L g1370 ( .A(n_1261), .B(n_1282), .Y(n_1370) );
NAND2xp5_ASAP7_75t_L g1378 ( .A(n_1261), .B(n_1379), .Y(n_1378) );
AND2x2_ASAP7_75t_L g1394 ( .A(n_1261), .B(n_1355), .Y(n_1394) );
NAND2xp5_ASAP7_75t_L g1430 ( .A(n_1261), .B(n_1282), .Y(n_1430) );
INVx1_ASAP7_75t_L g1443 ( .A(n_1261), .Y(n_1443) );
AND2x2_ASAP7_75t_L g1261 ( .A(n_1262), .B(n_1270), .Y(n_1261) );
INVx1_ASAP7_75t_L g1335 ( .A(n_1263), .Y(n_1335) );
AND2x4_ASAP7_75t_L g1263 ( .A(n_1264), .B(n_1267), .Y(n_1263) );
AND2x2_ASAP7_75t_L g1320 ( .A(n_1264), .B(n_1267), .Y(n_1320) );
HB1xp67_ASAP7_75t_L g1611 ( .A(n_1264), .Y(n_1611) );
INVx1_ASAP7_75t_L g1264 ( .A(n_1265), .Y(n_1264) );
AND2x4_ASAP7_75t_L g1269 ( .A(n_1265), .B(n_1267), .Y(n_1269) );
INVx1_ASAP7_75t_L g1265 ( .A(n_1266), .Y(n_1265) );
NAND2xp5_ASAP7_75t_L g1273 ( .A(n_1266), .B(n_1274), .Y(n_1273) );
INVx1_ASAP7_75t_L g1274 ( .A(n_1268), .Y(n_1274) );
INVx2_ASAP7_75t_L g1337 ( .A(n_1269), .Y(n_1337) );
AND2x4_ASAP7_75t_L g1271 ( .A(n_1272), .B(n_1275), .Y(n_1271) );
INVx1_ASAP7_75t_L g1272 ( .A(n_1273), .Y(n_1272) );
OR2x2_ASAP7_75t_L g1294 ( .A(n_1273), .B(n_1276), .Y(n_1294) );
HB1xp67_ASAP7_75t_L g1613 ( .A(n_1274), .Y(n_1613) );
AND2x4_ASAP7_75t_L g1277 ( .A(n_1275), .B(n_1278), .Y(n_1277) );
INVx1_ASAP7_75t_L g1275 ( .A(n_1276), .Y(n_1275) );
OR2x2_ASAP7_75t_L g1296 ( .A(n_1276), .B(n_1279), .Y(n_1296) );
INVx1_ASAP7_75t_L g1278 ( .A(n_1279), .Y(n_1278) );
AND2x2_ASAP7_75t_L g1280 ( .A(n_1281), .B(n_1289), .Y(n_1280) );
INVx1_ASAP7_75t_L g1325 ( .A(n_1281), .Y(n_1325) );
NAND2xp5_ASAP7_75t_L g1445 ( .A(n_1281), .B(n_1304), .Y(n_1445) );
AND2x2_ASAP7_75t_L g1457 ( .A(n_1281), .B(n_1314), .Y(n_1457) );
AND2x2_ASAP7_75t_L g1281 ( .A(n_1282), .B(n_1285), .Y(n_1281) );
INVx3_ASAP7_75t_L g1309 ( .A(n_1282), .Y(n_1309) );
INVx4_ASAP7_75t_L g1355 ( .A(n_1282), .Y(n_1355) );
NAND2xp5_ASAP7_75t_L g1413 ( .A(n_1282), .B(n_1304), .Y(n_1413) );
AND2x4_ASAP7_75t_L g1282 ( .A(n_1283), .B(n_1284), .Y(n_1282) );
NAND2xp5_ASAP7_75t_L g1391 ( .A(n_1285), .B(n_1366), .Y(n_1391) );
NAND2xp5_ASAP7_75t_L g1396 ( .A(n_1285), .B(n_1297), .Y(n_1396) );
OR2x2_ASAP7_75t_L g1417 ( .A(n_1285), .B(n_1418), .Y(n_1417) );
NOR2xp33_ASAP7_75t_L g1426 ( .A(n_1285), .B(n_1297), .Y(n_1426) );
OR2x2_ASAP7_75t_L g1475 ( .A(n_1285), .B(n_1386), .Y(n_1475) );
BUFx3_ASAP7_75t_L g1285 ( .A(n_1286), .Y(n_1285) );
AND2x2_ASAP7_75t_L g1303 ( .A(n_1286), .B(n_1304), .Y(n_1303) );
INVx2_ASAP7_75t_L g1307 ( .A(n_1286), .Y(n_1307) );
AND2x2_ASAP7_75t_L g1313 ( .A(n_1286), .B(n_1314), .Y(n_1313) );
AND2x2_ASAP7_75t_L g1357 ( .A(n_1286), .B(n_1358), .Y(n_1357) );
AND2x2_ASAP7_75t_L g1424 ( .A(n_1286), .B(n_1386), .Y(n_1424) );
OR2x2_ASAP7_75t_L g1433 ( .A(n_1286), .B(n_1422), .Y(n_1433) );
AND2x2_ASAP7_75t_L g1286 ( .A(n_1287), .B(n_1288), .Y(n_1286) );
NAND2xp5_ASAP7_75t_L g1308 ( .A(n_1289), .B(n_1309), .Y(n_1308) );
AOI21xp5_ASAP7_75t_L g1392 ( .A1(n_1289), .A2(n_1354), .B(n_1393), .Y(n_1392) );
INVx1_ASAP7_75t_L g1418 ( .A(n_1289), .Y(n_1418) );
NAND2xp5_ASAP7_75t_L g1461 ( .A(n_1289), .B(n_1380), .Y(n_1461) );
AND2x2_ASAP7_75t_L g1289 ( .A(n_1290), .B(n_1297), .Y(n_1289) );
INVx1_ASAP7_75t_L g1305 ( .A(n_1290), .Y(n_1305) );
AND2x2_ASAP7_75t_L g1314 ( .A(n_1290), .B(n_1298), .Y(n_1314) );
INVx1_ASAP7_75t_L g1386 ( .A(n_1290), .Y(n_1386) );
OAI22xp33_ASAP7_75t_L g1291 ( .A1(n_1292), .A2(n_1293), .B1(n_1295), .B2(n_1296), .Y(n_1291) );
OAI22xp5_ASAP7_75t_L g1299 ( .A1(n_1293), .A2(n_1296), .B1(n_1300), .B2(n_1301), .Y(n_1299) );
BUFx3_ASAP7_75t_L g1339 ( .A(n_1293), .Y(n_1339) );
OAI22xp33_ASAP7_75t_L g1346 ( .A1(n_1293), .A2(n_1347), .B1(n_1348), .B2(n_1349), .Y(n_1346) );
BUFx6f_ASAP7_75t_L g1293 ( .A(n_1294), .Y(n_1293) );
INVx1_ASAP7_75t_L g1342 ( .A(n_1296), .Y(n_1342) );
HB1xp67_ASAP7_75t_L g1349 ( .A(n_1296), .Y(n_1349) );
AND2x2_ASAP7_75t_L g1327 ( .A(n_1297), .B(n_1307), .Y(n_1327) );
AND2x2_ASAP7_75t_L g1358 ( .A(n_1297), .B(n_1305), .Y(n_1358) );
INVx2_ASAP7_75t_L g1366 ( .A(n_1297), .Y(n_1366) );
INVx2_ASAP7_75t_L g1297 ( .A(n_1298), .Y(n_1297) );
AND2x2_ASAP7_75t_L g1304 ( .A(n_1298), .B(n_1305), .Y(n_1304) );
AOI21xp33_ASAP7_75t_SL g1435 ( .A1(n_1302), .A2(n_1436), .B(n_1437), .Y(n_1435) );
INVx1_ASAP7_75t_L g1302 ( .A(n_1303), .Y(n_1302) );
AND2x2_ASAP7_75t_L g1379 ( .A(n_1304), .B(n_1380), .Y(n_1379) );
INVx1_ASAP7_75t_L g1422 ( .A(n_1304), .Y(n_1422) );
OR2x2_ASAP7_75t_L g1306 ( .A(n_1307), .B(n_1308), .Y(n_1306) );
NAND2xp5_ASAP7_75t_L g1375 ( .A(n_1307), .B(n_1358), .Y(n_1375) );
AND2x2_ASAP7_75t_L g1380 ( .A(n_1307), .B(n_1355), .Y(n_1380) );
NOR2x1_ASAP7_75t_L g1400 ( .A(n_1307), .B(n_1386), .Y(n_1400) );
NAND4xp25_ASAP7_75t_L g1401 ( .A(n_1307), .B(n_1330), .C(n_1360), .D(n_1402), .Y(n_1401) );
AND2x2_ASAP7_75t_L g1411 ( .A(n_1307), .B(n_1412), .Y(n_1411) );
AND2x2_ASAP7_75t_L g1467 ( .A(n_1307), .B(n_1314), .Y(n_1467) );
INVx2_ASAP7_75t_L g1330 ( .A(n_1309), .Y(n_1330) );
NAND2xp5_ASAP7_75t_L g1373 ( .A(n_1309), .B(n_1357), .Y(n_1373) );
AND2x2_ASAP7_75t_L g1415 ( .A(n_1309), .B(n_1313), .Y(n_1415) );
AND2x2_ASAP7_75t_L g1452 ( .A(n_1309), .B(n_1426), .Y(n_1452) );
OR2x2_ASAP7_75t_L g1469 ( .A(n_1309), .B(n_1375), .Y(n_1469) );
OAI221xp5_ASAP7_75t_L g1311 ( .A1(n_1312), .A2(n_1315), .B1(n_1322), .B2(n_1325), .C(n_1326), .Y(n_1311) );
INVx1_ASAP7_75t_L g1312 ( .A(n_1313), .Y(n_1312) );
NAND2xp5_ASAP7_75t_L g1352 ( .A(n_1314), .B(n_1353), .Y(n_1352) );
INVx1_ASAP7_75t_L g1403 ( .A(n_1314), .Y(n_1403) );
OAI321xp33_ASAP7_75t_L g1395 ( .A1(n_1315), .A2(n_1383), .A3(n_1396), .B1(n_1397), .B2(n_1398), .C(n_1401), .Y(n_1395) );
INVx1_ASAP7_75t_L g1315 ( .A(n_1316), .Y(n_1315) );
AND2x2_ASAP7_75t_L g1389 ( .A(n_1316), .B(n_1390), .Y(n_1389) );
AND2x2_ASAP7_75t_L g1316 ( .A(n_1317), .B(n_1318), .Y(n_1316) );
NAND2xp5_ASAP7_75t_L g1397 ( .A(n_1317), .B(n_1381), .Y(n_1397) );
CKINVDCx6p67_ASAP7_75t_R g1324 ( .A(n_1318), .Y(n_1324) );
AND2x2_ASAP7_75t_L g1360 ( .A(n_1318), .B(n_1361), .Y(n_1360) );
OAI221xp5_ASAP7_75t_L g1454 ( .A1(n_1318), .A2(n_1385), .B1(n_1451), .B2(n_1455), .C(n_1456), .Y(n_1454) );
NAND2xp5_ASAP7_75t_L g1470 ( .A(n_1318), .B(n_1471), .Y(n_1470) );
OR2x6_ASAP7_75t_L g1318 ( .A(n_1319), .B(n_1321), .Y(n_1318) );
NOR2xp33_ASAP7_75t_L g1374 ( .A(n_1322), .B(n_1375), .Y(n_1374) );
INVx1_ASAP7_75t_L g1322 ( .A(n_1323), .Y(n_1322) );
NAND2xp5_ASAP7_75t_L g1455 ( .A(n_1323), .B(n_1355), .Y(n_1455) );
NAND2xp5_ASAP7_75t_L g1456 ( .A(n_1323), .B(n_1457), .Y(n_1456) );
AND2x4_ASAP7_75t_SL g1368 ( .A(n_1324), .B(n_1361), .Y(n_1368) );
AND2x2_ASAP7_75t_L g1381 ( .A(n_1324), .B(n_1345), .Y(n_1381) );
OR2x2_ASAP7_75t_L g1408 ( .A(n_1324), .B(n_1361), .Y(n_1408) );
NAND2xp5_ASAP7_75t_L g1428 ( .A(n_1324), .B(n_1429), .Y(n_1428) );
AND2x2_ASAP7_75t_L g1434 ( .A(n_1324), .B(n_1365), .Y(n_1434) );
NOR2xp33_ASAP7_75t_L g1448 ( .A(n_1324), .B(n_1449), .Y(n_1448) );
NAND2xp5_ASAP7_75t_L g1465 ( .A(n_1324), .B(n_1438), .Y(n_1465) );
NAND2xp5_ASAP7_75t_L g1326 ( .A(n_1327), .B(n_1328), .Y(n_1326) );
INVx1_ASAP7_75t_L g1328 ( .A(n_1329), .Y(n_1328) );
NAND2xp5_ASAP7_75t_L g1329 ( .A(n_1330), .B(n_1331), .Y(n_1329) );
INVx1_ASAP7_75t_L g1437 ( .A(n_1331), .Y(n_1437) );
NOR2xp33_ASAP7_75t_L g1332 ( .A(n_1333), .B(n_1343), .Y(n_1332) );
OAI31xp33_ASAP7_75t_L g1350 ( .A1(n_1333), .A2(n_1351), .A3(n_1372), .B(n_1374), .Y(n_1350) );
AOI221xp5_ASAP7_75t_L g1376 ( .A1(n_1333), .A2(n_1377), .B1(n_1381), .B2(n_1382), .C(n_1395), .Y(n_1376) );
BUFx3_ASAP7_75t_L g1438 ( .A(n_1333), .Y(n_1438) );
NAND2xp5_ASAP7_75t_L g1459 ( .A(n_1333), .B(n_1343), .Y(n_1459) );
INVx1_ASAP7_75t_L g1471 ( .A(n_1333), .Y(n_1471) );
INVx1_ASAP7_75t_L g1334 ( .A(n_1335), .Y(n_1334) );
INVx2_ASAP7_75t_L g1336 ( .A(n_1337), .Y(n_1336) );
INVx1_ASAP7_75t_L g1478 ( .A(n_1337), .Y(n_1478) );
INVx1_ASAP7_75t_L g1341 ( .A(n_1342), .Y(n_1341) );
NOR3xp33_ASAP7_75t_L g1369 ( .A(n_1343), .B(n_1370), .C(n_1371), .Y(n_1369) );
NAND2xp5_ASAP7_75t_L g1420 ( .A(n_1343), .B(n_1387), .Y(n_1420) );
INVx2_ASAP7_75t_L g1343 ( .A(n_1344), .Y(n_1343) );
AND2x2_ASAP7_75t_L g1353 ( .A(n_1344), .B(n_1354), .Y(n_1353) );
OAI322xp33_ASAP7_75t_L g1382 ( .A1(n_1344), .A2(n_1383), .A3(n_1385), .B1(n_1387), .B2(n_1388), .C1(n_1391), .C2(n_1392), .Y(n_1382) );
INVx2_ASAP7_75t_L g1390 ( .A(n_1344), .Y(n_1390) );
NAND3xp33_ASAP7_75t_L g1466 ( .A(n_1344), .B(n_1394), .C(n_1467), .Y(n_1466) );
INVx2_ASAP7_75t_L g1344 ( .A(n_1345), .Y(n_1344) );
INVx2_ASAP7_75t_SL g1361 ( .A(n_1345), .Y(n_1361) );
OAI221xp5_ASAP7_75t_L g1351 ( .A1(n_1352), .A2(n_1355), .B1(n_1356), .B2(n_1359), .C(n_1362), .Y(n_1351) );
INVx1_ASAP7_75t_L g1450 ( .A(n_1353), .Y(n_1450) );
AND2x2_ASAP7_75t_L g1476 ( .A(n_1354), .B(n_1355), .Y(n_1476) );
INVx1_ASAP7_75t_L g1365 ( .A(n_1355), .Y(n_1365) );
NOR2xp33_ASAP7_75t_L g1384 ( .A(n_1355), .B(n_1361), .Y(n_1384) );
AND2x2_ASAP7_75t_L g1399 ( .A(n_1355), .B(n_1400), .Y(n_1399) );
NAND2xp5_ASAP7_75t_L g1432 ( .A(n_1356), .B(n_1433), .Y(n_1432) );
INVx1_ASAP7_75t_L g1356 ( .A(n_1357), .Y(n_1356) );
OAI21xp5_ASAP7_75t_L g1473 ( .A1(n_1357), .A2(n_1474), .B(n_1476), .Y(n_1473) );
INVx1_ASAP7_75t_L g1371 ( .A(n_1358), .Y(n_1371) );
AND2x2_ASAP7_75t_L g1393 ( .A(n_1358), .B(n_1394), .Y(n_1393) );
NAND2xp5_ASAP7_75t_L g1436 ( .A(n_1358), .B(n_1380), .Y(n_1436) );
INVx2_ASAP7_75t_L g1359 ( .A(n_1360), .Y(n_1359) );
NAND2xp5_ASAP7_75t_L g1463 ( .A(n_1361), .B(n_1387), .Y(n_1463) );
AOI21xp5_ASAP7_75t_L g1362 ( .A1(n_1363), .A2(n_1368), .B(n_1369), .Y(n_1362) );
INVxp67_ASAP7_75t_SL g1363 ( .A(n_1364), .Y(n_1363) );
NAND3xp33_ASAP7_75t_L g1364 ( .A(n_1365), .B(n_1366), .C(n_1367), .Y(n_1364) );
AND2x2_ASAP7_75t_L g1425 ( .A(n_1365), .B(n_1426), .Y(n_1425) );
NAND2xp5_ASAP7_75t_L g1402 ( .A(n_1371), .B(n_1403), .Y(n_1402) );
INVx1_ASAP7_75t_L g1446 ( .A(n_1373), .Y(n_1446) );
INVx1_ASAP7_75t_L g1377 ( .A(n_1378), .Y(n_1377) );
INVx1_ASAP7_75t_L g1464 ( .A(n_1379), .Y(n_1464) );
INVx1_ASAP7_75t_L g1427 ( .A(n_1381), .Y(n_1427) );
INVx1_ASAP7_75t_L g1383 ( .A(n_1384), .Y(n_1383) );
INVx1_ASAP7_75t_L g1385 ( .A(n_1386), .Y(n_1385) );
NOR2xp33_ASAP7_75t_L g1409 ( .A(n_1387), .B(n_1410), .Y(n_1409) );
O2A1O1Ixp33_ASAP7_75t_L g1462 ( .A1(n_1387), .A2(n_1407), .B(n_1438), .C(n_1463), .Y(n_1462) );
OAI221xp5_ASAP7_75t_L g1421 ( .A1(n_1388), .A2(n_1422), .B1(n_1423), .B2(n_1427), .C(n_1428), .Y(n_1421) );
INVx1_ASAP7_75t_L g1388 ( .A(n_1389), .Y(n_1388) );
NOR2xp33_ASAP7_75t_L g1429 ( .A(n_1396), .B(n_1430), .Y(n_1429) );
INVx1_ASAP7_75t_L g1398 ( .A(n_1399), .Y(n_1398) );
AOI31xp33_ASAP7_75t_L g1404 ( .A1(n_1405), .A2(n_1414), .A3(n_1431), .B(n_1438), .Y(n_1404) );
AOI21xp5_ASAP7_75t_L g1405 ( .A1(n_1406), .A2(n_1407), .B(n_1409), .Y(n_1405) );
INVx1_ASAP7_75t_L g1407 ( .A(n_1408), .Y(n_1407) );
INVx1_ASAP7_75t_L g1410 ( .A(n_1411), .Y(n_1410) );
INVx1_ASAP7_75t_L g1412 ( .A(n_1413), .Y(n_1412) );
O2A1O1Ixp33_ASAP7_75t_L g1414 ( .A1(n_1415), .A2(n_1416), .B(n_1419), .C(n_1421), .Y(n_1414) );
INVx1_ASAP7_75t_L g1416 ( .A(n_1417), .Y(n_1416) );
INVx1_ASAP7_75t_L g1419 ( .A(n_1420), .Y(n_1419) );
AOI21xp33_ASAP7_75t_L g1431 ( .A1(n_1432), .A2(n_1434), .B(n_1435), .Y(n_1431) );
OAI221xp5_ASAP7_75t_L g1468 ( .A1(n_1433), .A2(n_1469), .B1(n_1470), .B2(n_1472), .C(n_1473), .Y(n_1468) );
INVx2_ASAP7_75t_L g1449 ( .A(n_1438), .Y(n_1449) );
OAI221xp5_ASAP7_75t_SL g1439 ( .A1(n_1440), .A2(n_1447), .B1(n_1450), .B2(n_1451), .C(n_1453), .Y(n_1439) );
AND2x2_ASAP7_75t_L g1441 ( .A(n_1442), .B(n_1444), .Y(n_1441) );
INVx1_ASAP7_75t_L g1442 ( .A(n_1443), .Y(n_1442) );
INVx1_ASAP7_75t_L g1444 ( .A(n_1445), .Y(n_1444) );
INVxp67_ASAP7_75t_L g1447 ( .A(n_1448), .Y(n_1447) );
INVx1_ASAP7_75t_L g1451 ( .A(n_1452), .Y(n_1451) );
AOI21xp5_ASAP7_75t_SL g1453 ( .A1(n_1454), .A2(n_1458), .B(n_1460), .Y(n_1453) );
INVx1_ASAP7_75t_L g1458 ( .A(n_1459), .Y(n_1458) );
OAI221xp5_ASAP7_75t_L g1460 ( .A1(n_1461), .A2(n_1462), .B1(n_1464), .B2(n_1465), .C(n_1466), .Y(n_1460) );
INVx1_ASAP7_75t_L g1474 ( .A(n_1475), .Y(n_1474) );
INVx1_ASAP7_75t_L g1477 ( .A(n_1478), .Y(n_1477) );
INVx1_ASAP7_75t_L g1479 ( .A(n_1480), .Y(n_1479) );
INVx1_ASAP7_75t_L g1480 ( .A(n_1481), .Y(n_1480) );
AND3x1_ASAP7_75t_L g1482 ( .A(n_1483), .B(n_1506), .C(n_1508), .Y(n_1482) );
NOR2xp33_ASAP7_75t_L g1483 ( .A(n_1484), .B(n_1491), .Y(n_1483) );
NAND2xp5_ASAP7_75t_L g1484 ( .A(n_1485), .B(n_1488), .Y(n_1484) );
INVx1_ASAP7_75t_L g1503 ( .A(n_1504), .Y(n_1503) );
INVx2_ASAP7_75t_L g1511 ( .A(n_1512), .Y(n_1511) );
INVx2_ASAP7_75t_L g1512 ( .A(n_1513), .Y(n_1512) );
HB1xp67_ASAP7_75t_L g1517 ( .A(n_1518), .Y(n_1517) );
OAI22xp5_ASAP7_75t_SL g1520 ( .A1(n_1521), .A2(n_1522), .B1(n_1523), .B2(n_1524), .Y(n_1520) );
INVx1_ASAP7_75t_L g1524 ( .A(n_1525), .Y(n_1524) );
INVx1_ASAP7_75t_L g1525 ( .A(n_1526), .Y(n_1525) );
INVx2_ASAP7_75t_L g1530 ( .A(n_1531), .Y(n_1530) );
INVx1_ASAP7_75t_SL g1534 ( .A(n_1535), .Y(n_1534) );
INVx1_ASAP7_75t_L g1535 ( .A(n_1536), .Y(n_1535) );
INVx1_ASAP7_75t_L g1536 ( .A(n_1537), .Y(n_1536) );
INVx1_ASAP7_75t_L g1537 ( .A(n_1538), .Y(n_1537) );
INVx1_ASAP7_75t_L g1538 ( .A(n_1539), .Y(n_1538) );
INVx1_ASAP7_75t_L g1541 ( .A(n_1542), .Y(n_1541) );
CKINVDCx5p33_ASAP7_75t_R g1542 ( .A(n_1543), .Y(n_1542) );
A2O1A1Ixp33_ASAP7_75t_L g1609 ( .A1(n_1544), .A2(n_1610), .B(n_1612), .C(n_1614), .Y(n_1609) );
INVxp33_ASAP7_75t_SL g1545 ( .A(n_1546), .Y(n_1545) );
HB1xp67_ASAP7_75t_L g1547 ( .A(n_1548), .Y(n_1547) );
INVx1_ASAP7_75t_L g1548 ( .A(n_1549), .Y(n_1548) );
NOR3xp33_ASAP7_75t_L g1551 ( .A(n_1552), .B(n_1559), .C(n_1563), .Y(n_1551) );
NAND2xp5_ASAP7_75t_L g1552 ( .A(n_1553), .B(n_1556), .Y(n_1552) );
OAI221xp5_ASAP7_75t_L g1598 ( .A1(n_1554), .A2(n_1558), .B1(n_1588), .B2(n_1599), .C(n_1601), .Y(n_1598) );
INVx2_ASAP7_75t_L g1560 ( .A(n_1561), .Y(n_1560) );
INVx2_ASAP7_75t_SL g1566 ( .A(n_1567), .Y(n_1566) );
OAI221xp5_ASAP7_75t_L g1585 ( .A1(n_1568), .A2(n_1570), .B1(n_1586), .B2(n_1588), .C(n_1589), .Y(n_1585) );
INVx1_ASAP7_75t_L g1574 ( .A(n_1575), .Y(n_1574) );
INVx1_ASAP7_75t_L g1579 ( .A(n_1580), .Y(n_1579) );
OAI31xp33_ASAP7_75t_L g1582 ( .A1(n_1583), .A2(n_1592), .A3(n_1605), .B(n_1606), .Y(n_1582) );
INVx1_ASAP7_75t_L g1586 ( .A(n_1587), .Y(n_1586) );
INVx1_ASAP7_75t_L g1599 ( .A(n_1600), .Y(n_1599) );
INVx1_ASAP7_75t_L g1602 ( .A(n_1603), .Y(n_1602) );
BUFx2_ASAP7_75t_L g1607 ( .A(n_1608), .Y(n_1607) );
HB1xp67_ASAP7_75t_L g1608 ( .A(n_1609), .Y(n_1608) );
INVx1_ASAP7_75t_L g1610 ( .A(n_1611), .Y(n_1610) );
INVx1_ASAP7_75t_L g1612 ( .A(n_1613), .Y(n_1612) );
endmodule