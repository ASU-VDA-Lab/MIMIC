module fake_jpeg_17623_n_227 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_227);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_227;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx6_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx16f_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx6_ASAP7_75t_SL g30 ( 
.A(n_1),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

INVx3_ASAP7_75t_SL g34 ( 
.A(n_16),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_34),
.B(n_41),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx2_ASAP7_75t_SL g37 ( 
.A(n_30),
.Y(n_37)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

BUFx8_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

CKINVDCx16_ASAP7_75t_R g46 ( 
.A(n_38),
.Y(n_46)
);

BUFx16f_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_22),
.B(n_2),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_18),
.B(n_2),
.Y(n_42)
);

A2O1A1Ixp33_ASAP7_75t_L g58 ( 
.A1(n_42),
.A2(n_21),
.B(n_24),
.C(n_23),
.Y(n_58)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_38),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_49),
.B(n_54),
.Y(n_63)
);

CKINVDCx12_ASAP7_75t_R g50 ( 
.A(n_39),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_52),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_34),
.A2(n_18),
.B1(n_31),
.B2(n_16),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_53),
.A2(n_34),
.B1(n_37),
.B2(n_40),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_38),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_34),
.A2(n_31),
.B1(n_22),
.B2(n_30),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_56),
.A2(n_40),
.B1(n_37),
.B2(n_36),
.Y(n_87)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_57),
.Y(n_60)
);

OR2x4_ASAP7_75t_L g73 ( 
.A(n_58),
.B(n_39),
.Y(n_73)
);

A2O1A1Ixp33_ASAP7_75t_L g61 ( 
.A1(n_48),
.A2(n_41),
.B(n_42),
.C(n_39),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_61),
.B(n_67),
.Y(n_90)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_62),
.Y(n_93)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_55),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_64),
.B(n_72),
.Y(n_100)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_65),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_48),
.B(n_41),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_58),
.B(n_38),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_68),
.B(n_80),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_49),
.B(n_39),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_70),
.A2(n_85),
.B(n_86),
.Y(n_92)
);

OR2x2_ASAP7_75t_L g71 ( 
.A(n_58),
.B(n_25),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_71),
.B(n_76),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_47),
.Y(n_72)
);

NAND2xp33_ASAP7_75t_SL g91 ( 
.A(n_73),
.B(n_83),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_SL g74 ( 
.A1(n_46),
.A2(n_39),
.B(n_38),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_74),
.A2(n_27),
.B(n_51),
.Y(n_106)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_52),
.Y(n_75)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_75),
.Y(n_94)
);

OR2x2_ASAP7_75t_L g76 ( 
.A(n_44),
.B(n_25),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_50),
.Y(n_77)
);

HB1xp67_ASAP7_75t_L g98 ( 
.A(n_77),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_44),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_78),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_79),
.A2(n_87),
.B1(n_27),
.B2(n_28),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_54),
.B(n_38),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_47),
.Y(n_81)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_81),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_55),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_82),
.Y(n_97)
);

OR2x2_ASAP7_75t_L g83 ( 
.A(n_46),
.B(n_26),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_43),
.A2(n_34),
.B1(n_40),
.B2(n_17),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_84),
.A2(n_37),
.B1(n_36),
.B2(n_51),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_57),
.B(n_38),
.Y(n_85)
);

OR2x2_ASAP7_75t_L g86 ( 
.A(n_55),
.B(n_33),
.Y(n_86)
);

OA22x2_ASAP7_75t_L g88 ( 
.A1(n_73),
.A2(n_35),
.B1(n_37),
.B2(n_47),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_88),
.B(n_96),
.Y(n_123)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_62),
.Y(n_95)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_95),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_68),
.A2(n_36),
.B1(n_20),
.B2(n_32),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_101),
.B(n_108),
.Y(n_117)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_65),
.Y(n_102)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_102),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_67),
.B(n_3),
.Y(n_104)
);

XNOR2x1_ASAP7_75t_L g120 ( 
.A(n_104),
.B(n_106),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_61),
.B(n_51),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_105),
.B(n_71),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_74),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_87),
.A2(n_20),
.B1(n_32),
.B2(n_28),
.Y(n_109)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_109),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_70),
.A2(n_85),
.B1(n_86),
.B2(n_83),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_110),
.B(n_80),
.C(n_63),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_112),
.B(n_76),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_113),
.B(n_126),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_114),
.B(n_127),
.C(n_128),
.Y(n_159)
);

AND2x6_ASAP7_75t_L g115 ( 
.A(n_108),
.B(n_70),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_115),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_99),
.B(n_66),
.C(n_85),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_116),
.B(n_133),
.C(n_103),
.Y(n_149)
);

BUFx2_ASAP7_75t_L g118 ( 
.A(n_102),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_118),
.B(n_130),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_121),
.A2(n_104),
.B1(n_88),
.B2(n_91),
.Y(n_143)
);

OAI32xp33_ASAP7_75t_L g124 ( 
.A1(n_99),
.A2(n_78),
.A3(n_64),
.B1(n_33),
.B2(n_26),
.Y(n_124)
);

CKINVDCx14_ASAP7_75t_R g155 ( 
.A(n_124),
.Y(n_155)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_100),
.Y(n_125)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_125),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_90),
.B(n_75),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_90),
.B(n_92),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_92),
.B(n_69),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_94),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_129),
.B(n_131),
.Y(n_154)
);

INVx11_ASAP7_75t_L g130 ( 
.A(n_95),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_94),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_105),
.B(n_69),
.C(n_19),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_107),
.B(n_10),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_134),
.B(n_135),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_98),
.B(n_13),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_97),
.B(n_60),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_136),
.Y(n_137)
);

OAI22xp33_ASAP7_75t_L g138 ( 
.A1(n_122),
.A2(n_81),
.B1(n_106),
.B2(n_60),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_138),
.Y(n_160)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_132),
.Y(n_139)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_139),
.Y(n_173)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_132),
.Y(n_141)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_141),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_143),
.B(n_147),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_126),
.B(n_127),
.Y(n_144)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_144),
.Y(n_177)
);

AO22x1_ASAP7_75t_L g145 ( 
.A1(n_123),
.A2(n_88),
.B1(n_110),
.B2(n_109),
.Y(n_145)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_145),
.Y(n_170)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_119),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_113),
.B(n_104),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_148),
.B(n_124),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_149),
.B(n_150),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_128),
.B(n_89),
.C(n_93),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_125),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_151),
.B(n_152),
.Y(n_163)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_118),
.Y(n_152)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_130),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_157),
.B(n_111),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_116),
.B(n_89),
.C(n_111),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_158),
.B(n_133),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_156),
.A2(n_144),
.B(n_120),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_164),
.A2(n_172),
.B(n_176),
.Y(n_181)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_165),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_153),
.B(n_114),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_166),
.B(n_167),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_146),
.B(n_120),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_169),
.B(n_158),
.C(n_149),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_171),
.B(n_174),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_155),
.A2(n_123),
.B(n_117),
.Y(n_172)
);

NAND3xp33_ASAP7_75t_L g174 ( 
.A(n_148),
.B(n_115),
.C(n_88),
.Y(n_174)
);

MAJx2_ASAP7_75t_L g175 ( 
.A(n_159),
.B(n_123),
.C(n_122),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_175),
.B(n_159),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_138),
.B(n_97),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_164),
.A2(n_143),
.B(n_154),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_179),
.A2(n_176),
.B(n_170),
.Y(n_200)
);

MAJx2_ASAP7_75t_L g201 ( 
.A(n_180),
.B(n_177),
.C(n_170),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_162),
.B(n_150),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_182),
.B(n_183),
.C(n_184),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_162),
.B(n_169),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_163),
.B(n_146),
.Y(n_185)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_185),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_177),
.B(n_142),
.C(n_137),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_186),
.B(n_171),
.Y(n_195)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_168),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_188),
.Y(n_202)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_168),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_189),
.A2(n_191),
.B1(n_140),
.B2(n_139),
.Y(n_198)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_173),
.Y(n_191)
);

NOR2x1_ASAP7_75t_L g192 ( 
.A(n_181),
.B(n_161),
.Y(n_192)
);

OR2x2_ASAP7_75t_L g205 ( 
.A(n_192),
.B(n_190),
.Y(n_205)
);

XNOR2x1_ASAP7_75t_L g194 ( 
.A(n_181),
.B(n_175),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_194),
.B(n_200),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_195),
.B(n_197),
.C(n_201),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_182),
.B(n_172),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_198),
.B(n_178),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_187),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_199),
.B(n_186),
.Y(n_207)
);

AOI322xp5_ASAP7_75t_L g212 ( 
.A1(n_204),
.A2(n_196),
.A3(n_194),
.B1(n_199),
.B2(n_201),
.C1(n_145),
.C2(n_14),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_205),
.B(n_207),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_202),
.A2(n_160),
.B1(n_176),
.B2(n_141),
.Y(n_206)
);

A2O1A1Ixp33_ASAP7_75t_SL g214 ( 
.A1(n_206),
.A2(n_59),
.B(n_4),
.C(n_5),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_192),
.A2(n_142),
.B(n_180),
.Y(n_208)
);

MAJx2_ASAP7_75t_L g213 ( 
.A(n_208),
.B(n_15),
.C(n_13),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_193),
.B(n_184),
.C(n_183),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_210),
.B(n_211),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_193),
.B(n_19),
.C(n_145),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_212),
.A2(n_213),
.B1(n_214),
.B2(n_3),
.Y(n_221)
);

AOI322xp5_ASAP7_75t_L g215 ( 
.A1(n_207),
.A2(n_59),
.A3(n_4),
.B1(n_5),
.B2(n_6),
.C1(n_3),
.C2(n_8),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_215),
.B(n_216),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_218),
.A2(n_219),
.B1(n_221),
.B2(n_6),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_217),
.B(n_206),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_214),
.B(n_203),
.C(n_209),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_220),
.Y(n_223)
);

AOI21x1_ASAP7_75t_L g222 ( 
.A1(n_220),
.A2(n_5),
.B(n_6),
.Y(n_222)
);

AOI322xp5_ASAP7_75t_L g225 ( 
.A1(n_222),
.A2(n_7),
.A3(n_9),
.B1(n_223),
.B2(n_221),
.C1(n_224),
.C2(n_218),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_225),
.B(n_7),
.Y(n_226)
);

BUFx24_ASAP7_75t_SL g227 ( 
.A(n_226),
.Y(n_227)
);


endmodule