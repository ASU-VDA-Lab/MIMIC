module real_aes_6814_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_357;
wire n_287;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_555;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_545;
wire n_341;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_666;
wire n_320;
wire n_551;
wire n_537;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_656;
wire n_532;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_649;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_119;
wire n_310;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_417;
wire n_363;
wire n_754;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_756;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_728;
wire n_713;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_749;
wire n_162;
wire n_358;
wire n_275;
wire n_214;
wire n_385;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_481;
wire n_148;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_546;
wire n_151;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_424;
wire n_225;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g113 ( .A(n_0), .Y(n_113) );
A2O1A1Ixp33_ASAP7_75t_L g234 ( .A1(n_1), .A2(n_152), .B(n_155), .C(n_235), .Y(n_234) );
AOI21xp5_ASAP7_75t_L g201 ( .A1(n_2), .A2(n_181), .B(n_202), .Y(n_201) );
INVx1_ASAP7_75t_L g512 ( .A(n_3), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_4), .B(n_211), .Y(n_210) );
AOI21xp33_ASAP7_75t_L g495 ( .A1(n_5), .A2(n_181), .B(n_496), .Y(n_495) );
AND2x6_ASAP7_75t_L g152 ( .A(n_6), .B(n_153), .Y(n_152) );
INVx1_ASAP7_75t_L g248 ( .A(n_7), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g110 ( .A(n_8), .B(n_43), .Y(n_110) );
NOR2xp33_ASAP7_75t_L g447 ( .A(n_8), .B(n_43), .Y(n_447) );
AOI21xp5_ASAP7_75t_L g542 ( .A1(n_9), .A2(n_180), .B(n_543), .Y(n_542) );
NAND2xp5_ASAP7_75t_SL g237 ( .A(n_10), .B(n_164), .Y(n_237) );
INVx1_ASAP7_75t_L g500 ( .A(n_11), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_12), .B(n_205), .Y(n_535) );
OAI22xp5_ASAP7_75t_SL g454 ( .A1(n_13), .A2(n_455), .B1(n_456), .B2(n_462), .Y(n_454) );
CKINVDCx20_ASAP7_75t_R g462 ( .A(n_13), .Y(n_462) );
INVx1_ASAP7_75t_L g144 ( .A(n_14), .Y(n_144) );
INVx1_ASAP7_75t_L g547 ( .A(n_15), .Y(n_547) );
OAI22xp5_ASAP7_75t_L g459 ( .A1(n_16), .A2(n_80), .B1(n_460), .B2(n_461), .Y(n_459) );
CKINVDCx20_ASAP7_75t_R g460 ( .A(n_16), .Y(n_460) );
A2O1A1Ixp33_ASAP7_75t_L g269 ( .A1(n_17), .A2(n_189), .B(n_270), .C(n_272), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_18), .B(n_211), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_19), .B(n_478), .Y(n_557) );
NAND2xp5_ASAP7_75t_SL g521 ( .A(n_20), .B(n_181), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_21), .B(n_195), .Y(n_194) );
A2O1A1Ixp33_ASAP7_75t_L g255 ( .A1(n_22), .A2(n_205), .B(n_256), .C(n_258), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_23), .B(n_211), .Y(n_481) );
NAND2xp5_ASAP7_75t_SL g163 ( .A(n_24), .B(n_164), .Y(n_163) );
A2O1A1Ixp33_ASAP7_75t_L g545 ( .A1(n_25), .A2(n_191), .B(n_272), .C(n_546), .Y(n_545) );
NAND2xp5_ASAP7_75t_SL g219 ( .A(n_26), .B(n_164), .Y(n_219) );
CKINVDCx16_ASAP7_75t_R g146 ( .A(n_27), .Y(n_146) );
INVx1_ASAP7_75t_L g218 ( .A(n_28), .Y(n_218) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_29), .Y(n_151) );
CKINVDCx20_ASAP7_75t_R g233 ( .A(n_30), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_31), .B(n_164), .Y(n_513) );
NAND2xp5_ASAP7_75t_SL g448 ( .A(n_32), .B(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g187 ( .A(n_33), .Y(n_187) );
INVx1_ASAP7_75t_L g490 ( .A(n_34), .Y(n_490) );
AOI22xp5_ASAP7_75t_L g456 ( .A1(n_35), .A2(n_457), .B1(n_458), .B2(n_459), .Y(n_456) );
CKINVDCx20_ASAP7_75t_R g457 ( .A(n_35), .Y(n_457) );
INVx2_ASAP7_75t_L g150 ( .A(n_36), .Y(n_150) );
CKINVDCx20_ASAP7_75t_R g239 ( .A(n_37), .Y(n_239) );
A2O1A1Ixp33_ASAP7_75t_L g204 ( .A1(n_38), .A2(n_205), .B(n_206), .C(n_208), .Y(n_204) );
INVxp67_ASAP7_75t_L g190 ( .A(n_39), .Y(n_190) );
CKINVDCx14_ASAP7_75t_R g203 ( .A(n_40), .Y(n_203) );
A2O1A1Ixp33_ASAP7_75t_L g216 ( .A1(n_41), .A2(n_155), .B(n_217), .C(n_221), .Y(n_216) );
A2O1A1Ixp33_ASAP7_75t_L g522 ( .A1(n_42), .A2(n_152), .B(n_155), .C(n_523), .Y(n_522) );
INVx1_ASAP7_75t_L g489 ( .A(n_44), .Y(n_489) );
A2O1A1Ixp33_ASAP7_75t_L g245 ( .A1(n_45), .A2(n_166), .B(n_246), .C(n_247), .Y(n_245) );
NAND2xp5_ASAP7_75t_SL g556 ( .A(n_46), .B(n_164), .Y(n_556) );
CKINVDCx20_ASAP7_75t_R g223 ( .A(n_47), .Y(n_223) );
CKINVDCx20_ASAP7_75t_R g183 ( .A(n_48), .Y(n_183) );
INVx1_ASAP7_75t_L g254 ( .A(n_49), .Y(n_254) );
CKINVDCx16_ASAP7_75t_R g491 ( .A(n_50), .Y(n_491) );
AOI222xp33_ASAP7_75t_SL g452 ( .A1(n_51), .A2(n_453), .B1(n_454), .B2(n_463), .C1(n_749), .C2(n_752), .Y(n_452) );
OAI22xp5_ASAP7_75t_SL g435 ( .A1(n_52), .A2(n_61), .B1(n_436), .B2(n_437), .Y(n_435) );
CKINVDCx20_ASAP7_75t_R g436 ( .A(n_52), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_53), .B(n_181), .Y(n_537) );
AOI22xp5_ASAP7_75t_L g487 ( .A1(n_54), .A2(n_155), .B1(n_258), .B2(n_488), .Y(n_487) );
CKINVDCx20_ASAP7_75t_R g527 ( .A(n_55), .Y(n_527) );
CKINVDCx16_ASAP7_75t_R g509 ( .A(n_56), .Y(n_509) );
CKINVDCx14_ASAP7_75t_R g244 ( .A(n_57), .Y(n_244) );
A2O1A1Ixp33_ASAP7_75t_L g498 ( .A1(n_58), .A2(n_208), .B(n_246), .C(n_499), .Y(n_498) );
AOI22xp5_ASAP7_75t_L g125 ( .A1(n_59), .A2(n_126), .B1(n_127), .B2(n_440), .Y(n_125) );
CKINVDCx20_ASAP7_75t_R g440 ( .A(n_59), .Y(n_440) );
INVx1_ASAP7_75t_L g497 ( .A(n_60), .Y(n_497) );
CKINVDCx20_ASAP7_75t_R g437 ( .A(n_61), .Y(n_437) );
INVx1_ASAP7_75t_L g153 ( .A(n_62), .Y(n_153) );
INVx1_ASAP7_75t_L g143 ( .A(n_63), .Y(n_143) );
INVx1_ASAP7_75t_SL g207 ( .A(n_64), .Y(n_207) );
CKINVDCx20_ASAP7_75t_R g123 ( .A(n_65), .Y(n_123) );
OAI22xp5_ASAP7_75t_SL g434 ( .A1(n_66), .A2(n_435), .B1(n_438), .B2(n_439), .Y(n_434) );
CKINVDCx20_ASAP7_75t_R g438 ( .A(n_66), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_67), .B(n_211), .Y(n_260) );
INVx1_ASAP7_75t_L g159 ( .A(n_68), .Y(n_159) );
A2O1A1Ixp33_ASAP7_75t_SL g477 ( .A1(n_69), .A2(n_208), .B(n_478), .C(n_479), .Y(n_477) );
INVxp67_ASAP7_75t_L g480 ( .A(n_70), .Y(n_480) );
INVx1_ASAP7_75t_L g117 ( .A(n_71), .Y(n_117) );
AOI21xp5_ASAP7_75t_L g242 ( .A1(n_72), .A2(n_181), .B(n_243), .Y(n_242) );
CKINVDCx20_ASAP7_75t_R g171 ( .A(n_73), .Y(n_171) );
AOI21xp5_ASAP7_75t_L g266 ( .A1(n_74), .A2(n_181), .B(n_267), .Y(n_266) );
CKINVDCx20_ASAP7_75t_R g493 ( .A(n_75), .Y(n_493) );
INVx1_ASAP7_75t_L g553 ( .A(n_76), .Y(n_553) );
AOI21xp5_ASAP7_75t_L g179 ( .A1(n_77), .A2(n_180), .B(n_182), .Y(n_179) );
CKINVDCx16_ASAP7_75t_R g215 ( .A(n_78), .Y(n_215) );
INVx1_ASAP7_75t_L g268 ( .A(n_79), .Y(n_268) );
CKINVDCx20_ASAP7_75t_R g461 ( .A(n_80), .Y(n_461) );
A2O1A1Ixp33_ASAP7_75t_L g554 ( .A1(n_81), .A2(n_152), .B(n_155), .C(n_555), .Y(n_554) );
AOI21xp5_ASAP7_75t_L g252 ( .A1(n_82), .A2(n_181), .B(n_253), .Y(n_252) );
INVx1_ASAP7_75t_L g271 ( .A(n_83), .Y(n_271) );
NAND2xp5_ASAP7_75t_SL g524 ( .A(n_84), .B(n_188), .Y(n_524) );
INVx2_ASAP7_75t_L g141 ( .A(n_85), .Y(n_141) );
INVx1_ASAP7_75t_L g236 ( .A(n_86), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_87), .B(n_478), .Y(n_525) );
A2O1A1Ixp33_ASAP7_75t_L g510 ( .A1(n_88), .A2(n_152), .B(n_155), .C(n_511), .Y(n_510) );
INVx2_ASAP7_75t_L g114 ( .A(n_89), .Y(n_114) );
OR2x2_ASAP7_75t_L g444 ( .A(n_89), .B(n_445), .Y(n_444) );
OR2x2_ASAP7_75t_L g464 ( .A(n_89), .B(n_446), .Y(n_464) );
A2O1A1Ixp33_ASAP7_75t_L g154 ( .A1(n_90), .A2(n_155), .B(n_158), .C(n_168), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_91), .B(n_173), .Y(n_501) );
AOI22xp5_ASAP7_75t_L g104 ( .A1(n_92), .A2(n_105), .B1(n_118), .B2(n_756), .Y(n_104) );
CKINVDCx20_ASAP7_75t_R g516 ( .A(n_93), .Y(n_516) );
A2O1A1Ixp33_ASAP7_75t_L g532 ( .A1(n_94), .A2(n_152), .B(n_155), .C(n_533), .Y(n_532) );
CKINVDCx20_ASAP7_75t_R g539 ( .A(n_95), .Y(n_539) );
INVx1_ASAP7_75t_L g476 ( .A(n_96), .Y(n_476) );
CKINVDCx16_ASAP7_75t_R g544 ( .A(n_97), .Y(n_544) );
NAND2xp5_ASAP7_75t_SL g534 ( .A(n_98), .B(n_188), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_99), .B(n_139), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_100), .B(n_139), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g116 ( .A(n_101), .B(n_117), .Y(n_116) );
INVx2_ASAP7_75t_L g257 ( .A(n_102), .Y(n_257) );
AOI21xp5_ASAP7_75t_L g474 ( .A1(n_103), .A2(n_181), .B(n_475), .Y(n_474) );
INVx1_ASAP7_75t_SL g105 ( .A(n_106), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
INVx1_ASAP7_75t_SL g756 ( .A(n_107), .Y(n_756) );
CKINVDCx9p33_ASAP7_75t_R g107 ( .A(n_108), .Y(n_107) );
NAND2xp5_ASAP7_75t_L g108 ( .A(n_109), .B(n_111), .Y(n_108) );
CKINVDCx20_ASAP7_75t_R g109 ( .A(n_110), .Y(n_109) );
CKINVDCx14_ASAP7_75t_R g111 ( .A(n_112), .Y(n_111) );
NAND3xp33_ASAP7_75t_SL g112 ( .A(n_113), .B(n_114), .C(n_115), .Y(n_112) );
AND2x2_ASAP7_75t_L g446 ( .A(n_113), .B(n_447), .Y(n_446) );
OR2x2_ASAP7_75t_L g748 ( .A(n_114), .B(n_446), .Y(n_748) );
NOR2x2_ASAP7_75t_L g751 ( .A(n_114), .B(n_445), .Y(n_751) );
INVx1_ASAP7_75t_SL g115 ( .A(n_116), .Y(n_115) );
OA21x2_ASAP7_75t_L g118 ( .A1(n_119), .A2(n_124), .B(n_451), .Y(n_118) );
INVx1_ASAP7_75t_SL g119 ( .A(n_120), .Y(n_119) );
INVx1_ASAP7_75t_SL g120 ( .A(n_121), .Y(n_120) );
BUFx2_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
INVx2_ASAP7_75t_SL g755 ( .A(n_122), .Y(n_755) );
INVx2_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
OAI21xp5_ASAP7_75t_SL g124 ( .A1(n_125), .A2(n_441), .B(n_448), .Y(n_124) );
INVxp67_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
XOR2xp5_ASAP7_75t_L g127 ( .A(n_128), .B(n_434), .Y(n_127) );
OAI22xp5_ASAP7_75t_SL g463 ( .A1(n_128), .A2(n_464), .B1(n_465), .B2(n_746), .Y(n_463) );
INVx2_ASAP7_75t_L g753 ( .A(n_128), .Y(n_753) );
OR2x2_ASAP7_75t_L g128 ( .A(n_129), .B(n_368), .Y(n_128) );
NAND5xp2_ASAP7_75t_L g129 ( .A(n_130), .B(n_297), .C(n_327), .D(n_348), .E(n_354), .Y(n_129) );
AOI221xp5_ASAP7_75t_SL g130 ( .A1(n_131), .A2(n_227), .B1(n_261), .B2(n_263), .C(n_274), .Y(n_130) );
INVxp67_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
NOR2xp33_ASAP7_75t_L g132 ( .A(n_133), .B(n_224), .Y(n_132) );
NOR2xp33_ASAP7_75t_L g133 ( .A(n_134), .B(n_196), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
A2O1A1Ixp33_ASAP7_75t_SL g348 ( .A1(n_135), .A2(n_212), .B(n_349), .C(n_352), .Y(n_348) );
AND2x2_ASAP7_75t_L g418 ( .A(n_135), .B(n_213), .Y(n_418) );
AND2x2_ASAP7_75t_L g135 ( .A(n_136), .B(n_174), .Y(n_135) );
AND2x2_ASAP7_75t_L g276 ( .A(n_136), .B(n_277), .Y(n_276) );
OR2x2_ASAP7_75t_L g280 ( .A(n_136), .B(n_277), .Y(n_280) );
OR2x2_ASAP7_75t_L g306 ( .A(n_136), .B(n_213), .Y(n_306) );
AND2x2_ASAP7_75t_L g308 ( .A(n_136), .B(n_199), .Y(n_308) );
AND2x2_ASAP7_75t_L g326 ( .A(n_136), .B(n_198), .Y(n_326) );
INVx1_ASAP7_75t_L g359 ( .A(n_136), .Y(n_359) );
INVx2_ASAP7_75t_SL g136 ( .A(n_137), .Y(n_136) );
BUFx2_ASAP7_75t_L g226 ( .A(n_137), .Y(n_226) );
AND2x2_ASAP7_75t_L g262 ( .A(n_137), .B(n_199), .Y(n_262) );
AND2x2_ASAP7_75t_L g415 ( .A(n_137), .B(n_213), .Y(n_415) );
AO21x2_ASAP7_75t_L g137 ( .A1(n_138), .A2(n_145), .B(n_170), .Y(n_137) );
INVx3_ASAP7_75t_L g211 ( .A(n_138), .Y(n_211) );
NOR2xp33_ASAP7_75t_L g222 ( .A(n_138), .B(n_223), .Y(n_222) );
NOR2xp33_ASAP7_75t_L g238 ( .A(n_138), .B(n_239), .Y(n_238) );
NOR2xp33_ASAP7_75t_SL g526 ( .A(n_138), .B(n_527), .Y(n_526) );
INVx4_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
HB1xp67_ASAP7_75t_L g200 ( .A(n_139), .Y(n_200) );
OA21x2_ASAP7_75t_L g473 ( .A1(n_139), .A2(n_474), .B(n_481), .Y(n_473) );
BUFx6f_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
INVx1_ASAP7_75t_L g177 ( .A(n_140), .Y(n_177) );
AND2x2_ASAP7_75t_L g140 ( .A(n_141), .B(n_142), .Y(n_140) );
AND2x2_ASAP7_75t_SL g173 ( .A(n_141), .B(n_142), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_143), .B(n_144), .Y(n_142) );
OAI21xp5_ASAP7_75t_L g145 ( .A1(n_146), .A2(n_147), .B(n_154), .Y(n_145) );
O2A1O1Ixp33_ASAP7_75t_L g214 ( .A1(n_147), .A2(n_173), .B(n_215), .C(n_216), .Y(n_214) );
OAI21xp5_ASAP7_75t_L g232 ( .A1(n_147), .A2(n_233), .B(n_234), .Y(n_232) );
OAI22xp33_ASAP7_75t_L g486 ( .A1(n_147), .A2(n_169), .B1(n_487), .B2(n_491), .Y(n_486) );
OAI21xp5_ASAP7_75t_L g508 ( .A1(n_147), .A2(n_509), .B(n_510), .Y(n_508) );
OAI21xp5_ASAP7_75t_L g552 ( .A1(n_147), .A2(n_553), .B(n_554), .Y(n_552) );
NAND2x1p5_ASAP7_75t_L g147 ( .A(n_148), .B(n_152), .Y(n_147) );
AND2x4_ASAP7_75t_L g181 ( .A(n_148), .B(n_152), .Y(n_181) );
AND2x2_ASAP7_75t_L g148 ( .A(n_149), .B(n_151), .Y(n_148) );
INVx1_ASAP7_75t_L g192 ( .A(n_149), .Y(n_192) );
INVx1_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx2_ASAP7_75t_L g156 ( .A(n_150), .Y(n_156) );
INVx1_ASAP7_75t_L g259 ( .A(n_150), .Y(n_259) );
INVx1_ASAP7_75t_L g157 ( .A(n_151), .Y(n_157) );
BUFx6f_ASAP7_75t_L g162 ( .A(n_151), .Y(n_162) );
BUFx6f_ASAP7_75t_L g164 ( .A(n_151), .Y(n_164) );
INVx3_ASAP7_75t_L g189 ( .A(n_151), .Y(n_189) );
INVx1_ASAP7_75t_L g478 ( .A(n_151), .Y(n_478) );
INVx4_ASAP7_75t_SL g169 ( .A(n_152), .Y(n_169) );
BUFx3_ASAP7_75t_L g221 ( .A(n_152), .Y(n_221) );
INVx5_ASAP7_75t_L g184 ( .A(n_155), .Y(n_184) );
AND2x6_ASAP7_75t_L g155 ( .A(n_156), .B(n_157), .Y(n_155) );
BUFx3_ASAP7_75t_L g167 ( .A(n_156), .Y(n_167) );
BUFx6f_ASAP7_75t_L g209 ( .A(n_156), .Y(n_209) );
O2A1O1Ixp33_ASAP7_75t_L g158 ( .A1(n_159), .A2(n_160), .B(n_163), .C(n_165), .Y(n_158) );
O2A1O1Ixp5_ASAP7_75t_L g235 ( .A1(n_160), .A2(n_165), .B(n_236), .C(n_237), .Y(n_235) );
INVx2_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
OAI22xp5_ASAP7_75t_SL g488 ( .A1(n_161), .A2(n_162), .B1(n_489), .B2(n_490), .Y(n_488) );
INVx2_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
INVx4_ASAP7_75t_L g191 ( .A(n_162), .Y(n_191) );
INVx4_ASAP7_75t_L g205 ( .A(n_164), .Y(n_205) );
INVx2_ASAP7_75t_L g246 ( .A(n_164), .Y(n_246) );
AOI21xp5_ASAP7_75t_L g523 ( .A1(n_165), .A2(n_524), .B(n_525), .Y(n_523) );
AOI21xp5_ASAP7_75t_L g555 ( .A1(n_165), .A2(n_556), .B(n_557), .Y(n_555) );
INVx2_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
INVx2_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
INVx1_ASAP7_75t_L g272 ( .A(n_167), .Y(n_272) );
INVx1_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
O2A1O1Ixp33_ASAP7_75t_SL g182 ( .A1(n_169), .A2(n_183), .B(n_184), .C(n_185), .Y(n_182) );
O2A1O1Ixp33_ASAP7_75t_L g202 ( .A1(n_169), .A2(n_184), .B(n_203), .C(n_204), .Y(n_202) );
O2A1O1Ixp33_ASAP7_75t_SL g243 ( .A1(n_169), .A2(n_184), .B(n_244), .C(n_245), .Y(n_243) );
O2A1O1Ixp33_ASAP7_75t_SL g253 ( .A1(n_169), .A2(n_184), .B(n_254), .C(n_255), .Y(n_253) );
O2A1O1Ixp33_ASAP7_75t_SL g267 ( .A1(n_169), .A2(n_184), .B(n_268), .C(n_269), .Y(n_267) );
O2A1O1Ixp33_ASAP7_75t_L g475 ( .A1(n_169), .A2(n_184), .B(n_476), .C(n_477), .Y(n_475) );
O2A1O1Ixp33_ASAP7_75t_L g496 ( .A1(n_169), .A2(n_184), .B(n_497), .C(n_498), .Y(n_496) );
O2A1O1Ixp33_ASAP7_75t_L g543 ( .A1(n_169), .A2(n_184), .B(n_544), .C(n_545), .Y(n_543) );
NOR2xp33_ASAP7_75t_L g170 ( .A(n_171), .B(n_172), .Y(n_170) );
INVx1_ASAP7_75t_L g195 ( .A(n_172), .Y(n_195) );
AO21x2_ASAP7_75t_L g530 ( .A1(n_172), .A2(n_531), .B(n_538), .Y(n_530) );
INVx2_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
INVx1_ASAP7_75t_L g231 ( .A(n_173), .Y(n_231) );
OA21x2_ASAP7_75t_L g241 ( .A1(n_173), .A2(n_242), .B(n_249), .Y(n_241) );
OA21x2_ASAP7_75t_L g541 ( .A1(n_173), .A2(n_542), .B(n_548), .Y(n_541) );
AND2x2_ASAP7_75t_L g296 ( .A(n_174), .B(n_197), .Y(n_296) );
OR2x2_ASAP7_75t_L g300 ( .A(n_174), .B(n_213), .Y(n_300) );
AND2x2_ASAP7_75t_L g325 ( .A(n_174), .B(n_326), .Y(n_325) );
INVx1_ASAP7_75t_SL g372 ( .A(n_174), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_174), .B(n_334), .Y(n_420) );
AO21x2_ASAP7_75t_L g174 ( .A1(n_175), .A2(n_178), .B(n_193), .Y(n_174) );
INVx1_ASAP7_75t_L g278 ( .A(n_175), .Y(n_278) );
AO21x2_ASAP7_75t_L g551 ( .A1(n_175), .A2(n_552), .B(n_558), .Y(n_551) );
INVx1_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
AOI21xp5_ASAP7_75t_SL g520 ( .A1(n_176), .A2(n_521), .B(n_522), .Y(n_520) );
INVx2_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
AO21x2_ASAP7_75t_L g485 ( .A1(n_177), .A2(n_486), .B(n_492), .Y(n_485) );
NOR2xp33_ASAP7_75t_L g492 ( .A(n_177), .B(n_493), .Y(n_492) );
AO21x2_ASAP7_75t_L g507 ( .A1(n_177), .A2(n_508), .B(n_515), .Y(n_507) );
INVx1_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
OA21x2_ASAP7_75t_L g277 ( .A1(n_179), .A2(n_194), .B(n_278), .Y(n_277) );
BUFx2_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
NAND2xp5_ASAP7_75t_SL g185 ( .A(n_186), .B(n_192), .Y(n_185) );
OAI22xp33_ASAP7_75t_L g186 ( .A1(n_187), .A2(n_188), .B1(n_190), .B2(n_191), .Y(n_186) );
O2A1O1Ixp33_ASAP7_75t_L g217 ( .A1(n_188), .A2(n_218), .B(n_219), .C(n_220), .Y(n_217) );
O2A1O1Ixp33_ASAP7_75t_L g511 ( .A1(n_188), .A2(n_512), .B(n_513), .C(n_514), .Y(n_511) );
INVx5_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
NOR2xp33_ASAP7_75t_L g247 ( .A(n_189), .B(n_248), .Y(n_247) );
NOR2xp33_ASAP7_75t_L g479 ( .A(n_189), .B(n_480), .Y(n_479) );
NOR2xp33_ASAP7_75t_L g499 ( .A(n_189), .B(n_500), .Y(n_499) );
NOR2xp33_ASAP7_75t_L g256 ( .A(n_191), .B(n_257), .Y(n_256) );
NOR2xp33_ASAP7_75t_L g270 ( .A(n_191), .B(n_271), .Y(n_270) );
NOR2xp33_ASAP7_75t_L g546 ( .A(n_191), .B(n_547), .Y(n_546) );
INVx2_ASAP7_75t_L g220 ( .A(n_192), .Y(n_220) );
INVx1_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
OAI322xp33_ASAP7_75t_L g421 ( .A1(n_196), .A2(n_357), .A3(n_380), .B1(n_401), .B2(n_422), .C1(n_424), .C2(n_425), .Y(n_421) );
INVx1_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_197), .B(n_277), .Y(n_424) );
AND2x2_ASAP7_75t_L g197 ( .A(n_198), .B(n_212), .Y(n_197) );
AND2x2_ASAP7_75t_L g225 ( .A(n_198), .B(n_226), .Y(n_225) );
AND2x4_ASAP7_75t_L g293 ( .A(n_198), .B(n_213), .Y(n_293) );
INVx2_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
AND2x2_ASAP7_75t_L g334 ( .A(n_199), .B(n_213), .Y(n_334) );
AND2x2_ASAP7_75t_L g378 ( .A(n_199), .B(n_212), .Y(n_378) );
OA21x2_ASAP7_75t_L g199 ( .A1(n_200), .A2(n_201), .B(n_210), .Y(n_199) );
OA21x2_ASAP7_75t_L g251 ( .A1(n_200), .A2(n_252), .B(n_260), .Y(n_251) );
OA21x2_ASAP7_75t_L g265 ( .A1(n_200), .A2(n_266), .B(n_273), .Y(n_265) );
NOR2xp33_ASAP7_75t_L g206 ( .A(n_205), .B(n_207), .Y(n_206) );
INVx3_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
HB1xp67_ASAP7_75t_L g536 ( .A(n_209), .Y(n_536) );
OA21x2_ASAP7_75t_L g494 ( .A1(n_211), .A2(n_495), .B(n_501), .Y(n_494) );
AND2x2_ASAP7_75t_L g261 ( .A(n_212), .B(n_262), .Y(n_261) );
OR2x2_ASAP7_75t_L g279 ( .A(n_212), .B(n_280), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_212), .B(n_308), .Y(n_432) );
INVx3_ASAP7_75t_SL g212 ( .A(n_213), .Y(n_212) );
AND2x2_ASAP7_75t_L g224 ( .A(n_213), .B(n_225), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_213), .B(n_276), .Y(n_275) );
AND2x2_ASAP7_75t_L g346 ( .A(n_213), .B(n_277), .Y(n_346) );
AND2x2_ASAP7_75t_L g373 ( .A(n_213), .B(n_308), .Y(n_373) );
OR2x2_ASAP7_75t_L g429 ( .A(n_213), .B(n_280), .Y(n_429) );
OR2x6_ASAP7_75t_L g213 ( .A(n_214), .B(n_222), .Y(n_213) );
INVx1_ASAP7_75t_SL g315 ( .A(n_224), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_225), .B(n_346), .Y(n_347) );
AND2x2_ASAP7_75t_L g381 ( .A(n_225), .B(n_371), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_225), .B(n_304), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_225), .B(n_426), .Y(n_425) );
OAI31xp33_ASAP7_75t_L g399 ( .A1(n_227), .A2(n_261), .A3(n_400), .B(n_402), .Y(n_399) );
AND2x2_ASAP7_75t_L g227 ( .A(n_228), .B(n_240), .Y(n_227) );
NAND2xp5_ASAP7_75t_SL g366 ( .A(n_228), .B(n_367), .Y(n_366) );
AND2x2_ASAP7_75t_L g382 ( .A(n_228), .B(n_317), .Y(n_382) );
OR2x2_ASAP7_75t_L g389 ( .A(n_228), .B(n_390), .Y(n_389) );
OR2x2_ASAP7_75t_L g401 ( .A(n_228), .B(n_290), .Y(n_401) );
CKINVDCx16_ASAP7_75t_R g228 ( .A(n_229), .Y(n_228) );
OR2x2_ASAP7_75t_L g335 ( .A(n_229), .B(n_336), .Y(n_335) );
BUFx3_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
AND2x2_ASAP7_75t_L g263 ( .A(n_230), .B(n_264), .Y(n_263) );
INVx4_ASAP7_75t_L g284 ( .A(n_230), .Y(n_284) );
AND2x2_ASAP7_75t_L g321 ( .A(n_230), .B(n_265), .Y(n_321) );
AO21x2_ASAP7_75t_L g230 ( .A1(n_231), .A2(n_232), .B(n_238), .Y(n_230) );
NOR2xp33_ASAP7_75t_L g515 ( .A(n_231), .B(n_516), .Y(n_515) );
NOR2xp33_ASAP7_75t_L g538 ( .A(n_231), .B(n_539), .Y(n_538) );
NOR2xp33_ASAP7_75t_L g558 ( .A(n_231), .B(n_440), .Y(n_558) );
AND2x2_ASAP7_75t_L g320 ( .A(n_240), .B(n_321), .Y(n_320) );
INVx1_ASAP7_75t_SL g390 ( .A(n_240), .Y(n_390) );
AND2x2_ASAP7_75t_L g240 ( .A(n_241), .B(n_250), .Y(n_240) );
NOR2xp33_ASAP7_75t_L g283 ( .A(n_241), .B(n_284), .Y(n_283) );
OR2x2_ASAP7_75t_L g290 ( .A(n_241), .B(n_251), .Y(n_290) );
INVx2_ASAP7_75t_L g310 ( .A(n_241), .Y(n_310) );
AND2x2_ASAP7_75t_L g324 ( .A(n_241), .B(n_251), .Y(n_324) );
AND2x2_ASAP7_75t_L g331 ( .A(n_241), .B(n_287), .Y(n_331) );
BUFx3_ASAP7_75t_L g341 ( .A(n_241), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_241), .B(n_344), .Y(n_343) );
INVx2_ASAP7_75t_L g286 ( .A(n_250), .Y(n_286) );
AND2x2_ASAP7_75t_L g294 ( .A(n_250), .B(n_284), .Y(n_294) );
INVx2_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
AND2x2_ASAP7_75t_L g264 ( .A(n_251), .B(n_265), .Y(n_264) );
HB1xp67_ASAP7_75t_L g318 ( .A(n_251), .Y(n_318) );
INVx2_ASAP7_75t_L g514 ( .A(n_258), .Y(n_514) );
INVx3_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
INVx2_ASAP7_75t_SL g301 ( .A(n_262), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_262), .B(n_346), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_262), .B(n_371), .Y(n_392) );
NAND2xp5_ASAP7_75t_SL g394 ( .A(n_263), .B(n_341), .Y(n_394) );
INVx1_ASAP7_75t_SL g428 ( .A(n_263), .Y(n_428) );
INVx1_ASAP7_75t_SL g336 ( .A(n_264), .Y(n_336) );
INVx1_ASAP7_75t_SL g287 ( .A(n_265), .Y(n_287) );
HB1xp67_ASAP7_75t_L g298 ( .A(n_265), .Y(n_298) );
OR2x2_ASAP7_75t_L g309 ( .A(n_265), .B(n_284), .Y(n_309) );
AND2x2_ASAP7_75t_L g323 ( .A(n_265), .B(n_284), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_265), .B(n_313), .Y(n_375) );
A2O1A1Ixp33_ASAP7_75t_L g274 ( .A1(n_275), .A2(n_279), .B(n_281), .C(n_292), .Y(n_274) );
AOI31xp33_ASAP7_75t_L g391 ( .A1(n_275), .A2(n_392), .A3(n_393), .B(n_394), .Y(n_391) );
AND2x2_ASAP7_75t_L g364 ( .A(n_276), .B(n_293), .Y(n_364) );
BUFx3_ASAP7_75t_L g304 ( .A(n_277), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_277), .B(n_308), .Y(n_307) );
OR2x2_ASAP7_75t_L g340 ( .A(n_277), .B(n_341), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_277), .B(n_359), .Y(n_358) );
INVx1_ASAP7_75t_SL g295 ( .A(n_280), .Y(n_295) );
OAI222xp33_ASAP7_75t_L g404 ( .A1(n_280), .A2(n_405), .B1(n_408), .B2(n_409), .C1(n_410), .C2(n_411), .Y(n_404) );
NOR2xp33_ASAP7_75t_L g281 ( .A(n_282), .B(n_288), .Y(n_281) );
INVx1_ASAP7_75t_L g410 ( .A(n_282), .Y(n_410) );
AND2x2_ASAP7_75t_L g282 ( .A(n_283), .B(n_285), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_284), .B(n_287), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_284), .B(n_310), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_284), .B(n_285), .Y(n_380) );
INVx1_ASAP7_75t_L g431 ( .A(n_284), .Y(n_431) );
NAND2xp5_ASAP7_75t_SL g361 ( .A(n_285), .B(n_362), .Y(n_361) );
INVx1_ASAP7_75t_L g433 ( .A(n_285), .Y(n_433) );
AND2x2_ASAP7_75t_L g285 ( .A(n_286), .B(n_287), .Y(n_285) );
INVx2_ASAP7_75t_L g313 ( .A(n_286), .Y(n_313) );
HB1xp67_ASAP7_75t_L g356 ( .A(n_287), .Y(n_356) );
AOI32xp33_ASAP7_75t_L g292 ( .A1(n_288), .A2(n_293), .A3(n_294), .B1(n_295), .B2(n_296), .Y(n_292) );
INVx2_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
OR2x2_ASAP7_75t_L g289 ( .A(n_290), .B(n_291), .Y(n_289) );
NOR2xp33_ASAP7_75t_L g355 ( .A(n_290), .B(n_356), .Y(n_355) );
INVx1_ASAP7_75t_L g367 ( .A(n_290), .Y(n_367) );
OR2x2_ASAP7_75t_L g408 ( .A(n_290), .B(n_309), .Y(n_408) );
INVx1_ASAP7_75t_L g344 ( .A(n_291), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_293), .B(n_304), .Y(n_329) );
INVx3_ASAP7_75t_L g338 ( .A(n_293), .Y(n_338) );
AOI322xp5_ASAP7_75t_L g354 ( .A1(n_293), .A2(n_338), .A3(n_355), .B1(n_357), .B2(n_360), .C1(n_364), .C2(n_365), .Y(n_354) );
AND2x2_ASAP7_75t_L g330 ( .A(n_294), .B(n_331), .Y(n_330) );
INVxp67_ASAP7_75t_L g407 ( .A(n_294), .Y(n_407) );
A2O1A1O1Ixp25_ASAP7_75t_L g297 ( .A1(n_298), .A2(n_299), .B(n_302), .C(n_310), .D(n_311), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_298), .B(n_341), .Y(n_406) );
NOR2xp33_ASAP7_75t_L g299 ( .A(n_300), .B(n_301), .Y(n_299) );
OAI221xp5_ASAP7_75t_L g311 ( .A1(n_300), .A2(n_312), .B1(n_315), .B2(n_316), .C(n_319), .Y(n_311) );
INVx1_ASAP7_75t_SL g426 ( .A(n_300), .Y(n_426) );
AOI21xp33_ASAP7_75t_L g302 ( .A1(n_303), .A2(n_307), .B(n_309), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_304), .B(n_305), .Y(n_303) );
NAND2xp5_ASAP7_75t_SL g414 ( .A(n_304), .B(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
OAI221xp5_ASAP7_75t_SL g396 ( .A1(n_306), .A2(n_390), .B1(n_397), .B2(n_398), .C(n_399), .Y(n_396) );
OAI222xp33_ASAP7_75t_L g427 ( .A1(n_307), .A2(n_428), .B1(n_429), .B2(n_430), .C1(n_432), .C2(n_433), .Y(n_427) );
AND2x2_ASAP7_75t_L g385 ( .A(n_308), .B(n_371), .Y(n_385) );
AOI21xp5_ASAP7_75t_L g397 ( .A1(n_308), .A2(n_323), .B(n_370), .Y(n_397) );
INVx1_ASAP7_75t_L g411 ( .A(n_308), .Y(n_411) );
INVx2_ASAP7_75t_SL g314 ( .A(n_309), .Y(n_314) );
AND2x2_ASAP7_75t_L g317 ( .A(n_310), .B(n_318), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_313), .B(n_314), .Y(n_312) );
INVx1_ASAP7_75t_SL g351 ( .A(n_313), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_313), .B(n_323), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_314), .B(n_351), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_314), .B(n_324), .Y(n_353) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
OAI21xp5_ASAP7_75t_SL g319 ( .A1(n_320), .A2(n_322), .B(n_325), .Y(n_319) );
INVx1_ASAP7_75t_SL g337 ( .A(n_321), .Y(n_337) );
AND2x2_ASAP7_75t_L g384 ( .A(n_321), .B(n_367), .Y(n_384) );
AND2x2_ASAP7_75t_L g322 ( .A(n_323), .B(n_324), .Y(n_322) );
AND2x2_ASAP7_75t_L g423 ( .A(n_323), .B(n_341), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_324), .B(n_431), .Y(n_430) );
INVx1_ASAP7_75t_SL g409 ( .A(n_325), .Y(n_409) );
AOI221xp5_ASAP7_75t_L g327 ( .A1(n_328), .A2(n_330), .B1(n_332), .B2(n_339), .C(n_342), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
OAI22xp5_ASAP7_75t_L g332 ( .A1(n_333), .A2(n_335), .B1(n_337), .B2(n_338), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
OAI22xp33_ASAP7_75t_L g342 ( .A1(n_336), .A2(n_343), .B1(n_345), .B2(n_347), .Y(n_342) );
OR2x2_ASAP7_75t_L g413 ( .A(n_337), .B(n_341), .Y(n_413) );
OR2x2_ASAP7_75t_L g416 ( .A(n_337), .B(n_351), .Y(n_416) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
OAI221xp5_ASAP7_75t_L g412 ( .A1(n_358), .A2(n_413), .B1(n_414), .B2(n_416), .C(n_417), .Y(n_412) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVxp67_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
NAND3xp33_ASAP7_75t_SL g368 ( .A(n_369), .B(n_383), .C(n_395), .Y(n_368) );
AOI222xp33_ASAP7_75t_L g369 ( .A1(n_370), .A2(n_374), .B1(n_376), .B2(n_379), .C1(n_381), .C2(n_382), .Y(n_369) );
AND2x2_ASAP7_75t_L g370 ( .A(n_371), .B(n_373), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_371), .B(n_378), .Y(n_377) );
INVx2_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
INVx1_ASAP7_75t_L g393 ( .A(n_373), .Y(n_393) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVxp67_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
AOI221xp5_ASAP7_75t_L g383 ( .A1(n_384), .A2(n_385), .B1(n_386), .B2(n_388), .C(n_391), .Y(n_383) );
INVx1_ASAP7_75t_L g398 ( .A(n_384), .Y(n_398) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
OAI21xp33_ASAP7_75t_L g417 ( .A1(n_388), .A2(n_418), .B(n_419), .Y(n_417) );
INVx1_ASAP7_75t_SL g388 ( .A(n_389), .Y(n_388) );
NOR5xp2_ASAP7_75t_L g395 ( .A(n_396), .B(n_404), .C(n_412), .D(n_421), .E(n_427), .Y(n_395) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
OR2x2_ASAP7_75t_L g405 ( .A(n_406), .B(n_407), .Y(n_405) );
INVxp67_ASAP7_75t_SL g419 ( .A(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
CKINVDCx20_ASAP7_75t_R g439 ( .A(n_435), .Y(n_439) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx1_ASAP7_75t_SL g442 ( .A(n_443), .Y(n_442) );
INVx1_ASAP7_75t_SL g443 ( .A(n_444), .Y(n_443) );
BUFx2_ASAP7_75t_L g450 ( .A(n_444), .Y(n_450) );
INVx2_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
NAND3xp33_ASAP7_75t_L g451 ( .A(n_448), .B(n_452), .C(n_754), .Y(n_451) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
OAI22xp5_ASAP7_75t_SL g752 ( .A1(n_464), .A2(n_466), .B1(n_746), .B2(n_753), .Y(n_752) );
INVx1_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
AND2x2_ASAP7_75t_SL g466 ( .A(n_467), .B(n_683), .Y(n_466) );
NOR4xp25_ASAP7_75t_L g467 ( .A(n_468), .B(n_613), .C(n_644), .D(n_663), .Y(n_467) );
NAND4xp25_ASAP7_75t_L g468 ( .A(n_469), .B(n_571), .C(n_586), .D(n_604), .Y(n_468) );
AOI222xp33_ASAP7_75t_L g469 ( .A1(n_470), .A2(n_517), .B1(n_549), .B2(n_559), .C1(n_564), .C2(n_566), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_471), .B(n_502), .Y(n_470) );
INVx1_ASAP7_75t_L g627 ( .A(n_471), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_472), .B(n_482), .Y(n_471) );
AND2x2_ASAP7_75t_L g503 ( .A(n_472), .B(n_494), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_472), .B(n_506), .Y(n_656) );
INVx3_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
OR2x2_ASAP7_75t_L g563 ( .A(n_473), .B(n_484), .Y(n_563) );
AND2x2_ASAP7_75t_L g572 ( .A(n_473), .B(n_573), .Y(n_572) );
INVx1_ASAP7_75t_L g598 ( .A(n_473), .Y(n_598) );
AND2x2_ASAP7_75t_L g619 ( .A(n_473), .B(n_484), .Y(n_619) );
BUFx2_ASAP7_75t_L g642 ( .A(n_473), .Y(n_642) );
AND2x2_ASAP7_75t_L g666 ( .A(n_473), .B(n_485), .Y(n_666) );
AND2x2_ASAP7_75t_L g730 ( .A(n_473), .B(n_494), .Y(n_730) );
AND2x2_ASAP7_75t_L g631 ( .A(n_482), .B(n_562), .Y(n_631) );
INVx1_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
NOR2xp33_ASAP7_75t_L g655 ( .A(n_483), .B(n_656), .Y(n_655) );
OR2x2_ASAP7_75t_L g483 ( .A(n_484), .B(n_494), .Y(n_483) );
OR2x2_ASAP7_75t_L g591 ( .A(n_484), .B(n_507), .Y(n_591) );
AND2x2_ASAP7_75t_L g603 ( .A(n_484), .B(n_562), .Y(n_603) );
BUFx2_ASAP7_75t_L g735 ( .A(n_484), .Y(n_735) );
INVx3_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
OR2x2_ASAP7_75t_L g505 ( .A(n_485), .B(n_506), .Y(n_505) );
AND2x2_ASAP7_75t_L g585 ( .A(n_485), .B(n_507), .Y(n_585) );
AND2x2_ASAP7_75t_L g638 ( .A(n_485), .B(n_494), .Y(n_638) );
HB1xp67_ASAP7_75t_L g674 ( .A(n_485), .Y(n_674) );
AND2x2_ASAP7_75t_L g561 ( .A(n_494), .B(n_562), .Y(n_561) );
INVx1_ASAP7_75t_SL g573 ( .A(n_494), .Y(n_573) );
INVx2_ASAP7_75t_L g584 ( .A(n_494), .Y(n_584) );
BUFx2_ASAP7_75t_L g608 ( .A(n_494), .Y(n_608) );
AND2x2_ASAP7_75t_SL g665 ( .A(n_494), .B(n_666), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_503), .B(n_504), .Y(n_502) );
AOI332xp33_ASAP7_75t_L g586 ( .A1(n_503), .A2(n_587), .A3(n_591), .B1(n_592), .B2(n_596), .B3(n_599), .C1(n_600), .C2(n_602), .Y(n_586) );
NAND2x1_ASAP7_75t_L g671 ( .A(n_503), .B(n_562), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_503), .B(n_576), .Y(n_722) );
A2O1A1Ixp33_ASAP7_75t_SL g604 ( .A1(n_504), .A2(n_605), .B(n_608), .C(n_609), .Y(n_604) );
AND2x2_ASAP7_75t_L g743 ( .A(n_504), .B(n_584), .Y(n_743) );
INVx3_ASAP7_75t_SL g504 ( .A(n_505), .Y(n_504) );
OR2x2_ASAP7_75t_L g640 ( .A(n_505), .B(n_641), .Y(n_640) );
OR2x2_ASAP7_75t_L g645 ( .A(n_505), .B(n_642), .Y(n_645) );
INVx1_ASAP7_75t_L g576 ( .A(n_506), .Y(n_576) );
AND2x2_ASAP7_75t_L g679 ( .A(n_506), .B(n_638), .Y(n_679) );
AND2x2_ASAP7_75t_L g680 ( .A(n_506), .B(n_619), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_506), .B(n_690), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_506), .B(n_597), .Y(n_705) );
INVx3_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
INVx3_ASAP7_75t_L g562 ( .A(n_507), .Y(n_562) );
OAI31xp33_ASAP7_75t_L g744 ( .A1(n_517), .A2(n_665), .A3(n_672), .B(n_745), .Y(n_744) );
AND2x2_ASAP7_75t_L g517 ( .A(n_518), .B(n_528), .Y(n_517) );
AND2x2_ASAP7_75t_L g549 ( .A(n_518), .B(n_550), .Y(n_549) );
NAND2x1_ASAP7_75t_SL g567 ( .A(n_518), .B(n_568), .Y(n_567) );
HB1xp67_ASAP7_75t_L g654 ( .A(n_518), .Y(n_654) );
AND2x2_ASAP7_75t_L g659 ( .A(n_518), .B(n_570), .Y(n_659) );
INVx3_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
A2O1A1Ixp33_ASAP7_75t_L g571 ( .A1(n_519), .A2(n_572), .B(n_574), .C(n_577), .Y(n_571) );
OR2x2_ASAP7_75t_L g588 ( .A(n_519), .B(n_589), .Y(n_588) );
INVx1_ASAP7_75t_L g601 ( .A(n_519), .Y(n_601) );
AND2x2_ASAP7_75t_L g607 ( .A(n_519), .B(n_551), .Y(n_607) );
INVx2_ASAP7_75t_L g625 ( .A(n_519), .Y(n_625) );
AND2x2_ASAP7_75t_L g636 ( .A(n_519), .B(n_590), .Y(n_636) );
AND2x2_ASAP7_75t_L g668 ( .A(n_519), .B(n_626), .Y(n_668) );
AND2x2_ASAP7_75t_L g672 ( .A(n_519), .B(n_595), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_519), .B(n_528), .Y(n_677) );
AND2x2_ASAP7_75t_L g711 ( .A(n_519), .B(n_712), .Y(n_711) );
NOR2xp33_ASAP7_75t_L g745 ( .A(n_519), .B(n_614), .Y(n_745) );
OR2x6_ASAP7_75t_L g519 ( .A(n_520), .B(n_526), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_528), .B(n_576), .Y(n_575) );
INVx1_ASAP7_75t_L g653 ( .A(n_528), .Y(n_653) );
AND2x2_ASAP7_75t_L g715 ( .A(n_528), .B(n_636), .Y(n_715) );
AND2x2_ASAP7_75t_L g528 ( .A(n_529), .B(n_540), .Y(n_528) );
OR2x2_ASAP7_75t_L g569 ( .A(n_529), .B(n_570), .Y(n_569) );
AND2x2_ASAP7_75t_L g579 ( .A(n_529), .B(n_580), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_529), .B(n_590), .Y(n_589) );
INVx1_ASAP7_75t_L g687 ( .A(n_529), .Y(n_687) );
AND2x2_ASAP7_75t_L g704 ( .A(n_529), .B(n_551), .Y(n_704) );
INVx2_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
AND2x2_ASAP7_75t_L g595 ( .A(n_530), .B(n_540), .Y(n_595) );
AND2x2_ASAP7_75t_L g624 ( .A(n_530), .B(n_625), .Y(n_624) );
INVx1_ASAP7_75t_L g635 ( .A(n_530), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_530), .B(n_590), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_532), .B(n_537), .Y(n_531) );
AOI21xp5_ASAP7_75t_L g533 ( .A1(n_534), .A2(n_535), .B(n_536), .Y(n_533) );
INVx1_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
AND2x2_ASAP7_75t_L g550 ( .A(n_541), .B(n_551), .Y(n_550) );
INVx2_ASAP7_75t_L g570 ( .A(n_541), .Y(n_570) );
AND2x2_ASAP7_75t_L g626 ( .A(n_541), .B(n_590), .Y(n_626) );
INVx1_ASAP7_75t_L g728 ( .A(n_549), .Y(n_728) );
INVx1_ASAP7_75t_L g732 ( .A(n_550), .Y(n_732) );
INVx2_ASAP7_75t_L g590 ( .A(n_551), .Y(n_590) );
NOR2xp33_ASAP7_75t_L g559 ( .A(n_560), .B(n_563), .Y(n_559) );
INVx1_ASAP7_75t_SL g560 ( .A(n_561), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_561), .B(n_707), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_561), .B(n_666), .Y(n_724) );
OR2x2_ASAP7_75t_L g565 ( .A(n_562), .B(n_563), .Y(n_565) );
INVx1_ASAP7_75t_SL g617 ( .A(n_562), .Y(n_617) );
INVx1_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
INVx1_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
AOI221xp5_ASAP7_75t_L g620 ( .A1(n_568), .A2(n_621), .B1(n_623), .B2(n_627), .C(n_628), .Y(n_620) );
INVx2_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
OR2x2_ASAP7_75t_L g648 ( .A(n_569), .B(n_612), .Y(n_648) );
INVx2_ASAP7_75t_L g580 ( .A(n_570), .Y(n_580) );
INVx1_ASAP7_75t_L g606 ( .A(n_570), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_570), .B(n_590), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_570), .B(n_593), .Y(n_700) );
INVx1_ASAP7_75t_L g708 ( .A(n_570), .Y(n_708) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_572), .B(n_576), .Y(n_622) );
AND2x4_ASAP7_75t_L g597 ( .A(n_573), .B(n_598), .Y(n_597) );
INVx1_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
AND2x2_ASAP7_75t_L g710 ( .A(n_576), .B(n_666), .Y(n_710) );
NOR2xp33_ASAP7_75t_L g577 ( .A(n_578), .B(n_581), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_579), .B(n_611), .Y(n_610) );
INVxp67_ASAP7_75t_L g718 ( .A(n_580), .Y(n_718) );
INVxp67_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
AND2x2_ASAP7_75t_L g582 ( .A(n_583), .B(n_585), .Y(n_582) );
INVx1_ASAP7_75t_SL g583 ( .A(n_584), .Y(n_583) );
AND2x2_ASAP7_75t_L g618 ( .A(n_584), .B(n_619), .Y(n_618) );
AND2x2_ASAP7_75t_L g690 ( .A(n_584), .B(n_666), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_584), .B(n_603), .Y(n_696) );
AOI322xp5_ASAP7_75t_L g650 ( .A1(n_585), .A2(n_619), .A3(n_626), .B1(n_651), .B2(n_654), .C1(n_655), .C2(n_657), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_585), .B(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
OR2x2_ASAP7_75t_L g716 ( .A(n_588), .B(n_717), .Y(n_716) );
INVx1_ASAP7_75t_L g662 ( .A(n_589), .Y(n_662) );
INVx2_ASAP7_75t_L g593 ( .A(n_590), .Y(n_593) );
INVx1_ASAP7_75t_L g652 ( .A(n_590), .Y(n_652) );
CKINVDCx16_ASAP7_75t_R g599 ( .A(n_591), .Y(n_599) );
NOR2xp33_ASAP7_75t_L g592 ( .A(n_593), .B(n_594), .Y(n_592) );
AND2x2_ASAP7_75t_L g688 ( .A(n_593), .B(n_601), .Y(n_688) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
AND2x2_ASAP7_75t_L g600 ( .A(n_595), .B(n_601), .Y(n_600) );
AND2x2_ASAP7_75t_L g643 ( .A(n_595), .B(n_636), .Y(n_643) );
AND2x2_ASAP7_75t_L g647 ( .A(n_595), .B(n_607), .Y(n_647) );
OAI21xp33_ASAP7_75t_SL g657 ( .A1(n_596), .A2(n_658), .B(n_660), .Y(n_657) );
OAI22xp33_ASAP7_75t_L g727 ( .A1(n_596), .A2(n_728), .B1(n_729), .B2(n_731), .Y(n_727) );
INVx3_ASAP7_75t_SL g596 ( .A(n_597), .Y(n_596) );
AND2x2_ASAP7_75t_L g602 ( .A(n_597), .B(n_603), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_597), .B(n_617), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g736 ( .A(n_599), .B(n_737), .Y(n_736) );
AND2x2_ASAP7_75t_L g605 ( .A(n_606), .B(n_607), .Y(n_605) );
INVx1_ASAP7_75t_L g739 ( .A(n_606), .Y(n_739) );
INVx4_ASAP7_75t_L g612 ( .A(n_607), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_607), .B(n_634), .Y(n_682) );
INVx1_ASAP7_75t_SL g694 ( .A(n_608), .Y(n_694) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
NOR2xp67_ASAP7_75t_L g707 ( .A(n_612), .B(n_708), .Y(n_707) );
OAI211xp5_ASAP7_75t_SL g613 ( .A1(n_614), .A2(n_615), .B(n_620), .C(n_637), .Y(n_613) );
OAI221xp5_ASAP7_75t_SL g733 ( .A1(n_615), .A2(n_653), .B1(n_732), .B2(n_734), .C(n_736), .Y(n_733) );
INVx1_ASAP7_75t_SL g615 ( .A(n_616), .Y(n_615) );
AND2x2_ASAP7_75t_L g616 ( .A(n_617), .B(n_618), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_617), .B(n_730), .Y(n_729) );
OAI31xp33_ASAP7_75t_L g709 ( .A1(n_618), .A2(n_695), .A3(n_710), .B(n_711), .Y(n_709) );
INVx1_ASAP7_75t_L g649 ( .A(n_619), .Y(n_649) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
AND2x2_ASAP7_75t_L g623 ( .A(n_624), .B(n_626), .Y(n_623) );
INVx1_ASAP7_75t_L g699 ( .A(n_624), .Y(n_699) );
AND2x2_ASAP7_75t_L g712 ( .A(n_626), .B(n_635), .Y(n_712) );
AOI21xp33_ASAP7_75t_L g628 ( .A1(n_629), .A2(n_630), .B(n_632), .Y(n_628) );
INVx1_ASAP7_75t_SL g630 ( .A(n_631), .Y(n_630) );
INVxp67_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
AND2x2_ASAP7_75t_L g633 ( .A(n_634), .B(n_636), .Y(n_633) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g738 ( .A(n_636), .B(n_739), .Y(n_738) );
OAI21xp33_ASAP7_75t_L g637 ( .A1(n_638), .A2(n_639), .B(n_643), .Y(n_637) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
INVx1_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
OAI221xp5_ASAP7_75t_SL g644 ( .A1(n_645), .A2(n_646), .B1(n_648), .B2(n_649), .C(n_650), .Y(n_644) );
A2O1A1Ixp33_ASAP7_75t_L g713 ( .A1(n_645), .A2(n_714), .B(n_716), .C(n_719), .Y(n_713) );
CKINVDCx16_ASAP7_75t_R g646 ( .A(n_647), .Y(n_646) );
NAND2xp5_ASAP7_75t_SL g697 ( .A(n_648), .B(n_698), .Y(n_697) );
NOR2xp33_ASAP7_75t_L g651 ( .A(n_652), .B(n_653), .Y(n_651) );
INVx1_ASAP7_75t_L g675 ( .A(n_656), .Y(n_675) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
AND2x2_ASAP7_75t_L g661 ( .A(n_659), .B(n_662), .Y(n_661) );
AND2x2_ASAP7_75t_L g703 ( .A(n_659), .B(n_704), .Y(n_703) );
INVx2_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
OAI211xp5_ASAP7_75t_L g663 ( .A1(n_664), .A2(n_667), .B(n_669), .C(n_678), .Y(n_663) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
OAI221xp5_ASAP7_75t_L g740 ( .A1(n_667), .A2(n_677), .B1(n_741), .B2(n_742), .C(n_744), .Y(n_740) );
INVx1_ASAP7_75t_SL g667 ( .A(n_668), .Y(n_667) );
AOI22xp5_ASAP7_75t_L g669 ( .A1(n_670), .A2(n_672), .B1(n_673), .B2(n_676), .Y(n_669) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
AND2x2_ASAP7_75t_L g673 ( .A(n_674), .B(n_675), .Y(n_673) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
OAI21xp5_ASAP7_75t_SL g678 ( .A1(n_679), .A2(n_680), .B(n_681), .Y(n_678) );
INVx1_ASAP7_75t_SL g741 ( .A(n_680), .Y(n_741) );
INVxp67_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
NOR4xp25_ASAP7_75t_L g683 ( .A(n_684), .B(n_713), .C(n_733), .D(n_740), .Y(n_683) );
OAI211xp5_ASAP7_75t_L g684 ( .A1(n_685), .A2(n_689), .B(n_691), .C(n_709), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_686), .B(n_688), .Y(n_685) );
INVxp67_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
O2A1O1Ixp33_ASAP7_75t_L g691 ( .A1(n_692), .A2(n_695), .B(n_697), .C(n_701), .Y(n_691) );
INVx1_ASAP7_75t_SL g692 ( .A(n_693), .Y(n_692) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
INVx1_ASAP7_75t_SL g720 ( .A(n_698), .Y(n_720) );
OR2x2_ASAP7_75t_L g698 ( .A(n_699), .B(n_700), .Y(n_698) );
OR2x2_ASAP7_75t_L g731 ( .A(n_699), .B(n_732), .Y(n_731) );
OAI21xp33_ASAP7_75t_L g701 ( .A1(n_702), .A2(n_705), .B(n_706), .Y(n_701) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
INVx1_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
HB1xp67_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
AOI221xp5_ASAP7_75t_L g719 ( .A1(n_720), .A2(n_721), .B1(n_723), .B2(n_725), .C(n_727), .Y(n_719) );
INVx1_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVxp67_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_730), .B(n_735), .Y(n_734) );
INVx1_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
INVx1_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
INVx2_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
INVx1_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
INVx1_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
INVx2_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
INVx2_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
endmodule