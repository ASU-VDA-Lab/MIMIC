module fake_jpeg_17215_n_260 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_260);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_260;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_14;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_145;
wire n_20;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_93;
wire n_91;
wire n_54;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_96;

INVx1_ASAP7_75t_L g13 ( 
.A(n_9),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx10_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_26),
.B(n_0),
.Y(n_29)
);

AND2x2_ASAP7_75t_SL g38 ( 
.A(n_29),
.B(n_21),
.Y(n_38)
);

BUFx2_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_30),
.B(n_32),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_29),
.Y(n_53)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_39),
.B(n_44),
.Y(n_59)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_30),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_46),
.B(n_47),
.Y(n_60)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_31),
.Y(n_51)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_51),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_53),
.B(n_68),
.Y(n_74)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_56),
.Y(n_80)
);

AND2x2_ASAP7_75t_SL g57 ( 
.A(n_38),
.B(n_29),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_57),
.B(n_53),
.C(n_63),
.Y(n_83)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_58),
.Y(n_82)
);

BUFx12_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g73 ( 
.A(n_61),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_48),
.A2(n_33),
.B1(n_26),
.B2(n_37),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_62),
.A2(n_51),
.B1(n_52),
.B2(n_49),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_38),
.B(n_33),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_63),
.B(n_67),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_64),
.Y(n_84)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_65),
.Y(n_81)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_66),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_42),
.B(n_33),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_40),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_43),
.B(n_15),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_69),
.B(n_15),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_43),
.B(n_22),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_70),
.B(n_71),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_41),
.B(n_13),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_41),
.B(n_13),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_72),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_60),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_76),
.B(n_89),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_78),
.A2(n_93),
.B1(n_55),
.B2(n_58),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_83),
.B(n_28),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_67),
.A2(n_52),
.B1(n_35),
.B2(n_28),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_85),
.A2(n_90),
.B1(n_92),
.B2(n_89),
.Y(n_114)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_61),
.Y(n_87)
);

BUFx2_ASAP7_75t_L g105 ( 
.A(n_87),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_57),
.A2(n_50),
.B(n_18),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_88),
.A2(n_72),
.B(n_71),
.Y(n_106)
);

OA22x2_ASAP7_75t_L g90 ( 
.A1(n_65),
.A2(n_50),
.B1(n_31),
.B2(n_36),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_61),
.Y(n_91)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_91),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_68),
.A2(n_57),
.B1(n_69),
.B2(n_35),
.Y(n_92)
);

INVx1_ASAP7_75t_SL g93 ( 
.A(n_57),
.Y(n_93)
);

AO22x1_ASAP7_75t_SL g94 ( 
.A1(n_79),
.A2(n_36),
.B1(n_70),
.B2(n_54),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_94),
.A2(n_77),
.B1(n_79),
.B2(n_93),
.Y(n_119)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_81),
.Y(n_95)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_95),
.Y(n_121)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_87),
.Y(n_96)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_96),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_84),
.A2(n_55),
.B1(n_66),
.B2(n_54),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_97),
.A2(n_64),
.B(n_56),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_91),
.B(n_59),
.Y(n_98)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_98),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_99),
.B(n_102),
.Y(n_122)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_81),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_101),
.B(n_104),
.Y(n_117)
);

INVx13_ASAP7_75t_L g102 ( 
.A(n_73),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_75),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_106),
.A2(n_114),
.B(n_88),
.Y(n_120)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_75),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_107),
.B(n_109),
.Y(n_118)
);

INVx13_ASAP7_75t_L g108 ( 
.A(n_73),
.Y(n_108)
);

INVx1_ASAP7_75t_SL g126 ( 
.A(n_108),
.Y(n_126)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_80),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_82),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_110),
.B(n_111),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_86),
.B(n_61),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_112),
.B(n_78),
.Y(n_127)
);

INVx13_ASAP7_75t_L g113 ( 
.A(n_84),
.Y(n_113)
);

INVx1_ASAP7_75t_SL g131 ( 
.A(n_113),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_103),
.B(n_89),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_116),
.B(n_130),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_119),
.A2(n_123),
.B1(n_132),
.B2(n_134),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_120),
.A2(n_124),
.B(n_104),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_112),
.A2(n_77),
.B1(n_74),
.B2(n_83),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_112),
.B(n_92),
.C(n_85),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_125),
.B(n_127),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_106),
.B(n_64),
.C(n_32),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_129),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_114),
.B(n_90),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_94),
.A2(n_90),
.B1(n_37),
.B2(n_36),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_95),
.B(n_64),
.C(n_32),
.Y(n_133)
);

HB1xp67_ASAP7_75t_L g144 ( 
.A(n_133),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_94),
.A2(n_90),
.B1(n_37),
.B2(n_27),
.Y(n_134)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_100),
.Y(n_135)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_135),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_118),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_137),
.B(n_150),
.Y(n_171)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_117),
.Y(n_140)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_140),
.Y(n_172)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_135),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_141),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_142),
.A2(n_145),
.B(n_148),
.Y(n_167)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_121),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_143),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_127),
.B(n_94),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_120),
.A2(n_96),
.B(n_110),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_128),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_149),
.B(n_152),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_115),
.B(n_109),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_129),
.A2(n_101),
.B(n_14),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_151),
.A2(n_158),
.B(n_21),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_136),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_132),
.A2(n_107),
.B1(n_100),
.B2(n_113),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_153),
.A2(n_159),
.B1(n_131),
.B2(n_126),
.Y(n_166)
);

NOR2x1p5_ASAP7_75t_L g154 ( 
.A(n_130),
.B(n_24),
.Y(n_154)
);

AO21x1_ASAP7_75t_L g178 ( 
.A1(n_154),
.A2(n_124),
.B(n_24),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_134),
.A2(n_23),
.B1(n_14),
.B2(n_27),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_156),
.A2(n_157),
.B1(n_19),
.B2(n_16),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_122),
.A2(n_113),
.B1(n_102),
.B2(n_108),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_125),
.A2(n_13),
.B(n_27),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_119),
.A2(n_102),
.B1(n_14),
.B2(n_22),
.Y(n_159)
);

HB1xp67_ASAP7_75t_L g161 ( 
.A(n_139),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_161),
.B(n_170),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_145),
.B(n_123),
.Y(n_163)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_163),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_147),
.B(n_144),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_164),
.B(n_151),
.C(n_154),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_145),
.B(n_133),
.Y(n_165)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_165),
.Y(n_188)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_166),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_157),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_168),
.B(n_173),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_169),
.A2(n_158),
.B(n_23),
.Y(n_181)
);

INVx2_ASAP7_75t_SL g170 ( 
.A(n_153),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_159),
.B(n_126),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_148),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_174),
.B(n_177),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_147),
.B(n_142),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_175),
.B(n_155),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_138),
.B(n_131),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_178),
.B(n_25),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_179),
.A2(n_16),
.B1(n_20),
.B2(n_19),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_146),
.A2(n_105),
.B(n_1),
.Y(n_180)
);

A2O1A1Ixp33_ASAP7_75t_SL g191 ( 
.A1(n_180),
.A2(n_105),
.B(n_1),
.C(n_2),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_181),
.A2(n_191),
.B1(n_20),
.B2(n_176),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_184),
.B(n_185),
.C(n_187),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_164),
.B(n_146),
.C(n_154),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_SL g189 ( 
.A(n_163),
.B(n_105),
.C(n_11),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_189),
.A2(n_169),
.B(n_180),
.Y(n_200)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_190),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_194),
.B(n_186),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_160),
.B(n_10),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_195),
.B(n_171),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_172),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_196),
.B(n_176),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_175),
.B(n_165),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_197),
.B(n_177),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_182),
.A2(n_174),
.B1(n_170),
.B2(n_168),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_198),
.A2(n_202),
.B1(n_191),
.B2(n_1),
.Y(n_216)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_199),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_200),
.A2(n_204),
.B(n_9),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_201),
.B(n_203),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_193),
.A2(n_170),
.B1(n_172),
.B2(n_162),
.Y(n_202)
);

XOR2x2_ASAP7_75t_SL g204 ( 
.A(n_184),
.B(n_167),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_192),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_205),
.B(n_206),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_183),
.A2(n_185),
.B1(n_188),
.B2(n_187),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_208),
.B(n_212),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_209),
.B(n_178),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_197),
.B(n_167),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_211),
.B(n_191),
.C(n_18),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_194),
.B(n_166),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_213),
.B(n_215),
.Y(n_226)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_216),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_204),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_217),
.B(n_211),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_207),
.B(n_191),
.C(n_32),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_218),
.B(n_221),
.C(n_198),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_207),
.B(n_30),
.Y(n_221)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_222),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_205),
.A2(n_10),
.B(n_12),
.Y(n_224)
);

AO21x1_ASAP7_75t_L g231 ( 
.A1(n_224),
.A2(n_210),
.B(n_11),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_225),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_227),
.B(n_221),
.C(n_218),
.Y(n_236)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_219),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_230),
.B(n_231),
.Y(n_235)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_224),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_232),
.B(n_8),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_214),
.B(n_209),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_233),
.B(n_234),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_220),
.B(n_223),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_236),
.B(n_226),
.C(n_228),
.Y(n_244)
);

AOI31xp33_ASAP7_75t_L g237 ( 
.A1(n_229),
.A2(n_217),
.A3(n_213),
.B(n_215),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_237),
.A2(n_239),
.B(n_240),
.Y(n_243)
);

MAJx2_ASAP7_75t_L g239 ( 
.A(n_226),
.B(n_8),
.C(n_10),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g240 ( 
.A1(n_227),
.A2(n_8),
.B(n_4),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_242),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_L g249 ( 
.A1(n_244),
.A2(n_247),
.B(n_248),
.Y(n_249)
);

AOI31xp67_ASAP7_75t_SL g250 ( 
.A1(n_245),
.A2(n_237),
.A3(n_4),
.B(n_5),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_238),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_246),
.A2(n_12),
.B1(n_5),
.B2(n_6),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_241),
.B(n_231),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_235),
.B(n_25),
.Y(n_248)
);

CKINVDCx14_ASAP7_75t_R g254 ( 
.A(n_250),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_251),
.B(n_252),
.C(n_243),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_246),
.A2(n_7),
.B1(n_12),
.B2(n_3),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_253),
.Y(n_255)
);

AOI321xp33_ASAP7_75t_L g256 ( 
.A1(n_255),
.A2(n_249),
.A3(n_254),
.B1(n_30),
.B2(n_25),
.C(n_3),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_256),
.B(n_25),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_257),
.Y(n_258)
);

OAI21x1_ASAP7_75t_L g259 ( 
.A1(n_258),
.A2(n_18),
.B(n_17),
.Y(n_259)
);

NOR3xp33_ASAP7_75t_L g260 ( 
.A(n_259),
.B(n_17),
.C(n_18),
.Y(n_260)
);


endmodule