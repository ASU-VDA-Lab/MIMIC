module real_jpeg_15299_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_598;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_630;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_643;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_498;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_640;
wire n_160;
wire n_211;
wire n_574;
wire n_627;
wire n_595;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_578;
wire n_456;
wire n_620;
wire n_259;
wire n_556;
wire n_507;
wire n_57;
wire n_157;
wire n_560;
wire n_84;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_623;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_605;
wire n_483;
wire n_367;
wire n_639;
wire n_127;
wire n_365;
wire n_356;
wire n_464;
wire n_423;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_621;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_601;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_525;
wire n_221;
wire n_611;
wire n_489;
wire n_393;
wire n_104;
wire n_153;
wire n_634;
wire n_443;
wire n_599;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_607;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_378;
wire n_98;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_214;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_631;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_470;
wire n_372;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_593;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_590;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_612;
wire n_110;
wire n_195;
wire n_592;
wire n_533;
wire n_289;
wire n_117;
wire n_614;
wire n_193;
wire n_382;
wire n_411;
wire n_278;
wire n_314;
wire n_103;
wire n_559;
wire n_232;
wire n_582;
wire n_615;
wire n_448;
wire n_212;
wire n_579;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_583;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_589;
wire n_25;
wire n_542;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_632;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_633;
wire n_497;
wire n_638;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_596;
wire n_312;
wire n_617;
wire n_325;
wire n_316;
wire n_307;
wire n_594;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_604;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_572;
wire n_586;
wire n_548;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_637;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_613;
wire n_265;
wire n_231;
wire n_44;
wire n_635;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_642;
wire n_106;
wire n_172;
wire n_285;
wire n_546;
wire n_531;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_616;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_600;
wire n_392;
wire n_575;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_584;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_622;
wire n_183;
wire n_248;
wire n_192;
wire n_624;
wire n_318;
wire n_537;
wire n_603;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_628;
wire n_413;
wire n_585;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_581;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_587;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_608;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_602;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_610;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_636;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_606;
wire n_245;
wire n_451;
wire n_626;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_597;
wire n_618;
wire n_609;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_619;
wire n_116;
wire n_416;
wire n_513;
wire n_588;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_567;
wire n_51;
wire n_509;
wire n_519;
wire n_205;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_568;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_130;
wire n_641;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_629;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_625;
wire n_591;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_0),
.A2(n_21),
.B(n_642),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g642 ( 
.A(n_0),
.B(n_643),
.Y(n_642)
);

BUFx5_ASAP7_75t_L g244 ( 
.A(n_1),
.Y(n_244)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_1),
.Y(n_286)
);

BUFx3_ASAP7_75t_L g329 ( 
.A(n_1),
.Y(n_329)
);

BUFx5_ASAP7_75t_L g418 ( 
.A(n_1),
.Y(n_418)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_2),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_3),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_3),
.Y(n_90)
);

BUFx5_ASAP7_75t_L g92 ( 
.A(n_3),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g472 ( 
.A(n_3),
.Y(n_472)
);

OAI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_4),
.A2(n_110),
.B1(n_118),
.B2(n_119),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_4),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_4),
.A2(n_118),
.B1(n_196),
.B2(n_199),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_4),
.A2(n_118),
.B1(n_255),
.B2(n_259),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_4),
.A2(n_118),
.B1(n_298),
.B2(n_300),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_5),
.A2(n_186),
.B1(n_188),
.B2(n_190),
.Y(n_185)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_5),
.Y(n_190)
);

OAI22xp33_ASAP7_75t_SL g316 ( 
.A1(n_5),
.A2(n_190),
.B1(n_317),
.B2(n_321),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_5),
.A2(n_190),
.B1(n_336),
.B2(n_340),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_SL g386 ( 
.A1(n_5),
.A2(n_190),
.B1(n_387),
.B2(n_388),
.Y(n_386)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_6),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_6),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g252 ( 
.A(n_6),
.Y(n_252)
);

BUFx4f_ASAP7_75t_L g258 ( 
.A(n_6),
.Y(n_258)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_7),
.Y(n_643)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_8),
.A2(n_218),
.B1(n_220),
.B2(n_221),
.Y(n_217)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_8),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g362 ( 
.A1(n_8),
.A2(n_220),
.B1(n_363),
.B2(n_365),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_8),
.A2(n_63),
.B1(n_113),
.B2(n_220),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_SL g497 ( 
.A1(n_8),
.A2(n_220),
.B1(n_498),
.B2(n_501),
.Y(n_497)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_9),
.A2(n_109),
.B1(n_112),
.B2(n_115),
.Y(n_108)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_9),
.Y(n_115)
);

OAI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_9),
.A2(n_115),
.B1(n_247),
.B2(n_249),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_9),
.A2(n_115),
.B1(n_306),
.B2(n_310),
.Y(n_305)
);

AOI22xp33_ASAP7_75t_L g426 ( 
.A1(n_9),
.A2(n_115),
.B1(n_161),
.B2(n_427),
.Y(n_426)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_10),
.A2(n_46),
.B1(n_52),
.B2(n_56),
.Y(n_45)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_10),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_10),
.A2(n_56),
.B1(n_126),
.B2(n_130),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g280 ( 
.A1(n_10),
.A2(n_56),
.B1(n_281),
.B2(n_282),
.Y(n_280)
);

AOI22xp33_ASAP7_75t_SL g405 ( 
.A1(n_10),
.A2(n_56),
.B1(n_406),
.B2(n_409),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_11),
.A2(n_269),
.B1(n_273),
.B2(n_274),
.Y(n_268)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_11),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_11),
.A2(n_222),
.B1(n_273),
.B2(n_353),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_SL g506 ( 
.A1(n_11),
.A2(n_273),
.B1(n_507),
.B2(n_509),
.Y(n_506)
);

AOI22xp33_ASAP7_75t_SL g518 ( 
.A1(n_11),
.A2(n_273),
.B1(n_519),
.B2(n_522),
.Y(n_518)
);

OAI22xp33_ASAP7_75t_L g209 ( 
.A1(n_12),
.A2(n_210),
.B1(n_213),
.B2(n_214),
.Y(n_209)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_12),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_12),
.A2(n_110),
.B1(n_186),
.B2(n_213),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g489 ( 
.A1(n_12),
.A2(n_213),
.B1(n_259),
.B2(n_490),
.Y(n_489)
);

OAI22xp5_ASAP7_75t_L g584 ( 
.A1(n_12),
.A2(n_213),
.B1(n_585),
.B2(n_588),
.Y(n_584)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_13),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_13),
.Y(n_148)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_13),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_14),
.B(n_236),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g359 ( 
.A1(n_14),
.A2(n_186),
.B(n_235),
.Y(n_359)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_14),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_14),
.B(n_172),
.Y(n_503)
);

OAI22xp5_ASAP7_75t_SL g541 ( 
.A1(n_14),
.A2(n_242),
.B1(n_542),
.B2(n_544),
.Y(n_541)
);

OAI32xp33_ASAP7_75t_L g557 ( 
.A1(n_14),
.A2(n_558),
.A3(n_560),
.B1(n_563),
.B2(n_568),
.Y(n_557)
);

AOI22xp33_ASAP7_75t_SL g576 ( 
.A1(n_14),
.A2(n_394),
.B1(n_577),
.B2(n_579),
.Y(n_576)
);

AOI22xp33_ASAP7_75t_SL g266 ( 
.A1(n_15),
.A2(n_53),
.B1(n_188),
.B2(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_15),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_SL g377 ( 
.A1(n_15),
.A2(n_267),
.B1(n_378),
.B2(n_382),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_SL g483 ( 
.A1(n_15),
.A2(n_267),
.B1(n_484),
.B2(n_486),
.Y(n_483)
);

AOI22xp5_ASAP7_75t_SL g542 ( 
.A1(n_15),
.A2(n_267),
.B1(n_520),
.B2(n_543),
.Y(n_542)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_16),
.A2(n_59),
.B1(n_64),
.B2(n_67),
.Y(n_58)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_16),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_16),
.A2(n_67),
.B1(n_97),
.B2(n_102),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g160 ( 
.A1(n_16),
.A2(n_67),
.B1(n_161),
.B2(n_166),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g288 ( 
.A1(n_16),
.A2(n_67),
.B1(n_289),
.B2(n_292),
.Y(n_288)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_17),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_17),
.Y(n_95)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_17),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_17),
.Y(n_105)
);

BUFx5_ASAP7_75t_L g303 ( 
.A(n_17),
.Y(n_303)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_17),
.Y(n_320)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_17),
.Y(n_324)
);

BUFx3_ASAP7_75t_L g408 ( 
.A(n_17),
.Y(n_408)
);

BUFx3_ASAP7_75t_L g567 ( 
.A(n_17),
.Y(n_567)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

BUFx8_ASAP7_75t_L g31 ( 
.A(n_19),
.Y(n_31)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_19),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g111 ( 
.A(n_19),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_176),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_174),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_68),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_24),
.B(n_68),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_45),
.B1(n_57),
.B2(n_58),
.Y(n_24)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_25),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_25),
.A2(n_45),
.B1(n_57),
.B2(n_170),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_25),
.A2(n_57),
.B1(n_108),
.B2(n_185),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_25),
.A2(n_57),
.B1(n_266),
.B2(n_268),
.Y(n_265)
);

OAI22xp33_ASAP7_75t_L g331 ( 
.A1(n_25),
.A2(n_57),
.B1(n_268),
.B2(n_332),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_25),
.A2(n_57),
.B1(n_266),
.B2(n_359),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_L g423 ( 
.A1(n_25),
.A2(n_57),
.B1(n_332),
.B2(n_424),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_SL g450 ( 
.A1(n_25),
.A2(n_57),
.B1(n_185),
.B2(n_424),
.Y(n_450)
);

AO21x2_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_32),
.B(n_36),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_30),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_31),
.B(n_33),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_32),
.A2(n_226),
.B1(n_234),
.B2(n_237),
.Y(n_225)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_35),
.Y(n_230)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_36),
.A2(n_107),
.B1(n_116),
.B2(n_117),
.Y(n_106)
);

AO22x2_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_40),
.B1(n_41),
.B2(n_43),
.Y(n_36)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_37),
.Y(n_167)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_38),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_39),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_39),
.Y(n_151)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_39),
.Y(n_165)
);

BUFx5_ASAP7_75t_L g233 ( 
.A(n_39),
.Y(n_233)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_41),
.Y(n_223)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_41),
.Y(n_428)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_42),
.Y(n_129)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_42),
.Y(n_133)
);

INVx4_ASAP7_75t_L g198 ( 
.A(n_42),
.Y(n_198)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_42),
.Y(n_581)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_49),
.Y(n_63)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_50),
.Y(n_114)
);

INVx8_ASAP7_75t_L g121 ( 
.A(n_50),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_50),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_51),
.Y(n_272)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_55),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_55),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_57),
.B(n_394),
.Y(n_393)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

BUFx2_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_169),
.C(n_171),
.Y(n_68)
);

FAx1_ASAP7_75t_SL g179 ( 
.A(n_69),
.B(n_169),
.CI(n_171),
.CON(n_179),
.SN(n_179)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_106),
.C(n_122),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_70),
.A2(n_123),
.B1(n_124),
.B2(n_183),
.Y(n_182)
);

INVx1_ASAP7_75t_SL g183 ( 
.A(n_70),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_70),
.B(n_193),
.C(n_194),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g626 ( 
.A(n_70),
.B(n_194),
.Y(n_626)
);

OA21x2_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_82),
.B(n_96),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_71),
.B(n_296),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_71),
.A2(n_82),
.B1(n_305),
.B2(n_316),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_SL g442 ( 
.A1(n_71),
.A2(n_82),
.B1(n_96),
.B2(n_443),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_L g478 ( 
.A1(n_71),
.A2(n_82),
.B1(n_479),
.B2(n_483),
.Y(n_478)
);

AOI22xp5_ASAP7_75t_SL g505 ( 
.A1(n_71),
.A2(n_82),
.B1(n_483),
.B2(n_506),
.Y(n_505)
);

AOI22xp5_ASAP7_75t_L g583 ( 
.A1(n_71),
.A2(n_82),
.B1(n_506),
.B2(n_584),
.Y(n_583)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_72),
.A2(n_361),
.B1(n_362),
.B2(n_369),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g404 ( 
.A1(n_72),
.A2(n_297),
.B1(n_361),
.B2(n_405),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g549 ( 
.A(n_72),
.B(n_394),
.Y(n_549)
);

OAI22xp5_ASAP7_75t_SL g600 ( 
.A1(n_72),
.A2(n_361),
.B1(n_362),
.B2(n_601),
.Y(n_600)
);

BUFx2_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_73),
.B(n_83),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_75),
.B1(n_78),
.B2(n_81),
.Y(n_73)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_74),
.Y(n_81)
);

OR2x2_ASAP7_75t_L g242 ( 
.A(n_75),
.B(n_243),
.Y(n_242)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_75),
.Y(n_500)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_76),
.Y(n_283)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_76),
.Y(n_521)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_77),
.Y(n_263)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_80),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_82),
.B(n_305),
.Y(n_304)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_82),
.Y(n_361)
);

OAI22xp33_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_88),
.B1(n_91),
.B2(n_93),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_86),
.Y(n_562)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_92),
.Y(n_467)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_94),
.A2(n_153),
.B1(n_156),
.B2(n_157),
.Y(n_152)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_94),
.Y(n_299)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_100),
.Y(n_156)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_101),
.Y(n_309)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_101),
.Y(n_368)
);

BUFx3_ASAP7_75t_L g482 ( 
.A(n_101),
.Y(n_482)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_101),
.Y(n_512)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

BUFx12f_ASAP7_75t_L g311 ( 
.A(n_105),
.Y(n_311)
);

INVx4_ASAP7_75t_L g508 ( 
.A(n_105),
.Y(n_508)
);

BUFx3_ASAP7_75t_L g587 ( 
.A(n_105),
.Y(n_587)
);

XNOR2x1_ASAP7_75t_L g181 ( 
.A(n_106),
.B(n_182),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx8_ASAP7_75t_L g236 ( 
.A(n_111),
.Y(n_236)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx6_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_117),
.Y(n_170)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

HB1xp67_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_125),
.A2(n_134),
.B1(n_160),
.B2(n_168),
.Y(n_124)
);

OAI22x1_ASAP7_75t_L g194 ( 
.A1(n_125),
.A2(n_134),
.B1(n_168),
.B2(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_SL g126 ( 
.A(n_127),
.Y(n_126)
);

INVx6_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

HB1xp67_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_131),
.Y(n_383)
);

BUFx3_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_133),
.Y(n_339)
);

OAI22x1_ASAP7_75t_SL g333 ( 
.A1(n_134),
.A2(n_168),
.B1(n_334),
.B2(n_335),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_L g351 ( 
.A1(n_134),
.A2(n_168),
.B1(n_352),
.B2(n_357),
.Y(n_351)
);

OAI22xp33_ASAP7_75t_SL g376 ( 
.A1(n_134),
.A2(n_168),
.B1(n_352),
.B2(n_377),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_L g425 ( 
.A1(n_134),
.A2(n_168),
.B1(n_335),
.B2(n_426),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_SL g575 ( 
.A1(n_134),
.A2(n_168),
.B1(n_377),
.B2(n_576),
.Y(n_575)
);

INVx3_ASAP7_75t_SL g134 ( 
.A(n_135),
.Y(n_134)
);

OAI21xp33_ASAP7_75t_SL g171 ( 
.A1(n_135),
.A2(n_172),
.B(n_173),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_135),
.A2(n_172),
.B1(n_209),
.B2(n_217),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_135),
.A2(n_172),
.B1(n_440),
.B2(n_441),
.Y(n_439)
);

OA21x2_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_145),
.B(n_152),
.Y(n_135)
);

INVxp33_ASAP7_75t_L g568 ( 
.A(n_136),
.Y(n_568)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_142),
.Y(n_136)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

BUFx3_ASAP7_75t_L g201 ( 
.A(n_144),
.Y(n_201)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_144),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_149),
.Y(n_145)
);

INVx6_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_148),
.Y(n_155)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_151),
.Y(n_212)
);

INVx3_ASAP7_75t_L g343 ( 
.A(n_151),
.Y(n_343)
);

BUFx2_ASAP7_75t_L g168 ( 
.A(n_152),
.Y(n_168)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVxp33_ASAP7_75t_L g173 ( 
.A(n_160),
.Y(n_173)
);

INVx8_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_164),
.Y(n_356)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

BUFx2_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_168),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_202),
.B(n_640),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_180),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g641 ( 
.A(n_179),
.B(n_180),
.Y(n_641)
);

BUFx24_ASAP7_75t_SL g644 ( 
.A(n_179),
.Y(n_644)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_184),
.C(n_191),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g621 ( 
.A1(n_181),
.A2(n_184),
.B1(n_193),
.B2(n_622),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_181),
.Y(n_622)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_184),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g625 ( 
.A1(n_184),
.A2(n_193),
.B1(n_626),
.B2(n_627),
.Y(n_625)
);

INVx5_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx3_ASAP7_75t_SL g188 ( 
.A(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g620 ( 
.A(n_192),
.B(n_621),
.Y(n_620)
);

INVxp67_ASAP7_75t_L g441 ( 
.A(n_195),
.Y(n_441)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx6_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx6_ASAP7_75t_L g381 ( 
.A(n_198),
.Y(n_381)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_203),
.A2(n_616),
.B(n_637),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_204),
.A2(n_454),
.B(n_611),
.Y(n_203)
);

NAND3xp33_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_397),
.C(n_432),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_206),
.A2(n_344),
.B(n_370),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g612 ( 
.A(n_206),
.B(n_344),
.C(n_613),
.Y(n_612)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_275),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_207),
.B(n_276),
.C(n_312),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_224),
.C(n_264),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_208),
.A2(n_264),
.B1(n_265),
.B2(n_347),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_208),
.Y(n_347)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_209),
.Y(n_357)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

HB1xp67_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

BUFx2_ASAP7_75t_SL g215 ( 
.A(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_217),
.Y(n_334)
);

HB1xp67_ASAP7_75t_L g559 ( 
.A(n_218),
.Y(n_559)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_219),
.Y(n_578)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g345 ( 
.A(n_224),
.B(n_346),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_241),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_225),
.B(n_241),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_231),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx4_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx2_ASAP7_75t_SL g240 ( 
.A(n_233),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx3_ASAP7_75t_SL g274 ( 
.A(n_236),
.Y(n_274)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_242),
.A2(n_245),
.B1(n_253),
.B2(n_254),
.Y(n_241)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_242),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_242),
.A2(n_254),
.B1(n_280),
.B2(n_326),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_L g414 ( 
.A1(n_242),
.A2(n_288),
.B(n_415),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_L g488 ( 
.A1(n_242),
.A2(n_489),
.B1(n_494),
.B2(n_496),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_SL g547 ( 
.A1(n_242),
.A2(n_518),
.B1(n_542),
.B2(n_548),
.Y(n_547)
);

INVx6_ASAP7_75t_L g253 ( 
.A(n_243),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g516 ( 
.A1(n_243),
.A2(n_278),
.B1(n_517),
.B2(n_526),
.Y(n_516)
);

BUFx12f_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_246),
.A2(n_278),
.B1(n_386),
.B2(n_392),
.Y(n_385)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_247),
.Y(n_501)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_247),
.Y(n_543)
);

INVx5_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

OAI32xp33_ASAP7_75t_L g460 ( 
.A1(n_250),
.A2(n_461),
.A3(n_464),
.B1(n_468),
.B2(n_470),
.Y(n_460)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx4_ASAP7_75t_L g281 ( 
.A(n_252),
.Y(n_281)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_252),
.Y(n_291)
);

INVx5_ASAP7_75t_L g493 ( 
.A(n_252),
.Y(n_493)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_258),
.Y(n_476)
);

INVx3_ASAP7_75t_L g534 ( 
.A(n_258),
.Y(n_534)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx4_ASAP7_75t_L g391 ( 
.A(n_263),
.Y(n_391)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

BUFx2_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx4_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_312),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_294),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g421 ( 
.A1(n_277),
.A2(n_295),
.B(n_304),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_278),
.A2(n_279),
.B1(n_284),
.B2(n_287),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g569 ( 
.A1(n_278),
.A2(n_386),
.B1(n_497),
.B2(n_570),
.Y(n_569)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_281),
.Y(n_387)
);

BUFx2_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

BUFx3_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx6_ASAP7_75t_L g548 ( 
.A(n_285),
.Y(n_548)
);

INVx3_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_286),
.Y(n_540)
);

INVxp67_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_291),
.Y(n_293)
);

HB1xp67_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_304),
.Y(n_294)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx4_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

BUFx6f_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_303),
.Y(n_364)
);

BUFx2_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

INVx5_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx1_ASAP7_75t_SL g486 ( 
.A(n_311),
.Y(n_486)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_330),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g401 ( 
.A(n_313),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_314),
.B(n_325),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_314),
.A2(n_315),
.B1(n_325),
.B2(n_349),
.Y(n_348)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_316),
.Y(n_369)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_320),
.Y(n_412)
);

INVx4_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

BUFx6f_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

BUFx6f_ASAP7_75t_L g589 ( 
.A(n_324),
.Y(n_589)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_325),
.Y(n_349)
);

INVx5_ASAP7_75t_L g392 ( 
.A(n_326),
.Y(n_392)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_326),
.Y(n_570)
);

INVx6_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx5_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx3_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

BUFx3_ASAP7_75t_L g495 ( 
.A(n_329),
.Y(n_495)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_331),
.B(n_333),
.Y(n_330)
);

HB1xp67_ASAP7_75t_L g400 ( 
.A(n_331),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_333),
.B(n_400),
.C(n_401),
.Y(n_399)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_345),
.B(n_348),
.C(n_350),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_SL g395 ( 
.A(n_345),
.B(n_396),
.Y(n_395)
);

XNOR2x1_ASAP7_75t_L g396 ( 
.A(n_348),
.B(n_350),
.Y(n_396)
);

MAJx2_ASAP7_75t_L g350 ( 
.A(n_351),
.B(n_358),
.C(n_360),
.Y(n_350)
);

XOR2xp5_ASAP7_75t_L g373 ( 
.A(n_351),
.B(n_360),
.Y(n_373)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_SL g372 ( 
.A(n_358),
.B(n_373),
.Y(n_372)
);

BUFx2_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

INVx1_ASAP7_75t_SL g365 ( 
.A(n_366),
.Y(n_365)
);

BUFx3_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_371),
.B(n_395),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_371),
.B(n_395),
.Y(n_613)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_372),
.B(n_374),
.C(n_375),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_L g607 ( 
.A(n_372),
.B(n_608),
.Y(n_607)
);

XNOR2xp5_ASAP7_75t_L g608 ( 
.A(n_374),
.B(n_375),
.Y(n_608)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_376),
.B(n_384),
.C(n_393),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g594 ( 
.A(n_376),
.B(n_595),
.Y(n_594)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

INVx5_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

INVx4_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_SL g595 ( 
.A1(n_384),
.A2(n_385),
.B1(n_393),
.B2(n_596),
.Y(n_595)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

BUFx6f_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

BUFx6f_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

INVx3_ASAP7_75t_L g525 ( 
.A(n_391),
.Y(n_525)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_393),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_394),
.B(n_469),
.Y(n_468)
);

OAI21xp33_ASAP7_75t_SL g479 ( 
.A1(n_394),
.A2(n_468),
.B(n_480),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_SL g535 ( 
.A(n_394),
.B(n_536),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g563 ( 
.A(n_394),
.B(n_564),
.Y(n_563)
);

A2O1A1O1Ixp25_ASAP7_75t_L g611 ( 
.A1(n_397),
.A2(n_432),
.B(n_612),
.C(n_614),
.D(n_615),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_SL g397 ( 
.A(n_398),
.B(n_431),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g614 ( 
.A(n_398),
.B(n_431),
.Y(n_614)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_399),
.B(n_402),
.Y(n_398)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_399),
.Y(n_453)
);

AOI22xp5_ASAP7_75t_L g402 ( 
.A1(n_403),
.A2(n_420),
.B1(n_429),
.B2(n_430),
.Y(n_402)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_403),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_403),
.B(n_430),
.C(n_453),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_SL g403 ( 
.A1(n_404),
.A2(n_413),
.B1(n_414),
.B2(n_419),
.Y(n_403)
);

INVxp67_ASAP7_75t_L g419 ( 
.A(n_404),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_404),
.B(n_414),
.Y(n_446)
);

INVxp33_ASAP7_75t_SL g443 ( 
.A(n_405),
.Y(n_443)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_406),
.Y(n_469)
);

BUFx2_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

INVx3_ASAP7_75t_L g485 ( 
.A(n_408),
.Y(n_485)
);

BUFx3_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

INVx3_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

HB1xp67_ASAP7_75t_L g463 ( 
.A(n_412),
.Y(n_463)
);

AOI22xp5_ASAP7_75t_L g448 ( 
.A1(n_413),
.A2(n_414),
.B1(n_449),
.B2(n_450),
.Y(n_448)
);

OAI21xp5_ASAP7_75t_L g629 ( 
.A1(n_413),
.A2(n_450),
.B(n_451),
.Y(n_629)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

INVx3_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_420),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_L g420 ( 
.A(n_421),
.B(n_422),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_421),
.B(n_435),
.C(n_436),
.Y(n_434)
);

XOR2xp5_ASAP7_75t_L g422 ( 
.A(n_423),
.B(n_425),
.Y(n_422)
);

HB1xp67_ASAP7_75t_L g436 ( 
.A(n_423),
.Y(n_436)
);

HB1xp67_ASAP7_75t_L g435 ( 
.A(n_425),
.Y(n_435)
);

INVxp67_ASAP7_75t_L g440 ( 
.A(n_426),
.Y(n_440)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_SL g432 ( 
.A(n_433),
.B(n_452),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g615 ( 
.A(n_433),
.B(n_452),
.Y(n_615)
);

XNOR2xp5_ASAP7_75t_L g433 ( 
.A(n_434),
.B(n_437),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g631 ( 
.A(n_434),
.B(n_632),
.C(n_633),
.Y(n_631)
);

XNOR2xp5_ASAP7_75t_L g437 ( 
.A(n_438),
.B(n_445),
.Y(n_437)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_438),
.Y(n_633)
);

OAI21xp5_ASAP7_75t_SL g438 ( 
.A1(n_439),
.A2(n_442),
.B(n_444),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_439),
.B(n_442),
.Y(n_444)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_444),
.Y(n_628)
);

AOI22xp5_ASAP7_75t_L g635 ( 
.A1(n_444),
.A2(n_625),
.B1(n_628),
.B2(n_636),
.Y(n_635)
);

INVxp67_ASAP7_75t_L g632 ( 
.A(n_445),
.Y(n_632)
);

OAI22xp5_ASAP7_75t_SL g445 ( 
.A1(n_446),
.A2(n_447),
.B1(n_448),
.B2(n_451),
.Y(n_445)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_446),
.Y(n_451)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_450),
.Y(n_449)
);

AOI21x1_ASAP7_75t_L g454 ( 
.A1(n_455),
.A2(n_606),
.B(n_610),
.Y(n_454)
);

OAI21x1_ASAP7_75t_L g455 ( 
.A1(n_456),
.A2(n_591),
.B(n_605),
.Y(n_455)
);

AOI21xp5_ASAP7_75t_L g456 ( 
.A1(n_457),
.A2(n_553),
.B(n_590),
.Y(n_456)
);

OAI21x1_ASAP7_75t_L g457 ( 
.A1(n_458),
.A2(n_514),
.B(n_552),
.Y(n_457)
);

AND2x2_ASAP7_75t_L g458 ( 
.A(n_459),
.B(n_487),
.Y(n_458)
);

OR2x2_ASAP7_75t_L g552 ( 
.A(n_459),
.B(n_487),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_460),
.B(n_477),
.Y(n_459)
);

AOI22xp5_ASAP7_75t_L g527 ( 
.A1(n_460),
.A2(n_477),
.B1(n_478),
.B2(n_528),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_460),
.Y(n_528)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_462),
.Y(n_461)
);

HB1xp67_ASAP7_75t_L g462 ( 
.A(n_463),
.Y(n_462)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_465),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_466),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_467),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_471),
.B(n_473),
.Y(n_470)
);

INVx6_ASAP7_75t_L g471 ( 
.A(n_472),
.Y(n_471)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_474),
.Y(n_473)
);

BUFx3_ASAP7_75t_L g474 ( 
.A(n_475),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_476),
.Y(n_475)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_478),
.Y(n_477)
);

BUFx2_ASAP7_75t_L g480 ( 
.A(n_481),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_482),
.Y(n_481)
);

INVx3_ASAP7_75t_L g484 ( 
.A(n_485),
.Y(n_484)
);

XNOR2xp5_ASAP7_75t_L g487 ( 
.A(n_488),
.B(n_502),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g554 ( 
.A(n_488),
.B(n_504),
.C(n_513),
.Y(n_554)
);

INVxp67_ASAP7_75t_L g526 ( 
.A(n_489),
.Y(n_526)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_491),
.Y(n_490)
);

HB1xp67_ASAP7_75t_L g491 ( 
.A(n_492),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_493),
.Y(n_492)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_495),
.Y(n_494)
);

INVxp67_ASAP7_75t_L g496 ( 
.A(n_497),
.Y(n_496)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_499),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_500),
.Y(n_499)
);

OAI22xp5_ASAP7_75t_L g502 ( 
.A1(n_503),
.A2(n_504),
.B1(n_505),
.B2(n_513),
.Y(n_502)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_503),
.Y(n_513)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_505),
.Y(n_504)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_508),
.Y(n_507)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_510),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_511),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_512),
.Y(n_511)
);

AOI21xp5_ASAP7_75t_L g514 ( 
.A1(n_515),
.A2(n_529),
.B(n_551),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_516),
.B(n_527),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g551 ( 
.A(n_516),
.B(n_527),
.Y(n_551)
);

INVxp67_ASAP7_75t_L g517 ( 
.A(n_518),
.Y(n_517)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_520),
.Y(n_519)
);

HB1xp67_ASAP7_75t_L g520 ( 
.A(n_521),
.Y(n_520)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_523),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_524),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_525),
.Y(n_524)
);

OAI21xp5_ASAP7_75t_L g529 ( 
.A1(n_530),
.A2(n_546),
.B(n_550),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_531),
.B(n_541),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_532),
.B(n_535),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_533),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_534),
.Y(n_533)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_537),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_538),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_539),
.Y(n_538)
);

BUFx6f_ASAP7_75t_L g545 ( 
.A(n_539),
.Y(n_545)
);

BUFx6f_ASAP7_75t_L g539 ( 
.A(n_540),
.Y(n_539)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_545),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_547),
.B(n_549),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_547),
.B(n_549),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_554),
.B(n_555),
.Y(n_553)
);

NOR2xp33_ASAP7_75t_L g590 ( 
.A(n_554),
.B(n_555),
.Y(n_590)
);

XOR2xp5_ASAP7_75t_L g555 ( 
.A(n_556),
.B(n_573),
.Y(n_555)
);

MAJIxp5_ASAP7_75t_L g604 ( 
.A(n_556),
.B(n_574),
.C(n_583),
.Y(n_604)
);

AOI22xp5_ASAP7_75t_L g556 ( 
.A1(n_557),
.A2(n_569),
.B1(n_571),
.B2(n_572),
.Y(n_556)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_557),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_557),
.B(n_572),
.Y(n_599)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_559),
.Y(n_558)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_561),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_562),
.Y(n_561)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_565),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_566),
.Y(n_565)
);

INVx3_ASAP7_75t_L g566 ( 
.A(n_567),
.Y(n_566)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_569),
.Y(n_572)
);

OAI22xp5_ASAP7_75t_SL g573 ( 
.A1(n_574),
.A2(n_575),
.B1(n_582),
.B2(n_583),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_575),
.Y(n_574)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_578),
.Y(n_577)
);

BUFx3_ASAP7_75t_L g579 ( 
.A(n_580),
.Y(n_579)
);

INVx2_ASAP7_75t_SL g580 ( 
.A(n_581),
.Y(n_580)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_583),
.Y(n_582)
);

INVxp67_ASAP7_75t_L g601 ( 
.A(n_584),
.Y(n_601)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_586),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_587),
.Y(n_586)
);

BUFx6f_ASAP7_75t_L g588 ( 
.A(n_589),
.Y(n_588)
);

NOR2xp67_ASAP7_75t_L g591 ( 
.A(n_592),
.B(n_604),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_592),
.B(n_604),
.Y(n_605)
);

OAI22xp5_ASAP7_75t_SL g592 ( 
.A1(n_593),
.A2(n_594),
.B1(n_597),
.B2(n_598),
.Y(n_592)
);

MAJIxp5_ASAP7_75t_L g609 ( 
.A(n_593),
.B(n_600),
.C(n_602),
.Y(n_609)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_594),
.Y(n_593)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_598),
.Y(n_597)
);

OAI22xp5_ASAP7_75t_SL g598 ( 
.A1(n_599),
.A2(n_600),
.B1(n_602),
.B2(n_603),
.Y(n_598)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_599),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_600),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_SL g606 ( 
.A(n_607),
.B(n_609),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_L g610 ( 
.A(n_607),
.B(n_609),
.Y(n_610)
);

INVxp67_ASAP7_75t_L g616 ( 
.A(n_617),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_618),
.B(n_630),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_619),
.Y(n_618)
);

OAI21xp5_ASAP7_75t_L g637 ( 
.A1(n_619),
.A2(n_638),
.B(n_639),
.Y(n_637)
);

NOR2x1_ASAP7_75t_L g619 ( 
.A(n_620),
.B(n_623),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_620),
.B(n_623),
.Y(n_639)
);

MAJIxp5_ASAP7_75t_L g623 ( 
.A(n_624),
.B(n_628),
.C(n_629),
.Y(n_623)
);

HB1xp67_ASAP7_75t_L g624 ( 
.A(n_625),
.Y(n_624)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_625),
.Y(n_636)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_626),
.Y(n_627)
);

XOR2xp5_ASAP7_75t_L g634 ( 
.A(n_629),
.B(n_635),
.Y(n_634)
);

OR2x2_ASAP7_75t_L g630 ( 
.A(n_631),
.B(n_634),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_631),
.B(n_634),
.Y(n_638)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_641),
.Y(n_640)
);


endmodule