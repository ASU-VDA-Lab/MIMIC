module fake_jpeg_503_n_640 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_640);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_640;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_543;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_596;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_442;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_17),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx8_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_5),
.Y(n_29)
);

INVx1_ASAP7_75t_SL g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_17),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_1),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_12),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

BUFx24_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_3),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_16),
.Y(n_46)
);

INVx11_ASAP7_75t_SL g47 ( 
.A(n_6),
.Y(n_47)
);

CKINVDCx16_ASAP7_75t_R g48 ( 
.A(n_1),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_1),
.Y(n_49)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_10),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_13),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_15),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_15),
.Y(n_53)
);

BUFx12_ASAP7_75t_L g54 ( 
.A(n_12),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_0),
.B(n_10),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_14),
.Y(n_56)
);

BUFx10_ASAP7_75t_L g57 ( 
.A(n_4),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_7),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

BUFx10_ASAP7_75t_L g145 ( 
.A(n_59),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_55),
.B(n_8),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_60),
.B(n_74),
.Y(n_175)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_27),
.Y(n_61)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_61),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_62),
.Y(n_134)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_26),
.Y(n_63)
);

INVx5_ASAP7_75t_L g174 ( 
.A(n_63),
.Y(n_174)
);

BUFx5_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

INVx2_ASAP7_75t_SL g132 ( 
.A(n_64),
.Y(n_132)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_27),
.Y(n_65)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_65),
.Y(n_144)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_33),
.Y(n_66)
);

INVx4_ASAP7_75t_SL g137 ( 
.A(n_66),
.Y(n_137)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_26),
.Y(n_67)
);

INVx5_ASAP7_75t_L g176 ( 
.A(n_67),
.Y(n_176)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_68),
.Y(n_148)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_69),
.Y(n_151)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_33),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g178 ( 
.A(n_70),
.Y(n_178)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_26),
.Y(n_71)
);

INVx8_ASAP7_75t_L g140 ( 
.A(n_71),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_33),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g187 ( 
.A(n_72),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_42),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_73),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_55),
.B(n_8),
.Y(n_74)
);

BUFx8_ASAP7_75t_L g75 ( 
.A(n_26),
.Y(n_75)
);

BUFx2_ASAP7_75t_SL g198 ( 
.A(n_75),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_42),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_76),
.Y(n_177)
);

BUFx2_ASAP7_75t_L g77 ( 
.A(n_26),
.Y(n_77)
);

INVx2_ASAP7_75t_SL g142 ( 
.A(n_77),
.Y(n_142)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_35),
.Y(n_78)
);

INVx2_ASAP7_75t_SL g154 ( 
.A(n_78),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_42),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_79),
.Y(n_179)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_35),
.Y(n_80)
);

INVx2_ASAP7_75t_SL g159 ( 
.A(n_80),
.Y(n_159)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_35),
.Y(n_81)
);

INVx2_ASAP7_75t_SL g180 ( 
.A(n_81),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_43),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_82),
.Y(n_191)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_21),
.Y(n_83)
);

INVx5_ASAP7_75t_L g200 ( 
.A(n_83),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_43),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_84),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_19),
.B(n_8),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_85),
.B(n_93),
.Y(n_131)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_36),
.Y(n_86)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_86),
.Y(n_157)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_20),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g201 ( 
.A(n_87),
.Y(n_201)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_23),
.Y(n_88)
);

HB1xp67_ASAP7_75t_L g139 ( 
.A(n_88),
.Y(n_139)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_43),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_89),
.Y(n_206)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_20),
.Y(n_90)
);

BUFx2_ASAP7_75t_L g163 ( 
.A(n_90),
.Y(n_163)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_21),
.Y(n_91)
);

INVx3_ASAP7_75t_SL g171 ( 
.A(n_91),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_43),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_92),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g93 ( 
.A(n_57),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_36),
.Y(n_94)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_94),
.Y(n_161)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_21),
.Y(n_95)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_95),
.Y(n_196)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_23),
.Y(n_96)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_96),
.Y(n_172)
);

INVx3_ASAP7_75t_SL g97 ( 
.A(n_20),
.Y(n_97)
);

HB1xp67_ASAP7_75t_L g160 ( 
.A(n_97),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_48),
.B(n_8),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_98),
.B(n_30),
.Y(n_129)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_23),
.Y(n_99)
);

HB1xp67_ASAP7_75t_L g169 ( 
.A(n_99),
.Y(n_169)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_28),
.Y(n_100)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_100),
.Y(n_135)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_28),
.Y(n_101)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_101),
.Y(n_153)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_32),
.Y(n_102)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_102),
.Y(n_182)
);

CKINVDCx14_ASAP7_75t_R g103 ( 
.A(n_48),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_103),
.B(n_120),
.Y(n_133)
);

BUFx12_ASAP7_75t_L g104 ( 
.A(n_44),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_104),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_38),
.Y(n_105)
);

INVx6_ASAP7_75t_L g167 ( 
.A(n_105),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_38),
.Y(n_106)
);

INVx6_ASAP7_75t_L g203 ( 
.A(n_106),
.Y(n_203)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_21),
.Y(n_107)
);

INVx4_ASAP7_75t_L g219 ( 
.A(n_107),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_38),
.Y(n_108)
);

INVx6_ASAP7_75t_L g204 ( 
.A(n_108),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_19),
.B(n_9),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_109),
.B(n_115),
.Y(n_136)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_31),
.Y(n_110)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_110),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_28),
.Y(n_111)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_111),
.Y(n_166)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_31),
.Y(n_112)
);

INVx4_ASAP7_75t_L g205 ( 
.A(n_112),
.Y(n_205)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_32),
.Y(n_113)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_113),
.Y(n_190)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_32),
.Y(n_114)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_114),
.Y(n_195)
);

BUFx12_ASAP7_75t_L g115 ( 
.A(n_44),
.Y(n_115)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_22),
.Y(n_116)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_116),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_22),
.Y(n_117)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_117),
.Y(n_202)
);

INVx4_ASAP7_75t_SL g118 ( 
.A(n_44),
.Y(n_118)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_118),
.Y(n_141)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_31),
.Y(n_119)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_119),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_25),
.B(n_9),
.Y(n_120)
);

BUFx12f_ASAP7_75t_L g121 ( 
.A(n_54),
.Y(n_121)
);

INVx11_ASAP7_75t_L g138 ( 
.A(n_121),
.Y(n_138)
);

INVx8_ASAP7_75t_L g122 ( 
.A(n_22),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_122),
.B(n_123),
.Y(n_184)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_50),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_22),
.Y(n_124)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_124),
.Y(n_156)
);

BUFx5_ASAP7_75t_L g125 ( 
.A(n_44),
.Y(n_125)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_125),
.Y(n_165)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_34),
.Y(n_126)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_126),
.Y(n_194)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_50),
.Y(n_127)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_127),
.Y(n_212)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_34),
.Y(n_128)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_128),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_129),
.B(n_152),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_71),
.A2(n_30),
.B1(n_50),
.B2(n_49),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_130),
.A2(n_149),
.B1(n_162),
.B2(n_164),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_60),
.B(n_58),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_146),
.B(n_150),
.Y(n_285)
);

O2A1O1Ixp33_ASAP7_75t_SL g147 ( 
.A1(n_75),
.A2(n_44),
.B(n_30),
.C(n_56),
.Y(n_147)
);

A2O1A1Ixp33_ASAP7_75t_L g268 ( 
.A1(n_147),
.A2(n_130),
.B(n_164),
.C(n_162),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_74),
.A2(n_120),
.B1(n_98),
.B2(n_108),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_103),
.B(n_46),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_118),
.B(n_46),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_121),
.B(n_51),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_158),
.B(n_168),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_71),
.A2(n_40),
.B1(n_29),
.B2(n_25),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_77),
.A2(n_49),
.B1(n_40),
.B2(n_29),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_121),
.B(n_51),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_59),
.B(n_41),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_173),
.B(n_183),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_63),
.A2(n_58),
.B1(n_39),
.B2(n_56),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_181),
.A2(n_185),
.B1(n_186),
.B2(n_189),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_67),
.B(n_24),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_83),
.A2(n_39),
.B1(n_52),
.B2(n_53),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_L g186 ( 
.A1(n_105),
.A2(n_106),
.B1(n_124),
.B2(n_117),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_97),
.B(n_52),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_188),
.B(n_199),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_91),
.A2(n_53),
.B1(n_41),
.B2(n_37),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_89),
.A2(n_37),
.B1(n_24),
.B2(n_57),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_193),
.A2(n_217),
.B1(n_141),
.B2(n_92),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_62),
.B(n_10),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_73),
.B(n_9),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_209),
.B(n_210),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_76),
.B(n_9),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_79),
.B(n_11),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_211),
.B(n_215),
.Y(n_295)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_95),
.Y(n_214)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_214),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_107),
.B(n_11),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_122),
.B(n_11),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_216),
.B(n_7),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_82),
.A2(n_57),
.B1(n_54),
.B2(n_7),
.Y(n_217)
);

BUFx3_ASAP7_75t_L g220 ( 
.A(n_140),
.Y(n_220)
);

INVx4_ASAP7_75t_L g333 ( 
.A(n_220),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_133),
.B(n_0),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_221),
.B(n_256),
.Y(n_305)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_202),
.Y(n_222)
);

BUFx2_ASAP7_75t_L g327 ( 
.A(n_222),
.Y(n_327)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_198),
.Y(n_223)
);

INVx4_ASAP7_75t_L g338 ( 
.A(n_223),
.Y(n_338)
);

AND2x2_ASAP7_75t_L g322 ( 
.A(n_224),
.B(n_253),
.Y(n_322)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_219),
.Y(n_225)
);

INVx3_ASAP7_75t_L g301 ( 
.A(n_225),
.Y(n_301)
);

AOI22xp33_ASAP7_75t_L g227 ( 
.A1(n_194),
.A2(n_84),
.B1(n_57),
.B2(n_54),
.Y(n_227)
);

OAI22xp33_ASAP7_75t_SL g310 ( 
.A1(n_227),
.A2(n_240),
.B1(n_282),
.B2(n_288),
.Y(n_310)
);

INVx5_ASAP7_75t_L g229 ( 
.A(n_140),
.Y(n_229)
);

INVx1_ASAP7_75t_SL g336 ( 
.A(n_229),
.Y(n_336)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_208),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_230),
.B(n_234),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_160),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_231),
.B(n_246),
.Y(n_314)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_197),
.Y(n_233)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_233),
.Y(n_321)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_163),
.Y(n_234)
);

INVx8_ASAP7_75t_L g236 ( 
.A(n_208),
.Y(n_236)
);

INVx6_ASAP7_75t_L g345 ( 
.A(n_236),
.Y(n_345)
);

AOI22x1_ASAP7_75t_SL g237 ( 
.A1(n_147),
.A2(n_57),
.B1(n_104),
.B2(n_115),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g318 ( 
.A(n_237),
.Y(n_318)
);

INVxp67_ASAP7_75t_SL g238 ( 
.A(n_165),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g299 ( 
.A(n_238),
.Y(n_299)
);

INVx4_ASAP7_75t_L g239 ( 
.A(n_142),
.Y(n_239)
);

HB1xp67_ASAP7_75t_L g300 ( 
.A(n_239),
.Y(n_300)
);

AOI22xp33_ASAP7_75t_L g240 ( 
.A1(n_156),
.A2(n_57),
.B1(n_54),
.B2(n_7),
.Y(n_240)
);

INVx4_ASAP7_75t_L g241 ( 
.A(n_142),
.Y(n_241)
);

HB1xp67_ASAP7_75t_L g356 ( 
.A(n_241),
.Y(n_356)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_134),
.Y(n_242)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_242),
.Y(n_344)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_154),
.Y(n_243)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_243),
.Y(n_302)
);

AND2x2_ASAP7_75t_SL g245 ( 
.A(n_143),
.B(n_0),
.Y(n_245)
);

CKINVDCx14_ASAP7_75t_R g307 ( 
.A(n_245),
.Y(n_307)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_213),
.Y(n_247)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_247),
.Y(n_304)
);

OAI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_186),
.A2(n_54),
.B1(n_6),
.B2(n_13),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_248),
.A2(n_179),
.B1(n_192),
.B2(n_191),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_136),
.B(n_16),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_249),
.B(n_250),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_139),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_175),
.A2(n_18),
.B1(n_14),
.B2(n_13),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_251),
.A2(n_296),
.B1(n_204),
.B2(n_203),
.Y(n_308)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_154),
.Y(n_252)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_252),
.Y(n_311)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_157),
.B(n_161),
.Y(n_253)
);

INVx6_ASAP7_75t_L g254 ( 
.A(n_134),
.Y(n_254)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_254),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_169),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_255),
.B(n_262),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_144),
.B(n_0),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_159),
.Y(n_257)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_257),
.Y(n_329)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_132),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g347 ( 
.A(n_258),
.Y(n_347)
);

BUFx2_ASAP7_75t_L g259 ( 
.A(n_171),
.Y(n_259)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_259),
.Y(n_334)
);

INVx3_ASAP7_75t_L g261 ( 
.A(n_219),
.Y(n_261)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_261),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_131),
.B(n_14),
.Y(n_262)
);

HB1xp67_ASAP7_75t_L g264 ( 
.A(n_159),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_264),
.Y(n_309)
);

BUFx5_ASAP7_75t_L g265 ( 
.A(n_218),
.Y(n_265)
);

INVx13_ASAP7_75t_L g303 ( 
.A(n_265),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_148),
.B(n_0),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_266),
.B(n_272),
.Y(n_306)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_180),
.Y(n_267)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_267),
.Y(n_354)
);

O2A1O1Ixp33_ASAP7_75t_L g341 ( 
.A1(n_268),
.A2(n_178),
.B(n_187),
.C(n_145),
.Y(n_341)
);

INVx6_ASAP7_75t_L g269 ( 
.A(n_170),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_269),
.Y(n_352)
);

AND2x2_ASAP7_75t_L g270 ( 
.A(n_151),
.B(n_2),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_270),
.B(n_274),
.C(n_245),
.Y(n_312)
);

BUFx3_ASAP7_75t_L g271 ( 
.A(n_174),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_271),
.B(n_273),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_172),
.B(n_2),
.Y(n_272)
);

INVx3_ASAP7_75t_L g273 ( 
.A(n_174),
.Y(n_273)
);

AND2x2_ASAP7_75t_L g274 ( 
.A(n_180),
.B(n_2),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_184),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_275),
.B(n_278),
.Y(n_343)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_185),
.A2(n_181),
.B(n_189),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g330 ( 
.A1(n_276),
.A2(n_135),
.B(n_153),
.Y(n_330)
);

BUFx6f_ASAP7_75t_L g277 ( 
.A(n_170),
.Y(n_277)
);

AOI22xp33_ASAP7_75t_SL g298 ( 
.A1(n_277),
.A2(n_284),
.B1(n_289),
.B2(n_290),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_184),
.Y(n_278)
);

BUFx2_ASAP7_75t_L g279 ( 
.A(n_171),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_279),
.B(n_283),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_163),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_280),
.B(n_281),
.Y(n_351)
);

INVx3_ASAP7_75t_L g281 ( 
.A(n_176),
.Y(n_281)
);

AOI22xp33_ASAP7_75t_L g282 ( 
.A1(n_182),
.A2(n_18),
.B1(n_4),
.B2(n_5),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_167),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_167),
.Y(n_284)
);

INVx3_ASAP7_75t_L g286 ( 
.A(n_176),
.Y(n_286)
);

AOI22xp33_ASAP7_75t_SL g350 ( 
.A1(n_286),
.A2(n_293),
.B1(n_223),
.B2(n_259),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_166),
.A2(n_18),
.B1(n_4),
.B2(n_5),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_L g319 ( 
.A1(n_287),
.A2(n_205),
.B(n_155),
.Y(n_319)
);

AOI22xp33_ASAP7_75t_L g288 ( 
.A1(n_190),
.A2(n_3),
.B1(n_5),
.B2(n_195),
.Y(n_288)
);

INVx1_ASAP7_75t_SL g289 ( 
.A(n_137),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_212),
.Y(n_290)
);

AOI22xp33_ASAP7_75t_SL g291 ( 
.A1(n_132),
.A2(n_3),
.B1(n_5),
.B2(n_166),
.Y(n_291)
);

AOI22xp33_ASAP7_75t_SL g346 ( 
.A1(n_291),
.A2(n_294),
.B1(n_145),
.B2(n_289),
.Y(n_346)
);

HB1xp67_ASAP7_75t_L g293 ( 
.A(n_135),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_203),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_206),
.A2(n_3),
.B1(n_196),
.B2(n_207),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_196),
.B(n_3),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_297),
.B(n_137),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_308),
.A2(n_316),
.B1(n_337),
.B2(n_258),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_312),
.B(n_315),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_224),
.A2(n_204),
.B1(n_206),
.B2(n_207),
.Y(n_316)
);

OR2x2_ASAP7_75t_L g378 ( 
.A(n_319),
.B(n_271),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_L g400 ( 
.A1(n_320),
.A2(n_323),
.B1(n_254),
.B2(n_269),
.Y(n_400)
);

AOI22xp33_ASAP7_75t_L g323 ( 
.A1(n_292),
.A2(n_200),
.B1(n_179),
.B2(n_192),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_263),
.B(n_200),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_326),
.B(n_348),
.Y(n_384)
);

AOI21xp5_ASAP7_75t_L g401 ( 
.A1(n_330),
.A2(n_341),
.B(n_322),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_295),
.B(n_205),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_SL g377 ( 
.A(n_331),
.B(n_339),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_226),
.B(n_138),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_332),
.B(n_340),
.C(n_342),
.Y(n_365)
);

AO22x1_ASAP7_75t_SL g335 ( 
.A1(n_235),
.A2(n_153),
.B1(n_191),
.B2(n_177),
.Y(n_335)
);

OA21x2_ASAP7_75t_L g363 ( 
.A1(n_335),
.A2(n_349),
.B(n_274),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_L g337 ( 
.A1(n_276),
.A2(n_177),
.B1(n_201),
.B2(n_155),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_260),
.B(n_201),
.Y(n_339)
);

MAJx2_ASAP7_75t_L g340 ( 
.A(n_221),
.B(n_138),
.C(n_178),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_232),
.B(n_187),
.C(n_145),
.Y(n_342)
);

INVxp67_ASAP7_75t_L g358 ( 
.A(n_346),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_245),
.B(n_256),
.Y(n_348)
);

OA22x2_ASAP7_75t_SL g349 ( 
.A1(n_237),
.A2(n_268),
.B1(n_287),
.B2(n_274),
.Y(n_349)
);

INVx1_ASAP7_75t_SL g366 ( 
.A(n_350),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_317),
.B(n_285),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_SL g406 ( 
.A(n_357),
.B(n_362),
.Y(n_406)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_355),
.Y(n_359)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_359),
.Y(n_405)
);

AOI22xp33_ASAP7_75t_SL g360 ( 
.A1(n_337),
.A2(n_286),
.B1(n_281),
.B2(n_273),
.Y(n_360)
);

INVx1_ASAP7_75t_SL g430 ( 
.A(n_360),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_318),
.A2(n_297),
.B1(n_272),
.B2(n_266),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_361),
.A2(n_363),
.B1(n_367),
.B2(n_374),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_324),
.B(n_314),
.Y(n_362)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_304),
.Y(n_364)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_364),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_318),
.A2(n_296),
.B1(n_270),
.B2(n_244),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_328),
.Y(n_368)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_368),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_327),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_369),
.B(n_370),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_327),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_304),
.Y(n_371)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_371),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_326),
.B(n_253),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_372),
.B(n_376),
.Y(n_413)
);

OAI21xp5_ASAP7_75t_L g373 ( 
.A1(n_330),
.A2(n_251),
.B(n_270),
.Y(n_373)
);

OAI21xp5_ASAP7_75t_L g403 ( 
.A1(n_373),
.A2(n_378),
.B(n_382),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_322),
.A2(n_253),
.B1(n_294),
.B2(n_284),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_302),
.Y(n_375)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_375),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_327),
.Y(n_376)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_302),
.Y(n_379)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_379),
.Y(n_431)
);

INVxp67_ASAP7_75t_L g380 ( 
.A(n_313),
.Y(n_380)
);

INVxp67_ASAP7_75t_L g420 ( 
.A(n_380),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_351),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_381),
.Y(n_407)
);

OR2x2_ASAP7_75t_L g382 ( 
.A(n_319),
.B(n_241),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_311),
.Y(n_383)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_383),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_L g434 ( 
.A1(n_385),
.A2(n_400),
.B1(n_316),
.B2(n_308),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_309),
.B(n_228),
.Y(n_387)
);

INVxp67_ASAP7_75t_L g421 ( 
.A(n_387),
.Y(n_421)
);

AOI22xp33_ASAP7_75t_SL g388 ( 
.A1(n_341),
.A2(n_225),
.B1(n_261),
.B2(n_220),
.Y(n_388)
);

INVxp67_ASAP7_75t_L g436 ( 
.A(n_388),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_332),
.B(n_233),
.C(n_222),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_389),
.B(n_390),
.C(n_399),
.Y(n_426)
);

XOR2xp5_ASAP7_75t_L g390 ( 
.A(n_306),
.B(n_243),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_328),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_391),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_L g392 ( 
.A1(n_322),
.A2(n_283),
.B1(n_257),
.B2(n_252),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_SL g409 ( 
.A1(n_392),
.A2(n_320),
.B1(n_352),
.B2(n_309),
.Y(n_409)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_311),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_SL g404 ( 
.A(n_393),
.B(n_394),
.Y(n_404)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_329),
.Y(n_394)
);

CKINVDCx14_ASAP7_75t_R g395 ( 
.A(n_313),
.Y(n_395)
);

CKINVDCx16_ASAP7_75t_R g412 ( 
.A(n_395),
.Y(n_412)
);

INVxp67_ASAP7_75t_L g396 ( 
.A(n_343),
.Y(n_396)
);

CKINVDCx16_ASAP7_75t_R g414 ( 
.A(n_396),
.Y(n_414)
);

INVx4_ASAP7_75t_L g397 ( 
.A(n_345),
.Y(n_397)
);

CKINVDCx16_ASAP7_75t_R g429 ( 
.A(n_397),
.Y(n_429)
);

INVxp67_ASAP7_75t_L g398 ( 
.A(n_300),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_L g411 ( 
.A(n_398),
.B(n_342),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_306),
.B(n_267),
.C(n_230),
.Y(n_399)
);

AOI21xp5_ASAP7_75t_L g427 ( 
.A1(n_401),
.A2(n_312),
.B(n_325),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_340),
.B(n_239),
.C(n_279),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_402),
.B(n_353),
.C(n_335),
.Y(n_428)
);

AND2x2_ASAP7_75t_L g463 ( 
.A(n_409),
.B(n_382),
.Y(n_463)
);

INVx1_ASAP7_75t_SL g447 ( 
.A(n_411),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_SL g415 ( 
.A1(n_385),
.A2(n_349),
.B1(n_307),
.B2(n_335),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_415),
.A2(n_422),
.B1(n_434),
.B2(n_438),
.Y(n_441)
);

XOR2xp5_ASAP7_75t_L g416 ( 
.A(n_365),
.B(n_339),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_416),
.B(n_418),
.C(n_365),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_L g418 ( 
.A(n_386),
.B(n_305),
.Y(n_418)
);

OAI32xp33_ASAP7_75t_L g419 ( 
.A1(n_384),
.A2(n_349),
.A3(n_315),
.B1(n_348),
.B2(n_305),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_419),
.B(n_433),
.Y(n_474)
);

OAI22xp5_ASAP7_75t_SL g422 ( 
.A1(n_401),
.A2(n_384),
.B1(n_373),
.B2(n_349),
.Y(n_422)
);

OAI21xp5_ASAP7_75t_SL g449 ( 
.A1(n_427),
.A2(n_381),
.B(n_362),
.Y(n_449)
);

XOR2xp5_ASAP7_75t_L g459 ( 
.A(n_428),
.B(n_402),
.Y(n_459)
);

OAI32xp33_ASAP7_75t_L g433 ( 
.A1(n_377),
.A2(n_335),
.A3(n_331),
.B1(n_353),
.B2(n_329),
.Y(n_433)
);

AOI21xp5_ASAP7_75t_L g435 ( 
.A1(n_378),
.A2(n_298),
.B(n_347),
.Y(n_435)
);

AOI21xp5_ASAP7_75t_L g443 ( 
.A1(n_435),
.A2(n_378),
.B(n_382),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_363),
.A2(n_310),
.B1(n_352),
.B2(n_344),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_363),
.A2(n_277),
.B1(n_242),
.B2(n_344),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_L g461 ( 
.A1(n_439),
.A2(n_440),
.B1(n_374),
.B2(n_392),
.Y(n_461)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_363),
.A2(n_336),
.B1(n_301),
.B2(n_354),
.Y(n_440)
);

OAI32xp33_ASAP7_75t_L g442 ( 
.A1(n_413),
.A2(n_377),
.A3(n_372),
.B1(n_365),
.B2(n_359),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_442),
.B(n_458),
.Y(n_493)
);

AOI21xp5_ASAP7_75t_L g484 ( 
.A1(n_443),
.A2(n_456),
.B(n_468),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_444),
.B(n_445),
.C(n_448),
.Y(n_490)
);

XNOR2xp5_ASAP7_75t_L g445 ( 
.A(n_416),
.B(n_386),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_404),
.Y(n_446)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_446),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_426),
.B(n_390),
.C(n_389),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_SL g509 ( 
.A(n_449),
.B(n_451),
.Y(n_509)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_404),
.Y(n_450)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_450),
.Y(n_488)
);

CKINVDCx20_ASAP7_75t_R g451 ( 
.A(n_437),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_437),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_452),
.B(n_464),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_426),
.B(n_390),
.C(n_389),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_453),
.B(n_459),
.C(n_462),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_SL g454 ( 
.A(n_406),
.B(n_357),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_SL g501 ( 
.A(n_454),
.B(n_460),
.Y(n_501)
);

AOI22x1_ASAP7_75t_L g455 ( 
.A1(n_422),
.A2(n_367),
.B1(n_400),
.B2(n_358),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_L g478 ( 
.A1(n_455),
.A2(n_461),
.B1(n_466),
.B2(n_473),
.Y(n_478)
);

AOI21xp5_ASAP7_75t_L g456 ( 
.A1(n_403),
.A2(n_388),
.B(n_366),
.Y(n_456)
);

INVx4_ASAP7_75t_L g457 ( 
.A(n_408),
.Y(n_457)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_457),
.Y(n_479)
);

INVxp33_ASAP7_75t_SL g458 ( 
.A(n_406),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_407),
.B(n_395),
.Y(n_460)
);

XNOR2xp5_ASAP7_75t_L g462 ( 
.A(n_418),
.B(n_399),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_463),
.B(n_432),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_407),
.B(n_387),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_414),
.B(n_399),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_465),
.B(n_469),
.Y(n_492)
);

AOI22xp5_ASAP7_75t_L g466 ( 
.A1(n_415),
.A2(n_439),
.B1(n_425),
.B2(n_428),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_417),
.Y(n_467)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_467),
.Y(n_491)
);

AOI21x1_ASAP7_75t_L g468 ( 
.A1(n_403),
.A2(n_402),
.B(n_360),
.Y(n_468)
);

OAI21xp5_ASAP7_75t_L g469 ( 
.A1(n_435),
.A2(n_427),
.B(n_413),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_405),
.B(n_364),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_470),
.B(n_376),
.Y(n_504)
);

XNOR2xp5_ASAP7_75t_L g471 ( 
.A(n_411),
.B(n_361),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_471),
.B(n_475),
.C(n_375),
.Y(n_506)
);

BUFx6f_ASAP7_75t_L g472 ( 
.A(n_405),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g499 ( 
.A(n_472),
.Y(n_499)
);

AOI22xp5_ASAP7_75t_L g473 ( 
.A1(n_425),
.A2(n_438),
.B1(n_434),
.B2(n_409),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_L g475 ( 
.A(n_419),
.B(n_420),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_L g476 ( 
.A1(n_473),
.A2(n_440),
.B1(n_436),
.B2(n_430),
.Y(n_476)
);

OAI22xp5_ASAP7_75t_L g512 ( 
.A1(n_476),
.A2(n_480),
.B1(n_482),
.B2(n_485),
.Y(n_512)
);

XNOR2xp5_ASAP7_75t_SL g477 ( 
.A(n_445),
.B(n_433),
.Y(n_477)
);

XNOR2xp5_ASAP7_75t_SL g522 ( 
.A(n_477),
.B(n_394),
.Y(n_522)
);

OAI22xp5_ASAP7_75t_L g480 ( 
.A1(n_441),
.A2(n_421),
.B1(n_414),
.B2(n_412),
.Y(n_480)
);

AOI22xp5_ASAP7_75t_L g482 ( 
.A1(n_441),
.A2(n_430),
.B1(n_412),
.B2(n_366),
.Y(n_482)
);

AOI22xp5_ASAP7_75t_L g485 ( 
.A1(n_466),
.A2(n_430),
.B1(n_366),
.B2(n_410),
.Y(n_485)
);

AOI22xp5_ASAP7_75t_L g486 ( 
.A1(n_468),
.A2(n_410),
.B1(n_417),
.B2(n_423),
.Y(n_486)
);

AOI22xp5_ASAP7_75t_L g510 ( 
.A1(n_486),
.A2(n_489),
.B1(n_497),
.B2(n_443),
.Y(n_510)
);

OAI22xp5_ASAP7_75t_L g487 ( 
.A1(n_455),
.A2(n_423),
.B1(n_431),
.B2(n_424),
.Y(n_487)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_487),
.Y(n_514)
);

OAI22xp5_ASAP7_75t_SL g489 ( 
.A1(n_474),
.A2(n_432),
.B1(n_431),
.B2(n_424),
.Y(n_489)
);

OAI21xp5_ASAP7_75t_L g531 ( 
.A1(n_494),
.A2(n_391),
.B(n_321),
.Y(n_531)
);

XNOR2xp5_ASAP7_75t_L g496 ( 
.A(n_444),
.B(n_371),
.Y(n_496)
);

XOR2xp5_ASAP7_75t_L g532 ( 
.A(n_496),
.B(n_498),
.Y(n_532)
);

AOI22xp5_ASAP7_75t_L g497 ( 
.A1(n_463),
.A2(n_429),
.B1(n_408),
.B2(n_397),
.Y(n_497)
);

XNOR2xp5_ASAP7_75t_L g498 ( 
.A(n_459),
.B(n_471),
.Y(n_498)
);

XNOR2xp5_ASAP7_75t_L g500 ( 
.A(n_462),
.B(n_379),
.Y(n_500)
);

XNOR2xp5_ASAP7_75t_L g515 ( 
.A(n_500),
.B(n_506),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_474),
.B(n_429),
.Y(n_502)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_502),
.Y(n_516)
);

CKINVDCx16_ASAP7_75t_R g503 ( 
.A(n_472),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_503),
.B(n_449),
.Y(n_511)
);

CKINVDCx14_ASAP7_75t_R g525 ( 
.A(n_504),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_475),
.B(n_463),
.Y(n_505)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_505),
.Y(n_528)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_457),
.Y(n_507)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_507),
.Y(n_529)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_461),
.Y(n_508)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_508),
.Y(n_533)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_510),
.Y(n_546)
);

CKINVDCx16_ASAP7_75t_R g550 ( 
.A(n_511),
.Y(n_550)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_495),
.B(n_453),
.C(n_448),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g553 ( 
.A(n_513),
.B(n_524),
.C(n_534),
.Y(n_553)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_501),
.B(n_447),
.Y(n_517)
);

CKINVDCx16_ASAP7_75t_R g556 ( 
.A(n_517),
.Y(n_556)
);

XNOR2xp5_ASAP7_75t_L g518 ( 
.A(n_490),
.B(n_447),
.Y(n_518)
);

XNOR2xp5_ASAP7_75t_L g540 ( 
.A(n_518),
.B(n_522),
.Y(n_540)
);

AOI22xp5_ASAP7_75t_L g519 ( 
.A1(n_508),
.A2(n_456),
.B1(n_469),
.B2(n_455),
.Y(n_519)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_519),
.Y(n_549)
);

AOI22xp5_ASAP7_75t_SL g520 ( 
.A1(n_478),
.A2(n_442),
.B1(n_397),
.B2(n_369),
.Y(n_520)
);

OAI21xp5_ASAP7_75t_SL g548 ( 
.A1(n_520),
.A2(n_521),
.B(n_530),
.Y(n_548)
);

AOI21xp5_ASAP7_75t_L g521 ( 
.A1(n_484),
.A2(n_370),
.B(n_333),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_SL g523 ( 
.A(n_501),
.B(n_393),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_SL g544 ( 
.A(n_523),
.B(n_526),
.Y(n_544)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_495),
.B(n_333),
.C(n_383),
.Y(n_524)
);

CKINVDCx16_ASAP7_75t_R g526 ( 
.A(n_509),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_SL g527 ( 
.A(n_481),
.B(n_354),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_SL g560 ( 
.A(n_527),
.B(n_491),
.Y(n_560)
);

AOI21xp5_ASAP7_75t_L g530 ( 
.A1(n_484),
.A2(n_336),
.B(n_368),
.Y(n_530)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_531),
.Y(n_557)
);

MAJIxp5_ASAP7_75t_L g534 ( 
.A(n_490),
.B(n_301),
.C(n_356),
.Y(n_534)
);

AND2x2_ASAP7_75t_L g535 ( 
.A(n_476),
.B(n_345),
.Y(n_535)
);

INVx1_ASAP7_75t_SL g551 ( 
.A(n_535),
.Y(n_551)
);

AOI22xp5_ASAP7_75t_SL g536 ( 
.A1(n_492),
.A2(n_229),
.B1(n_299),
.B2(n_334),
.Y(n_536)
);

INVxp67_ASAP7_75t_L g542 ( 
.A(n_536),
.Y(n_542)
);

XNOR2xp5_ASAP7_75t_L g537 ( 
.A(n_496),
.B(n_299),
.Y(n_537)
);

XNOR2xp5_ASAP7_75t_L g559 ( 
.A(n_537),
.B(n_505),
.Y(n_559)
);

INVxp67_ASAP7_75t_L g538 ( 
.A(n_486),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_538),
.B(n_497),
.Y(n_547)
);

AOI21xp5_ASAP7_75t_L g539 ( 
.A1(n_493),
.A2(n_338),
.B(n_334),
.Y(n_539)
);

OAI21xp5_ASAP7_75t_L g555 ( 
.A1(n_539),
.A2(n_494),
.B(n_482),
.Y(n_555)
);

XOR2x2_ASAP7_75t_L g541 ( 
.A(n_519),
.B(n_493),
.Y(n_541)
);

INVx1_ASAP7_75t_SL g580 ( 
.A(n_541),
.Y(n_580)
);

XOR2xp5_ASAP7_75t_L g543 ( 
.A(n_532),
.B(n_498),
.Y(n_543)
);

XOR2xp5_ASAP7_75t_L g564 ( 
.A(n_543),
.B(n_545),
.Y(n_564)
);

XOR2xp5_ASAP7_75t_L g545 ( 
.A(n_532),
.B(n_506),
.Y(n_545)
);

NAND2xp33_ASAP7_75t_SL g582 ( 
.A(n_547),
.B(n_555),
.Y(n_582)
);

AOI22xp33_ASAP7_75t_SL g552 ( 
.A1(n_535),
.A2(n_488),
.B1(n_483),
.B2(n_499),
.Y(n_552)
);

OAI22xp5_ASAP7_75t_SL g573 ( 
.A1(n_552),
.A2(n_485),
.B1(n_539),
.B2(n_510),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_525),
.B(n_489),
.Y(n_554)
);

CKINVDCx20_ASAP7_75t_R g571 ( 
.A(n_554),
.Y(n_571)
);

MAJIxp5_ASAP7_75t_L g558 ( 
.A(n_513),
.B(n_500),
.C(n_477),
.Y(n_558)
);

MAJIxp5_ASAP7_75t_L g565 ( 
.A(n_558),
.B(n_534),
.C(n_524),
.Y(n_565)
);

XOR2xp5_ASAP7_75t_L g569 ( 
.A(n_559),
.B(n_562),
.Y(n_569)
);

AOI22xp5_ASAP7_75t_L g566 ( 
.A1(n_560),
.A2(n_561),
.B1(n_563),
.B2(n_483),
.Y(n_566)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_529),
.Y(n_561)
);

XOR2xp5_ASAP7_75t_L g562 ( 
.A(n_515),
.B(n_518),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_529),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_SL g598 ( 
.A(n_565),
.B(n_570),
.Y(n_598)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_566),
.Y(n_584)
);

AOI22xp5_ASAP7_75t_L g567 ( 
.A1(n_546),
.A2(n_512),
.B1(n_514),
.B2(n_535),
.Y(n_567)
);

OAI22xp5_ASAP7_75t_SL g591 ( 
.A1(n_567),
.A2(n_575),
.B1(n_551),
.B2(n_549),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_L g568 ( 
.A(n_556),
.B(n_488),
.Y(n_568)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_568),
.Y(n_587)
);

MAJIxp5_ASAP7_75t_L g570 ( 
.A(n_553),
.B(n_515),
.C(n_538),
.Y(n_570)
);

MAJIxp5_ASAP7_75t_L g572 ( 
.A(n_553),
.B(n_537),
.C(n_520),
.Y(n_572)
);

MAJIxp5_ASAP7_75t_L g589 ( 
.A(n_572),
.B(n_576),
.C(n_570),
.Y(n_589)
);

AOI22xp5_ASAP7_75t_L g590 ( 
.A1(n_573),
.A2(n_542),
.B1(n_551),
.B2(n_549),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_SL g574 ( 
.A(n_544),
.B(n_528),
.Y(n_574)
);

NOR3xp33_ASAP7_75t_L g596 ( 
.A(n_574),
.B(n_563),
.C(n_561),
.Y(n_596)
);

AOI22xp5_ASAP7_75t_L g575 ( 
.A1(n_546),
.A2(n_514),
.B1(n_533),
.B2(n_516),
.Y(n_575)
);

MAJIxp5_ASAP7_75t_L g576 ( 
.A(n_562),
.B(n_528),
.C(n_521),
.Y(n_576)
);

FAx1_ASAP7_75t_SL g577 ( 
.A(n_541),
.B(n_522),
.CI(n_516),
.CON(n_577),
.SN(n_577)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_577),
.B(n_559),
.Y(n_585)
);

XNOR2xp5_ASAP7_75t_L g578 ( 
.A(n_545),
.B(n_502),
.Y(n_578)
);

XOR2xp5_ASAP7_75t_L g588 ( 
.A(n_578),
.B(n_579),
.Y(n_588)
);

XOR2xp5_ASAP7_75t_L g579 ( 
.A(n_543),
.B(n_533),
.Y(n_579)
);

XNOR2xp5_ASAP7_75t_L g581 ( 
.A(n_558),
.B(n_536),
.Y(n_581)
);

XOR2xp5_ASAP7_75t_L g592 ( 
.A(n_581),
.B(n_540),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_L g583 ( 
.A(n_550),
.B(n_491),
.Y(n_583)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_583),
.Y(n_597)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_585),
.Y(n_601)
);

AOI21xp5_ASAP7_75t_L g586 ( 
.A1(n_580),
.A2(n_548),
.B(n_555),
.Y(n_586)
);

AOI21xp5_ASAP7_75t_L g606 ( 
.A1(n_586),
.A2(n_593),
.B(n_576),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_589),
.B(n_595),
.Y(n_612)
);

OAI22xp5_ASAP7_75t_SL g609 ( 
.A1(n_590),
.A2(n_599),
.B1(n_600),
.B2(n_586),
.Y(n_609)
);

AOI22xp5_ASAP7_75t_L g608 ( 
.A1(n_591),
.A2(n_577),
.B1(n_578),
.B2(n_581),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_592),
.B(n_596),
.Y(n_604)
);

OAI21xp5_ASAP7_75t_L g593 ( 
.A1(n_580),
.A2(n_547),
.B(n_554),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_575),
.Y(n_594)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_594),
.Y(n_607)
);

MAJIxp5_ASAP7_75t_L g595 ( 
.A(n_565),
.B(n_579),
.C(n_564),
.Y(n_595)
);

AOI22xp5_ASAP7_75t_L g599 ( 
.A1(n_571),
.A2(n_542),
.B1(n_550),
.B2(n_557),
.Y(n_599)
);

AOI22xp5_ASAP7_75t_L g600 ( 
.A1(n_567),
.A2(n_557),
.B1(n_530),
.B2(n_548),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_L g602 ( 
.A(n_598),
.B(n_582),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_602),
.B(n_603),
.Y(n_617)
);

MAJIxp5_ASAP7_75t_L g603 ( 
.A(n_595),
.B(n_564),
.C(n_569),
.Y(n_603)
);

MAJIxp5_ASAP7_75t_L g605 ( 
.A(n_589),
.B(n_569),
.C(n_572),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_605),
.B(n_608),
.Y(n_623)
);

AOI21xp33_ASAP7_75t_L g618 ( 
.A1(n_606),
.A2(n_599),
.B(n_593),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_L g621 ( 
.A(n_609),
.B(n_610),
.Y(n_621)
);

AOI22xp5_ASAP7_75t_L g610 ( 
.A1(n_584),
.A2(n_577),
.B1(n_499),
.B2(n_531),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_597),
.B(n_507),
.Y(n_611)
);

CKINVDCx20_ASAP7_75t_R g615 ( 
.A(n_611),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_L g613 ( 
.A(n_587),
.B(n_479),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_SL g614 ( 
.A(n_613),
.B(n_611),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_614),
.B(n_616),
.Y(n_625)
);

NOR2xp33_ASAP7_75t_SL g616 ( 
.A(n_612),
.B(n_604),
.Y(n_616)
);

OAI21xp5_ASAP7_75t_L g629 ( 
.A1(n_618),
.A2(n_609),
.B(n_594),
.Y(n_629)
);

NOR2x1_ASAP7_75t_L g619 ( 
.A(n_604),
.B(n_585),
.Y(n_619)
);

AOI21x1_ASAP7_75t_L g626 ( 
.A1(n_619),
.A2(n_620),
.B(n_622),
.Y(n_626)
);

AOI21xp5_ASAP7_75t_L g620 ( 
.A1(n_606),
.A2(n_605),
.B(n_603),
.Y(n_620)
);

AOI21xp5_ASAP7_75t_L g622 ( 
.A1(n_608),
.A2(n_588),
.B(n_592),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g624 ( 
.A(n_617),
.B(n_601),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_624),
.B(n_627),
.Y(n_634)
);

INVxp67_ASAP7_75t_L g627 ( 
.A(n_623),
.Y(n_627)
);

OAI21xp5_ASAP7_75t_SL g628 ( 
.A1(n_619),
.A2(n_607),
.B(n_610),
.Y(n_628)
);

NAND3xp33_ASAP7_75t_SL g631 ( 
.A(n_628),
.B(n_629),
.C(n_630),
.Y(n_631)
);

O2A1O1Ixp33_ASAP7_75t_SL g630 ( 
.A1(n_621),
.A2(n_591),
.B(n_600),
.C(n_590),
.Y(n_630)
);

MAJIxp5_ASAP7_75t_L g632 ( 
.A(n_626),
.B(n_615),
.C(n_588),
.Y(n_632)
);

OAI21xp5_ASAP7_75t_L g636 ( 
.A1(n_632),
.A2(n_633),
.B(n_631),
.Y(n_636)
);

OAI21xp5_ASAP7_75t_SL g633 ( 
.A1(n_625),
.A2(n_618),
.B(n_479),
.Y(n_633)
);

OAI21x1_ASAP7_75t_L g635 ( 
.A1(n_634),
.A2(n_540),
.B(n_321),
.Y(n_635)
);

MAJIxp5_ASAP7_75t_L g637 ( 
.A(n_635),
.B(n_636),
.C(n_338),
.Y(n_637)
);

AOI21xp33_ASAP7_75t_SL g638 ( 
.A1(n_637),
.A2(n_303),
.B(n_236),
.Y(n_638)
);

MAJIxp5_ASAP7_75t_L g639 ( 
.A(n_638),
.B(n_347),
.C(n_303),
.Y(n_639)
);

AOI21xp5_ASAP7_75t_L g640 ( 
.A1(n_639),
.A2(n_303),
.B(n_265),
.Y(n_640)
);


endmodule