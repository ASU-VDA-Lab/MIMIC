module fake_jpeg_29530_n_539 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_539);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_539;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

HB1xp67_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_11),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

HB1xp67_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

CKINVDCx16_ASAP7_75t_R g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_14),
.B(n_13),
.Y(n_30)
);

INVx11_ASAP7_75t_SL g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_11),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_7),
.B(n_3),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

BUFx16f_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_9),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_8),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_8),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_9),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_8),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_3),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_1),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_13),
.Y(n_50)
);

CKINVDCx16_ASAP7_75t_R g51 ( 
.A(n_6),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_10),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_7),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_54),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_29),
.Y(n_55)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_55),
.Y(n_112)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_26),
.Y(n_56)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_56),
.Y(n_108)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_26),
.Y(n_57)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_57),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_30),
.B(n_16),
.C(n_15),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_58),
.B(n_61),
.Y(n_107)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_29),
.Y(n_59)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_59),
.Y(n_118)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_29),
.Y(n_60)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_60),
.Y(n_145)
);

INVx6_ASAP7_75t_SL g61 ( 
.A(n_42),
.Y(n_61)
);

INVx3_ASAP7_75t_SL g62 ( 
.A(n_49),
.Y(n_62)
);

INVx2_ASAP7_75t_SL g158 ( 
.A(n_62),
.Y(n_158)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_49),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_63),
.Y(n_124)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_64),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_30),
.B(n_16),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_65),
.B(n_67),
.Y(n_114)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_66),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_38),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_31),
.Y(n_68)
);

BUFx5_ASAP7_75t_L g128 ( 
.A(n_68),
.Y(n_128)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_69),
.Y(n_115)
);

INVx4_ASAP7_75t_SL g70 ( 
.A(n_26),
.Y(n_70)
);

INVx4_ASAP7_75t_SL g110 ( 
.A(n_70),
.Y(n_110)
);

INVxp67_ASAP7_75t_SL g71 ( 
.A(n_31),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_71),
.B(n_82),
.Y(n_159)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_38),
.Y(n_72)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_72),
.Y(n_153)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_73),
.Y(n_125)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_36),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_74),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_36),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_75),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_36),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_76),
.Y(n_150)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_42),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_77),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_37),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_78),
.Y(n_166)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_37),
.Y(n_79)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_79),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_37),
.Y(n_80)
);

INVx6_ASAP7_75t_L g147 ( 
.A(n_80),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_37),
.Y(n_81)
);

INVx6_ASAP7_75t_L g160 ( 
.A(n_81),
.Y(n_160)
);

INVx1_ASAP7_75t_SL g82 ( 
.A(n_42),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_52),
.Y(n_83)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_83),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_19),
.Y(n_84)
);

INVx6_ASAP7_75t_L g164 ( 
.A(n_84),
.Y(n_164)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_38),
.Y(n_85)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_85),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_19),
.Y(n_86)
);

INVx5_ASAP7_75t_L g144 ( 
.A(n_86),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_40),
.B(n_16),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_87),
.B(n_95),
.Y(n_152)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_52),
.Y(n_88)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_88),
.Y(n_143)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_19),
.Y(n_89)
);

INVx5_ASAP7_75t_L g149 ( 
.A(n_89),
.Y(n_149)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_52),
.Y(n_90)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_90),
.Y(n_146)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_22),
.Y(n_91)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_91),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_40),
.B(n_15),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_92),
.B(n_105),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_25),
.Y(n_93)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_93),
.Y(n_111)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_22),
.Y(n_94)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_94),
.Y(n_121)
);

INVx2_ASAP7_75t_SL g95 ( 
.A(n_42),
.Y(n_95)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_48),
.Y(n_96)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_96),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_25),
.Y(n_97)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_97),
.Y(n_131)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_48),
.Y(n_98)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_98),
.Y(n_165)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_45),
.Y(n_99)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_99),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_25),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g139 ( 
.A(n_100),
.Y(n_139)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_25),
.Y(n_101)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_101),
.Y(n_122)
);

BUFx5_ASAP7_75t_L g102 ( 
.A(n_42),
.Y(n_102)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_102),
.Y(n_123)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_32),
.Y(n_103)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_103),
.Y(n_132)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_45),
.Y(n_104)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_104),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_18),
.B(n_15),
.Y(n_105)
);

AOI21xp33_ASAP7_75t_L g106 ( 
.A1(n_70),
.A2(n_39),
.B(n_50),
.Y(n_106)
);

AOI21xp33_ASAP7_75t_L g202 ( 
.A1(n_106),
.A2(n_137),
.B(n_28),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_62),
.A2(n_17),
.B1(n_20),
.B2(n_35),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_109),
.A2(n_127),
.B1(n_140),
.B2(n_161),
.Y(n_171)
);

OAI22xp33_ASAP7_75t_L g117 ( 
.A1(n_74),
.A2(n_45),
.B1(n_35),
.B2(n_32),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_117),
.A2(n_120),
.B1(n_134),
.B2(n_51),
.Y(n_186)
);

OAI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_84),
.A2(n_20),
.B1(n_17),
.B2(n_35),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_103),
.A2(n_55),
.B1(n_82),
.B2(n_89),
.Y(n_127)
);

AO22x1_ASAP7_75t_L g134 ( 
.A1(n_95),
.A2(n_51),
.B1(n_28),
.B2(n_21),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_68),
.B(n_18),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_136),
.B(n_141),
.Y(n_168)
);

A2O1A1Ixp33_ASAP7_75t_L g137 ( 
.A1(n_94),
.A2(n_41),
.B(n_50),
.C(n_34),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_86),
.A2(n_33),
.B1(n_43),
.B2(n_32),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_56),
.Y(n_141)
);

BUFx4f_ASAP7_75t_L g151 ( 
.A(n_79),
.Y(n_151)
);

INVx2_ASAP7_75t_SL g211 ( 
.A(n_151),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_57),
.B(n_43),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_157),
.B(n_163),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_59),
.A2(n_35),
.B1(n_32),
.B2(n_41),
.Y(n_161)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_77),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_139),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_167),
.B(n_170),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_114),
.B(n_33),
.Y(n_170)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_154),
.Y(n_172)
);

INVx4_ASAP7_75t_SL g260 ( 
.A(n_172),
.Y(n_260)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_155),
.Y(n_173)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_173),
.Y(n_255)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_126),
.Y(n_174)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_174),
.Y(n_258)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_142),
.Y(n_175)
);

BUFx2_ASAP7_75t_L g230 ( 
.A(n_175),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_119),
.Y(n_176)
);

INVx11_ASAP7_75t_L g250 ( 
.A(n_176),
.Y(n_250)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_143),
.Y(n_177)
);

INVx4_ASAP7_75t_L g245 ( 
.A(n_177),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_134),
.A2(n_85),
.B1(n_72),
.B2(n_34),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g232 ( 
.A1(n_178),
.A2(n_200),
.B1(n_215),
.B2(n_216),
.Y(n_232)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_146),
.Y(n_179)
);

INVx4_ASAP7_75t_L g252 ( 
.A(n_179),
.Y(n_252)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_153),
.Y(n_180)
);

HB1xp67_ASAP7_75t_L g261 ( 
.A(n_180),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_139),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_181),
.B(n_188),
.Y(n_238)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_148),
.Y(n_182)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_182),
.Y(n_221)
);

INVx6_ASAP7_75t_L g183 ( 
.A(n_119),
.Y(n_183)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_183),
.Y(n_225)
);

BUFx3_ASAP7_75t_L g184 ( 
.A(n_128),
.Y(n_184)
);

INVx3_ASAP7_75t_L g226 ( 
.A(n_184),
.Y(n_226)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_156),
.Y(n_185)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_185),
.Y(n_222)
);

OR2x2_ASAP7_75t_L g246 ( 
.A(n_186),
.B(n_198),
.Y(n_246)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_113),
.Y(n_187)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_187),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_159),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_135),
.Y(n_189)
);

INVx3_ASAP7_75t_L g263 ( 
.A(n_189),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_135),
.Y(n_190)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_190),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_151),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_191),
.B(n_192),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_152),
.Y(n_192)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_122),
.Y(n_193)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_193),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_107),
.B(n_21),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_194),
.B(n_201),
.Y(n_243)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_162),
.Y(n_195)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_195),
.Y(n_254)
);

HB1xp67_ASAP7_75t_L g196 ( 
.A(n_129),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_196),
.Y(n_229)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_162),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_197),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_161),
.Y(n_198)
);

OAI22xp33_ASAP7_75t_L g199 ( 
.A1(n_164),
.A2(n_54),
.B1(n_76),
.B2(n_78),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_199),
.A2(n_212),
.B1(n_120),
.B2(n_111),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_110),
.A2(n_158),
.B1(n_165),
.B2(n_130),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_115),
.B(n_24),
.Y(n_201)
);

OAI21xp33_ASAP7_75t_L g240 ( 
.A1(n_202),
.A2(n_204),
.B(n_123),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_116),
.A2(n_81),
.B1(n_80),
.B2(n_75),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_L g247 ( 
.A1(n_203),
.A2(n_205),
.B1(n_214),
.B2(n_133),
.Y(n_247)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_138),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_109),
.A2(n_100),
.B1(n_97),
.B2(n_93),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_127),
.Y(n_206)
);

NOR3xp33_ASAP7_75t_L g233 ( 
.A(n_206),
.B(n_217),
.C(n_23),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_L g207 ( 
.A1(n_164),
.A2(n_101),
.B1(n_39),
.B2(n_79),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_207),
.A2(n_160),
.B1(n_147),
.B2(n_131),
.Y(n_224)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_121),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_208),
.Y(n_228)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_121),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_209),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_130),
.B(n_24),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_210),
.B(n_213),
.Y(n_249)
);

OAI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_144),
.A2(n_73),
.B1(n_63),
.B2(n_53),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_165),
.B(n_23),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_147),
.A2(n_160),
.B1(n_166),
.B2(n_150),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_110),
.A2(n_68),
.B1(n_53),
.B2(n_47),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_158),
.A2(n_47),
.B1(n_44),
.B2(n_27),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_108),
.B(n_44),
.C(n_27),
.Y(n_217)
);

BUFx3_ASAP7_75t_L g218 ( 
.A(n_112),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_SL g237 ( 
.A1(n_218),
.A2(n_219),
.B1(n_220),
.B2(n_166),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_150),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_111),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_223),
.A2(n_224),
.B1(n_242),
.B2(n_256),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_233),
.B(n_213),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_192),
.B(n_145),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g298 ( 
.A(n_236),
.B(n_251),
.Y(n_298)
);

INVxp67_ASAP7_75t_SL g267 ( 
.A(n_237),
.Y(n_267)
);

CKINVDCx16_ASAP7_75t_R g266 ( 
.A(n_240),
.Y(n_266)
);

A2O1A1Ixp33_ASAP7_75t_L g241 ( 
.A1(n_194),
.A2(n_132),
.B(n_117),
.C(n_14),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_241),
.B(n_12),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_198),
.A2(n_133),
.B1(n_131),
.B2(n_149),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_206),
.A2(n_188),
.B1(n_171),
.B2(n_118),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_244),
.A2(n_253),
.B1(n_259),
.B2(n_211),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_247),
.A2(n_219),
.B1(n_176),
.B2(n_189),
.Y(n_290)
);

AO22x1_ASAP7_75t_SL g248 ( 
.A1(n_186),
.A2(n_125),
.B1(n_124),
.B2(n_71),
.Y(n_248)
);

OA22x2_ASAP7_75t_SL g273 ( 
.A1(n_248),
.A2(n_179),
.B1(n_175),
.B2(n_177),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_168),
.B(n_15),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_SL g253 ( 
.A1(n_187),
.A2(n_125),
.B1(n_124),
.B2(n_14),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_201),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_256)
);

OAI21xp33_ASAP7_75t_L g259 ( 
.A1(n_210),
.A2(n_13),
.B(n_12),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_264),
.B(n_275),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_257),
.B(n_169),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_265),
.B(n_268),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_249),
.B(n_217),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_249),
.B(n_173),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_269),
.B(n_274),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_246),
.A2(n_182),
.B1(n_183),
.B2(n_199),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_270),
.A2(n_292),
.B1(n_224),
.B2(n_260),
.Y(n_303)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_260),
.Y(n_272)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_272),
.Y(n_302)
);

OAI21xp33_ASAP7_75t_SL g321 ( 
.A1(n_273),
.A2(n_252),
.B(n_245),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_257),
.B(n_174),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_230),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_236),
.B(n_204),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_276),
.B(n_277),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_235),
.B(n_193),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_223),
.A2(n_167),
.B1(n_181),
.B2(n_208),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_278),
.A2(n_279),
.B1(n_260),
.B2(n_221),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_246),
.A2(n_209),
.B1(n_220),
.B2(n_185),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_227),
.Y(n_280)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_280),
.Y(n_312)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_227),
.Y(n_281)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_281),
.Y(n_314)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_239),
.Y(n_282)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_282),
.Y(n_320)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_250),
.Y(n_283)
);

BUFx3_ASAP7_75t_L g306 ( 
.A(n_283),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_243),
.B(n_180),
.C(n_218),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_284),
.B(n_294),
.C(n_234),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_285),
.A2(n_261),
.B1(n_226),
.B2(n_234),
.Y(n_315)
);

BUFx3_ASAP7_75t_L g286 ( 
.A(n_226),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_286),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_243),
.B(n_191),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_287),
.B(n_288),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_238),
.B(n_195),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_230),
.Y(n_289)
);

OR2x2_ASAP7_75t_L g318 ( 
.A(n_289),
.B(n_291),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_290),
.A2(n_250),
.B1(n_255),
.B2(n_258),
.Y(n_336)
);

O2A1O1Ixp33_ASAP7_75t_L g291 ( 
.A1(n_246),
.A2(n_211),
.B(n_197),
.C(n_172),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_232),
.A2(n_190),
.B1(n_211),
.B2(n_184),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_239),
.Y(n_293)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_293),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_238),
.B(n_190),
.C(n_1),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_242),
.A2(n_13),
.B(n_12),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g317 ( 
.A1(n_295),
.A2(n_9),
.B(n_231),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_296),
.A2(n_241),
.B(n_251),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_230),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_297),
.Y(n_329)
);

INVx3_ASAP7_75t_L g299 ( 
.A(n_225),
.Y(n_299)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_299),
.Y(n_331)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_221),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_300),
.B(n_228),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_268),
.B(n_235),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_301),
.B(n_316),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_303),
.A2(n_304),
.B1(n_310),
.B2(n_278),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_270),
.A2(n_248),
.B1(n_233),
.B2(n_241),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_305),
.B(n_298),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_308),
.A2(n_276),
.B1(n_273),
.B2(n_292),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_SL g309 ( 
.A1(n_296),
.A2(n_248),
.B(n_229),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_SL g338 ( 
.A1(n_309),
.A2(n_311),
.B(n_317),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_290),
.A2(n_248),
.B1(n_256),
.B2(n_254),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_SL g311 ( 
.A1(n_264),
.A2(n_261),
.B(n_262),
.Y(n_311)
);

INVxp67_ASAP7_75t_L g366 ( 
.A(n_315),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_287),
.B(n_222),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_321),
.A2(n_322),
.B1(n_332),
.B2(n_273),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_271),
.A2(n_231),
.B1(n_254),
.B2(n_225),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_326),
.B(n_284),
.Y(n_345)
);

OAI21xp5_ASAP7_75t_SL g327 ( 
.A1(n_288),
.A2(n_222),
.B(n_252),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_SL g349 ( 
.A1(n_327),
.A2(n_333),
.B(n_335),
.Y(n_349)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_269),
.B(n_228),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_328),
.B(n_258),
.C(n_289),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_L g332 ( 
.A1(n_271),
.A2(n_263),
.B1(n_252),
.B2(n_245),
.Y(n_332)
);

AOI22xp33_ASAP7_75t_SL g333 ( 
.A1(n_267),
.A2(n_286),
.B1(n_285),
.B2(n_299),
.Y(n_333)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_334),
.Y(n_350)
);

AOI22xp33_ASAP7_75t_SL g335 ( 
.A1(n_267),
.A2(n_263),
.B1(n_245),
.B2(n_255),
.Y(n_335)
);

AOI22xp33_ASAP7_75t_L g341 ( 
.A1(n_336),
.A2(n_272),
.B1(n_297),
.B2(n_275),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_337),
.A2(n_347),
.B1(n_353),
.B2(n_354),
.Y(n_400)
);

CKINVDCx16_ASAP7_75t_R g339 ( 
.A(n_334),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_339),
.B(n_368),
.Y(n_376)
);

OA22x2_ASAP7_75t_L g395 ( 
.A1(n_340),
.A2(n_321),
.B1(n_336),
.B2(n_332),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_341),
.A2(n_343),
.B1(n_340),
.B2(n_303),
.Y(n_389)
);

INVxp67_ASAP7_75t_SL g342 ( 
.A(n_308),
.Y(n_342)
);

INVxp67_ASAP7_75t_L g373 ( 
.A(n_342),
.Y(n_373)
);

OAI21xp5_ASAP7_75t_SL g372 ( 
.A1(n_344),
.A2(n_362),
.B(n_369),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_345),
.B(n_370),
.C(n_326),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_306),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_346),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_304),
.A2(n_279),
.B1(n_273),
.B2(n_266),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_325),
.B(n_274),
.Y(n_348)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_348),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_325),
.B(n_277),
.Y(n_352)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_352),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_L g353 ( 
.A1(n_318),
.A2(n_295),
.B1(n_266),
.B2(n_265),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_318),
.A2(n_294),
.B1(n_291),
.B2(n_281),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_306),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_355),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_306),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_356),
.Y(n_394)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_312),
.Y(n_357)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_357),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_313),
.B(n_298),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_358),
.Y(n_396)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_312),
.Y(n_359)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_359),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_323),
.B(n_280),
.Y(n_360)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_360),
.Y(n_387)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_314),
.Y(n_361)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_361),
.Y(n_391)
);

AOI21xp5_ASAP7_75t_SL g362 ( 
.A1(n_318),
.A2(n_291),
.B(n_293),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_314),
.Y(n_363)
);

CKINVDCx16_ASAP7_75t_R g375 ( 
.A(n_363),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_323),
.B(n_282),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_364),
.B(n_365),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g365 ( 
.A(n_319),
.B(n_300),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_367),
.B(n_326),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_313),
.Y(n_368)
);

OAI21xp5_ASAP7_75t_SL g369 ( 
.A1(n_333),
.A2(n_299),
.B(n_286),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_301),
.B(n_283),
.C(n_250),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_378),
.B(n_381),
.C(n_382),
.Y(n_409)
);

OAI21xp5_ASAP7_75t_SL g379 ( 
.A1(n_366),
.A2(n_335),
.B(n_315),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_SL g410 ( 
.A(n_379),
.B(n_388),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_345),
.B(n_328),
.C(n_307),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_370),
.B(n_328),
.C(n_307),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_383),
.B(n_403),
.C(n_367),
.Y(n_421)
);

OAI21xp5_ASAP7_75t_SL g388 ( 
.A1(n_362),
.A2(n_317),
.B(n_311),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_389),
.A2(n_398),
.B1(n_402),
.B2(n_339),
.Y(n_408)
);

OAI21xp5_ASAP7_75t_SL g390 ( 
.A1(n_362),
.A2(n_305),
.B(n_309),
.Y(n_390)
);

CKINVDCx14_ASAP7_75t_R g423 ( 
.A(n_390),
.Y(n_423)
);

INVxp67_ASAP7_75t_L g392 ( 
.A(n_341),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_392),
.B(n_337),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_L g393 ( 
.A1(n_358),
.A2(n_310),
.B1(n_319),
.B2(n_329),
.Y(n_393)
);

INVxp67_ASAP7_75t_L g413 ( 
.A(n_393),
.Y(n_413)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_395),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_368),
.B(n_316),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_397),
.B(n_351),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_343),
.A2(n_322),
.B1(n_329),
.B2(n_327),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_L g399 ( 
.A(n_351),
.B(n_330),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g426 ( 
.A(n_399),
.B(n_351),
.Y(n_426)
);

OAI21x1_ASAP7_75t_L g401 ( 
.A1(n_360),
.A2(n_330),
.B(n_320),
.Y(n_401)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_401),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_SL g402 ( 
.A1(n_340),
.A2(n_320),
.B1(n_302),
.B2(n_324),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_370),
.B(n_302),
.C(n_331),
.Y(n_403)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_405),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_376),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_406),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_L g437 ( 
.A1(n_408),
.A2(n_412),
.B1(n_418),
.B2(n_428),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_SL g411 ( 
.A1(n_400),
.A2(n_350),
.B1(n_344),
.B2(n_365),
.Y(n_411)
);

AOI22xp5_ASAP7_75t_L g439 ( 
.A1(n_411),
.A2(n_430),
.B1(n_373),
.B2(n_402),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_L g412 ( 
.A1(n_389),
.A2(n_354),
.B1(n_353),
.B2(n_347),
.Y(n_412)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_377),
.Y(n_414)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_414),
.Y(n_444)
);

CKINVDCx16_ASAP7_75t_R g415 ( 
.A(n_377),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_415),
.B(n_419),
.Y(n_450)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_384),
.Y(n_416)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_416),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_396),
.B(n_364),
.Y(n_417)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_417),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_SL g418 ( 
.A(n_396),
.B(n_352),
.Y(n_418)
);

AOI32xp33_ASAP7_75t_L g419 ( 
.A1(n_372),
.A2(n_338),
.A3(n_349),
.B1(n_350),
.B2(n_369),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_386),
.B(n_348),
.Y(n_420)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_420),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_421),
.B(n_381),
.C(n_378),
.Y(n_433)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_384),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_422),
.B(n_424),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_386),
.B(n_363),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_L g434 ( 
.A(n_425),
.B(n_427),
.Y(n_434)
);

XOR2xp5_ASAP7_75t_L g440 ( 
.A(n_426),
.B(n_383),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_387),
.B(n_361),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_391),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_391),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_L g448 ( 
.A1(n_429),
.A2(n_431),
.B1(n_394),
.B2(n_380),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_L g430 ( 
.A1(n_400),
.A2(n_349),
.B1(n_342),
.B2(n_367),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_401),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_387),
.B(n_357),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_L g438 ( 
.A(n_432),
.B(n_398),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_433),
.B(n_441),
.C(n_451),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_438),
.B(n_445),
.Y(n_469)
);

OAI22xp5_ASAP7_75t_SL g467 ( 
.A1(n_439),
.A2(n_412),
.B1(n_413),
.B2(n_408),
.Y(n_467)
);

XOR2xp5_ASAP7_75t_L g459 ( 
.A(n_440),
.B(n_443),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_409),
.B(n_403),
.C(n_382),
.Y(n_441)
);

OAI21xp5_ASAP7_75t_L g442 ( 
.A1(n_410),
.A2(n_372),
.B(n_373),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_442),
.B(n_410),
.Y(n_460)
);

XNOR2xp5_ASAP7_75t_SL g443 ( 
.A(n_426),
.B(n_399),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_SL g445 ( 
.A(n_406),
.B(n_374),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_SL g447 ( 
.A(n_411),
.B(n_390),
.Y(n_447)
);

XOR2xp5_ASAP7_75t_L g466 ( 
.A(n_447),
.B(n_419),
.Y(n_466)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_448),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_409),
.B(n_388),
.C(n_338),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_421),
.B(n_374),
.C(n_371),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_453),
.B(n_454),
.C(n_455),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_423),
.B(n_371),
.C(n_395),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_430),
.B(n_395),
.C(n_394),
.Y(n_455)
);

INVx1_ASAP7_75t_SL g458 ( 
.A(n_444),
.Y(n_458)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_458),
.Y(n_477)
);

XOR2xp5_ASAP7_75t_L g484 ( 
.A(n_460),
.B(n_466),
.Y(n_484)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_440),
.B(n_441),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g481 ( 
.A(n_461),
.B(n_474),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_446),
.B(n_418),
.Y(n_462)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_462),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_SL g463 ( 
.A(n_450),
.B(n_417),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_463),
.B(n_464),
.Y(n_478)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_449),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_452),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_465),
.B(n_467),
.Y(n_487)
);

INVx1_ASAP7_75t_SL g470 ( 
.A(n_452),
.Y(n_470)
);

OR2x2_ASAP7_75t_L g490 ( 
.A(n_470),
.B(n_380),
.Y(n_490)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_456),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_471),
.B(n_473),
.Y(n_491)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_456),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_434),
.B(n_385),
.Y(n_474)
);

XOR2xp5_ASAP7_75t_L g475 ( 
.A(n_443),
.B(n_424),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_L g489 ( 
.A(n_475),
.B(n_435),
.Y(n_489)
);

OAI22xp33_ASAP7_75t_SL g476 ( 
.A1(n_457),
.A2(n_404),
.B1(n_436),
.B2(n_407),
.Y(n_476)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_476),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_468),
.B(n_433),
.C(n_453),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_479),
.B(n_480),
.Y(n_500)
);

OAI22xp5_ASAP7_75t_SL g480 ( 
.A1(n_462),
.A2(n_439),
.B1(n_455),
.B2(n_404),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_468),
.B(n_451),
.C(n_454),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_482),
.B(n_483),
.C(n_486),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_472),
.B(n_437),
.C(n_438),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_472),
.B(n_447),
.C(n_442),
.Y(n_486)
);

OAI22x1_ASAP7_75t_L g488 ( 
.A1(n_466),
.A2(n_395),
.B1(n_405),
.B2(n_379),
.Y(n_488)
);

OR2x2_ASAP7_75t_L g499 ( 
.A(n_488),
.B(n_493),
.Y(n_499)
);

XNOR2xp5_ASAP7_75t_L g495 ( 
.A(n_489),
.B(n_475),
.Y(n_495)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_490),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_461),
.B(n_434),
.C(n_432),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_492),
.B(n_474),
.C(n_470),
.Y(n_505)
);

OAI321xp33_ASAP7_75t_L g493 ( 
.A1(n_469),
.A2(n_420),
.A3(n_425),
.B1(n_427),
.B2(n_431),
.C(n_407),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_481),
.B(n_460),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_494),
.B(n_495),
.Y(n_513)
);

XNOR2xp5_ASAP7_75t_L g496 ( 
.A(n_484),
.B(n_459),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g520 ( 
.A(n_496),
.B(n_503),
.C(n_505),
.Y(n_520)
);

AND2x2_ASAP7_75t_L g502 ( 
.A(n_486),
.B(n_467),
.Y(n_502)
);

OR2x2_ASAP7_75t_L g511 ( 
.A(n_502),
.B(n_482),
.Y(n_511)
);

XNOR2xp5_ASAP7_75t_L g503 ( 
.A(n_484),
.B(n_459),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_478),
.B(n_458),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_504),
.B(n_506),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_492),
.B(n_385),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_485),
.B(n_415),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_507),
.B(n_508),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_483),
.B(n_392),
.C(n_428),
.Y(n_508)
);

BUFx4f_ASAP7_75t_SL g509 ( 
.A(n_501),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_509),
.B(n_510),
.Y(n_521)
);

AO22x1_ASAP7_75t_L g510 ( 
.A1(n_497),
.A2(n_488),
.B1(n_490),
.B2(n_476),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_511),
.B(n_512),
.Y(n_522)
);

OAI22xp5_ASAP7_75t_SL g512 ( 
.A1(n_499),
.A2(n_487),
.B1(n_491),
.B2(n_477),
.Y(n_512)
);

AOI321xp33_ASAP7_75t_L g514 ( 
.A1(n_499),
.A2(n_375),
.A3(n_422),
.B1(n_416),
.B2(n_414),
.C(n_429),
.Y(n_514)
);

AOI21xp5_ASAP7_75t_L g524 ( 
.A1(n_514),
.A2(n_517),
.B(n_505),
.Y(n_524)
);

XOR2xp5_ASAP7_75t_L g516 ( 
.A(n_502),
.B(n_359),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_516),
.B(n_519),
.Y(n_523)
);

AOI321xp33_ASAP7_75t_L g517 ( 
.A1(n_498),
.A2(n_356),
.A3(n_355),
.B1(n_346),
.B2(n_324),
.C(n_331),
.Y(n_517)
);

OAI22xp5_ASAP7_75t_L g519 ( 
.A1(n_500),
.A2(n_283),
.B1(n_1),
.B2(n_2),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_524),
.B(n_509),
.Y(n_529)
);

OAI21xp5_ASAP7_75t_L g525 ( 
.A1(n_511),
.A2(n_498),
.B(n_508),
.Y(n_525)
);

OAI21xp5_ASAP7_75t_L g528 ( 
.A1(n_525),
.A2(n_526),
.B(n_527),
.Y(n_528)
);

OAI21xp5_ASAP7_75t_L g526 ( 
.A1(n_513),
.A2(n_0),
.B(n_1),
.Y(n_526)
);

AOI21xp5_ASAP7_75t_L g527 ( 
.A1(n_515),
.A2(n_7),
.B(n_2),
.Y(n_527)
);

AOI21xp5_ASAP7_75t_L g533 ( 
.A1(n_529),
.A2(n_530),
.B(n_531),
.Y(n_533)
);

OAI21xp5_ASAP7_75t_L g530 ( 
.A1(n_522),
.A2(n_509),
.B(n_520),
.Y(n_530)
);

MAJIxp5_ASAP7_75t_L g531 ( 
.A(n_521),
.B(n_518),
.C(n_516),
.Y(n_531)
);

OAI321xp33_ASAP7_75t_L g532 ( 
.A1(n_528),
.A2(n_510),
.A3(n_523),
.B1(n_3),
.B2(n_4),
.C(n_0),
.Y(n_532)
);

OAI21xp5_ASAP7_75t_L g534 ( 
.A1(n_532),
.A2(n_2),
.B(n_3),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_534),
.Y(n_535)
);

MAJIxp5_ASAP7_75t_L g536 ( 
.A(n_535),
.B(n_533),
.C(n_5),
.Y(n_536)
);

MAJIxp5_ASAP7_75t_L g537 ( 
.A(n_536),
.B(n_7),
.C(n_4),
.Y(n_537)
);

OAI22xp5_ASAP7_75t_L g538 ( 
.A1(n_537),
.A2(n_4),
.B1(n_6),
.B2(n_501),
.Y(n_538)
);

AO21x1_ASAP7_75t_L g539 ( 
.A1(n_538),
.A2(n_4),
.B(n_6),
.Y(n_539)
);


endmodule