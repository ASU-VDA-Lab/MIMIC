module fake_netlist_6_1261_n_180 (n_16, n_1, n_9, n_8, n_18, n_10, n_21, n_24, n_6, n_15, n_27, n_3, n_14, n_0, n_4, n_22, n_26, n_13, n_11, n_28, n_17, n_23, n_12, n_20, n_7, n_30, n_2, n_5, n_19, n_29, n_31, n_25, n_180);

input n_16;
input n_1;
input n_9;
input n_8;
input n_18;
input n_10;
input n_21;
input n_24;
input n_6;
input n_15;
input n_27;
input n_3;
input n_14;
input n_0;
input n_4;
input n_22;
input n_26;
input n_13;
input n_11;
input n_28;
input n_17;
input n_23;
input n_12;
input n_20;
input n_7;
input n_30;
input n_2;
input n_5;
input n_19;
input n_29;
input n_31;
input n_25;

output n_180;

wire n_52;
wire n_119;
wire n_146;
wire n_46;
wire n_163;
wire n_91;
wire n_147;
wire n_154;
wire n_88;
wire n_98;
wire n_113;
wire n_39;
wire n_63;
wire n_73;
wire n_148;
wire n_138;
wire n_161;
wire n_68;
wire n_166;
wire n_50;
wire n_158;
wire n_49;
wire n_83;
wire n_101;
wire n_167;
wire n_144;
wire n_174;
wire n_127;
wire n_125;
wire n_153;
wire n_168;
wire n_178;
wire n_77;
wire n_156;
wire n_149;
wire n_152;
wire n_106;
wire n_145;
wire n_92;
wire n_42;
wire n_133;
wire n_96;
wire n_90;
wire n_160;
wire n_131;
wire n_105;
wire n_54;
wire n_132;
wire n_102;
wire n_87;
wire n_32;
wire n_66;
wire n_85;
wire n_130;
wire n_78;
wire n_99;
wire n_84;
wire n_164;
wire n_100;
wire n_129;
wire n_121;
wire n_137;
wire n_142;
wire n_143;
wire n_47;
wire n_62;
wire n_155;
wire n_75;
wire n_109;
wire n_150;
wire n_122;
wire n_45;
wire n_34;
wire n_140;
wire n_70;
wire n_120;
wire n_37;
wire n_67;
wire n_33;
wire n_82;
wire n_38;
wire n_110;
wire n_151;
wire n_61;
wire n_112;
wire n_172;
wire n_81;
wire n_59;
wire n_76;
wire n_36;
wire n_124;
wire n_55;
wire n_126;
wire n_97;
wire n_94;
wire n_108;
wire n_58;
wire n_116;
wire n_64;
wire n_117;
wire n_118;
wire n_175;
wire n_48;
wire n_65;
wire n_40;
wire n_93;
wire n_141;
wire n_80;
wire n_135;
wire n_165;
wire n_139;
wire n_41;
wire n_134;
wire n_177;
wire n_176;
wire n_114;
wire n_86;
wire n_104;
wire n_95;
wire n_179;
wire n_107;
wire n_71;
wire n_74;
wire n_123;
wire n_136;
wire n_72;
wire n_89;
wire n_173;
wire n_103;
wire n_111;
wire n_60;
wire n_159;
wire n_157;
wire n_162;
wire n_170;
wire n_35;
wire n_115;
wire n_69;
wire n_128;
wire n_79;
wire n_43;
wire n_171;
wire n_57;
wire n_169;
wire n_53;
wire n_51;
wire n_44;
wire n_56;

INVx1_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

CKINVDCx5p33_ASAP7_75t_R g33 ( 
.A(n_1),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_0),
.Y(n_35)
);

CKINVDCx5p33_ASAP7_75t_R g36 ( 
.A(n_29),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_26),
.Y(n_37)
);

CKINVDCx5p33_ASAP7_75t_R g38 ( 
.A(n_16),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_23),
.Y(n_39)
);

CKINVDCx5p33_ASAP7_75t_R g40 ( 
.A(n_19),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_28),
.B(n_12),
.Y(n_42)
);

CKINVDCx5p33_ASAP7_75t_R g43 ( 
.A(n_3),
.Y(n_43)
);

CKINVDCx5p33_ASAP7_75t_R g44 ( 
.A(n_27),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_4),
.B(n_3),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_11),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_1),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_7),
.B(n_14),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_2),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_9),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_4),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_52),
.Y(n_53)
);

AND2x6_ASAP7_75t_L g54 ( 
.A(n_34),
.B(n_31),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_32),
.B(n_0),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_51),
.Y(n_57)
);

AND2x4_ASAP7_75t_L g58 ( 
.A(n_47),
.B(n_30),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_41),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_59)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_48),
.B(n_5),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_33),
.B(n_6),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_38),
.B(n_8),
.Y(n_65)
);

OR2x6_ASAP7_75t_L g66 ( 
.A(n_42),
.B(n_49),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_33),
.Y(n_67)
);

OR2x2_ASAP7_75t_L g68 ( 
.A(n_43),
.B(n_8),
.Y(n_68)
);

INVx1_ASAP7_75t_SL g69 ( 
.A(n_35),
.Y(n_69)
);

OR2x6_ASAP7_75t_L g70 ( 
.A(n_43),
.B(n_10),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_38),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_40),
.B(n_10),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_40),
.Y(n_73)
);

AOI21x1_ASAP7_75t_L g74 ( 
.A1(n_58),
.A2(n_44),
.B(n_17),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_L g75 ( 
.A1(n_64),
.A2(n_44),
.B(n_39),
.Y(n_75)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_54),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_60),
.B(n_37),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_71),
.B(n_13),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_60),
.B(n_50),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_63),
.A2(n_18),
.B(n_20),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g81 ( 
.A1(n_66),
.A2(n_64),
.B(n_63),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_53),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_53),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_71),
.B(n_21),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_L g85 ( 
.A1(n_58),
.A2(n_22),
.B(n_25),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_69),
.Y(n_86)
);

HB1xp67_ASAP7_75t_L g87 ( 
.A(n_67),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_73),
.A2(n_66),
.B(n_71),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_71),
.B(n_73),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_66),
.A2(n_68),
.B1(n_59),
.B2(n_70),
.Y(n_90)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_74),
.Y(n_91)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_74),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_89),
.B(n_60),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_82),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_78),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_81),
.B(n_56),
.Y(n_96)
);

OR2x2_ASAP7_75t_L g97 ( 
.A(n_86),
.B(n_71),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_85),
.A2(n_66),
.B1(n_58),
.B2(n_54),
.Y(n_98)
);

O2A1O1Ixp33_ASAP7_75t_L g99 ( 
.A1(n_90),
.A2(n_57),
.B(n_72),
.C(n_61),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_82),
.B(n_56),
.Y(n_100)
);

BUFx2_ASAP7_75t_L g101 ( 
.A(n_75),
.Y(n_101)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_83),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_102),
.Y(n_103)
);

HB1xp67_ASAP7_75t_L g104 ( 
.A(n_97),
.Y(n_104)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_102),
.Y(n_105)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_102),
.Y(n_106)
);

HB1xp67_ASAP7_75t_L g107 ( 
.A(n_97),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_94),
.Y(n_108)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_94),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_100),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_110),
.B(n_96),
.Y(n_111)
);

OA21x2_ASAP7_75t_L g112 ( 
.A1(n_108),
.A2(n_98),
.B(n_85),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_110),
.A2(n_98),
.B1(n_101),
.B2(n_75),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_104),
.B(n_107),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_109),
.B(n_96),
.Y(n_115)
);

NAND3xp33_ASAP7_75t_L g116 ( 
.A(n_106),
.B(n_79),
.C(n_77),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_103),
.B(n_97),
.Y(n_117)
);

OR2x2_ASAP7_75t_L g118 ( 
.A(n_111),
.B(n_101),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_117),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_115),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_114),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_113),
.B(n_96),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_119),
.Y(n_123)
);

INVx2_ASAP7_75t_SL g124 ( 
.A(n_121),
.Y(n_124)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_120),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_122),
.A2(n_76),
.B(n_112),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_118),
.B(n_113),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_L g128 ( 
.A1(n_118),
.A2(n_116),
.B1(n_93),
.B2(n_112),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_119),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_120),
.B(n_112),
.Y(n_130)
);

OR2x2_ASAP7_75t_L g131 ( 
.A(n_118),
.B(n_88),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_119),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_121),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_124),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_125),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_127),
.B(n_125),
.Y(n_136)
);

NOR2x1_ASAP7_75t_L g137 ( 
.A(n_131),
.B(n_132),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_127),
.B(n_58),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_130),
.B(n_70),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_133),
.B(n_87),
.Y(n_140)
);

AND2x4_ASAP7_75t_L g141 ( 
.A(n_123),
.B(n_105),
.Y(n_141)
);

NOR2xp67_ASAP7_75t_L g142 ( 
.A(n_135),
.B(n_131),
.Y(n_142)
);

INVx2_ASAP7_75t_SL g143 ( 
.A(n_135),
.Y(n_143)
);

NAND5xp2_ASAP7_75t_L g144 ( 
.A(n_140),
.B(n_99),
.C(n_65),
.D(n_128),
.E(n_62),
.Y(n_144)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_136),
.Y(n_145)
);

AND3x2_ASAP7_75t_L g146 ( 
.A(n_134),
.B(n_132),
.C(n_123),
.Y(n_146)
);

NAND5xp2_ASAP7_75t_L g147 ( 
.A(n_138),
.B(n_99),
.C(n_62),
.D(n_61),
.E(n_55),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_136),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_137),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_139),
.B(n_130),
.Y(n_150)
);

HB1xp67_ASAP7_75t_L g151 ( 
.A(n_141),
.Y(n_151)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_145),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_143),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_149),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_144),
.A2(n_138),
.B1(n_139),
.B2(n_124),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_149),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_150),
.B(n_129),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_151),
.A2(n_142),
.B1(n_146),
.B2(n_150),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_145),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_155),
.B(n_148),
.Y(n_160)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_154),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_156),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_155),
.A2(n_147),
.B(n_126),
.Y(n_163)
);

XOR2x1_ASAP7_75t_L g164 ( 
.A(n_153),
.B(n_141),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_158),
.A2(n_141),
.B(n_147),
.Y(n_165)
);

OA22x2_ASAP7_75t_L g166 ( 
.A1(n_157),
.A2(n_148),
.B1(n_145),
.B2(n_70),
.Y(n_166)
);

NAND4xp75_ASAP7_75t_L g167 ( 
.A(n_159),
.B(n_55),
.C(n_57),
.D(n_80),
.Y(n_167)
);

AOI211xp5_ASAP7_75t_SL g168 ( 
.A1(n_165),
.A2(n_68),
.B(n_152),
.C(n_84),
.Y(n_168)
);

NAND4xp25_ASAP7_75t_L g169 ( 
.A(n_163),
.B(n_83),
.C(n_100),
.D(n_70),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_162),
.B(n_95),
.Y(n_170)
);

OAI221xp5_ASAP7_75t_L g171 ( 
.A1(n_166),
.A2(n_95),
.B1(n_91),
.B2(n_92),
.C(n_54),
.Y(n_171)
);

NOR3xp33_ASAP7_75t_L g172 ( 
.A(n_167),
.B(n_91),
.C(n_92),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_161),
.Y(n_173)
);

AND3x2_ASAP7_75t_L g174 ( 
.A(n_166),
.B(n_54),
.C(n_91),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_173),
.B(n_164),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_170),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_172),
.B(n_160),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_171),
.A2(n_168),
.B1(n_169),
.B2(n_174),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_178),
.A2(n_54),
.B(n_91),
.Y(n_179)
);

OAI221xp5_ASAP7_75t_R g180 ( 
.A1(n_179),
.A2(n_177),
.B1(n_175),
.B2(n_176),
.C(n_54),
.Y(n_180)
);


endmodule