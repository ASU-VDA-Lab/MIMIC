module fake_jpeg_858_n_71 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_71);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_71;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_10;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_47;
wire n_22;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_62;
wire n_25;
wire n_31;
wire n_17;
wire n_56;
wire n_67;
wire n_37;
wire n_43;
wire n_50;
wire n_29;
wire n_12;
wire n_32;
wire n_70;
wire n_15;
wire n_66;

NAND2xp5_ASAP7_75t_SL g9 ( 
.A(n_0),
.B(n_2),
.Y(n_9)
);

INVx5_ASAP7_75t_L g10 ( 
.A(n_2),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_4),
.Y(n_11)
);

BUFx24_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

INVx3_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_8),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_7),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_1),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_9),
.B(n_3),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_19),
.B(n_11),
.Y(n_31)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_20),
.Y(n_30)
);

CKINVDCx9p33_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g27 ( 
.A(n_21),
.Y(n_27)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_24),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_25),
.A2(n_23),
.B1(n_24),
.B2(n_10),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_31),
.B(n_33),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g32 ( 
.A(n_20),
.B(n_13),
.C(n_14),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g40 ( 
.A(n_32),
.B(n_22),
.Y(n_40)
);

O2A1O1Ixp33_ASAP7_75t_L g33 ( 
.A1(n_21),
.A2(n_18),
.B(n_15),
.C(n_11),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_34),
.B(n_27),
.Y(n_35)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_33),
.B(n_19),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_41),
.Y(n_45)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_L g39 ( 
.A1(n_30),
.A2(n_23),
.B1(n_17),
.B2(n_18),
.Y(n_39)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_40),
.B(n_43),
.C(n_28),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_32),
.B(n_15),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_26),
.B(n_16),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_42),
.B(n_44),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_26),
.B(n_25),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_28),
.A2(n_17),
.B1(n_25),
.B2(n_22),
.Y(n_44)
);

INVx13_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

INVx13_ASAP7_75t_L g52 ( 
.A(n_47),
.Y(n_52)
);

XNOR2xp5_ASAP7_75t_L g54 ( 
.A(n_50),
.B(n_40),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_48),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_53),
.B(n_55),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_54),
.Y(n_57)
);

NOR4xp25_ASAP7_75t_L g55 ( 
.A(n_45),
.B(n_36),
.C(n_3),
.D(n_4),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_45),
.B(n_39),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g58 ( 
.A(n_56),
.Y(n_58)
);

OA21x2_ASAP7_75t_L g60 ( 
.A1(n_56),
.A2(n_46),
.B(n_51),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_60),
.A2(n_46),
.B1(n_49),
.B2(n_50),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_SL g64 ( 
.A1(n_61),
.A2(n_60),
.B(n_49),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_59),
.B(n_57),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_62),
.B(n_63),
.C(n_29),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_58),
.B(n_48),
.C(n_47),
.Y(n_63)
);

AO21x1_ASAP7_75t_L g66 ( 
.A1(n_64),
.A2(n_63),
.B(n_52),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_65),
.B(n_29),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_66),
.B(n_67),
.Y(n_68)
);

AO21x1_ASAP7_75t_L g69 ( 
.A1(n_68),
.A2(n_51),
.B(n_44),
.Y(n_69)
);

OAI321xp33_ASAP7_75t_L g70 ( 
.A1(n_69),
.A2(n_0),
.A3(n_6),
.B1(n_7),
.B2(n_25),
.C(n_68),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_70),
.B(n_6),
.Y(n_71)
);


endmodule