module real_jpeg_6669_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_498;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_128;
wire n_202;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_470;
wire n_372;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_215;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_502;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx8_ASAP7_75t_L g170 ( 
.A(n_0),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_0),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_0),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_0),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g306 ( 
.A(n_0),
.Y(n_306)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_0),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_1),
.A2(n_234),
.B1(n_236),
.B2(n_237),
.Y(n_233)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_1),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_L g286 ( 
.A1(n_1),
.A2(n_236),
.B1(n_287),
.B2(n_289),
.Y(n_286)
);

OAI22xp33_ASAP7_75t_SL g394 ( 
.A1(n_1),
.A2(n_178),
.B1(n_236),
.B2(n_395),
.Y(n_394)
);

AOI22xp33_ASAP7_75t_SL g455 ( 
.A1(n_1),
.A2(n_236),
.B1(n_456),
.B2(n_458),
.Y(n_455)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_2),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_2),
.Y(n_54)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_2),
.Y(n_56)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_2),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_2),
.Y(n_235)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_2),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_3),
.A2(n_87),
.B1(n_89),
.B2(n_90),
.Y(n_86)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_3),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_3),
.A2(n_90),
.B1(n_135),
.B2(n_136),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_3),
.A2(n_90),
.B1(n_178),
.B2(n_180),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_4),
.A2(n_34),
.B1(n_235),
.B2(n_282),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_4),
.Y(n_282)
);

AOI22xp33_ASAP7_75t_SL g321 ( 
.A1(n_4),
.A2(n_231),
.B1(n_282),
.B2(n_322),
.Y(n_321)
);

AOI22xp33_ASAP7_75t_L g406 ( 
.A1(n_4),
.A2(n_282),
.B1(n_407),
.B2(n_408),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_L g428 ( 
.A1(n_4),
.A2(n_282),
.B1(n_429),
.B2(n_432),
.Y(n_428)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

INVx3_ASAP7_75t_L g501 ( 
.A(n_6),
.Y(n_501)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_7),
.Y(n_70)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_7),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g389 ( 
.A(n_7),
.Y(n_389)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_8),
.Y(n_67)
);

OAI22xp33_ASAP7_75t_L g46 ( 
.A1(n_9),
.A2(n_47),
.B1(n_48),
.B2(n_49),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_9),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_9),
.A2(n_47),
.B1(n_230),
.B2(n_231),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g298 ( 
.A1(n_9),
.A2(n_47),
.B1(n_299),
.B2(n_300),
.Y(n_298)
);

AOI22xp33_ASAP7_75t_L g351 ( 
.A1(n_9),
.A2(n_47),
.B1(n_274),
.B2(n_352),
.Y(n_351)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_10),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_10),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g173 ( 
.A(n_10),
.Y(n_173)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_11),
.Y(n_99)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_12),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_SL g382 ( 
.A1(n_12),
.A2(n_262),
.B1(n_300),
.B2(n_383),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_12),
.B(n_389),
.C(n_390),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_SL g411 ( 
.A(n_12),
.B(n_106),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_12),
.B(n_423),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_12),
.B(n_85),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_12),
.B(n_294),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g504 ( 
.A(n_13),
.Y(n_504)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_14),
.A2(n_114),
.B1(n_115),
.B2(n_116),
.Y(n_113)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_14),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_14),
.A2(n_115),
.B1(n_139),
.B2(n_140),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_14),
.A2(n_115),
.B1(n_185),
.B2(n_186),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_L g272 ( 
.A1(n_14),
.A2(n_115),
.B1(n_273),
.B2(n_275),
.Y(n_272)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_16),
.A2(n_53),
.B1(n_55),
.B2(n_57),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_16),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_16),
.A2(n_57),
.B1(n_159),
.B2(n_161),
.Y(n_158)
);

OAI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_16),
.A2(n_57),
.B1(n_223),
.B2(n_224),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g266 ( 
.A1(n_16),
.A2(n_57),
.B1(n_171),
.B2(n_267),
.Y(n_266)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_17),
.A2(n_122),
.B1(n_124),
.B2(n_126),
.Y(n_121)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_17),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_17),
.A2(n_126),
.B1(n_149),
.B2(n_152),
.Y(n_148)
);

OAI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_17),
.A2(n_126),
.B1(n_171),
.B2(n_216),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_18),
.A2(n_194),
.B1(n_195),
.B2(n_196),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_18),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_18),
.A2(n_159),
.B1(n_194),
.B2(n_293),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_18),
.A2(n_150),
.B1(n_194),
.B2(n_311),
.Y(n_310)
);

AOI22xp33_ASAP7_75t_L g401 ( 
.A1(n_18),
.A2(n_194),
.B1(n_353),
.B2(n_402),
.Y(n_401)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_499),
.B(n_502),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_200),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_199),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_142),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_24),
.B(n_142),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_26),
.B1(n_127),
.B2(n_128),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_58),
.C(n_91),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_27),
.A2(n_129),
.B1(n_130),
.B2(n_141),
.Y(n_128)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_27),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_27),
.A2(n_141),
.B1(n_144),
.B2(n_145),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g27 ( 
.A1(n_28),
.A2(n_45),
.B1(n_50),
.B2(n_52),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_28),
.A2(n_50),
.B1(n_52),
.B2(n_138),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_28),
.A2(n_233),
.B(n_240),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g333 ( 
.A1(n_28),
.A2(n_38),
.B1(n_233),
.B2(n_281),
.Y(n_333)
);

INVx1_ASAP7_75t_SL g28 ( 
.A(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_29),
.B(n_193),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_29),
.A2(n_315),
.B(n_319),
.Y(n_314)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_38),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_31),
.A2(n_34),
.B1(n_35),
.B2(n_36),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx5_ASAP7_75t_L g256 ( 
.A(n_33),
.Y(n_256)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_34),
.Y(n_140)
);

INVx8_ASAP7_75t_L g195 ( 
.A(n_34),
.Y(n_195)
);

INVx3_ASAP7_75t_L g253 ( 
.A(n_35),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_35),
.B(n_262),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_36),
.A2(n_39),
.B1(n_40),
.B2(n_43),
.Y(n_38)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_37),
.Y(n_39)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_38),
.B(n_262),
.Y(n_357)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_42),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g101 ( 
.A(n_42),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_42),
.Y(n_105)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_42),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g252 ( 
.A(n_42),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_44),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_44),
.Y(n_163)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_44),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_44),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_44),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_46),
.B(n_51),
.Y(n_191)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_48),
.Y(n_49)
);

OAI21xp5_ASAP7_75t_L g280 ( 
.A1(n_50),
.A2(n_192),
.B(n_281),
.Y(n_280)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_51),
.B(n_193),
.Y(n_240)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx8_ASAP7_75t_L g139 ( 
.A(n_54),
.Y(n_139)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_58),
.A2(n_59),
.B1(n_132),
.B2(n_133),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_58),
.A2(n_59),
.B1(n_91),
.B2(n_92),
.Y(n_144)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

AOI21xp5_ASAP7_75t_SL g59 ( 
.A1(n_60),
.A2(n_84),
.B(n_86),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_60),
.A2(n_84),
.B1(n_298),
.B2(n_302),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_SL g381 ( 
.A1(n_60),
.A2(n_382),
.B(n_384),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_SL g454 ( 
.A1(n_60),
.A2(n_84),
.B1(n_406),
.B2(n_455),
.Y(n_454)
);

OAI21xp5_ASAP7_75t_SL g480 ( 
.A1(n_60),
.A2(n_384),
.B(n_455),
.Y(n_480)
);

INVx2_ASAP7_75t_SL g60 ( 
.A(n_61),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_61),
.A2(n_85),
.B1(n_148),
.B2(n_154),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_61),
.A2(n_85),
.B1(n_148),
.B2(n_184),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_61),
.A2(n_85),
.B1(n_184),
.B2(n_222),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_61),
.B(n_310),
.Y(n_309)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_75),
.Y(n_61)
);

OAI22xp33_ASAP7_75t_L g62 ( 
.A1(n_63),
.A2(n_68),
.B1(n_71),
.B2(n_74),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_65),
.Y(n_89)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_66),
.Y(n_74)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_66),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_66),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_66),
.Y(n_227)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

BUFx5_ASAP7_75t_L g109 ( 
.A(n_67),
.Y(n_109)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_67),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g312 ( 
.A(n_67),
.Y(n_312)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_67),
.Y(n_409)
);

INVx3_ASAP7_75t_L g472 ( 
.A(n_67),
.Y(n_472)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_70),
.Y(n_76)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_73),
.Y(n_83)
);

AO22x2_ASAP7_75t_L g106 ( 
.A1(n_74),
.A2(n_107),
.B1(n_109),
.B2(n_110),
.Y(n_106)
);

INVx11_ASAP7_75t_L g407 ( 
.A(n_74),
.Y(n_407)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_75),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_SL g405 ( 
.A1(n_75),
.A2(n_309),
.B(n_406),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_77),
.B1(n_81),
.B2(n_83),
.Y(n_75)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_78),
.Y(n_274)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_79),
.Y(n_355)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_80),
.Y(n_217)
);

BUFx3_ASAP7_75t_L g277 ( 
.A(n_80),
.Y(n_277)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_82),
.Y(n_179)
);

BUFx5_ASAP7_75t_L g433 ( 
.A(n_82),
.Y(n_433)
);

OAI21xp5_ASAP7_75t_SL g308 ( 
.A1(n_84),
.A2(n_298),
.B(n_309),
.Y(n_308)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g384 ( 
.A(n_85),
.B(n_310),
.Y(n_384)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_86),
.Y(n_154)
);

BUFx2_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_88),
.Y(n_153)
);

INVx5_ASAP7_75t_L g457 ( 
.A(n_88),
.Y(n_457)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_93),
.A2(n_112),
.B1(n_120),
.B2(n_121),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_93),
.A2(n_120),
.B1(n_121),
.B2(n_134),
.Y(n_133)
);

INVx3_ASAP7_75t_SL g156 ( 
.A(n_93),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_93),
.A2(n_120),
.B1(n_158),
.B2(n_229),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_93),
.A2(n_120),
.B1(n_286),
.B2(n_321),
.Y(n_320)
);

OR2x2_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_106),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_95),
.A2(n_100),
.B1(n_102),
.B2(n_103),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_97),
.Y(n_102)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g469 ( 
.A(n_98),
.Y(n_469)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_99),
.Y(n_108)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_99),
.Y(n_111)
);

INVx3_ASAP7_75t_L g294 ( 
.A(n_100),
.Y(n_294)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_101),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g135 ( 
.A(n_101),
.Y(n_135)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

BUFx2_ASAP7_75t_L g114 ( 
.A(n_104),
.Y(n_114)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_105),
.Y(n_125)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_105),
.Y(n_136)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_105),
.Y(n_288)
);

INVx3_ASAP7_75t_L g323 ( 
.A(n_105),
.Y(n_323)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_106),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_106),
.A2(n_113),
.B1(n_156),
.B2(n_157),
.Y(n_155)
);

AOI22x1_ASAP7_75t_L g330 ( 
.A1(n_106),
.A2(n_156),
.B1(n_331),
.B2(n_332),
.Y(n_330)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx5_ASAP7_75t_L g185 ( 
.A(n_109),
.Y(n_185)
);

INVx4_ASAP7_75t_L g473 ( 
.A(n_110),
.Y(n_473)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_120),
.B(n_292),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_SL g348 ( 
.A1(n_120),
.A2(n_321),
.B(n_349),
.Y(n_348)
);

INVx6_ASAP7_75t_L g231 ( 
.A(n_122),
.Y(n_231)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx5_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_SL g130 ( 
.A(n_131),
.B(n_137),
.Y(n_130)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_146),
.C(n_164),
.Y(n_142)
);

FAx1_ASAP7_75t_SL g202 ( 
.A(n_143),
.B(n_146),
.CI(n_164),
.CON(n_202),
.SN(n_202)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_144),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_146),
.A2(n_210),
.B(n_211),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_155),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_147),
.Y(n_211)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_151),
.Y(n_301)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_155),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_156),
.A2(n_285),
.B(n_291),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_156),
.B(n_331),
.Y(n_349)
);

AOI21xp5_ASAP7_75t_L g460 ( 
.A1(n_156),
.A2(n_291),
.B(n_461),
.Y(n_460)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

OAI21xp33_ASAP7_75t_SL g461 ( 
.A1(n_161),
.A2(n_262),
.B(n_462),
.Y(n_461)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_165),
.A2(n_166),
.B(n_190),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_165),
.B(n_206),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_183),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_166),
.A2(n_190),
.B1(n_207),
.B2(n_208),
.Y(n_206)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_166),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_166),
.A2(n_183),
.B1(n_208),
.B2(n_367),
.Y(n_366)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_167),
.A2(n_174),
.B(n_177),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_167),
.A2(n_177),
.B1(n_215),
.B2(n_218),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_167),
.A2(n_265),
.B1(n_268),
.B2(n_271),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g393 ( 
.A1(n_167),
.A2(n_394),
.B(n_398),
.Y(n_393)
);

AOI21xp5_ASAP7_75t_L g425 ( 
.A1(n_167),
.A2(n_262),
.B(n_398),
.Y(n_425)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_168),
.A2(n_272),
.B1(n_304),
.B2(n_305),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_168),
.A2(n_266),
.B1(n_351),
.B2(n_356),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_168),
.B(n_401),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_SL g441 ( 
.A1(n_168),
.A2(n_442),
.B1(n_443),
.B2(n_444),
.Y(n_441)
);

OR2x2_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_171),
.Y(n_168)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_170),
.Y(n_400)
);

BUFx6f_ASAP7_75t_L g424 ( 
.A(n_170),
.Y(n_424)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_170),
.Y(n_436)
);

INVx8_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

BUFx2_ASAP7_75t_L g267 ( 
.A(n_172),
.Y(n_267)
);

BUFx8_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

BUFx5_ASAP7_75t_L g182 ( 
.A(n_173),
.Y(n_182)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_173),
.Y(n_421)
);

BUFx3_ASAP7_75t_L g431 ( 
.A(n_173),
.Y(n_431)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

BUFx2_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g367 ( 
.A(n_183),
.Y(n_367)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_185),
.Y(n_299)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_186),
.Y(n_223)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx4_ASAP7_75t_SL g187 ( 
.A(n_188),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

BUFx3_ASAP7_75t_L g387 ( 
.A(n_189),
.Y(n_387)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_190),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_192),
.Y(n_190)
);

INVx5_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_201),
.A2(n_241),
.B(n_498),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_202),
.B(n_203),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_202),
.B(n_203),
.Y(n_498)
);

BUFx24_ASAP7_75t_SL g505 ( 
.A(n_202),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_209),
.C(n_212),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_204),
.A2(n_205),
.B1(n_209),
.B2(n_371),
.Y(n_370)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_209),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_L g369 ( 
.A(n_212),
.B(n_370),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_228),
.C(n_232),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_213),
.B(n_365),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_221),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_214),
.B(n_221),
.Y(n_336)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_215),
.Y(n_304)
);

INVx4_ASAP7_75t_L g402 ( 
.A(n_216),
.Y(n_402)
);

INVx8_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

HB1xp67_ASAP7_75t_L g391 ( 
.A(n_217),
.Y(n_391)
);

BUFx3_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_222),
.Y(n_302)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_227),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_228),
.B(n_232),
.Y(n_365)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_229),
.Y(n_332)
);

AOI32xp33_ASAP7_75t_L g467 ( 
.A1(n_231),
.A2(n_312),
.A3(n_463),
.B1(n_468),
.B2(n_470),
.Y(n_467)
);

INVx4_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_239),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_240),
.Y(n_319)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

HB1xp67_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

OAI311xp33_ASAP7_75t_L g243 ( 
.A1(n_244),
.A2(n_361),
.A3(n_375),
.B1(n_492),
.C1(n_497),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_245),
.B(n_339),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_L g493 ( 
.A1(n_246),
.A2(n_494),
.B(n_495),
.Y(n_493)
);

NOR2x1_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_324),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_247),
.B(n_324),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_295),
.C(n_307),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g358 ( 
.A(n_248),
.B(n_359),
.Y(n_358)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_278),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_249),
.B(n_279),
.C(n_284),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_263),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g345 ( 
.A1(n_250),
.A2(n_263),
.B1(n_264),
.B2(n_346),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_250),
.Y(n_346)
);

OAI32xp33_ASAP7_75t_L g250 ( 
.A1(n_251),
.A2(n_253),
.A3(n_254),
.B1(n_257),
.B2(n_261),
.Y(n_250)
);

INVx4_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_255),
.B(n_258),
.Y(n_257)
);

INVx6_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

OAI21xp33_ASAP7_75t_SL g315 ( 
.A1(n_261),
.A2(n_262),
.B(n_316),
.Y(n_315)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx3_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

BUFx3_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g397 ( 
.A(n_277),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_279),
.A2(n_280),
.B1(n_283),
.B2(n_284),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx3_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

BUFx12f_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_292),
.Y(n_331)
);

INVx4_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_295),
.A2(n_296),
.B1(n_307),
.B2(n_360),
.Y(n_359)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_303),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_297),
.B(n_303),
.Y(n_328)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx4_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_307),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_313),
.C(n_320),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_SL g342 ( 
.A(n_308),
.B(n_320),
.Y(n_342)
);

INVx5_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_313),
.A2(n_314),
.B1(n_342),
.B2(n_343),
.Y(n_341)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx3_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx4_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_326),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_325),
.B(n_336),
.C(n_337),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_327),
.A2(n_336),
.B1(n_337),
.B2(n_338),
.Y(n_326)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_327),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_329),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_328),
.B(n_330),
.C(n_335),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_330),
.A2(n_333),
.B1(n_334),
.B2(n_335),
.Y(n_329)
);

INVx1_ASAP7_75t_SL g334 ( 
.A(n_330),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_333),
.Y(n_335)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_336),
.Y(n_338)
);

OR2x2_ASAP7_75t_L g339 ( 
.A(n_340),
.B(n_358),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_340),
.B(n_358),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_341),
.B(n_344),
.C(n_347),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g488 ( 
.A(n_341),
.B(n_489),
.Y(n_488)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_342),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g489 ( 
.A1(n_344),
.A2(n_345),
.B1(n_347),
.B2(n_490),
.Y(n_489)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_347),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_348),
.B(n_350),
.C(n_357),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_SL g482 ( 
.A(n_348),
.B(n_483),
.Y(n_482)
);

XOR2xp5_ASAP7_75t_L g483 ( 
.A(n_350),
.B(n_357),
.Y(n_483)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_351),
.Y(n_466)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

INVx4_ASAP7_75t_SL g353 ( 
.A(n_354),
.Y(n_353)
);

INVx4_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

NAND2xp33_ASAP7_75t_SL g361 ( 
.A(n_362),
.B(n_372),
.Y(n_361)
);

A2O1A1Ixp33_ASAP7_75t_SL g492 ( 
.A1(n_362),
.A2(n_372),
.B(n_493),
.C(n_496),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_363),
.B(n_369),
.Y(n_362)
);

OR2x2_ASAP7_75t_L g497 ( 
.A(n_363),
.B(n_369),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_364),
.B(n_366),
.C(n_368),
.Y(n_363)
);

FAx1_ASAP7_75t_SL g374 ( 
.A(n_364),
.B(n_366),
.CI(n_368),
.CON(n_374),
.SN(n_374)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_373),
.B(n_374),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_373),
.B(n_374),
.Y(n_496)
);

BUFx24_ASAP7_75t_SL g507 ( 
.A(n_374),
.Y(n_507)
);

AOI21xp5_ASAP7_75t_SL g375 ( 
.A1(n_376),
.A2(n_486),
.B(n_491),
.Y(n_375)
);

AO21x1_ASAP7_75t_SL g376 ( 
.A1(n_377),
.A2(n_475),
.B(n_485),
.Y(n_376)
);

OAI21xp5_ASAP7_75t_SL g377 ( 
.A1(n_378),
.A2(n_449),
.B(n_474),
.Y(n_377)
);

AOI21xp5_ASAP7_75t_L g378 ( 
.A1(n_379),
.A2(n_412),
.B(n_448),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_380),
.B(n_392),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_380),
.B(n_392),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_SL g380 ( 
.A(n_381),
.B(n_385),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_SL g445 ( 
.A1(n_381),
.A2(n_385),
.B1(n_386),
.B2(n_446),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_381),
.Y(n_446)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_387),
.B(n_388),
.Y(n_386)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_393),
.B(n_403),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_393),
.B(n_404),
.C(n_411),
.Y(n_450)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_394),
.Y(n_443)
);

INVx6_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

INVx4_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_399),
.B(n_401),
.Y(n_398)
);

INVx4_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_SL g403 ( 
.A1(n_404),
.A2(n_405),
.B1(n_410),
.B2(n_411),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_407),
.Y(n_458)
);

BUFx3_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

OAI21xp5_ASAP7_75t_L g412 ( 
.A1(n_413),
.A2(n_440),
.B(n_447),
.Y(n_412)
);

AOI21xp5_ASAP7_75t_L g413 ( 
.A1(n_414),
.A2(n_426),
.B(n_439),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_415),
.B(n_425),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_416),
.B(n_422),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

INVx1_ASAP7_75t_SL g417 ( 
.A(n_418),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_423),
.Y(n_444)
);

INVx8_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_SL g426 ( 
.A(n_427),
.B(n_438),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_427),
.B(n_438),
.Y(n_439)
);

AOI21xp5_ASAP7_75t_L g427 ( 
.A1(n_428),
.A2(n_434),
.B(n_437),
.Y(n_427)
);

INVxp67_ASAP7_75t_L g442 ( 
.A(n_428),
.Y(n_442)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

INVx5_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

INVx5_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

INVx3_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

AOI21xp5_ASAP7_75t_L g465 ( 
.A1(n_436),
.A2(n_437),
.B(n_466),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_441),
.B(n_445),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_441),
.B(n_445),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_450),
.B(n_451),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_450),
.B(n_451),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_L g451 ( 
.A(n_452),
.B(n_464),
.Y(n_451)
);

AOI22xp5_ASAP7_75t_L g452 ( 
.A1(n_453),
.A2(n_454),
.B1(n_459),
.B2(n_460),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_454),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_454),
.B(n_459),
.C(n_464),
.Y(n_476)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_457),
.Y(n_456)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_460),
.Y(n_459)
);

INVxp33_ASAP7_75t_L g462 ( 
.A(n_463),
.Y(n_462)
);

XOR2xp5_ASAP7_75t_L g464 ( 
.A(n_465),
.B(n_467),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_465),
.B(n_467),
.Y(n_481)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_469),
.Y(n_468)
);

NAND2xp33_ASAP7_75t_SL g470 ( 
.A(n_471),
.B(n_473),
.Y(n_470)
);

BUFx6f_ASAP7_75t_L g471 ( 
.A(n_472),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_476),
.B(n_477),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_SL g485 ( 
.A(n_476),
.B(n_477),
.Y(n_485)
);

AOI22xp5_ASAP7_75t_L g477 ( 
.A1(n_478),
.A2(n_479),
.B1(n_482),
.B2(n_484),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_479),
.Y(n_478)
);

XNOR2xp5_ASAP7_75t_SL g479 ( 
.A(n_480),
.B(n_481),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_480),
.B(n_481),
.C(n_484),
.Y(n_487)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_482),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_487),
.B(n_488),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_SL g491 ( 
.A(n_487),
.B(n_488),
.Y(n_491)
);

BUFx6f_ASAP7_75t_L g499 ( 
.A(n_500),
.Y(n_499)
);

BUFx6f_ASAP7_75t_L g503 ( 
.A(n_500),
.Y(n_503)
);

INVx13_ASAP7_75t_L g500 ( 
.A(n_501),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_503),
.B(n_504),
.Y(n_502)
);


endmodule