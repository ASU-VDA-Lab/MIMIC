module fake_jpeg_2229_n_425 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_425);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_425;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_260;
wire n_199;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_9),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_15),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx8_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_2),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

BUFx10_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_16),
.Y(n_37)
);

INVx13_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

INVx13_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_16),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

CKINVDCx16_ASAP7_75t_R g43 ( 
.A(n_8),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_17),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_17),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_7),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_12),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_12),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_11),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_3),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_5),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_13),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_10),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_37),
.B(n_0),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_55),
.B(n_70),
.Y(n_123)
);

INVx6_ASAP7_75t_SL g56 ( 
.A(n_31),
.Y(n_56)
);

CKINVDCx9p33_ASAP7_75t_R g117 ( 
.A(n_56),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_57),
.Y(n_116)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_32),
.Y(n_58)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_58),
.Y(n_136)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_31),
.Y(n_59)
);

INVx2_ASAP7_75t_SL g151 ( 
.A(n_59),
.Y(n_151)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_31),
.Y(n_60)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_60),
.Y(n_131)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_61),
.Y(n_142)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_32),
.Y(n_62)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_62),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_63),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_37),
.B(n_0),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_64),
.B(n_66),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_65),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_31),
.Y(n_66)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_35),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g172 ( 
.A(n_67),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_41),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_68),
.B(n_71),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_35),
.Y(n_69)
);

INVx6_ASAP7_75t_L g169 ( 
.A(n_69),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_41),
.B(n_0),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_46),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_46),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_72),
.B(n_77),
.Y(n_126)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_20),
.Y(n_73)
);

INVx1_ASAP7_75t_SL g154 ( 
.A(n_73),
.Y(n_154)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_74),
.Y(n_156)
);

BUFx4f_ASAP7_75t_SL g75 ( 
.A(n_20),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_75),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_35),
.Y(n_76)
);

INVx3_ASAP7_75t_SL g127 ( 
.A(n_76),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_27),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_50),
.Y(n_78)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_78),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_49),
.Y(n_79)
);

INVx3_ASAP7_75t_SL g148 ( 
.A(n_79),
.Y(n_148)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_49),
.Y(n_80)
);

INVx5_ASAP7_75t_L g157 ( 
.A(n_80),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_54),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_81),
.B(n_93),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_49),
.Y(n_82)
);

INVx8_ASAP7_75t_L g174 ( 
.A(n_82),
.Y(n_174)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_49),
.Y(n_83)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_83),
.Y(n_130)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_53),
.Y(n_84)
);

INVx5_ASAP7_75t_L g143 ( 
.A(n_84),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_53),
.Y(n_85)
);

BUFx12f_ASAP7_75t_L g115 ( 
.A(n_85),
.Y(n_115)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_53),
.Y(n_86)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_86),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_45),
.B(n_1),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_87),
.B(n_88),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_27),
.B(n_3),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_23),
.Y(n_89)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_89),
.Y(n_139)
);

BUFx12f_ASAP7_75t_L g90 ( 
.A(n_20),
.Y(n_90)
);

INVx5_ASAP7_75t_L g159 ( 
.A(n_90),
.Y(n_159)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_23),
.Y(n_91)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_91),
.Y(n_140)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_53),
.Y(n_92)
);

HB1xp67_ASAP7_75t_L g184 ( 
.A(n_92),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_54),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_18),
.Y(n_94)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_94),
.Y(n_161)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_18),
.Y(n_95)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_95),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_52),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_96),
.B(n_100),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_19),
.B(n_4),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_97),
.B(n_114),
.Y(n_153)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_38),
.Y(n_98)
);

INVx5_ASAP7_75t_L g185 ( 
.A(n_98),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_20),
.Y(n_99)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_99),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_38),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_19),
.Y(n_101)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_101),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_28),
.B(n_4),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_102),
.B(n_106),
.Y(n_173)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_21),
.Y(n_103)
);

BUFx24_ASAP7_75t_L g122 ( 
.A(n_103),
.Y(n_122)
);

INVx11_ASAP7_75t_L g104 ( 
.A(n_40),
.Y(n_104)
);

INVx5_ASAP7_75t_SL g128 ( 
.A(n_104),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_21),
.Y(n_105)
);

BUFx2_ASAP7_75t_SL g162 ( 
.A(n_105),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_52),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_22),
.Y(n_107)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_107),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_28),
.B(n_5),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_108),
.B(n_111),
.Y(n_178)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_22),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_109),
.B(n_110),
.Y(n_158)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_36),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_29),
.B(n_6),
.Y(n_111)
);

INVx8_ASAP7_75t_L g112 ( 
.A(n_40),
.Y(n_112)
);

BUFx12_ASAP7_75t_L g121 ( 
.A(n_112),
.Y(n_121)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_24),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_113),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_51),
.B(n_7),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_103),
.B(n_51),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_118),
.B(n_119),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_101),
.B(n_29),
.Y(n_119)
);

AND2x2_ASAP7_75t_SL g120 ( 
.A(n_59),
.B(n_33),
.Y(n_120)
);

CKINVDCx14_ASAP7_75t_R g233 ( 
.A(n_120),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_105),
.B(n_48),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_132),
.B(n_141),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_57),
.A2(n_33),
.B1(n_47),
.B2(n_42),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_133),
.A2(n_137),
.B1(n_152),
.B2(n_170),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_61),
.A2(n_34),
.B1(n_48),
.B2(n_30),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_134),
.A2(n_167),
.B1(n_168),
.B2(n_177),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_63),
.A2(n_47),
.B1(n_42),
.B2(n_39),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_83),
.B(n_34),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_98),
.B(n_30),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_147),
.B(n_160),
.Y(n_231)
);

OR2x2_ASAP7_75t_L g150 ( 
.A(n_92),
.B(n_25),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_150),
.B(n_155),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_L g152 ( 
.A1(n_60),
.A2(n_25),
.B1(n_39),
.B2(n_26),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_86),
.B(n_24),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_65),
.Y(n_160)
);

CKINVDCx12_ASAP7_75t_R g163 ( 
.A(n_75),
.Y(n_163)
);

BUFx12f_ASAP7_75t_L g229 ( 
.A(n_163),
.Y(n_229)
);

OR2x2_ASAP7_75t_L g165 ( 
.A(n_69),
.B(n_26),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_165),
.B(n_182),
.Y(n_230)
);

OAI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_76),
.A2(n_79),
.B1(n_85),
.B2(n_82),
.Y(n_167)
);

OAI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_110),
.A2(n_43),
.B1(n_36),
.B2(n_45),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_67),
.A2(n_36),
.B1(n_43),
.B2(n_12),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_80),
.A2(n_84),
.B1(n_104),
.B2(n_90),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_175),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_99),
.A2(n_36),
.B1(n_11),
.B2(n_15),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_L g181 ( 
.A1(n_112),
.A2(n_8),
.B1(n_15),
.B2(n_73),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_181),
.A2(n_168),
.B1(n_167),
.B2(n_179),
.Y(n_213)
);

OR2x2_ASAP7_75t_SL g182 ( 
.A(n_73),
.B(n_90),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_88),
.B(n_114),
.Y(n_186)
);

NOR2x1_ASAP7_75t_L g205 ( 
.A(n_186),
.B(n_153),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_144),
.B(n_126),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_187),
.B(n_189),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_125),
.B(n_124),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_146),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_190),
.B(n_203),
.Y(n_261)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_176),
.Y(n_191)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_191),
.Y(n_259)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_161),
.Y(n_192)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_192),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_173),
.B(n_171),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_193),
.B(n_197),
.Y(n_256)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_166),
.Y(n_194)
);

INVxp67_ASAP7_75t_SL g250 ( 
.A(n_194),
.Y(n_250)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_183),
.Y(n_195)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_195),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_123),
.B(n_135),
.Y(n_197)
);

OR2x2_ASAP7_75t_SL g198 ( 
.A(n_120),
.B(n_117),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g263 ( 
.A(n_198),
.Y(n_263)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_157),
.Y(n_200)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_200),
.Y(n_286)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_162),
.Y(n_201)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_201),
.Y(n_273)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_136),
.Y(n_202)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_202),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_146),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_156),
.Y(n_204)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_204),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_205),
.B(n_208),
.Y(n_269)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_158),
.Y(n_206)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_206),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_184),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_158),
.Y(n_209)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_209),
.Y(n_292)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_151),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_210),
.Y(n_257)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_142),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_211),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_150),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_212),
.B(n_217),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_213),
.A2(n_216),
.B1(n_236),
.B2(n_243),
.Y(n_268)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_142),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_214),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_178),
.B(n_129),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_151),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_218),
.B(n_220),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_138),
.B(n_165),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_219),
.B(n_234),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_130),
.B(n_140),
.Y(n_220)
);

INVx8_ASAP7_75t_L g221 ( 
.A(n_115),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_SL g287 ( 
.A1(n_221),
.A2(n_239),
.B1(n_241),
.B2(n_245),
.Y(n_287)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_139),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_222),
.B(n_223),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_149),
.B(n_185),
.Y(n_223)
);

AND2x2_ASAP7_75t_SL g224 ( 
.A(n_149),
.B(n_154),
.Y(n_224)
);

CKINVDCx16_ASAP7_75t_R g276 ( 
.A(n_224),
.Y(n_276)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_157),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g275 ( 
.A(n_225),
.Y(n_275)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_152),
.Y(n_226)
);

NAND2xp33_ASAP7_75t_SL g252 ( 
.A(n_226),
.B(n_227),
.Y(n_252)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_127),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_116),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_228),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_172),
.B(n_154),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_232),
.A2(n_235),
.B1(n_240),
.B2(n_247),
.Y(n_280)
);

AO22x1_ASAP7_75t_SL g234 ( 
.A1(n_116),
.A2(n_164),
.B1(n_145),
.B2(n_127),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_172),
.B(n_143),
.Y(n_235)
);

HAxp5_ASAP7_75t_SL g236 ( 
.A(n_122),
.B(n_181),
.CON(n_236),
.SN(n_236)
);

NOR3xp33_ASAP7_75t_SL g255 ( 
.A(n_236),
.B(n_237),
.C(n_242),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_169),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_164),
.B(n_169),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_238),
.B(n_243),
.Y(n_251)
);

INVx1_ASAP7_75t_SL g239 ( 
.A(n_159),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_128),
.B(n_174),
.Y(n_240)
);

INVx1_ASAP7_75t_SL g241 ( 
.A(n_131),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_180),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_180),
.B(n_148),
.Y(n_243)
);

AND2x2_ASAP7_75t_L g244 ( 
.A(n_131),
.B(n_148),
.Y(n_244)
);

AND2x2_ASAP7_75t_SL g260 ( 
.A(n_244),
.B(n_121),
.Y(n_260)
);

BUFx12f_ASAP7_75t_L g245 ( 
.A(n_121),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_115),
.B(n_170),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_246),
.B(n_213),
.Y(n_270)
);

BUFx2_ASAP7_75t_L g247 ( 
.A(n_174),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_196),
.A2(n_175),
.B1(n_115),
.B2(n_122),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_248),
.A2(n_254),
.B1(n_285),
.B2(n_221),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_196),
.A2(n_122),
.B1(n_128),
.B2(n_121),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_206),
.B(n_209),
.C(n_233),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_258),
.B(n_288),
.C(n_244),
.Y(n_293)
);

AND2x2_ASAP7_75t_L g306 ( 
.A(n_260),
.B(n_268),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_226),
.A2(n_207),
.B1(n_219),
.B2(n_246),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_265),
.A2(n_280),
.B1(n_251),
.B2(n_260),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_216),
.A2(n_230),
.B(n_198),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_L g317 ( 
.A1(n_266),
.A2(n_289),
.B(n_252),
.Y(n_317)
);

FAx1_ASAP7_75t_SL g267 ( 
.A(n_205),
.B(n_215),
.CI(n_199),
.CON(n_267),
.SN(n_267)
);

OAI32xp33_ASAP7_75t_L g314 ( 
.A1(n_267),
.A2(n_292),
.A3(n_251),
.B1(n_255),
.B2(n_262),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g320 ( 
.A(n_270),
.Y(n_320)
);

AOI22xp33_ASAP7_75t_L g271 ( 
.A1(n_202),
.A2(n_191),
.B1(n_234),
.B2(n_238),
.Y(n_271)
);

INVxp33_ASAP7_75t_L g299 ( 
.A(n_271),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_234),
.A2(n_214),
.B1(n_211),
.B2(n_224),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_224),
.B(n_218),
.C(n_200),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_201),
.A2(n_241),
.B(n_231),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_188),
.B(n_225),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_290),
.B(n_267),
.Y(n_304)
);

OAI22xp33_ASAP7_75t_SL g291 ( 
.A1(n_247),
.A2(n_227),
.B1(n_228),
.B2(n_239),
.Y(n_291)
);

AOI22xp33_ASAP7_75t_L g310 ( 
.A1(n_291),
.A2(n_273),
.B1(n_279),
.B2(n_249),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_293),
.B(n_301),
.C(n_305),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_277),
.B(n_244),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_294),
.B(n_300),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_295),
.A2(n_316),
.B1(n_248),
.B2(n_264),
.Y(n_327)
);

NAND3xp33_ASAP7_75t_L g296 ( 
.A(n_263),
.B(n_229),
.C(n_245),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_296),
.B(n_312),
.Y(n_328)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_274),
.Y(n_297)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_297),
.Y(n_329)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_274),
.Y(n_298)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_298),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_256),
.B(n_253),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_258),
.B(n_229),
.C(n_245),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_265),
.A2(n_229),
.B1(n_270),
.B2(n_249),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_L g345 ( 
.A1(n_302),
.A2(n_305),
.B1(n_293),
.B2(n_309),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_290),
.B(n_272),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_303),
.B(n_304),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_276),
.B(n_283),
.C(n_288),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_269),
.B(n_261),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_SL g344 ( 
.A(n_307),
.B(n_311),
.Y(n_344)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_262),
.Y(n_308)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_308),
.Y(n_347)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_283),
.B(n_292),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_SL g336 ( 
.A(n_309),
.B(n_314),
.Y(n_336)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_310),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_282),
.B(n_278),
.Y(n_311)
);

AND2x6_ASAP7_75t_L g312 ( 
.A(n_267),
.B(n_266),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_250),
.B(n_289),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_SL g346 ( 
.A(n_313),
.B(n_315),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_281),
.B(n_257),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_SL g343 ( 
.A1(n_317),
.A2(n_322),
.B(n_306),
.Y(n_343)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_280),
.B(n_260),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_318),
.B(n_319),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_281),
.B(n_259),
.Y(n_319)
);

INVx13_ASAP7_75t_L g321 ( 
.A(n_287),
.Y(n_321)
);

CKINVDCx16_ASAP7_75t_R g331 ( 
.A(n_321),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_259),
.B(n_255),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_322),
.B(n_325),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_257),
.B(n_286),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g348 ( 
.A(n_323),
.B(n_298),
.Y(n_348)
);

INVx11_ASAP7_75t_L g324 ( 
.A(n_286),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_324),
.B(n_326),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_254),
.B(n_285),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_273),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_L g360 ( 
.A1(n_327),
.A2(n_332),
.B1(n_339),
.B2(n_341),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_316),
.A2(n_275),
.B1(n_264),
.B2(n_284),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_319),
.B(n_275),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_334),
.B(n_337),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_302),
.B(n_284),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_320),
.A2(n_325),
.B1(n_295),
.B2(n_299),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_320),
.A2(n_299),
.B1(n_306),
.B2(n_318),
.Y(n_341)
);

AOI21xp5_ASAP7_75t_L g352 ( 
.A1(n_343),
.A2(n_301),
.B(n_314),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_345),
.A2(n_333),
.B1(n_341),
.B2(n_350),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_348),
.B(n_350),
.Y(n_357)
);

OR2x2_ASAP7_75t_L g350 ( 
.A(n_317),
.B(n_306),
.Y(n_350)
);

INVxp67_ASAP7_75t_L g382 ( 
.A(n_352),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_351),
.B(n_312),
.C(n_324),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_353),
.B(n_354),
.C(n_361),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_351),
.B(n_321),
.C(n_345),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_344),
.B(n_346),
.Y(n_355)
);

INVxp33_ASAP7_75t_L g377 ( 
.A(n_355),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_338),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_358),
.Y(n_385)
);

AND2x2_ASAP7_75t_L g359 ( 
.A(n_350),
.B(n_337),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_359),
.Y(n_380)
);

BUFx24_ASAP7_75t_SL g362 ( 
.A(n_344),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_SL g376 ( 
.A(n_362),
.B(n_365),
.Y(n_376)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_348),
.Y(n_363)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_363),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_334),
.B(n_349),
.Y(n_364)
);

HB1xp67_ASAP7_75t_L g378 ( 
.A(n_364),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_SL g365 ( 
.A(n_342),
.B(n_335),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_329),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_L g372 ( 
.A1(n_366),
.A2(n_368),
.B1(n_369),
.B2(n_370),
.Y(n_372)
);

XOR2xp5_ASAP7_75t_L g367 ( 
.A(n_333),
.B(n_336),
.Y(n_367)
);

XOR2xp5_ASAP7_75t_SL g374 ( 
.A(n_367),
.B(n_343),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_349),
.B(n_330),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_346),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_SL g370 ( 
.A(n_330),
.B(n_347),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_L g390 ( 
.A(n_374),
.B(n_367),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_360),
.A2(n_327),
.B1(n_339),
.B2(n_332),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_375),
.B(n_379),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_364),
.A2(n_328),
.B1(n_331),
.B2(n_336),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_352),
.A2(n_331),
.B1(n_329),
.B2(n_347),
.Y(n_381)
);

INVxp67_ASAP7_75t_L g388 ( 
.A(n_381),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_368),
.A2(n_340),
.B1(n_356),
.B2(n_359),
.Y(n_383)
);

INVxp67_ASAP7_75t_L g392 ( 
.A(n_383),
.Y(n_392)
);

AO22x1_ASAP7_75t_L g384 ( 
.A1(n_359),
.A2(n_340),
.B1(n_363),
.B2(n_357),
.Y(n_384)
);

OAI21xp5_ASAP7_75t_L g394 ( 
.A1(n_384),
.A2(n_357),
.B(n_356),
.Y(n_394)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_372),
.Y(n_386)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_386),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_385),
.B(n_369),
.Y(n_387)
);

INVxp67_ASAP7_75t_SL g406 ( 
.A(n_387),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_378),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_389),
.B(n_391),
.Y(n_399)
);

XOR2xp5_ASAP7_75t_L g398 ( 
.A(n_390),
.B(n_397),
.Y(n_398)
);

CKINVDCx16_ASAP7_75t_R g391 ( 
.A(n_383),
.Y(n_391)
);

INVx11_ASAP7_75t_L g393 ( 
.A(n_385),
.Y(n_393)
);

AO21x1_ASAP7_75t_L g403 ( 
.A1(n_393),
.A2(n_394),
.B(n_395),
.Y(n_403)
);

AOI321xp33_ASAP7_75t_L g395 ( 
.A1(n_380),
.A2(n_353),
.A3(n_354),
.B1(n_361),
.B2(n_358),
.C(n_366),
.Y(n_395)
);

XOR2x2_ASAP7_75t_L g397 ( 
.A(n_379),
.B(n_371),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_397),
.B(n_371),
.C(n_382),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_400),
.B(n_401),
.C(n_392),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_390),
.B(n_382),
.C(n_377),
.Y(n_401)
);

BUFx24_ASAP7_75t_SL g402 ( 
.A(n_395),
.Y(n_402)
);

OAI21xp5_ASAP7_75t_L g408 ( 
.A1(n_402),
.A2(n_405),
.B(n_406),
.Y(n_408)
);

A2O1A1Ixp33_ASAP7_75t_SL g405 ( 
.A1(n_396),
.A2(n_381),
.B(n_384),
.C(n_373),
.Y(n_405)
);

AOI21xp5_ASAP7_75t_L g407 ( 
.A1(n_403),
.A2(n_388),
.B(n_392),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_407),
.B(n_408),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g416 ( 
.A(n_409),
.B(n_412),
.Y(n_416)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_399),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_SL g414 ( 
.A(n_410),
.B(n_411),
.Y(n_414)
);

OAI21xp5_ASAP7_75t_L g411 ( 
.A1(n_404),
.A2(n_388),
.B(n_394),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_405),
.Y(n_412)
);

XOR2xp5_ASAP7_75t_L g413 ( 
.A(n_398),
.B(n_374),
.Y(n_413)
);

INVxp67_ASAP7_75t_L g418 ( 
.A(n_413),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_SL g417 ( 
.A1(n_409),
.A2(n_384),
.B1(n_373),
.B2(n_405),
.Y(n_417)
);

HB1xp67_ASAP7_75t_L g419 ( 
.A(n_417),
.Y(n_419)
);

NOR2xp67_ASAP7_75t_SL g420 ( 
.A(n_416),
.B(n_415),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_420),
.B(n_421),
.C(n_418),
.Y(n_423)
);

NAND2xp33_ASAP7_75t_R g421 ( 
.A(n_414),
.B(n_413),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_419),
.B(n_376),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_L g424 ( 
.A(n_422),
.B(n_423),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_424),
.B(n_418),
.Y(n_425)
);


endmodule