module fake_ariane_1886_n_1685 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_18, n_86, n_75, n_89, n_67, n_34, n_69, n_95, n_92, n_143, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_148, n_52, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_136, n_28, n_80, n_146, n_97, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_127, n_35, n_54, n_25, n_1685);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_34;
input n_69;
input n_95;
input n_92;
input n_143;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_52;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1685;

wire n_913;
wire n_1681;
wire n_1507;
wire n_1486;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_524;
wire n_634;
wire n_1214;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_1682;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_829;
wire n_1062;
wire n_339;
wire n_738;
wire n_672;
wire n_740;
wire n_1283;
wire n_167;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_495;
wire n_267;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_206;
wire n_899;
wire n_611;
wire n_1295;
wire n_238;
wire n_365;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1597;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_149;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_209;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1594;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_150;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_824;
wire n_428;
wire n_159;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_155;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_162;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1163;
wire n_186;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_158;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1304;
wire n_1608;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_545;
wire n_1015;
wire n_1614;
wire n_1162;
wire n_536;
wire n_1377;
wire n_325;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_163;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_321;
wire n_221;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_710;
wire n_534;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1572;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_769;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_430;
wire n_1206;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_521;
wire n_873;
wire n_1301;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_157;
wire n_1161;
wire n_811;
wire n_624;
wire n_876;
wire n_791;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_151;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_154;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_152;
wire n_169;
wire n_1288;
wire n_1201;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_166;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_168;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_683;
wire n_601;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_284;
wire n_593;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_820;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_161;
wire n_532;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_164;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_1536;
wire n_1471;
wire n_160;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_443;
wire n_1412;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1093;
wire n_1551;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_153;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_709;
wire n_809;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_896;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1670;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_156;
wire n_174;
wire n_275;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1313;
wire n_1001;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_165;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1233;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g149 ( 
.A(n_73),
.Y(n_149)
);

CKINVDCx5p33_ASAP7_75t_R g150 ( 
.A(n_135),
.Y(n_150)
);

CKINVDCx5p33_ASAP7_75t_R g151 ( 
.A(n_72),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_117),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_40),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_96),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_58),
.Y(n_155)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_58),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_123),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_23),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_66),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_16),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_74),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_114),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_69),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_29),
.Y(n_164)
);

BUFx3_ASAP7_75t_L g165 ( 
.A(n_147),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_16),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_137),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_44),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_111),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_62),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_134),
.Y(n_171)
);

BUFx10_ASAP7_75t_L g172 ( 
.A(n_146),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_46),
.Y(n_173)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_98),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_97),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_119),
.Y(n_176)
);

BUFx2_ASAP7_75t_L g177 ( 
.A(n_143),
.Y(n_177)
);

BUFx2_ASAP7_75t_L g178 ( 
.A(n_26),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_19),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_46),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_129),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_89),
.Y(n_182)
);

BUFx3_ASAP7_75t_L g183 ( 
.A(n_51),
.Y(n_183)
);

BUFx8_ASAP7_75t_SL g184 ( 
.A(n_115),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_118),
.Y(n_185)
);

BUFx5_ASAP7_75t_L g186 ( 
.A(n_145),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_107),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_100),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_40),
.Y(n_189)
);

BUFx3_ASAP7_75t_L g190 ( 
.A(n_103),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_104),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_64),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_22),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_63),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_101),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_108),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_24),
.Y(n_197)
);

INVx1_ASAP7_75t_SL g198 ( 
.A(n_148),
.Y(n_198)
);

BUFx10_ASAP7_75t_L g199 ( 
.A(n_21),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_124),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_90),
.Y(n_201)
);

BUFx2_ASAP7_75t_SL g202 ( 
.A(n_133),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_49),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_20),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_99),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_22),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_1),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_32),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_93),
.Y(n_209)
);

CKINVDCx14_ASAP7_75t_R g210 ( 
.A(n_79),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_10),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_81),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_50),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_0),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_35),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_139),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_32),
.Y(n_217)
);

INVx2_ASAP7_75t_SL g218 ( 
.A(n_142),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_8),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_67),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_3),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_80),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_52),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_77),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_1),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_41),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_12),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_49),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_94),
.Y(n_229)
);

INVx2_ASAP7_75t_SL g230 ( 
.A(n_6),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_50),
.Y(n_231)
);

BUFx10_ASAP7_75t_L g232 ( 
.A(n_127),
.Y(n_232)
);

BUFx2_ASAP7_75t_L g233 ( 
.A(n_30),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_8),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_109),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_43),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_113),
.Y(n_237)
);

BUFx2_ASAP7_75t_R g238 ( 
.A(n_43),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_29),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_83),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_14),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_130),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_84),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_59),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_128),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_2),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_138),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_12),
.Y(n_248)
);

BUFx10_ASAP7_75t_L g249 ( 
.A(n_54),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_54),
.Y(n_250)
);

BUFx2_ASAP7_75t_L g251 ( 
.A(n_27),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_37),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_26),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_36),
.Y(n_254)
);

INVx2_ASAP7_75t_SL g255 ( 
.A(n_60),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_4),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_132),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_57),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_48),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_0),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_136),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_63),
.Y(n_262)
);

INVx2_ASAP7_75t_SL g263 ( 
.A(n_144),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_41),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_62),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_17),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_75),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_33),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_85),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_10),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_6),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_106),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_11),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_17),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_11),
.Y(n_275)
);

INVx1_ASAP7_75t_SL g276 ( 
.A(n_25),
.Y(n_276)
);

BUFx10_ASAP7_75t_L g277 ( 
.A(n_86),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_42),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_45),
.Y(n_279)
);

INVx2_ASAP7_75t_SL g280 ( 
.A(n_3),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_141),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_87),
.Y(n_282)
);

INVx1_ASAP7_75t_SL g283 ( 
.A(n_9),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_24),
.Y(n_284)
);

CKINVDCx16_ASAP7_75t_R g285 ( 
.A(n_44),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_91),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_9),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_39),
.Y(n_288)
);

BUFx3_ASAP7_75t_L g289 ( 
.A(n_60),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_59),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_110),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_51),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_56),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_20),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_55),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_122),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_42),
.Y(n_297)
);

INVx1_ASAP7_75t_SL g298 ( 
.A(n_45),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_177),
.B(n_2),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_184),
.Y(n_300)
);

HB1xp67_ASAP7_75t_L g301 ( 
.A(n_178),
.Y(n_301)
);

INVxp33_ASAP7_75t_SL g302 ( 
.A(n_178),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_177),
.B(n_4),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_159),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_163),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_159),
.Y(n_306)
);

BUFx2_ASAP7_75t_L g307 ( 
.A(n_233),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_169),
.Y(n_308)
);

CKINVDCx16_ASAP7_75t_R g309 ( 
.A(n_217),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_285),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_182),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_176),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_182),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_188),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_188),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_191),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_222),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_191),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_153),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_192),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_217),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_238),
.B(n_5),
.Y(n_322)
);

HB1xp67_ASAP7_75t_L g323 ( 
.A(n_233),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_158),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_192),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_155),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_160),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_195),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_164),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_195),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_220),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_220),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_229),
.B(n_5),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_229),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_245),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_245),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_247),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_197),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_247),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_261),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_261),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_281),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_R g343 ( 
.A(n_210),
.B(n_102),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_281),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_282),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_166),
.Y(n_346)
);

INVxp67_ASAP7_75t_L g347 ( 
.A(n_251),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_282),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_286),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_286),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_296),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_296),
.Y(n_352)
);

HB1xp67_ASAP7_75t_L g353 ( 
.A(n_251),
.Y(n_353)
);

INVxp67_ASAP7_75t_L g354 ( 
.A(n_170),
.Y(n_354)
);

INVxp67_ASAP7_75t_L g355 ( 
.A(n_170),
.Y(n_355)
);

CKINVDCx14_ASAP7_75t_R g356 ( 
.A(n_172),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_253),
.Y(n_357)
);

CKINVDCx16_ASAP7_75t_R g358 ( 
.A(n_172),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_168),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_253),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_253),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_179),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_215),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_241),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_189),
.Y(n_365)
);

CKINVDCx16_ASAP7_75t_R g366 ( 
.A(n_199),
.Y(n_366)
);

HB1xp67_ASAP7_75t_L g367 ( 
.A(n_183),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_204),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_253),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_207),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_230),
.B(n_255),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_253),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_180),
.Y(n_373)
);

INVxp67_ASAP7_75t_L g374 ( 
.A(n_180),
.Y(n_374)
);

AND2x2_ASAP7_75t_L g375 ( 
.A(n_304),
.B(n_183),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_361),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_304),
.B(n_218),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_357),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_306),
.B(n_218),
.Y(n_379)
);

XOR2xp5_ASAP7_75t_L g380 ( 
.A(n_322),
.B(n_259),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_357),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_361),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_360),
.Y(n_383)
);

INVx3_ASAP7_75t_L g384 ( 
.A(n_360),
.Y(n_384)
);

INVx4_ASAP7_75t_L g385 ( 
.A(n_306),
.Y(n_385)
);

AND2x2_ASAP7_75t_L g386 ( 
.A(n_311),
.B(n_289),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_369),
.Y(n_387)
);

BUFx2_ASAP7_75t_L g388 ( 
.A(n_321),
.Y(n_388)
);

AND2x2_ASAP7_75t_L g389 ( 
.A(n_311),
.B(n_289),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_371),
.B(n_263),
.Y(n_390)
);

BUFx6f_ASAP7_75t_L g391 ( 
.A(n_369),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_SL g392 ( 
.A(n_343),
.B(n_172),
.Y(n_392)
);

NOR2x1_ASAP7_75t_L g393 ( 
.A(n_313),
.B(n_165),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_372),
.Y(n_394)
);

INVx4_ASAP7_75t_L g395 ( 
.A(n_313),
.Y(n_395)
);

INVx3_ASAP7_75t_L g396 ( 
.A(n_372),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_314),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_314),
.Y(n_398)
);

BUFx6f_ASAP7_75t_L g399 ( 
.A(n_315),
.Y(n_399)
);

AND2x4_ASAP7_75t_L g400 ( 
.A(n_315),
.B(n_230),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_316),
.Y(n_401)
);

BUFx6f_ASAP7_75t_L g402 ( 
.A(n_316),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_318),
.B(n_263),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_318),
.Y(n_404)
);

BUFx8_ASAP7_75t_L g405 ( 
.A(n_307),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_320),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_320),
.Y(n_407)
);

INVx4_ASAP7_75t_L g408 ( 
.A(n_325),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_325),
.B(n_198),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_328),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_328),
.Y(n_411)
);

BUFx6f_ASAP7_75t_L g412 ( 
.A(n_330),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_SL g413 ( 
.A(n_358),
.B(n_172),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_SL g414 ( 
.A(n_358),
.B(n_232),
.Y(n_414)
);

BUFx6f_ASAP7_75t_L g415 ( 
.A(n_330),
.Y(n_415)
);

BUFx2_ASAP7_75t_L g416 ( 
.A(n_310),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_331),
.Y(n_417)
);

INVx4_ASAP7_75t_L g418 ( 
.A(n_331),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_332),
.B(n_149),
.Y(n_419)
);

INVx4_ASAP7_75t_L g420 ( 
.A(n_332),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_334),
.Y(n_421)
);

NAND2xp33_ASAP7_75t_L g422 ( 
.A(n_334),
.B(n_186),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_SL g423 ( 
.A1(n_322),
.A2(n_294),
.B1(n_270),
.B2(n_283),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_335),
.B(n_150),
.Y(n_424)
);

AND2x2_ASAP7_75t_L g425 ( 
.A(n_335),
.B(n_156),
.Y(n_425)
);

INVx3_ASAP7_75t_L g426 ( 
.A(n_336),
.Y(n_426)
);

INVx5_ASAP7_75t_L g427 ( 
.A(n_366),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_299),
.B(n_232),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_336),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_SL g430 ( 
.A1(n_319),
.A2(n_298),
.B1(n_276),
.B2(n_295),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_302),
.B(n_174),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_337),
.Y(n_432)
);

AND2x4_ASAP7_75t_L g433 ( 
.A(n_337),
.B(n_255),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_339),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_339),
.B(n_151),
.Y(n_435)
);

BUFx6f_ASAP7_75t_L g436 ( 
.A(n_340),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_340),
.B(n_152),
.Y(n_437)
);

BUFx6f_ASAP7_75t_L g438 ( 
.A(n_341),
.Y(n_438)
);

BUFx8_ASAP7_75t_L g439 ( 
.A(n_307),
.Y(n_439)
);

BUFx6f_ASAP7_75t_L g440 ( 
.A(n_341),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_342),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_342),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_344),
.B(n_154),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_428),
.B(n_356),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_399),
.Y(n_445)
);

BUFx6f_ASAP7_75t_SL g446 ( 
.A(n_400),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_399),
.Y(n_447)
);

INVx3_ASAP7_75t_L g448 ( 
.A(n_399),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_399),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_384),
.Y(n_450)
);

NAND3xp33_ASAP7_75t_L g451 ( 
.A(n_390),
.B(n_333),
.C(n_303),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_399),
.Y(n_452)
);

INVx4_ASAP7_75t_L g453 ( 
.A(n_399),
.Y(n_453)
);

NAND3xp33_ASAP7_75t_L g454 ( 
.A(n_390),
.B(n_345),
.C(n_344),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_384),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_384),
.Y(n_456)
);

AND2x4_ASAP7_75t_L g457 ( 
.A(n_400),
.B(n_354),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_384),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g459 ( 
.A(n_427),
.B(n_324),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_399),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_419),
.B(n_345),
.Y(n_461)
);

HB1xp67_ASAP7_75t_L g462 ( 
.A(n_416),
.Y(n_462)
);

AND2x6_ASAP7_75t_L g463 ( 
.A(n_400),
.B(n_174),
.Y(n_463)
);

NAND2xp33_ASAP7_75t_L g464 ( 
.A(n_427),
.B(n_327),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_402),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_SL g466 ( 
.A(n_427),
.B(n_329),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_428),
.B(n_346),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_384),
.Y(n_468)
);

INVx4_ASAP7_75t_L g469 ( 
.A(n_402),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_396),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_SL g471 ( 
.A(n_427),
.B(n_359),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_402),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_392),
.B(n_362),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_419),
.B(n_424),
.Y(n_474)
);

BUFx6f_ASAP7_75t_L g475 ( 
.A(n_402),
.Y(n_475)
);

INVx2_ASAP7_75t_SL g476 ( 
.A(n_427),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_392),
.B(n_365),
.Y(n_477)
);

INVx5_ASAP7_75t_L g478 ( 
.A(n_402),
.Y(n_478)
);

INVx4_ASAP7_75t_L g479 ( 
.A(n_402),
.Y(n_479)
);

AND2x4_ASAP7_75t_L g480 ( 
.A(n_400),
.B(n_355),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_424),
.B(n_348),
.Y(n_481)
);

AOI22xp5_ASAP7_75t_L g482 ( 
.A1(n_431),
.A2(n_280),
.B1(n_227),
.B2(n_173),
.Y(n_482)
);

BUFx6f_ASAP7_75t_L g483 ( 
.A(n_402),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_SL g484 ( 
.A(n_427),
.B(n_368),
.Y(n_484)
);

AND2x2_ASAP7_75t_L g485 ( 
.A(n_425),
.B(n_373),
.Y(n_485)
);

OAI22xp33_ASAP7_75t_L g486 ( 
.A1(n_431),
.A2(n_309),
.B1(n_347),
.B2(n_409),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_396),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_412),
.Y(n_488)
);

OR2x2_ASAP7_75t_L g489 ( 
.A(n_416),
.B(n_309),
.Y(n_489)
);

AND2x2_ASAP7_75t_L g490 ( 
.A(n_425),
.B(n_373),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_413),
.B(n_370),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_396),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_412),
.Y(n_493)
);

NAND2xp33_ASAP7_75t_L g494 ( 
.A(n_427),
.B(n_300),
.Y(n_494)
);

INVx3_ASAP7_75t_L g495 ( 
.A(n_412),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_413),
.B(n_301),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_396),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_412),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_412),
.Y(n_499)
);

INVx3_ASAP7_75t_L g500 ( 
.A(n_412),
.Y(n_500)
);

INVx2_ASAP7_75t_SL g501 ( 
.A(n_427),
.Y(n_501)
);

AOI22xp33_ASAP7_75t_L g502 ( 
.A1(n_400),
.A2(n_323),
.B1(n_353),
.B2(n_350),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_412),
.Y(n_503)
);

INVxp33_ASAP7_75t_L g504 ( 
.A(n_380),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_396),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_414),
.B(n_348),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_415),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_387),
.Y(n_508)
);

INVxp33_ASAP7_75t_L g509 ( 
.A(n_380),
.Y(n_509)
);

AOI22xp33_ASAP7_75t_L g510 ( 
.A1(n_433),
.A2(n_352),
.B1(n_351),
.B2(n_350),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_415),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_387),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_414),
.B(n_349),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_387),
.Y(n_514)
);

AOI22xp33_ASAP7_75t_L g515 ( 
.A1(n_433),
.A2(n_280),
.B1(n_213),
.B2(n_156),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_415),
.Y(n_516)
);

BUFx6f_ASAP7_75t_SL g517 ( 
.A(n_433),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_435),
.B(n_374),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_376),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_376),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_SL g521 ( 
.A(n_409),
.B(n_312),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_376),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_382),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_415),
.Y(n_524)
);

NAND2xp33_ASAP7_75t_L g525 ( 
.A(n_435),
.B(n_157),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_382),
.Y(n_526)
);

AND2x4_ASAP7_75t_L g527 ( 
.A(n_433),
.B(n_367),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_382),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_415),
.Y(n_529)
);

INVx2_ASAP7_75t_SL g530 ( 
.A(n_375),
.Y(n_530)
);

CKINVDCx20_ASAP7_75t_R g531 ( 
.A(n_405),
.Y(n_531)
);

OR2x6_ASAP7_75t_L g532 ( 
.A(n_425),
.B(n_213),
.Y(n_532)
);

BUFx3_ASAP7_75t_L g533 ( 
.A(n_426),
.Y(n_533)
);

BUFx10_ASAP7_75t_L g534 ( 
.A(n_397),
.Y(n_534)
);

INVx5_ASAP7_75t_L g535 ( 
.A(n_415),
.Y(n_535)
);

INVx3_ASAP7_75t_L g536 ( 
.A(n_415),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_437),
.B(n_161),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_437),
.B(n_162),
.Y(n_538)
);

OR2x2_ASAP7_75t_L g539 ( 
.A(n_388),
.B(n_317),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_L g540 ( 
.A(n_443),
.B(n_305),
.Y(n_540)
);

BUFx6f_ASAP7_75t_SL g541 ( 
.A(n_405),
.Y(n_541)
);

INVx2_ASAP7_75t_SL g542 ( 
.A(n_375),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_443),
.B(n_167),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_436),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_385),
.B(n_171),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_385),
.B(n_175),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_436),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_436),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_SL g549 ( 
.A(n_388),
.B(n_385),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_SL g550 ( 
.A(n_388),
.B(n_199),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_385),
.B(n_185),
.Y(n_551)
);

INVx3_ASAP7_75t_L g552 ( 
.A(n_436),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_L g553 ( 
.A(n_385),
.B(n_308),
.Y(n_553)
);

BUFx3_ASAP7_75t_L g554 ( 
.A(n_426),
.Y(n_554)
);

OAI22xp5_ASAP7_75t_L g555 ( 
.A1(n_377),
.A2(n_246),
.B1(n_228),
.B2(n_226),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_436),
.Y(n_556)
);

AND2x2_ASAP7_75t_L g557 ( 
.A(n_386),
.B(n_199),
.Y(n_557)
);

AOI22xp5_ASAP7_75t_L g558 ( 
.A1(n_430),
.A2(n_208),
.B1(n_214),
.B2(n_211),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_436),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_436),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_438),
.Y(n_561)
);

NAND3xp33_ASAP7_75t_L g562 ( 
.A(n_395),
.B(n_248),
.C(n_297),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_438),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_SL g564 ( 
.A(n_395),
.B(n_199),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_438),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_438),
.Y(n_566)
);

HB1xp67_ASAP7_75t_L g567 ( 
.A(n_405),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_438),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_438),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_438),
.Y(n_570)
);

OR2x2_ASAP7_75t_L g571 ( 
.A(n_386),
.B(n_193),
.Y(n_571)
);

INVxp33_ASAP7_75t_L g572 ( 
.A(n_423),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_SL g573 ( 
.A(n_395),
.B(n_249),
.Y(n_573)
);

OR2x2_ASAP7_75t_L g574 ( 
.A(n_386),
.B(n_193),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_395),
.B(n_187),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_395),
.B(n_196),
.Y(n_576)
);

BUFx6f_ASAP7_75t_L g577 ( 
.A(n_440),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_440),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_440),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_405),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_440),
.Y(n_581)
);

OR2x6_ASAP7_75t_L g582 ( 
.A(n_389),
.B(n_430),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_440),
.Y(n_583)
);

BUFx2_ASAP7_75t_L g584 ( 
.A(n_405),
.Y(n_584)
);

INVx4_ASAP7_75t_L g585 ( 
.A(n_440),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_SL g586 ( 
.A(n_408),
.B(n_249),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_440),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_391),
.Y(n_588)
);

AND2x2_ASAP7_75t_L g589 ( 
.A(n_389),
.B(n_249),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_408),
.B(n_200),
.Y(n_590)
);

NOR3xp33_ASAP7_75t_L g591 ( 
.A(n_451),
.B(n_423),
.C(n_203),
.Y(n_591)
);

A2O1A1Ixp33_ASAP7_75t_L g592 ( 
.A1(n_506),
.A2(n_426),
.B(n_406),
.C(n_434),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_SL g593 ( 
.A(n_467),
.B(n_408),
.Y(n_593)
);

OAI22xp5_ASAP7_75t_L g594 ( 
.A1(n_451),
.A2(n_408),
.B1(n_418),
.B2(n_420),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_513),
.B(n_408),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_474),
.B(n_418),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_508),
.Y(n_597)
);

NOR2xp33_ASAP7_75t_L g598 ( 
.A(n_491),
.B(n_439),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_518),
.B(n_418),
.Y(n_599)
);

A2O1A1Ixp33_ASAP7_75t_L g600 ( 
.A1(n_473),
.A2(n_426),
.B(n_406),
.C(n_434),
.Y(n_600)
);

NAND2xp33_ASAP7_75t_L g601 ( 
.A(n_475),
.B(n_483),
.Y(n_601)
);

INVx2_ASAP7_75t_SL g602 ( 
.A(n_534),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_508),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_461),
.B(n_418),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_580),
.Y(n_605)
);

NOR2xp33_ASAP7_75t_L g606 ( 
.A(n_477),
.B(n_439),
.Y(n_606)
);

NAND2xp33_ASAP7_75t_L g607 ( 
.A(n_475),
.B(n_426),
.Y(n_607)
);

AOI221xp5_ASAP7_75t_L g608 ( 
.A1(n_486),
.A2(n_231),
.B1(n_236),
.B2(n_221),
.C(n_219),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_512),
.Y(n_609)
);

INVx2_ASAP7_75t_SL g610 ( 
.A(n_534),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_512),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_514),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_481),
.B(n_418),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_528),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_444),
.B(n_420),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_454),
.B(n_420),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_528),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_454),
.B(n_420),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_519),
.Y(n_619)
);

AOI21xp5_ASAP7_75t_L g620 ( 
.A1(n_545),
.A2(n_551),
.B(n_546),
.Y(n_620)
);

BUFx3_ASAP7_75t_L g621 ( 
.A(n_533),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_557),
.B(n_589),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_SL g623 ( 
.A(n_541),
.B(n_439),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_L g624 ( 
.A(n_521),
.B(n_439),
.Y(n_624)
);

INVx2_ASAP7_75t_SL g625 ( 
.A(n_534),
.Y(n_625)
);

AOI221xp5_ASAP7_75t_L g626 ( 
.A1(n_482),
.A2(n_231),
.B1(n_221),
.B2(n_219),
.C(n_236),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_557),
.B(n_589),
.Y(n_627)
);

INVx3_ASAP7_75t_L g628 ( 
.A(n_533),
.Y(n_628)
);

NAND2xp33_ASAP7_75t_L g629 ( 
.A(n_475),
.B(n_397),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_520),
.Y(n_630)
);

OAI221xp5_ASAP7_75t_L g631 ( 
.A1(n_482),
.A2(n_278),
.B1(n_206),
.B2(n_203),
.C(n_194),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_SL g632 ( 
.A(n_534),
.B(n_420),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_530),
.B(n_398),
.Y(n_633)
);

HB1xp67_ASAP7_75t_L g634 ( 
.A(n_462),
.Y(n_634)
);

OAI22xp5_ASAP7_75t_L g635 ( 
.A1(n_530),
.A2(n_442),
.B1(n_398),
.B2(n_401),
.Y(n_635)
);

NAND2xp33_ASAP7_75t_L g636 ( 
.A(n_475),
.B(n_401),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_542),
.B(n_407),
.Y(n_637)
);

NOR3xp33_ASAP7_75t_L g638 ( 
.A(n_553),
.B(n_206),
.C(n_194),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_542),
.B(n_407),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_520),
.Y(n_640)
);

NOR2xp33_ASAP7_75t_L g641 ( 
.A(n_496),
.B(n_439),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_522),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_SL g643 ( 
.A(n_457),
.B(n_379),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_522),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_485),
.B(n_410),
.Y(n_645)
);

AOI22xp33_ASAP7_75t_L g646 ( 
.A1(n_582),
.A2(n_393),
.B1(n_422),
.B2(n_403),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_523),
.Y(n_647)
);

AND2x4_ASAP7_75t_L g648 ( 
.A(n_532),
.B(n_584),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_L g649 ( 
.A(n_540),
.B(n_326),
.Y(n_649)
);

HB1xp67_ASAP7_75t_L g650 ( 
.A(n_489),
.Y(n_650)
);

AOI22xp5_ASAP7_75t_L g651 ( 
.A1(n_446),
.A2(n_422),
.B1(n_379),
.B2(n_403),
.Y(n_651)
);

NOR2xp33_ASAP7_75t_L g652 ( 
.A(n_549),
.B(n_338),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_514),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_523),
.Y(n_654)
);

AND2x4_ASAP7_75t_L g655 ( 
.A(n_532),
.B(n_417),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_526),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_490),
.B(n_417),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_526),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_SL g659 ( 
.A(n_457),
.B(n_429),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_487),
.Y(n_660)
);

BUFx3_ASAP7_75t_L g661 ( 
.A(n_533),
.Y(n_661)
);

INVxp67_ASAP7_75t_L g662 ( 
.A(n_539),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_487),
.Y(n_663)
);

HB1xp67_ASAP7_75t_L g664 ( 
.A(n_539),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_510),
.B(n_442),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_457),
.B(n_404),
.Y(n_666)
);

NOR3xp33_ASAP7_75t_L g667 ( 
.A(n_550),
.B(n_244),
.C(n_297),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_554),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_SL g669 ( 
.A(n_457),
.B(n_441),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_480),
.B(n_537),
.Y(n_670)
);

AOI22xp33_ASAP7_75t_L g671 ( 
.A1(n_582),
.A2(n_393),
.B1(n_432),
.B2(n_421),
.Y(n_671)
);

INVx3_ASAP7_75t_L g672 ( 
.A(n_554),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_554),
.Y(n_673)
);

INVxp67_ASAP7_75t_L g674 ( 
.A(n_527),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_487),
.Y(n_675)
);

INVxp67_ASAP7_75t_L g676 ( 
.A(n_527),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_580),
.Y(n_677)
);

NAND2xp33_ASAP7_75t_L g678 ( 
.A(n_475),
.B(n_483),
.Y(n_678)
);

NOR2xp33_ASAP7_75t_L g679 ( 
.A(n_538),
.B(n_363),
.Y(n_679)
);

NOR2xp33_ASAP7_75t_L g680 ( 
.A(n_543),
.B(n_364),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_450),
.Y(n_681)
);

AOI22xp5_ASAP7_75t_L g682 ( 
.A1(n_446),
.A2(n_517),
.B1(n_463),
.B2(n_532),
.Y(n_682)
);

INVx2_ASAP7_75t_SL g683 ( 
.A(n_480),
.Y(n_683)
);

BUFx6f_ASAP7_75t_L g684 ( 
.A(n_483),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_480),
.B(n_411),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_492),
.Y(n_686)
);

NOR2xp33_ASAP7_75t_L g687 ( 
.A(n_564),
.B(n_411),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_SL g688 ( 
.A(n_527),
.B(n_441),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_492),
.Y(n_689)
);

O2A1O1Ixp33_ASAP7_75t_L g690 ( 
.A1(n_555),
.A2(n_574),
.B(n_571),
.C(n_573),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_532),
.B(n_421),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_492),
.Y(n_692)
);

AND2x6_ASAP7_75t_L g693 ( 
.A(n_497),
.B(n_421),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_532),
.B(n_432),
.Y(n_694)
);

AOI22xp33_ASAP7_75t_L g695 ( 
.A1(n_582),
.A2(n_441),
.B1(n_432),
.B2(n_277),
.Y(n_695)
);

NOR2xp33_ASAP7_75t_SL g696 ( 
.A(n_541),
.B(n_232),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_497),
.Y(n_697)
);

OAI221xp5_ASAP7_75t_L g698 ( 
.A1(n_515),
.A2(n_502),
.B1(n_558),
.B2(n_571),
.C(n_574),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_497),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_SL g700 ( 
.A(n_476),
.B(n_249),
.Y(n_700)
);

AND2x2_ASAP7_75t_L g701 ( 
.A(n_582),
.B(n_244),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_455),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_455),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_SL g704 ( 
.A(n_476),
.B(n_501),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_SL g705 ( 
.A(n_501),
.B(n_223),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_456),
.Y(n_706)
);

HB1xp67_ASAP7_75t_L g707 ( 
.A(n_446),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_SL g708 ( 
.A(n_586),
.B(n_225),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_456),
.Y(n_709)
);

INVx2_ASAP7_75t_SL g710 ( 
.A(n_463),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_463),
.B(n_378),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_458),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_SL g713 ( 
.A(n_584),
.B(n_234),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_458),
.Y(n_714)
);

NOR2xp33_ASAP7_75t_L g715 ( 
.A(n_517),
.B(n_239),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_463),
.B(n_378),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_463),
.B(n_381),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_463),
.B(n_381),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_468),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_463),
.B(n_383),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_468),
.B(n_383),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_470),
.B(n_394),
.Y(n_722)
);

O2A1O1Ixp33_ASAP7_75t_L g723 ( 
.A1(n_525),
.A2(n_271),
.B(n_295),
.C(n_290),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_470),
.Y(n_724)
);

BUFx8_ASAP7_75t_L g725 ( 
.A(n_541),
.Y(n_725)
);

NOR2xp33_ASAP7_75t_L g726 ( 
.A(n_517),
.B(n_252),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_505),
.B(n_394),
.Y(n_727)
);

AOI22xp5_ASAP7_75t_L g728 ( 
.A1(n_464),
.A2(n_202),
.B1(n_242),
.B2(n_243),
.Y(n_728)
);

AND2x2_ASAP7_75t_L g729 ( 
.A(n_582),
.B(n_248),
.Y(n_729)
);

NAND2xp33_ASAP7_75t_L g730 ( 
.A(n_483),
.B(n_186),
.Y(n_730)
);

AO22x2_ASAP7_75t_L g731 ( 
.A1(n_572),
.A2(n_266),
.B1(n_290),
.B2(n_278),
.Y(n_731)
);

NOR3xp33_ASAP7_75t_L g732 ( 
.A(n_562),
.B(n_274),
.C(n_273),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_SL g733 ( 
.A(n_575),
.B(n_254),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_505),
.Y(n_734)
);

INVx2_ASAP7_75t_SL g735 ( 
.A(n_448),
.Y(n_735)
);

NOR2xp33_ASAP7_75t_SL g736 ( 
.A(n_567),
.B(n_232),
.Y(n_736)
);

INVx2_ASAP7_75t_SL g737 ( 
.A(n_448),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_576),
.B(n_590),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_529),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_448),
.B(n_495),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_448),
.B(n_250),
.Y(n_741)
);

OAI22xp5_ASAP7_75t_SL g742 ( 
.A1(n_531),
.A2(n_275),
.B1(n_256),
.B2(n_293),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_445),
.Y(n_743)
);

AOI22xp5_ASAP7_75t_L g744 ( 
.A1(n_494),
.A2(n_202),
.B1(n_205),
.B2(n_291),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_558),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_495),
.B(n_250),
.Y(n_746)
);

AND2x4_ASAP7_75t_L g747 ( 
.A(n_562),
.B(n_266),
.Y(n_747)
);

AOI22xp5_ASAP7_75t_L g748 ( 
.A1(n_459),
.A2(n_209),
.B1(n_212),
.B2(n_201),
.Y(n_748)
);

BUFx6f_ASAP7_75t_L g749 ( 
.A(n_483),
.Y(n_749)
);

AOI22xp33_ASAP7_75t_L g750 ( 
.A1(n_529),
.A2(n_569),
.B1(n_587),
.B2(n_570),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_445),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_SL g752 ( 
.A(n_577),
.B(n_258),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_495),
.B(n_500),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_L g754 ( 
.A(n_641),
.B(n_453),
.Y(n_754)
);

AOI21xp5_ASAP7_75t_L g755 ( 
.A1(n_738),
.A2(n_471),
.B(n_466),
.Y(n_755)
);

AND2x4_ASAP7_75t_L g756 ( 
.A(n_683),
.B(n_453),
.Y(n_756)
);

INVx4_ASAP7_75t_L g757 ( 
.A(n_648),
.Y(n_757)
);

NOR2xp33_ASAP7_75t_L g758 ( 
.A(n_745),
.B(n_453),
.Y(n_758)
);

AOI21xp5_ASAP7_75t_L g759 ( 
.A1(n_620),
.A2(n_484),
.B(n_449),
.Y(n_759)
);

O2A1O1Ixp33_ASAP7_75t_L g760 ( 
.A1(n_670),
.A2(n_273),
.B(n_274),
.C(n_271),
.Y(n_760)
);

AOI21xp5_ASAP7_75t_L g761 ( 
.A1(n_740),
.A2(n_449),
.B(n_447),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_SL g762 ( 
.A(n_602),
.B(n_577),
.Y(n_762)
);

AOI21xp5_ASAP7_75t_L g763 ( 
.A1(n_753),
.A2(n_447),
.B(n_499),
.Y(n_763)
);

AOI21xp5_ASAP7_75t_L g764 ( 
.A1(n_596),
.A2(n_452),
.B(n_460),
.Y(n_764)
);

NOR2xp33_ASAP7_75t_SL g765 ( 
.A(n_598),
.B(n_504),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_622),
.B(n_495),
.Y(n_766)
);

INVx3_ASAP7_75t_L g767 ( 
.A(n_621),
.Y(n_767)
);

BUFx6f_ASAP7_75t_L g768 ( 
.A(n_684),
.Y(n_768)
);

AOI21xp5_ASAP7_75t_L g769 ( 
.A1(n_593),
.A2(n_452),
.B(n_460),
.Y(n_769)
);

NOR2xp33_ASAP7_75t_L g770 ( 
.A(n_745),
.B(n_453),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_614),
.Y(n_771)
);

AO21x1_ASAP7_75t_L g772 ( 
.A1(n_606),
.A2(n_479),
.B(n_469),
.Y(n_772)
);

AOI21xp5_ASAP7_75t_L g773 ( 
.A1(n_604),
.A2(n_548),
.B(n_472),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_627),
.B(n_500),
.Y(n_774)
);

AOI21xp5_ASAP7_75t_L g775 ( 
.A1(n_613),
.A2(n_548),
.B(n_472),
.Y(n_775)
);

BUFx2_ASAP7_75t_L g776 ( 
.A(n_634),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_617),
.Y(n_777)
);

AND2x4_ASAP7_75t_L g778 ( 
.A(n_683),
.B(n_469),
.Y(n_778)
);

AOI21xp5_ASAP7_75t_L g779 ( 
.A1(n_599),
.A2(n_465),
.B(n_499),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_SL g780 ( 
.A(n_602),
.B(n_577),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_617),
.Y(n_781)
);

NOR2x1_ASAP7_75t_R g782 ( 
.A(n_605),
.B(n_260),
.Y(n_782)
);

AOI21xp5_ASAP7_75t_L g783 ( 
.A1(n_595),
.A2(n_465),
.B(n_498),
.Y(n_783)
);

AOI21xp5_ASAP7_75t_L g784 ( 
.A1(n_615),
.A2(n_556),
.B(n_524),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_643),
.B(n_500),
.Y(n_785)
);

A2O1A1Ixp33_ASAP7_75t_L g786 ( 
.A1(n_690),
.A2(n_608),
.B(n_638),
.C(n_723),
.Y(n_786)
);

OAI22xp5_ASAP7_75t_L g787 ( 
.A1(n_610),
.A2(n_469),
.B1(n_479),
.B2(n_585),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_645),
.B(n_536),
.Y(n_788)
);

INVx2_ASAP7_75t_SL g789 ( 
.A(n_664),
.Y(n_789)
);

O2A1O1Ixp5_ASAP7_75t_L g790 ( 
.A1(n_733),
.A2(n_469),
.B(n_479),
.C(n_585),
.Y(n_790)
);

AOI21xp5_ASAP7_75t_L g791 ( 
.A1(n_632),
.A2(n_561),
.B(n_503),
.Y(n_791)
);

NOR2xp33_ASAP7_75t_R g792 ( 
.A(n_605),
.B(n_552),
.Y(n_792)
);

OAI321xp33_ASAP7_75t_L g793 ( 
.A1(n_631),
.A2(n_181),
.A3(n_216),
.B1(n_235),
.B2(n_511),
.C(n_579),
.Y(n_793)
);

AND2x6_ASAP7_75t_L g794 ( 
.A(n_648),
.B(n_559),
.Y(n_794)
);

CKINVDCx10_ASAP7_75t_R g795 ( 
.A(n_742),
.Y(n_795)
);

AOI21xp5_ASAP7_75t_L g796 ( 
.A1(n_675),
.A2(n_561),
.B(n_503),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_706),
.Y(n_797)
);

NAND2xp33_ASAP7_75t_L g798 ( 
.A(n_610),
.B(n_577),
.Y(n_798)
);

O2A1O1Ixp33_ASAP7_75t_L g799 ( 
.A1(n_662),
.A2(n_516),
.B(n_493),
.C(n_583),
.Y(n_799)
);

CKINVDCx8_ASAP7_75t_R g800 ( 
.A(n_677),
.Y(n_800)
);

A2O1A1Ixp33_ASAP7_75t_L g801 ( 
.A1(n_666),
.A2(n_552),
.B(n_559),
.C(n_563),
.Y(n_801)
);

OAI21xp5_ASAP7_75t_L g802 ( 
.A1(n_600),
.A2(n_493),
.B(n_556),
.Y(n_802)
);

AOI21xp5_ASAP7_75t_L g803 ( 
.A1(n_686),
.A2(n_524),
.B(n_511),
.Y(n_803)
);

O2A1O1Ixp33_ASAP7_75t_L g804 ( 
.A1(n_616),
.A2(n_560),
.B(n_507),
.C(n_583),
.Y(n_804)
);

AOI21xp5_ASAP7_75t_L g805 ( 
.A1(n_689),
.A2(n_488),
.B(n_498),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_SL g806 ( 
.A(n_625),
.B(n_577),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_657),
.B(n_552),
.Y(n_807)
);

BUFx4f_ASAP7_75t_L g808 ( 
.A(n_648),
.Y(n_808)
);

AND2x2_ASAP7_75t_L g809 ( 
.A(n_649),
.B(n_509),
.Y(n_809)
);

AOI22xp33_ASAP7_75t_L g810 ( 
.A1(n_591),
.A2(n_277),
.B1(n_587),
.B2(n_570),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_SL g811 ( 
.A(n_625),
.B(n_479),
.Y(n_811)
);

OAI22xp5_ASAP7_75t_L g812 ( 
.A1(n_674),
.A2(n_676),
.B1(n_621),
.B2(n_661),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_685),
.B(n_585),
.Y(n_813)
);

AOI21xp5_ASAP7_75t_L g814 ( 
.A1(n_735),
.A2(n_507),
.B(n_488),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_SL g815 ( 
.A(n_655),
.B(n_478),
.Y(n_815)
);

AOI21xp5_ASAP7_75t_L g816 ( 
.A1(n_735),
.A2(n_547),
.B(n_560),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_709),
.Y(n_817)
);

BUFx6f_ASAP7_75t_L g818 ( 
.A(n_684),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_709),
.Y(n_819)
);

AOI21xp5_ASAP7_75t_L g820 ( 
.A1(n_737),
.A2(n_547),
.B(n_516),
.Y(n_820)
);

NOR3xp33_ASAP7_75t_L g821 ( 
.A(n_679),
.B(n_268),
.C(n_264),
.Y(n_821)
);

OAI21x1_ASAP7_75t_L g822 ( 
.A1(n_619),
.A2(n_566),
.B(n_565),
.Y(n_822)
);

AOI21xp5_ASAP7_75t_L g823 ( 
.A1(n_737),
.A2(n_579),
.B(n_563),
.Y(n_823)
);

BUFx6f_ASAP7_75t_L g824 ( 
.A(n_684),
.Y(n_824)
);

AOI21xp5_ASAP7_75t_L g825 ( 
.A1(n_660),
.A2(n_566),
.B(n_568),
.Y(n_825)
);

AOI21xp5_ASAP7_75t_L g826 ( 
.A1(n_660),
.A2(n_566),
.B(n_568),
.Y(n_826)
);

A2O1A1Ixp33_ASAP7_75t_L g827 ( 
.A1(n_680),
.A2(n_568),
.B(n_565),
.C(n_578),
.Y(n_827)
);

AOI21x1_ASAP7_75t_L g828 ( 
.A1(n_704),
.A2(n_581),
.B(n_578),
.Y(n_828)
);

BUFx4f_ASAP7_75t_SL g829 ( 
.A(n_725),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_724),
.Y(n_830)
);

AOI21xp5_ASAP7_75t_L g831 ( 
.A1(n_663),
.A2(n_565),
.B(n_581),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_633),
.B(n_544),
.Y(n_832)
);

HB1xp67_ASAP7_75t_L g833 ( 
.A(n_650),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_637),
.B(n_588),
.Y(n_834)
);

OAI21xp5_ASAP7_75t_L g835 ( 
.A1(n_592),
.A2(n_588),
.B(n_535),
.Y(n_835)
);

OAI21xp5_ASAP7_75t_L g836 ( 
.A1(n_594),
.A2(n_588),
.B(n_535),
.Y(n_836)
);

NOR2xp33_ASAP7_75t_L g837 ( 
.A(n_698),
.B(n_478),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_639),
.B(n_478),
.Y(n_838)
);

HB1xp67_ASAP7_75t_L g839 ( 
.A(n_691),
.Y(n_839)
);

AO21x1_ASAP7_75t_L g840 ( 
.A1(n_635),
.A2(n_181),
.B(n_235),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_724),
.Y(n_841)
);

O2A1O1Ixp33_ASAP7_75t_L g842 ( 
.A1(n_618),
.A2(n_216),
.B(n_165),
.C(n_190),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_701),
.B(n_478),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_SL g844 ( 
.A(n_628),
.B(n_478),
.Y(n_844)
);

NOR2xp33_ASAP7_75t_L g845 ( 
.A(n_624),
.B(n_535),
.Y(n_845)
);

AOI21xp5_ASAP7_75t_L g846 ( 
.A1(n_692),
.A2(n_535),
.B(n_240),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_697),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_701),
.B(n_535),
.Y(n_848)
);

O2A1O1Ixp33_ASAP7_75t_L g849 ( 
.A1(n_659),
.A2(n_190),
.B(n_262),
.C(n_265),
.Y(n_849)
);

OAI21xp5_ASAP7_75t_L g850 ( 
.A1(n_697),
.A2(n_279),
.B(n_292),
.Y(n_850)
);

INVx11_ASAP7_75t_L g851 ( 
.A(n_725),
.Y(n_851)
);

NOR2xp33_ASAP7_75t_L g852 ( 
.A(n_652),
.B(n_284),
.Y(n_852)
);

AOI21xp5_ASAP7_75t_L g853 ( 
.A1(n_699),
.A2(n_257),
.B(n_237),
.Y(n_853)
);

HB1xp67_ASAP7_75t_SL g854 ( 
.A(n_725),
.Y(n_854)
);

A2O1A1Ixp33_ASAP7_75t_L g855 ( 
.A1(n_651),
.A2(n_288),
.B(n_287),
.C(n_391),
.Y(n_855)
);

NOR2xp33_ASAP7_75t_L g856 ( 
.A(n_736),
.B(n_729),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_729),
.B(n_267),
.Y(n_857)
);

AND2x2_ASAP7_75t_L g858 ( 
.A(n_677),
.B(n_277),
.Y(n_858)
);

A2O1A1Ixp33_ASAP7_75t_L g859 ( 
.A1(n_626),
.A2(n_391),
.B(n_224),
.C(n_272),
.Y(n_859)
);

NOR2xp33_ASAP7_75t_L g860 ( 
.A(n_688),
.B(n_7),
.Y(n_860)
);

INVx4_ASAP7_75t_L g861 ( 
.A(n_661),
.Y(n_861)
);

AND2x2_ASAP7_75t_L g862 ( 
.A(n_715),
.B(n_277),
.Y(n_862)
);

BUFx4f_ASAP7_75t_L g863 ( 
.A(n_747),
.Y(n_863)
);

AND2x6_ASAP7_75t_L g864 ( 
.A(n_682),
.B(n_224),
.Y(n_864)
);

HB1xp67_ASAP7_75t_L g865 ( 
.A(n_694),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_646),
.B(n_747),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_681),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_747),
.B(n_671),
.Y(n_868)
);

INVx3_ASAP7_75t_L g869 ( 
.A(n_628),
.Y(n_869)
);

BUFx12f_ASAP7_75t_L g870 ( 
.A(n_684),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_669),
.B(n_269),
.Y(n_871)
);

NAND2xp33_ASAP7_75t_L g872 ( 
.A(n_693),
.B(n_391),
.Y(n_872)
);

OAI21xp5_ASAP7_75t_L g873 ( 
.A1(n_702),
.A2(n_391),
.B(n_186),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_695),
.B(n_391),
.Y(n_874)
);

NOR2xp33_ASAP7_75t_L g875 ( 
.A(n_668),
.B(n_7),
.Y(n_875)
);

INVx3_ASAP7_75t_L g876 ( 
.A(n_628),
.Y(n_876)
);

AND2x2_ASAP7_75t_L g877 ( 
.A(n_726),
.B(n_391),
.Y(n_877)
);

NOR2xp33_ASAP7_75t_L g878 ( 
.A(n_673),
.B(n_13),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_702),
.Y(n_879)
);

INVx3_ASAP7_75t_L g880 ( 
.A(n_672),
.Y(n_880)
);

INVx2_ASAP7_75t_SL g881 ( 
.A(n_707),
.Y(n_881)
);

AOI21xp5_ASAP7_75t_L g882 ( 
.A1(n_703),
.A2(n_224),
.B(n_186),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_665),
.B(n_13),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_672),
.B(n_14),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_SL g885 ( 
.A(n_672),
.B(n_186),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_712),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_712),
.Y(n_887)
);

OAI21xp33_ASAP7_75t_L g888 ( 
.A1(n_732),
.A2(n_741),
.B(n_746),
.Y(n_888)
);

AND2x2_ASAP7_75t_L g889 ( 
.A(n_731),
.B(n_15),
.Y(n_889)
);

INVxp67_ASAP7_75t_L g890 ( 
.A(n_731),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_731),
.B(n_15),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_SL g892 ( 
.A(n_684),
.B(n_186),
.Y(n_892)
);

AO21x1_ASAP7_75t_L g893 ( 
.A1(n_601),
.A2(n_186),
.B(n_224),
.Y(n_893)
);

NOR2xp33_ASAP7_75t_L g894 ( 
.A(n_713),
.B(n_18),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_714),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_731),
.B(n_18),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_719),
.Y(n_897)
);

OAI22xp33_ASAP7_75t_L g898 ( 
.A1(n_623),
.A2(n_19),
.B1(n_21),
.B2(n_23),
.Y(n_898)
);

OAI21xp5_ASAP7_75t_L g899 ( 
.A1(n_734),
.A2(n_140),
.B(n_131),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_SL g900 ( 
.A(n_749),
.B(n_27),
.Y(n_900)
);

OAI21xp5_ASAP7_75t_L g901 ( 
.A1(n_743),
.A2(n_126),
.B(n_125),
.Y(n_901)
);

AOI21xp5_ASAP7_75t_L g902 ( 
.A1(n_601),
.A2(n_121),
.B(n_120),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_597),
.Y(n_903)
);

O2A1O1Ixp5_ASAP7_75t_L g904 ( 
.A1(n_752),
.A2(n_28),
.B(n_30),
.C(n_31),
.Y(n_904)
);

A2O1A1Ixp33_ASAP7_75t_L g905 ( 
.A1(n_687),
.A2(n_28),
.B(n_31),
.C(n_33),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_597),
.B(n_603),
.Y(n_906)
);

AOI22xp5_ASAP7_75t_L g907 ( 
.A1(n_667),
.A2(n_34),
.B1(n_35),
.B2(n_36),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_603),
.B(n_34),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_609),
.Y(n_909)
);

CKINVDCx10_ASAP7_75t_R g910 ( 
.A(n_696),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_SL g911 ( 
.A(n_749),
.B(n_710),
.Y(n_911)
);

BUFx2_ASAP7_75t_L g912 ( 
.A(n_693),
.Y(n_912)
);

AOI21xp5_ASAP7_75t_L g913 ( 
.A1(n_678),
.A2(n_68),
.B(n_112),
.Y(n_913)
);

NOR2xp33_ASAP7_75t_L g914 ( 
.A(n_708),
.B(n_37),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_609),
.B(n_38),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_611),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_611),
.B(n_38),
.Y(n_917)
);

OAI21xp5_ASAP7_75t_L g918 ( 
.A1(n_751),
.A2(n_70),
.B(n_105),
.Y(n_918)
);

AND2x2_ASAP7_75t_L g919 ( 
.A(n_833),
.B(n_612),
.Y(n_919)
);

AOI21xp5_ASAP7_75t_L g920 ( 
.A1(n_754),
.A2(n_678),
.B(n_607),
.Y(n_920)
);

AOI21xp5_ASAP7_75t_L g921 ( 
.A1(n_754),
.A2(n_607),
.B(n_636),
.Y(n_921)
);

BUFx3_ASAP7_75t_L g922 ( 
.A(n_800),
.Y(n_922)
);

AOI22x1_ASAP7_75t_L g923 ( 
.A1(n_755),
.A2(n_749),
.B1(n_739),
.B2(n_653),
.Y(n_923)
);

AND2x2_ASAP7_75t_L g924 ( 
.A(n_833),
.B(n_612),
.Y(n_924)
);

O2A1O1Ixp5_ASAP7_75t_SL g925 ( 
.A1(n_900),
.A2(n_705),
.B(n_700),
.C(n_653),
.Y(n_925)
);

AOI21xp5_ASAP7_75t_L g926 ( 
.A1(n_798),
.A2(n_629),
.B(n_636),
.Y(n_926)
);

BUFx5_ASAP7_75t_L g927 ( 
.A(n_870),
.Y(n_927)
);

BUFx3_ASAP7_75t_L g928 ( 
.A(n_776),
.Y(n_928)
);

OAI21xp33_ASAP7_75t_SL g929 ( 
.A1(n_914),
.A2(n_728),
.B(n_722),
.Y(n_929)
);

NOR2xp33_ASAP7_75t_L g930 ( 
.A(n_852),
.B(n_739),
.Y(n_930)
);

BUFx2_ASAP7_75t_L g931 ( 
.A(n_789),
.Y(n_931)
);

AOI21xp5_ASAP7_75t_L g932 ( 
.A1(n_872),
.A2(n_629),
.B(n_749),
.Y(n_932)
);

OAI22xp5_ASAP7_75t_L g933 ( 
.A1(n_786),
.A2(n_744),
.B1(n_721),
.B2(n_727),
.Y(n_933)
);

AOI21xp5_ASAP7_75t_L g934 ( 
.A1(n_759),
.A2(n_730),
.B(n_711),
.Y(n_934)
);

OAI22x1_ASAP7_75t_L g935 ( 
.A1(n_852),
.A2(n_658),
.B1(n_640),
.B2(n_642),
.Y(n_935)
);

OR2x2_ASAP7_75t_L g936 ( 
.A(n_809),
.B(n_656),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_758),
.B(n_658),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_758),
.B(n_630),
.Y(n_938)
);

NOR2xp33_ASAP7_75t_L g939 ( 
.A(n_770),
.B(n_748),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_770),
.B(n_640),
.Y(n_940)
);

OAI22xp5_ASAP7_75t_L g941 ( 
.A1(n_863),
.A2(n_720),
.B1(n_718),
.B2(n_717),
.Y(n_941)
);

INVx3_ASAP7_75t_L g942 ( 
.A(n_757),
.Y(n_942)
);

BUFx3_ASAP7_75t_L g943 ( 
.A(n_829),
.Y(n_943)
);

NOR2xp33_ASAP7_75t_L g944 ( 
.A(n_856),
.B(n_656),
.Y(n_944)
);

OR2x2_ASAP7_75t_L g945 ( 
.A(n_857),
.B(n_654),
.Y(n_945)
);

AOI222xp33_ASAP7_75t_L g946 ( 
.A1(n_889),
.A2(n_856),
.B1(n_863),
.B2(n_890),
.C1(n_896),
.C2(n_891),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_862),
.B(n_757),
.Y(n_947)
);

OAI21xp5_ASAP7_75t_L g948 ( 
.A1(n_801),
.A2(n_693),
.B(n_750),
.Y(n_948)
);

INVx3_ASAP7_75t_SL g949 ( 
.A(n_854),
.Y(n_949)
);

NOR2xp33_ASAP7_75t_L g950 ( 
.A(n_765),
.B(n_654),
.Y(n_950)
);

OAI22xp5_ASAP7_75t_L g951 ( 
.A1(n_866),
.A2(n_716),
.B1(n_644),
.B2(n_647),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_868),
.B(n_647),
.Y(n_952)
);

INVxp67_ASAP7_75t_L g953 ( 
.A(n_894),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_867),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_839),
.B(n_644),
.Y(n_955)
);

AOI21xp5_ASAP7_75t_L g956 ( 
.A1(n_845),
.A2(n_693),
.B(n_65),
.Y(n_956)
);

BUFx6f_ASAP7_75t_L g957 ( 
.A(n_808),
.Y(n_957)
);

CKINVDCx20_ASAP7_75t_R g958 ( 
.A(n_829),
.Y(n_958)
);

AOI21xp5_ASAP7_75t_L g959 ( 
.A1(n_784),
.A2(n_693),
.B(n_71),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_839),
.B(n_693),
.Y(n_960)
);

A2O1A1Ixp33_ASAP7_75t_L g961 ( 
.A1(n_837),
.A2(n_39),
.B(n_47),
.C(n_48),
.Y(n_961)
);

AOI21xp5_ASAP7_75t_L g962 ( 
.A1(n_783),
.A2(n_76),
.B(n_95),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_SL g963 ( 
.A(n_808),
.B(n_47),
.Y(n_963)
);

INVx2_ASAP7_75t_SL g964 ( 
.A(n_851),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_865),
.B(n_52),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_865),
.B(n_53),
.Y(n_966)
);

AND2x2_ASAP7_75t_L g967 ( 
.A(n_858),
.B(n_53),
.Y(n_967)
);

AOI21xp5_ASAP7_75t_L g968 ( 
.A1(n_836),
.A2(n_78),
.B(n_92),
.Y(n_968)
);

O2A1O1Ixp33_ASAP7_75t_L g969 ( 
.A1(n_821),
.A2(n_905),
.B(n_914),
.C(n_894),
.Y(n_969)
);

AOI21xp5_ASAP7_75t_L g970 ( 
.A1(n_764),
.A2(n_82),
.B(n_88),
.Y(n_970)
);

NOR2xp33_ASAP7_75t_L g971 ( 
.A(n_821),
.B(n_55),
.Y(n_971)
);

NOR3xp33_ASAP7_75t_L g972 ( 
.A(n_905),
.B(n_56),
.C(n_57),
.Y(n_972)
);

INVx4_ASAP7_75t_R g973 ( 
.A(n_881),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_837),
.B(n_61),
.Y(n_974)
);

OAI21xp33_ASAP7_75t_SL g975 ( 
.A1(n_901),
.A2(n_61),
.B(n_116),
.Y(n_975)
);

NOR2xp33_ASAP7_75t_L g976 ( 
.A(n_910),
.B(n_782),
.Y(n_976)
);

AOI21xp5_ASAP7_75t_L g977 ( 
.A1(n_834),
.A2(n_779),
.B(n_775),
.Y(n_977)
);

BUFx10_ASAP7_75t_L g978 ( 
.A(n_860),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_794),
.B(n_860),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_SL g980 ( 
.A(n_792),
.B(n_812),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_797),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_817),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_819),
.Y(n_983)
);

NOR2xp33_ASAP7_75t_R g984 ( 
.A(n_795),
.B(n_767),
.Y(n_984)
);

AO32x1_ASAP7_75t_L g985 ( 
.A1(n_877),
.A2(n_841),
.A3(n_830),
.B1(n_909),
.B2(n_903),
.Y(n_985)
);

AO32x1_ASAP7_75t_L g986 ( 
.A1(n_916),
.A2(n_847),
.A3(n_879),
.B1(n_886),
.B2(n_887),
.Y(n_986)
);

AOI21xp5_ASAP7_75t_L g987 ( 
.A1(n_773),
.A2(n_823),
.B(n_814),
.Y(n_987)
);

INVx6_ASAP7_75t_L g988 ( 
.A(n_861),
.Y(n_988)
);

INVx4_ASAP7_75t_L g989 ( 
.A(n_794),
.Y(n_989)
);

AND2x4_ASAP7_75t_L g990 ( 
.A(n_794),
.B(n_815),
.Y(n_990)
);

NOR3xp33_ASAP7_75t_L g991 ( 
.A(n_898),
.B(n_900),
.C(n_850),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_766),
.B(n_774),
.Y(n_992)
);

OAI22xp5_ASAP7_75t_L g993 ( 
.A1(n_883),
.A2(n_907),
.B1(n_875),
.B2(n_878),
.Y(n_993)
);

AND2x4_ASAP7_75t_L g994 ( 
.A(n_794),
.B(n_815),
.Y(n_994)
);

AOI21xp5_ASAP7_75t_L g995 ( 
.A1(n_816),
.A2(n_820),
.B(n_761),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_792),
.B(n_810),
.Y(n_996)
);

NOR2xp67_ASAP7_75t_L g997 ( 
.A(n_861),
.B(n_767),
.Y(n_997)
);

INVx4_ASAP7_75t_L g998 ( 
.A(n_768),
.Y(n_998)
);

AOI22xp33_ASAP7_75t_L g999 ( 
.A1(n_810),
.A2(n_864),
.B1(n_843),
.B2(n_848),
.Y(n_999)
);

OAI21xp33_ASAP7_75t_L g1000 ( 
.A1(n_875),
.A2(n_878),
.B(n_888),
.Y(n_1000)
);

AOI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_763),
.A2(n_807),
.B(n_788),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_SL g1002 ( 
.A(n_756),
.B(n_778),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_SL g1003 ( 
.A(n_756),
.B(n_778),
.Y(n_1003)
);

NAND3xp33_ASAP7_75t_SL g1004 ( 
.A(n_760),
.B(n_849),
.C(n_918),
.Y(n_1004)
);

INVx6_ASAP7_75t_SL g1005 ( 
.A(n_898),
.Y(n_1005)
);

NOR2xp33_ASAP7_75t_L g1006 ( 
.A(n_869),
.B(n_876),
.Y(n_1006)
);

OAI22xp5_ASAP7_75t_L g1007 ( 
.A1(n_859),
.A2(n_917),
.B1(n_915),
.B2(n_908),
.Y(n_1007)
);

O2A1O1Ixp33_ASAP7_75t_L g1008 ( 
.A1(n_799),
.A2(n_855),
.B(n_827),
.C(n_884),
.Y(n_1008)
);

INVx1_ASAP7_75t_SL g1009 ( 
.A(n_768),
.Y(n_1009)
);

O2A1O1Ixp33_ASAP7_75t_L g1010 ( 
.A1(n_904),
.A2(n_859),
.B(n_785),
.C(n_804),
.Y(n_1010)
);

BUFx3_ASAP7_75t_L g1011 ( 
.A(n_818),
.Y(n_1011)
);

AOI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_762),
.A2(n_780),
.B(n_806),
.Y(n_1012)
);

AOI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_762),
.A2(n_780),
.B(n_832),
.Y(n_1013)
);

NOR3xp33_ASAP7_75t_L g1014 ( 
.A(n_793),
.B(n_790),
.C(n_811),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_895),
.Y(n_1015)
);

NOR2xp33_ASAP7_75t_L g1016 ( 
.A(n_869),
.B(n_880),
.Y(n_1016)
);

AOI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_831),
.A2(n_838),
.B(n_885),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_897),
.Y(n_1018)
);

OAI21xp33_ASAP7_75t_L g1019 ( 
.A1(n_813),
.A2(n_871),
.B(n_853),
.Y(n_1019)
);

AO32x1_ASAP7_75t_L g1020 ( 
.A1(n_771),
.A2(n_777),
.A3(n_781),
.B1(n_787),
.B2(n_840),
.Y(n_1020)
);

OAI22xp5_ASAP7_75t_L g1021 ( 
.A1(n_906),
.A2(n_912),
.B1(n_876),
.B2(n_880),
.Y(n_1021)
);

INVx3_ASAP7_75t_SL g1022 ( 
.A(n_818),
.Y(n_1022)
);

BUFx6f_ASAP7_75t_L g1023 ( 
.A(n_818),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_SL g1024 ( 
.A(n_824),
.B(n_772),
.Y(n_1024)
);

O2A1O1Ixp33_ASAP7_75t_L g1025 ( 
.A1(n_802),
.A2(n_811),
.B(n_844),
.C(n_835),
.Y(n_1025)
);

CKINVDCx20_ASAP7_75t_R g1026 ( 
.A(n_824),
.Y(n_1026)
);

CKINVDCx20_ASAP7_75t_R g1027 ( 
.A(n_824),
.Y(n_1027)
);

NOR2xp33_ASAP7_75t_L g1028 ( 
.A(n_911),
.B(n_892),
.Y(n_1028)
);

AND2x4_ASAP7_75t_L g1029 ( 
.A(n_864),
.B(n_844),
.Y(n_1029)
);

OAI22xp5_ASAP7_75t_L g1030 ( 
.A1(n_874),
.A2(n_899),
.B1(n_825),
.B2(n_826),
.Y(n_1030)
);

AO32x1_ASAP7_75t_L g1031 ( 
.A1(n_893),
.A2(n_842),
.A3(n_828),
.B1(n_892),
.B2(n_822),
.Y(n_1031)
);

A2O1A1Ixp33_ASAP7_75t_L g1032 ( 
.A1(n_796),
.A2(n_803),
.B(n_805),
.C(n_913),
.Y(n_1032)
);

OAI22xp5_ASAP7_75t_L g1033 ( 
.A1(n_791),
.A2(n_902),
.B1(n_769),
.B2(n_846),
.Y(n_1033)
);

AOI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_873),
.A2(n_882),
.B(n_754),
.Y(n_1034)
);

AOI22xp5_ASAP7_75t_L g1035 ( 
.A1(n_852),
.A2(n_649),
.B1(n_606),
.B2(n_598),
.Y(n_1035)
);

OAI22xp5_ASAP7_75t_L g1036 ( 
.A1(n_786),
.A2(n_451),
.B1(n_606),
.B2(n_670),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_SL g1037 ( 
.A(n_758),
.B(n_605),
.Y(n_1037)
);

HB1xp67_ASAP7_75t_L g1038 ( 
.A(n_776),
.Y(n_1038)
);

AOI222xp33_ASAP7_75t_L g1039 ( 
.A1(n_889),
.A2(n_608),
.B1(n_626),
.B2(n_423),
.C1(n_698),
.C2(n_745),
.Y(n_1039)
);

INVxp67_ASAP7_75t_L g1040 ( 
.A(n_776),
.Y(n_1040)
);

NOR2xp33_ASAP7_75t_L g1041 ( 
.A(n_852),
.B(n_649),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_SL g1042 ( 
.A(n_758),
.B(n_605),
.Y(n_1042)
);

AND2x2_ASAP7_75t_L g1043 ( 
.A(n_833),
.B(n_662),
.Y(n_1043)
);

AOI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_754),
.A2(n_738),
.B(n_610),
.Y(n_1044)
);

AND2x2_ASAP7_75t_L g1045 ( 
.A(n_833),
.B(n_662),
.Y(n_1045)
);

AOI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_754),
.A2(n_738),
.B(n_610),
.Y(n_1046)
);

O2A1O1Ixp33_ASAP7_75t_L g1047 ( 
.A1(n_1041),
.A2(n_969),
.B(n_1036),
.C(n_993),
.Y(n_1047)
);

O2A1O1Ixp33_ASAP7_75t_SL g1048 ( 
.A1(n_1036),
.A2(n_993),
.B(n_1037),
.C(n_1042),
.Y(n_1048)
);

AOI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_1044),
.A2(n_1046),
.B(n_920),
.Y(n_1049)
);

A2O1A1Ixp33_ASAP7_75t_L g1050 ( 
.A1(n_1035),
.A2(n_939),
.B(n_1000),
.C(n_929),
.Y(n_1050)
);

AO31x2_ASAP7_75t_L g1051 ( 
.A1(n_935),
.A2(n_1007),
.A3(n_1030),
.B(n_951),
.Y(n_1051)
);

OAI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_974),
.A2(n_1025),
.B(n_933),
.Y(n_1052)
);

A2O1A1Ixp33_ASAP7_75t_L g1053 ( 
.A1(n_991),
.A2(n_930),
.B(n_953),
.C(n_971),
.Y(n_1053)
);

AOI21x1_ASAP7_75t_L g1054 ( 
.A1(n_1024),
.A2(n_1030),
.B(n_977),
.Y(n_1054)
);

AOI22xp33_ASAP7_75t_L g1055 ( 
.A1(n_1039),
.A2(n_1005),
.B1(n_946),
.B2(n_972),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_944),
.B(n_992),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_992),
.B(n_937),
.Y(n_1057)
);

AOI22xp5_ASAP7_75t_L g1058 ( 
.A1(n_1039),
.A2(n_978),
.B1(n_1043),
.B2(n_1045),
.Y(n_1058)
);

BUFx6f_ASAP7_75t_L g1059 ( 
.A(n_957),
.Y(n_1059)
);

AO31x2_ASAP7_75t_L g1060 ( 
.A1(n_1007),
.A2(n_951),
.A3(n_1032),
.B(n_1033),
.Y(n_1060)
);

NOR2x1_ASAP7_75t_SL g1061 ( 
.A(n_989),
.B(n_980),
.Y(n_1061)
);

OAI21xp5_ASAP7_75t_L g1062 ( 
.A1(n_933),
.A2(n_1010),
.B(n_921),
.Y(n_1062)
);

AOI21xp5_ASAP7_75t_L g1063 ( 
.A1(n_1001),
.A2(n_1034),
.B(n_995),
.Y(n_1063)
);

AOI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_987),
.A2(n_926),
.B(n_932),
.Y(n_1064)
);

A2O1A1Ixp33_ASAP7_75t_L g1065 ( 
.A1(n_975),
.A2(n_1004),
.B(n_947),
.C(n_1008),
.Y(n_1065)
);

BUFx2_ASAP7_75t_L g1066 ( 
.A(n_928),
.Y(n_1066)
);

AOI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_1033),
.A2(n_1017),
.B(n_956),
.Y(n_1067)
);

NOR2xp33_ASAP7_75t_L g1068 ( 
.A(n_978),
.B(n_1040),
.Y(n_1068)
);

AOI21xp5_ASAP7_75t_L g1069 ( 
.A1(n_968),
.A2(n_934),
.B(n_940),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_919),
.Y(n_1070)
);

A2O1A1Ixp33_ASAP7_75t_L g1071 ( 
.A1(n_979),
.A2(n_950),
.B(n_1028),
.C(n_1019),
.Y(n_1071)
);

OAI21xp5_ASAP7_75t_L g1072 ( 
.A1(n_1013),
.A2(n_925),
.B(n_1012),
.Y(n_1072)
);

AOI21xp5_ASAP7_75t_L g1073 ( 
.A1(n_938),
.A2(n_959),
.B(n_1021),
.Y(n_1073)
);

OAI21x1_ASAP7_75t_SL g1074 ( 
.A1(n_948),
.A2(n_996),
.B(n_966),
.Y(n_1074)
);

OAI21x1_ASAP7_75t_L g1075 ( 
.A1(n_948),
.A2(n_962),
.B(n_970),
.Y(n_1075)
);

OAI21xp5_ASAP7_75t_L g1076 ( 
.A1(n_1014),
.A2(n_966),
.B(n_965),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_955),
.B(n_952),
.Y(n_1077)
);

OR2x2_ASAP7_75t_L g1078 ( 
.A(n_1038),
.B(n_936),
.Y(n_1078)
);

AOI21x1_ASAP7_75t_SL g1079 ( 
.A1(n_967),
.A2(n_965),
.B(n_924),
.Y(n_1079)
);

CKINVDCx11_ASAP7_75t_R g1080 ( 
.A(n_958),
.Y(n_1080)
);

BUFx3_ASAP7_75t_L g1081 ( 
.A(n_943),
.Y(n_1081)
);

NOR2xp33_ASAP7_75t_L g1082 ( 
.A(n_931),
.B(n_922),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_955),
.B(n_1002),
.Y(n_1083)
);

AOI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_985),
.A2(n_941),
.B(n_1031),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_954),
.Y(n_1085)
);

NAND3x1_ASAP7_75t_L g1086 ( 
.A(n_976),
.B(n_1005),
.C(n_983),
.Y(n_1086)
);

A2O1A1Ixp33_ASAP7_75t_L g1087 ( 
.A1(n_961),
.A2(n_999),
.B(n_960),
.C(n_945),
.Y(n_1087)
);

HB1xp67_ASAP7_75t_L g1088 ( 
.A(n_1026),
.Y(n_1088)
);

BUFx6f_ASAP7_75t_L g1089 ( 
.A(n_957),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_1003),
.B(n_946),
.Y(n_1090)
);

INVx3_ASAP7_75t_SL g1091 ( 
.A(n_949),
.Y(n_1091)
);

OAI21xp5_ASAP7_75t_L g1092 ( 
.A1(n_941),
.A2(n_1006),
.B(n_1016),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_981),
.B(n_982),
.Y(n_1093)
);

OR2x2_ASAP7_75t_L g1094 ( 
.A(n_1015),
.B(n_1018),
.Y(n_1094)
);

AOI22xp5_ASAP7_75t_L g1095 ( 
.A1(n_990),
.A2(n_994),
.B1(n_963),
.B2(n_1027),
.Y(n_1095)
);

BUFx6f_ASAP7_75t_L g1096 ( 
.A(n_957),
.Y(n_1096)
);

INVx3_ASAP7_75t_L g1097 ( 
.A(n_989),
.Y(n_1097)
);

AOI22xp5_ASAP7_75t_L g1098 ( 
.A1(n_990),
.A2(n_994),
.B1(n_1029),
.B2(n_964),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_1009),
.B(n_942),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_986),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_986),
.Y(n_1101)
);

AO31x2_ASAP7_75t_L g1102 ( 
.A1(n_1020),
.A2(n_986),
.A3(n_985),
.B(n_1031),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_988),
.Y(n_1103)
);

OR2x2_ASAP7_75t_L g1104 ( 
.A(n_1022),
.B(n_1011),
.Y(n_1104)
);

CKINVDCx20_ASAP7_75t_R g1105 ( 
.A(n_984),
.Y(n_1105)
);

AOI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_985),
.A2(n_1031),
.B(n_1020),
.Y(n_1106)
);

AND2x4_ASAP7_75t_L g1107 ( 
.A(n_997),
.B(n_998),
.Y(n_1107)
);

INVx4_ASAP7_75t_L g1108 ( 
.A(n_927),
.Y(n_1108)
);

OAI21x1_ASAP7_75t_L g1109 ( 
.A1(n_998),
.A2(n_1023),
.B(n_927),
.Y(n_1109)
);

INVx2_ASAP7_75t_SL g1110 ( 
.A(n_973),
.Y(n_1110)
);

A2O1A1Ixp33_ASAP7_75t_L g1111 ( 
.A1(n_1023),
.A2(n_1041),
.B(n_1035),
.C(n_969),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_988),
.Y(n_1112)
);

AOI221x1_ASAP7_75t_L g1113 ( 
.A1(n_927),
.A2(n_1041),
.B1(n_972),
.B2(n_991),
.C(n_993),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_919),
.Y(n_1114)
);

A2O1A1Ixp33_ASAP7_75t_L g1115 ( 
.A1(n_1041),
.A2(n_1035),
.B(n_969),
.C(n_939),
.Y(n_1115)
);

AOI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_1044),
.A2(n_1046),
.B(n_920),
.Y(n_1116)
);

OAI21xp5_ASAP7_75t_L g1117 ( 
.A1(n_1036),
.A2(n_929),
.B(n_1041),
.Y(n_1117)
);

OAI21x1_ASAP7_75t_L g1118 ( 
.A1(n_1017),
.A2(n_923),
.B(n_987),
.Y(n_1118)
);

AOI21xp5_ASAP7_75t_L g1119 ( 
.A1(n_1044),
.A2(n_1046),
.B(n_920),
.Y(n_1119)
);

NAND2xp33_ASAP7_75t_R g1120 ( 
.A(n_1041),
.B(n_580),
.Y(n_1120)
);

OAI22xp5_ASAP7_75t_L g1121 ( 
.A1(n_1035),
.A2(n_1041),
.B1(n_939),
.B2(n_1036),
.Y(n_1121)
);

AOI21xp5_ASAP7_75t_L g1122 ( 
.A1(n_1044),
.A2(n_1046),
.B(n_920),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_919),
.Y(n_1123)
);

NOR2xp33_ASAP7_75t_L g1124 ( 
.A(n_1041),
.B(n_649),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_919),
.Y(n_1125)
);

AOI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_1044),
.A2(n_1046),
.B(n_920),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_1036),
.B(n_1035),
.Y(n_1127)
);

BUFx2_ASAP7_75t_L g1128 ( 
.A(n_928),
.Y(n_1128)
);

AO31x2_ASAP7_75t_L g1129 ( 
.A1(n_935),
.A2(n_1007),
.A3(n_1030),
.B(n_951),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_919),
.Y(n_1130)
);

OA21x2_ASAP7_75t_L g1131 ( 
.A1(n_977),
.A2(n_987),
.B(n_995),
.Y(n_1131)
);

OAI21x1_ASAP7_75t_SL g1132 ( 
.A1(n_969),
.A2(n_974),
.B(n_993),
.Y(n_1132)
);

A2O1A1Ixp33_ASAP7_75t_L g1133 ( 
.A1(n_1041),
.A2(n_1035),
.B(n_969),
.C(n_939),
.Y(n_1133)
);

OAI21x1_ASAP7_75t_L g1134 ( 
.A1(n_1017),
.A2(n_923),
.B(n_987),
.Y(n_1134)
);

OAI21x1_ASAP7_75t_L g1135 ( 
.A1(n_1017),
.A2(n_923),
.B(n_987),
.Y(n_1135)
);

CKINVDCx6p67_ASAP7_75t_R g1136 ( 
.A(n_949),
.Y(n_1136)
);

AO31x2_ASAP7_75t_L g1137 ( 
.A1(n_935),
.A2(n_1007),
.A3(n_1030),
.B(n_951),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_919),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_919),
.Y(n_1139)
);

OAI21xp5_ASAP7_75t_L g1140 ( 
.A1(n_1036),
.A2(n_929),
.B(n_1041),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_SL g1141 ( 
.A(n_1035),
.B(n_1041),
.Y(n_1141)
);

OAI21x1_ASAP7_75t_L g1142 ( 
.A1(n_1017),
.A2(n_923),
.B(n_987),
.Y(n_1142)
);

A2O1A1Ixp33_ASAP7_75t_L g1143 ( 
.A1(n_1041),
.A2(n_1035),
.B(n_969),
.C(n_939),
.Y(n_1143)
);

AO31x2_ASAP7_75t_L g1144 ( 
.A1(n_935),
.A2(n_1007),
.A3(n_1030),
.B(n_951),
.Y(n_1144)
);

INVx1_ASAP7_75t_SL g1145 ( 
.A(n_928),
.Y(n_1145)
);

AOI22xp5_ASAP7_75t_L g1146 ( 
.A1(n_1041),
.A2(n_1035),
.B1(n_649),
.B2(n_939),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_919),
.Y(n_1147)
);

AOI21x1_ASAP7_75t_L g1148 ( 
.A1(n_1024),
.A2(n_1030),
.B(n_977),
.Y(n_1148)
);

INVx2_ASAP7_75t_SL g1149 ( 
.A(n_943),
.Y(n_1149)
);

AOI21xp5_ASAP7_75t_L g1150 ( 
.A1(n_1044),
.A2(n_1046),
.B(n_920),
.Y(n_1150)
);

CKINVDCx5p33_ASAP7_75t_R g1151 ( 
.A(n_958),
.Y(n_1151)
);

INVx1_ASAP7_75t_SL g1152 ( 
.A(n_928),
.Y(n_1152)
);

OR2x2_ASAP7_75t_L g1153 ( 
.A(n_1043),
.B(n_833),
.Y(n_1153)
);

OAI21xp5_ASAP7_75t_L g1154 ( 
.A1(n_1036),
.A2(n_929),
.B(n_1041),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_1036),
.B(n_1035),
.Y(n_1155)
);

AO22x2_ASAP7_75t_L g1156 ( 
.A1(n_993),
.A2(n_890),
.B1(n_991),
.B2(n_889),
.Y(n_1156)
);

INVx3_ASAP7_75t_L g1157 ( 
.A(n_989),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_919),
.Y(n_1158)
);

OAI22xp33_ASAP7_75t_L g1159 ( 
.A1(n_1035),
.A2(n_1041),
.B1(n_745),
.B2(n_1005),
.Y(n_1159)
);

AO31x2_ASAP7_75t_L g1160 ( 
.A1(n_935),
.A2(n_1007),
.A3(n_1030),
.B(n_951),
.Y(n_1160)
);

OAI21x1_ASAP7_75t_L g1161 ( 
.A1(n_1017),
.A2(n_923),
.B(n_987),
.Y(n_1161)
);

BUFx3_ASAP7_75t_L g1162 ( 
.A(n_958),
.Y(n_1162)
);

AOI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_1044),
.A2(n_1046),
.B(n_920),
.Y(n_1163)
);

OR2x6_ASAP7_75t_L g1164 ( 
.A(n_989),
.B(n_757),
.Y(n_1164)
);

AND2x2_ASAP7_75t_L g1165 ( 
.A(n_1043),
.B(n_1045),
.Y(n_1165)
);

AOI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_1044),
.A2(n_1046),
.B(n_920),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_919),
.Y(n_1167)
);

BUFx4_ASAP7_75t_SL g1168 ( 
.A(n_958),
.Y(n_1168)
);

A2O1A1Ixp33_ASAP7_75t_L g1169 ( 
.A1(n_1041),
.A2(n_1035),
.B(n_969),
.C(n_939),
.Y(n_1169)
);

O2A1O1Ixp33_ASAP7_75t_SL g1170 ( 
.A1(n_1041),
.A2(n_1036),
.B(n_993),
.C(n_1037),
.Y(n_1170)
);

A2O1A1Ixp33_ASAP7_75t_L g1171 ( 
.A1(n_1041),
.A2(n_1035),
.B(n_969),
.C(n_939),
.Y(n_1171)
);

OAI21xp5_ASAP7_75t_L g1172 ( 
.A1(n_1036),
.A2(n_929),
.B(n_1041),
.Y(n_1172)
);

AOI211x1_ASAP7_75t_L g1173 ( 
.A1(n_1000),
.A2(n_451),
.B(n_898),
.C(n_631),
.Y(n_1173)
);

NOR2xp33_ASAP7_75t_L g1174 ( 
.A(n_1041),
.B(n_649),
.Y(n_1174)
);

OAI222xp33_ASAP7_75t_L g1175 ( 
.A1(n_1035),
.A2(n_558),
.B1(n_745),
.B2(n_380),
.C1(n_322),
.C2(n_582),
.Y(n_1175)
);

INVx3_ASAP7_75t_L g1176 ( 
.A(n_989),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_919),
.Y(n_1177)
);

AOI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_1044),
.A2(n_1046),
.B(n_920),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_1036),
.B(n_1035),
.Y(n_1179)
);

OAI21x1_ASAP7_75t_L g1180 ( 
.A1(n_1017),
.A2(n_923),
.B(n_987),
.Y(n_1180)
);

AND2x4_ASAP7_75t_L g1181 ( 
.A(n_1098),
.B(n_1095),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_1094),
.Y(n_1182)
);

INVx1_ASAP7_75t_SL g1183 ( 
.A(n_1145),
.Y(n_1183)
);

AOI22xp33_ASAP7_75t_SL g1184 ( 
.A1(n_1121),
.A2(n_1090),
.B1(n_1156),
.B2(n_1124),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_1093),
.Y(n_1185)
);

AOI21xp5_ASAP7_75t_L g1186 ( 
.A1(n_1121),
.A2(n_1140),
.B(n_1117),
.Y(n_1186)
);

AOI22xp33_ASAP7_75t_L g1187 ( 
.A1(n_1055),
.A2(n_1174),
.B1(n_1090),
.B2(n_1146),
.Y(n_1187)
);

OAI21xp5_ASAP7_75t_SL g1188 ( 
.A1(n_1115),
.A2(n_1143),
.B(n_1133),
.Y(n_1188)
);

BUFx6f_ASAP7_75t_SL g1189 ( 
.A(n_1081),
.Y(n_1189)
);

OAI22xp33_ASAP7_75t_L g1190 ( 
.A1(n_1058),
.A2(n_1155),
.B1(n_1179),
.B2(n_1127),
.Y(n_1190)
);

AOI22xp33_ASAP7_75t_L g1191 ( 
.A1(n_1141),
.A2(n_1159),
.B1(n_1156),
.B2(n_1154),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_1056),
.B(n_1165),
.Y(n_1192)
);

AOI22xp33_ASAP7_75t_SL g1193 ( 
.A1(n_1117),
.A2(n_1140),
.B1(n_1154),
.B2(n_1172),
.Y(n_1193)
);

OAI22xp5_ASAP7_75t_L g1194 ( 
.A1(n_1169),
.A2(n_1171),
.B1(n_1155),
.B2(n_1127),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_1093),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_1085),
.Y(n_1196)
);

OAI22xp33_ASAP7_75t_L g1197 ( 
.A1(n_1179),
.A2(n_1172),
.B1(n_1113),
.B2(n_1120),
.Y(n_1197)
);

AOI22xp33_ASAP7_75t_L g1198 ( 
.A1(n_1132),
.A2(n_1076),
.B1(n_1052),
.B2(n_1056),
.Y(n_1198)
);

BUFx2_ASAP7_75t_SL g1199 ( 
.A(n_1105),
.Y(n_1199)
);

BUFx10_ASAP7_75t_L g1200 ( 
.A(n_1151),
.Y(n_1200)
);

CKINVDCx20_ASAP7_75t_R g1201 ( 
.A(n_1080),
.Y(n_1201)
);

CKINVDCx20_ASAP7_75t_R g1202 ( 
.A(n_1136),
.Y(n_1202)
);

CKINVDCx11_ASAP7_75t_R g1203 ( 
.A(n_1091),
.Y(n_1203)
);

AOI22xp33_ASAP7_75t_SL g1204 ( 
.A1(n_1052),
.A2(n_1076),
.B1(n_1175),
.B2(n_1074),
.Y(n_1204)
);

INVx6_ASAP7_75t_L g1205 ( 
.A(n_1059),
.Y(n_1205)
);

OAI22xp5_ASAP7_75t_L g1206 ( 
.A1(n_1050),
.A2(n_1111),
.B1(n_1053),
.B2(n_1047),
.Y(n_1206)
);

AOI22xp5_ASAP7_75t_L g1207 ( 
.A1(n_1086),
.A2(n_1068),
.B1(n_1170),
.B2(n_1082),
.Y(n_1207)
);

INVx6_ASAP7_75t_L g1208 ( 
.A(n_1089),
.Y(n_1208)
);

OAI22xp33_ASAP7_75t_L g1209 ( 
.A1(n_1153),
.A2(n_1057),
.B1(n_1078),
.B2(n_1125),
.Y(n_1209)
);

AOI22xp33_ASAP7_75t_SL g1210 ( 
.A1(n_1062),
.A2(n_1061),
.B1(n_1057),
.B2(n_1130),
.Y(n_1210)
);

INVx6_ASAP7_75t_L g1211 ( 
.A(n_1089),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1070),
.Y(n_1212)
);

INVx3_ASAP7_75t_L g1213 ( 
.A(n_1108),
.Y(n_1213)
);

BUFx10_ASAP7_75t_L g1214 ( 
.A(n_1110),
.Y(n_1214)
);

OAI22xp5_ASAP7_75t_L g1215 ( 
.A1(n_1173),
.A2(n_1065),
.B1(n_1062),
.B2(n_1152),
.Y(n_1215)
);

OAI21xp5_ASAP7_75t_SL g1216 ( 
.A1(n_1092),
.A2(n_1048),
.B(n_1084),
.Y(n_1216)
);

BUFx2_ASAP7_75t_SL g1217 ( 
.A(n_1162),
.Y(n_1217)
);

BUFx6f_ASAP7_75t_L g1218 ( 
.A(n_1089),
.Y(n_1218)
);

BUFx10_ASAP7_75t_L g1219 ( 
.A(n_1149),
.Y(n_1219)
);

CKINVDCx11_ASAP7_75t_R g1220 ( 
.A(n_1145),
.Y(n_1220)
);

BUFx10_ASAP7_75t_L g1221 ( 
.A(n_1168),
.Y(n_1221)
);

AOI21xp5_ASAP7_75t_L g1222 ( 
.A1(n_1067),
.A2(n_1063),
.B(n_1178),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1114),
.Y(n_1223)
);

AOI22xp33_ASAP7_75t_L g1224 ( 
.A1(n_1123),
.A2(n_1139),
.B1(n_1177),
.B2(n_1138),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_1147),
.B(n_1158),
.Y(n_1225)
);

OAI22xp33_ASAP7_75t_L g1226 ( 
.A1(n_1167),
.A2(n_1083),
.B1(n_1152),
.B2(n_1077),
.Y(n_1226)
);

OAI22xp33_ASAP7_75t_L g1227 ( 
.A1(n_1083),
.A2(n_1077),
.B1(n_1088),
.B2(n_1164),
.Y(n_1227)
);

INVx6_ASAP7_75t_L g1228 ( 
.A(n_1096),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1099),
.Y(n_1229)
);

BUFx3_ASAP7_75t_L g1230 ( 
.A(n_1066),
.Y(n_1230)
);

BUFx12f_ASAP7_75t_L g1231 ( 
.A(n_1128),
.Y(n_1231)
);

AOI22xp33_ASAP7_75t_SL g1232 ( 
.A1(n_1075),
.A2(n_1106),
.B1(n_1073),
.B2(n_1100),
.Y(n_1232)
);

CKINVDCx8_ASAP7_75t_R g1233 ( 
.A(n_1096),
.Y(n_1233)
);

OAI22xp5_ASAP7_75t_L g1234 ( 
.A1(n_1087),
.A2(n_1071),
.B1(n_1164),
.B2(n_1176),
.Y(n_1234)
);

OAI22xp5_ASAP7_75t_L g1235 ( 
.A1(n_1164),
.A2(n_1176),
.B1(n_1157),
.B2(n_1097),
.Y(n_1235)
);

AOI22xp33_ASAP7_75t_L g1236 ( 
.A1(n_1096),
.A2(n_1112),
.B1(n_1103),
.B2(n_1101),
.Y(n_1236)
);

OAI22xp33_ASAP7_75t_L g1237 ( 
.A1(n_1104),
.A2(n_1069),
.B1(n_1072),
.B2(n_1079),
.Y(n_1237)
);

OAI22xp33_ASAP7_75t_L g1238 ( 
.A1(n_1072),
.A2(n_1148),
.B1(n_1054),
.B2(n_1126),
.Y(n_1238)
);

INVx6_ASAP7_75t_L g1239 ( 
.A(n_1107),
.Y(n_1239)
);

CKINVDCx20_ASAP7_75t_R g1240 ( 
.A(n_1131),
.Y(n_1240)
);

HB1xp67_ASAP7_75t_L g1241 ( 
.A(n_1051),
.Y(n_1241)
);

BUFx12f_ASAP7_75t_L g1242 ( 
.A(n_1109),
.Y(n_1242)
);

AOI22xp33_ASAP7_75t_L g1243 ( 
.A1(n_1049),
.A2(n_1166),
.B1(n_1163),
.B2(n_1119),
.Y(n_1243)
);

AOI22xp33_ASAP7_75t_SL g1244 ( 
.A1(n_1060),
.A2(n_1051),
.B1(n_1137),
.B2(n_1160),
.Y(n_1244)
);

AOI22xp33_ASAP7_75t_L g1245 ( 
.A1(n_1116),
.A2(n_1150),
.B1(n_1122),
.B2(n_1064),
.Y(n_1245)
);

OAI21xp5_ASAP7_75t_L g1246 ( 
.A1(n_1118),
.A2(n_1180),
.B(n_1161),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1060),
.Y(n_1247)
);

INVx3_ASAP7_75t_L g1248 ( 
.A(n_1129),
.Y(n_1248)
);

CKINVDCx20_ASAP7_75t_R g1249 ( 
.A(n_1160),
.Y(n_1249)
);

INVx3_ASAP7_75t_L g1250 ( 
.A(n_1137),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_SL g1251 ( 
.A(n_1134),
.B(n_1135),
.Y(n_1251)
);

AOI22xp33_ASAP7_75t_L g1252 ( 
.A1(n_1142),
.A2(n_1055),
.B1(n_1041),
.B2(n_1005),
.Y(n_1252)
);

AOI22xp33_ASAP7_75t_L g1253 ( 
.A1(n_1144),
.A2(n_1055),
.B1(n_1041),
.B2(n_1005),
.Y(n_1253)
);

INVx1_ASAP7_75t_SL g1254 ( 
.A(n_1102),
.Y(n_1254)
);

INVx6_ASAP7_75t_L g1255 ( 
.A(n_1102),
.Y(n_1255)
);

BUFx2_ASAP7_75t_L g1256 ( 
.A(n_1102),
.Y(n_1256)
);

CKINVDCx20_ASAP7_75t_R g1257 ( 
.A(n_1080),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1094),
.Y(n_1258)
);

AOI22xp33_ASAP7_75t_L g1259 ( 
.A1(n_1055),
.A2(n_1041),
.B1(n_1005),
.B2(n_1039),
.Y(n_1259)
);

INVx6_ASAP7_75t_L g1260 ( 
.A(n_1059),
.Y(n_1260)
);

CKINVDCx20_ASAP7_75t_R g1261 ( 
.A(n_1080),
.Y(n_1261)
);

OAI22xp33_ASAP7_75t_L g1262 ( 
.A1(n_1146),
.A2(n_1121),
.B1(n_1035),
.B2(n_1005),
.Y(n_1262)
);

OAI22xp33_ASAP7_75t_L g1263 ( 
.A1(n_1146),
.A2(n_1121),
.B1(n_1035),
.B2(n_1005),
.Y(n_1263)
);

AOI22xp33_ASAP7_75t_L g1264 ( 
.A1(n_1055),
.A2(n_1039),
.B1(n_1041),
.B2(n_1005),
.Y(n_1264)
);

OAI22xp5_ASAP7_75t_L g1265 ( 
.A1(n_1146),
.A2(n_1124),
.B1(n_1174),
.B2(n_1133),
.Y(n_1265)
);

AOI22xp33_ASAP7_75t_L g1266 ( 
.A1(n_1055),
.A2(n_1039),
.B1(n_1041),
.B2(n_1005),
.Y(n_1266)
);

AOI22xp33_ASAP7_75t_L g1267 ( 
.A1(n_1055),
.A2(n_1039),
.B1(n_1041),
.B2(n_1005),
.Y(n_1267)
);

BUFx3_ASAP7_75t_L g1268 ( 
.A(n_1091),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1094),
.Y(n_1269)
);

AOI22xp33_ASAP7_75t_SL g1270 ( 
.A1(n_1121),
.A2(n_1090),
.B1(n_889),
.B2(n_1041),
.Y(n_1270)
);

INVx1_ASAP7_75t_SL g1271 ( 
.A(n_1145),
.Y(n_1271)
);

AOI22xp33_ASAP7_75t_L g1272 ( 
.A1(n_1055),
.A2(n_1039),
.B1(n_1041),
.B2(n_1005),
.Y(n_1272)
);

CKINVDCx11_ASAP7_75t_R g1273 ( 
.A(n_1105),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1094),
.Y(n_1274)
);

INVx6_ASAP7_75t_L g1275 ( 
.A(n_1059),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1094),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1094),
.Y(n_1277)
);

AOI22xp33_ASAP7_75t_L g1278 ( 
.A1(n_1055),
.A2(n_1039),
.B1(n_1041),
.B2(n_1005),
.Y(n_1278)
);

BUFx8_ASAP7_75t_L g1279 ( 
.A(n_1066),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_L g1280 ( 
.A(n_1124),
.B(n_1174),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1094),
.Y(n_1281)
);

INVx2_ASAP7_75t_SL g1282 ( 
.A(n_1168),
.Y(n_1282)
);

AOI22xp33_ASAP7_75t_L g1283 ( 
.A1(n_1055),
.A2(n_1039),
.B1(n_1041),
.B2(n_1005),
.Y(n_1283)
);

INVx1_ASAP7_75t_SL g1284 ( 
.A(n_1145),
.Y(n_1284)
);

BUFx3_ASAP7_75t_L g1285 ( 
.A(n_1091),
.Y(n_1285)
);

AOI22xp5_ASAP7_75t_L g1286 ( 
.A1(n_1124),
.A2(n_1041),
.B1(n_1174),
.B2(n_1146),
.Y(n_1286)
);

CKINVDCx11_ASAP7_75t_R g1287 ( 
.A(n_1105),
.Y(n_1287)
);

BUFx6f_ASAP7_75t_L g1288 ( 
.A(n_1059),
.Y(n_1288)
);

CKINVDCx6p67_ASAP7_75t_R g1289 ( 
.A(n_1091),
.Y(n_1289)
);

INVx4_ASAP7_75t_L g1290 ( 
.A(n_1091),
.Y(n_1290)
);

OAI22xp5_ASAP7_75t_L g1291 ( 
.A1(n_1146),
.A2(n_1124),
.B1(n_1174),
.B2(n_1133),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1241),
.Y(n_1292)
);

OAI21x1_ASAP7_75t_L g1293 ( 
.A1(n_1222),
.A2(n_1246),
.B(n_1245),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1241),
.Y(n_1294)
);

OAI21x1_ASAP7_75t_L g1295 ( 
.A1(n_1222),
.A2(n_1243),
.B(n_1251),
.Y(n_1295)
);

INVx4_ASAP7_75t_L g1296 ( 
.A(n_1242),
.Y(n_1296)
);

OAI21x1_ASAP7_75t_L g1297 ( 
.A1(n_1186),
.A2(n_1250),
.B(n_1248),
.Y(n_1297)
);

AOI22xp33_ASAP7_75t_L g1298 ( 
.A1(n_1264),
.A2(n_1272),
.B1(n_1278),
.B2(n_1267),
.Y(n_1298)
);

AND2x2_ASAP7_75t_L g1299 ( 
.A(n_1193),
.B(n_1186),
.Y(n_1299)
);

AOI22xp33_ASAP7_75t_L g1300 ( 
.A1(n_1264),
.A2(n_1272),
.B1(n_1278),
.B2(n_1267),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1247),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1229),
.Y(n_1302)
);

AND2x2_ASAP7_75t_L g1303 ( 
.A(n_1193),
.B(n_1256),
.Y(n_1303)
);

OR2x2_ASAP7_75t_SL g1304 ( 
.A(n_1184),
.B(n_1255),
.Y(n_1304)
);

BUFx2_ASAP7_75t_L g1305 ( 
.A(n_1240),
.Y(n_1305)
);

BUFx2_ASAP7_75t_L g1306 ( 
.A(n_1255),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1196),
.Y(n_1307)
);

AND2x2_ASAP7_75t_L g1308 ( 
.A(n_1244),
.B(n_1254),
.Y(n_1308)
);

INVx3_ASAP7_75t_L g1309 ( 
.A(n_1213),
.Y(n_1309)
);

BUFx3_ASAP7_75t_L g1310 ( 
.A(n_1230),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1185),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1195),
.Y(n_1312)
);

HB1xp67_ASAP7_75t_L g1313 ( 
.A(n_1215),
.Y(n_1313)
);

AOI22xp33_ASAP7_75t_SL g1314 ( 
.A1(n_1265),
.A2(n_1291),
.B1(n_1206),
.B2(n_1194),
.Y(n_1314)
);

AND2x2_ASAP7_75t_L g1315 ( 
.A(n_1244),
.B(n_1232),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1212),
.Y(n_1316)
);

NOR2x1_ASAP7_75t_R g1317 ( 
.A(n_1203),
.B(n_1273),
.Y(n_1317)
);

AND2x2_ASAP7_75t_L g1318 ( 
.A(n_1232),
.B(n_1198),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1223),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1249),
.Y(n_1320)
);

AO21x2_ASAP7_75t_L g1321 ( 
.A1(n_1238),
.A2(n_1237),
.B(n_1190),
.Y(n_1321)
);

BUFx2_ASAP7_75t_L g1322 ( 
.A(n_1227),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1226),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_L g1324 ( 
.A(n_1226),
.B(n_1198),
.Y(n_1324)
);

AO21x1_ASAP7_75t_SL g1325 ( 
.A1(n_1191),
.A2(n_1236),
.B(n_1252),
.Y(n_1325)
);

AND2x2_ASAP7_75t_L g1326 ( 
.A(n_1224),
.B(n_1191),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1182),
.Y(n_1327)
);

INVx1_ASAP7_75t_SL g1328 ( 
.A(n_1183),
.Y(n_1328)
);

BUFx2_ASAP7_75t_L g1329 ( 
.A(n_1227),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1258),
.Y(n_1330)
);

INVx3_ASAP7_75t_L g1331 ( 
.A(n_1213),
.Y(n_1331)
);

AND2x4_ASAP7_75t_L g1332 ( 
.A(n_1181),
.B(n_1269),
.Y(n_1332)
);

AND2x4_ASAP7_75t_L g1333 ( 
.A(n_1181),
.B(n_1274),
.Y(n_1333)
);

OR2x2_ASAP7_75t_L g1334 ( 
.A(n_1192),
.B(n_1209),
.Y(n_1334)
);

BUFx2_ASAP7_75t_L g1335 ( 
.A(n_1231),
.Y(n_1335)
);

AND2x2_ASAP7_75t_L g1336 ( 
.A(n_1216),
.B(n_1184),
.Y(n_1336)
);

CKINVDCx6p67_ASAP7_75t_R g1337 ( 
.A(n_1189),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1276),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1277),
.Y(n_1339)
);

NOR2x1_ASAP7_75t_SL g1340 ( 
.A(n_1188),
.B(n_1234),
.Y(n_1340)
);

OA21x2_ASAP7_75t_L g1341 ( 
.A1(n_1253),
.A2(n_1224),
.B(n_1225),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1281),
.Y(n_1342)
);

BUFx2_ASAP7_75t_L g1343 ( 
.A(n_1237),
.Y(n_1343)
);

OR2x2_ASAP7_75t_L g1344 ( 
.A(n_1209),
.B(n_1190),
.Y(n_1344)
);

AND2x2_ASAP7_75t_L g1345 ( 
.A(n_1204),
.B(n_1270),
.Y(n_1345)
);

AOI21xp5_ASAP7_75t_L g1346 ( 
.A1(n_1262),
.A2(n_1263),
.B(n_1238),
.Y(n_1346)
);

OR2x6_ASAP7_75t_L g1347 ( 
.A(n_1239),
.B(n_1235),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1197),
.Y(n_1348)
);

AND2x4_ASAP7_75t_L g1349 ( 
.A(n_1218),
.B(n_1288),
.Y(n_1349)
);

NAND2x1p5_ASAP7_75t_L g1350 ( 
.A(n_1207),
.B(n_1288),
.Y(n_1350)
);

BUFx6f_ASAP7_75t_L g1351 ( 
.A(n_1288),
.Y(n_1351)
);

BUFx3_ASAP7_75t_L g1352 ( 
.A(n_1279),
.Y(n_1352)
);

HB1xp67_ASAP7_75t_L g1353 ( 
.A(n_1197),
.Y(n_1353)
);

OR2x2_ASAP7_75t_L g1354 ( 
.A(n_1271),
.B(n_1284),
.Y(n_1354)
);

CKINVDCx20_ASAP7_75t_R g1355 ( 
.A(n_1287),
.Y(n_1355)
);

BUFx3_ASAP7_75t_L g1356 ( 
.A(n_1279),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1210),
.Y(n_1357)
);

NOR2xp33_ASAP7_75t_R g1358 ( 
.A(n_1201),
.B(n_1257),
.Y(n_1358)
);

OAI21xp5_ASAP7_75t_L g1359 ( 
.A1(n_1286),
.A2(n_1262),
.B(n_1263),
.Y(n_1359)
);

BUFx3_ASAP7_75t_L g1360 ( 
.A(n_1233),
.Y(n_1360)
);

NAND2xp5_ASAP7_75t_L g1361 ( 
.A(n_1187),
.B(n_1270),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1210),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1204),
.Y(n_1363)
);

AO21x1_ASAP7_75t_L g1364 ( 
.A1(n_1280),
.A2(n_1283),
.B(n_1266),
.Y(n_1364)
);

AND2x2_ASAP7_75t_L g1365 ( 
.A(n_1303),
.B(n_1217),
.Y(n_1365)
);

OAI21xp5_ASAP7_75t_L g1366 ( 
.A1(n_1314),
.A2(n_1283),
.B(n_1266),
.Y(n_1366)
);

AND2x6_ASAP7_75t_L g1367 ( 
.A(n_1299),
.B(n_1285),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1307),
.Y(n_1368)
);

OR2x2_ASAP7_75t_L g1369 ( 
.A(n_1305),
.B(n_1259),
.Y(n_1369)
);

BUFx2_ASAP7_75t_L g1370 ( 
.A(n_1306),
.Y(n_1370)
);

OAI22xp5_ASAP7_75t_L g1371 ( 
.A1(n_1314),
.A2(n_1289),
.B1(n_1282),
.B2(n_1290),
.Y(n_1371)
);

OAI22xp5_ASAP7_75t_L g1372 ( 
.A1(n_1359),
.A2(n_1290),
.B1(n_1268),
.B2(n_1261),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_SL g1373 ( 
.A(n_1359),
.B(n_1219),
.Y(n_1373)
);

OAI22xp5_ASAP7_75t_L g1374 ( 
.A1(n_1298),
.A2(n_1202),
.B1(n_1199),
.B2(n_1260),
.Y(n_1374)
);

INVxp67_ASAP7_75t_L g1375 ( 
.A(n_1354),
.Y(n_1375)
);

AND2x2_ASAP7_75t_L g1376 ( 
.A(n_1303),
.B(n_1220),
.Y(n_1376)
);

AO32x2_ASAP7_75t_L g1377 ( 
.A1(n_1296),
.A2(n_1189),
.A3(n_1219),
.B1(n_1205),
.B2(n_1208),
.Y(n_1377)
);

OAI22xp5_ASAP7_75t_L g1378 ( 
.A1(n_1300),
.A2(n_1275),
.B1(n_1205),
.B2(n_1208),
.Y(n_1378)
);

INVx1_ASAP7_75t_SL g1379 ( 
.A(n_1354),
.Y(n_1379)
);

AOI22xp33_ASAP7_75t_L g1380 ( 
.A1(n_1364),
.A2(n_1275),
.B1(n_1205),
.B2(n_1208),
.Y(n_1380)
);

AO32x2_ASAP7_75t_L g1381 ( 
.A1(n_1296),
.A2(n_1211),
.A3(n_1228),
.B1(n_1260),
.B2(n_1214),
.Y(n_1381)
);

AND2x2_ASAP7_75t_L g1382 ( 
.A(n_1303),
.B(n_1221),
.Y(n_1382)
);

AND2x2_ASAP7_75t_L g1383 ( 
.A(n_1315),
.B(n_1221),
.Y(n_1383)
);

OR2x2_ASAP7_75t_L g1384 ( 
.A(n_1305),
.B(n_1200),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_L g1385 ( 
.A(n_1299),
.B(n_1211),
.Y(n_1385)
);

OAI21xp5_ASAP7_75t_L g1386 ( 
.A1(n_1346),
.A2(n_1324),
.B(n_1353),
.Y(n_1386)
);

NOR2xp33_ASAP7_75t_L g1387 ( 
.A(n_1355),
.B(n_1200),
.Y(n_1387)
);

HB1xp67_ASAP7_75t_L g1388 ( 
.A(n_1328),
.Y(n_1388)
);

AOI21xp5_ASAP7_75t_L g1389 ( 
.A1(n_1346),
.A2(n_1214),
.B(n_1321),
.Y(n_1389)
);

AOI22xp33_ASAP7_75t_L g1390 ( 
.A1(n_1364),
.A2(n_1345),
.B1(n_1363),
.B2(n_1336),
.Y(n_1390)
);

AO32x2_ASAP7_75t_L g1391 ( 
.A1(n_1296),
.A2(n_1353),
.A3(n_1334),
.B1(n_1329),
.B2(n_1322),
.Y(n_1391)
);

NOR2xp33_ASAP7_75t_L g1392 ( 
.A(n_1310),
.B(n_1335),
.Y(n_1392)
);

AND2x2_ASAP7_75t_L g1393 ( 
.A(n_1318),
.B(n_1308),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_L g1394 ( 
.A(n_1328),
.B(n_1334),
.Y(n_1394)
);

AND2x2_ASAP7_75t_L g1395 ( 
.A(n_1318),
.B(n_1308),
.Y(n_1395)
);

AND2x2_ASAP7_75t_L g1396 ( 
.A(n_1318),
.B(n_1308),
.Y(n_1396)
);

A2O1A1Ixp33_ASAP7_75t_L g1397 ( 
.A1(n_1345),
.A2(n_1336),
.B(n_1344),
.C(n_1361),
.Y(n_1397)
);

AND2x2_ASAP7_75t_L g1398 ( 
.A(n_1321),
.B(n_1316),
.Y(n_1398)
);

BUFx2_ASAP7_75t_SL g1399 ( 
.A(n_1360),
.Y(n_1399)
);

AOI22xp33_ASAP7_75t_L g1400 ( 
.A1(n_1363),
.A2(n_1336),
.B1(n_1325),
.B2(n_1320),
.Y(n_1400)
);

AND2x2_ASAP7_75t_L g1401 ( 
.A(n_1321),
.B(n_1316),
.Y(n_1401)
);

AND2x2_ASAP7_75t_L g1402 ( 
.A(n_1321),
.B(n_1319),
.Y(n_1402)
);

OR2x2_ASAP7_75t_L g1403 ( 
.A(n_1344),
.B(n_1292),
.Y(n_1403)
);

AND2x2_ASAP7_75t_L g1404 ( 
.A(n_1319),
.B(n_1343),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_L g1405 ( 
.A(n_1313),
.B(n_1311),
.Y(n_1405)
);

AND2x2_ASAP7_75t_L g1406 ( 
.A(n_1297),
.B(n_1311),
.Y(n_1406)
);

OR2x2_ASAP7_75t_L g1407 ( 
.A(n_1292),
.B(n_1294),
.Y(n_1407)
);

A2O1A1Ixp33_ASAP7_75t_L g1408 ( 
.A1(n_1361),
.A2(n_1324),
.B(n_1322),
.C(n_1329),
.Y(n_1408)
);

AND2x2_ASAP7_75t_L g1409 ( 
.A(n_1312),
.B(n_1332),
.Y(n_1409)
);

NOR2xp33_ASAP7_75t_L g1410 ( 
.A(n_1310),
.B(n_1335),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1301),
.Y(n_1411)
);

OAI21xp5_ASAP7_75t_L g1412 ( 
.A1(n_1313),
.A2(n_1348),
.B(n_1357),
.Y(n_1412)
);

OAI22xp5_ASAP7_75t_SL g1413 ( 
.A1(n_1304),
.A2(n_1352),
.B1(n_1356),
.B2(n_1357),
.Y(n_1413)
);

OR2x2_ASAP7_75t_L g1414 ( 
.A(n_1403),
.B(n_1327),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_L g1415 ( 
.A(n_1398),
.B(n_1401),
.Y(n_1415)
);

INVxp67_ASAP7_75t_SL g1416 ( 
.A(n_1398),
.Y(n_1416)
);

INVx2_ASAP7_75t_L g1417 ( 
.A(n_1406),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1407),
.Y(n_1418)
);

INVxp67_ASAP7_75t_SL g1419 ( 
.A(n_1401),
.Y(n_1419)
);

OAI222xp33_ASAP7_75t_L g1420 ( 
.A1(n_1390),
.A2(n_1326),
.B1(n_1362),
.B2(n_1323),
.C1(n_1320),
.C2(n_1333),
.Y(n_1420)
);

NOR2x1_ASAP7_75t_L g1421 ( 
.A(n_1399),
.B(n_1405),
.Y(n_1421)
);

BUFx2_ASAP7_75t_L g1422 ( 
.A(n_1367),
.Y(n_1422)
);

AOI22xp33_ASAP7_75t_L g1423 ( 
.A1(n_1366),
.A2(n_1326),
.B1(n_1325),
.B2(n_1362),
.Y(n_1423)
);

OR2x2_ASAP7_75t_L g1424 ( 
.A(n_1403),
.B(n_1327),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_L g1425 ( 
.A(n_1402),
.B(n_1302),
.Y(n_1425)
);

INVx2_ASAP7_75t_L g1426 ( 
.A(n_1411),
.Y(n_1426)
);

INVx2_ASAP7_75t_L g1427 ( 
.A(n_1411),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_L g1428 ( 
.A(n_1402),
.B(n_1302),
.Y(n_1428)
);

AND2x2_ASAP7_75t_L g1429 ( 
.A(n_1393),
.B(n_1293),
.Y(n_1429)
);

AND2x2_ASAP7_75t_L g1430 ( 
.A(n_1393),
.B(n_1293),
.Y(n_1430)
);

OAI22xp5_ASAP7_75t_L g1431 ( 
.A1(n_1397),
.A2(n_1340),
.B1(n_1347),
.B2(n_1332),
.Y(n_1431)
);

HB1xp67_ASAP7_75t_L g1432 ( 
.A(n_1404),
.Y(n_1432)
);

AND2x2_ASAP7_75t_L g1433 ( 
.A(n_1395),
.B(n_1293),
.Y(n_1433)
);

AND2x2_ASAP7_75t_L g1434 ( 
.A(n_1395),
.B(n_1295),
.Y(n_1434)
);

AND2x2_ASAP7_75t_L g1435 ( 
.A(n_1396),
.B(n_1295),
.Y(n_1435)
);

OR2x2_ASAP7_75t_L g1436 ( 
.A(n_1396),
.B(n_1330),
.Y(n_1436)
);

AOI22xp33_ASAP7_75t_L g1437 ( 
.A1(n_1386),
.A2(n_1341),
.B1(n_1333),
.B2(n_1332),
.Y(n_1437)
);

INVx4_ASAP7_75t_L g1438 ( 
.A(n_1367),
.Y(n_1438)
);

HB1xp67_ASAP7_75t_L g1439 ( 
.A(n_1388),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_L g1440 ( 
.A(n_1394),
.B(n_1368),
.Y(n_1440)
);

INVx2_ASAP7_75t_L g1441 ( 
.A(n_1417),
.Y(n_1441)
);

AND2x2_ASAP7_75t_L g1442 ( 
.A(n_1434),
.B(n_1391),
.Y(n_1442)
);

AOI21xp5_ASAP7_75t_L g1443 ( 
.A1(n_1416),
.A2(n_1340),
.B(n_1389),
.Y(n_1443)
);

INVx4_ASAP7_75t_L g1444 ( 
.A(n_1438),
.Y(n_1444)
);

NAND3xp33_ASAP7_75t_L g1445 ( 
.A(n_1439),
.B(n_1408),
.C(n_1371),
.Y(n_1445)
);

AOI22xp33_ASAP7_75t_SL g1446 ( 
.A1(n_1431),
.A2(n_1376),
.B1(n_1367),
.B2(n_1413),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1426),
.Y(n_1447)
);

NOR2xp33_ASAP7_75t_L g1448 ( 
.A(n_1439),
.B(n_1317),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1426),
.Y(n_1449)
);

INVx4_ASAP7_75t_L g1450 ( 
.A(n_1438),
.Y(n_1450)
);

NAND2xp5_ASAP7_75t_L g1451 ( 
.A(n_1425),
.B(n_1385),
.Y(n_1451)
);

OAI33xp33_ASAP7_75t_L g1452 ( 
.A1(n_1415),
.A2(n_1375),
.A3(n_1372),
.B1(n_1338),
.B2(n_1342),
.B3(n_1339),
.Y(n_1452)
);

OAI321xp33_ASAP7_75t_L g1453 ( 
.A1(n_1423),
.A2(n_1400),
.A3(n_1412),
.B1(n_1369),
.B2(n_1374),
.C(n_1376),
.Y(n_1453)
);

OAI221xp5_ASAP7_75t_L g1454 ( 
.A1(n_1423),
.A2(n_1369),
.B1(n_1380),
.B2(n_1373),
.C(n_1383),
.Y(n_1454)
);

AOI221xp5_ASAP7_75t_SL g1455 ( 
.A1(n_1416),
.A2(n_1383),
.B1(n_1365),
.B2(n_1382),
.C(n_1384),
.Y(n_1455)
);

AOI33xp33_ASAP7_75t_L g1456 ( 
.A1(n_1429),
.A2(n_1382),
.A3(n_1365),
.B1(n_1379),
.B2(n_1330),
.B3(n_1339),
.Y(n_1456)
);

AND2x4_ASAP7_75t_L g1457 ( 
.A(n_1422),
.B(n_1438),
.Y(n_1457)
);

AND2x2_ASAP7_75t_L g1458 ( 
.A(n_1432),
.B(n_1370),
.Y(n_1458)
);

INVx2_ASAP7_75t_L g1459 ( 
.A(n_1417),
.Y(n_1459)
);

NOR2xp33_ASAP7_75t_L g1460 ( 
.A(n_1436),
.B(n_1317),
.Y(n_1460)
);

INVx2_ASAP7_75t_L g1461 ( 
.A(n_1417),
.Y(n_1461)
);

INVx3_ASAP7_75t_L g1462 ( 
.A(n_1422),
.Y(n_1462)
);

BUFx6f_ASAP7_75t_L g1463 ( 
.A(n_1422),
.Y(n_1463)
);

OAI31xp33_ASAP7_75t_L g1464 ( 
.A1(n_1431),
.A2(n_1391),
.A3(n_1333),
.B(n_1350),
.Y(n_1464)
);

AND2x2_ASAP7_75t_L g1465 ( 
.A(n_1434),
.B(n_1435),
.Y(n_1465)
);

AND2x2_ASAP7_75t_L g1466 ( 
.A(n_1434),
.B(n_1391),
.Y(n_1466)
);

NAND2xp5_ASAP7_75t_L g1467 ( 
.A(n_1425),
.B(n_1409),
.Y(n_1467)
);

HB1xp67_ASAP7_75t_L g1468 ( 
.A(n_1427),
.Y(n_1468)
);

HB1xp67_ASAP7_75t_L g1469 ( 
.A(n_1427),
.Y(n_1469)
);

AND2x2_ASAP7_75t_L g1470 ( 
.A(n_1432),
.B(n_1370),
.Y(n_1470)
);

INVx4_ASAP7_75t_L g1471 ( 
.A(n_1438),
.Y(n_1471)
);

AND2x2_ASAP7_75t_L g1472 ( 
.A(n_1435),
.B(n_1391),
.Y(n_1472)
);

NOR2xp33_ASAP7_75t_L g1473 ( 
.A(n_1436),
.B(n_1387),
.Y(n_1473)
);

OR2x2_ASAP7_75t_L g1474 ( 
.A(n_1451),
.B(n_1442),
.Y(n_1474)
);

BUFx2_ASAP7_75t_L g1475 ( 
.A(n_1457),
.Y(n_1475)
);

INVx1_ASAP7_75t_SL g1476 ( 
.A(n_1448),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1468),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1468),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1469),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1469),
.Y(n_1480)
);

AND2x4_ASAP7_75t_L g1481 ( 
.A(n_1457),
.B(n_1438),
.Y(n_1481)
);

BUFx3_ASAP7_75t_L g1482 ( 
.A(n_1463),
.Y(n_1482)
);

OR2x2_ASAP7_75t_L g1483 ( 
.A(n_1451),
.B(n_1428),
.Y(n_1483)
);

NOR2xp33_ASAP7_75t_L g1484 ( 
.A(n_1473),
.B(n_1352),
.Y(n_1484)
);

NOR2xp67_ASAP7_75t_L g1485 ( 
.A(n_1462),
.B(n_1435),
.Y(n_1485)
);

NAND2xp5_ASAP7_75t_SL g1486 ( 
.A(n_1455),
.B(n_1421),
.Y(n_1486)
);

INVx2_ASAP7_75t_L g1487 ( 
.A(n_1441),
.Y(n_1487)
);

NAND2x1p5_ASAP7_75t_SL g1488 ( 
.A(n_1442),
.B(n_1421),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1447),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1447),
.Y(n_1490)
);

OR2x2_ASAP7_75t_L g1491 ( 
.A(n_1442),
.B(n_1428),
.Y(n_1491)
);

AND2x2_ASAP7_75t_L g1492 ( 
.A(n_1466),
.B(n_1429),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_L g1493 ( 
.A(n_1456),
.B(n_1440),
.Y(n_1493)
);

AND2x2_ASAP7_75t_L g1494 ( 
.A(n_1466),
.B(n_1429),
.Y(n_1494)
);

NAND2xp33_ASAP7_75t_R g1495 ( 
.A(n_1462),
.B(n_1358),
.Y(n_1495)
);

INVx2_ASAP7_75t_L g1496 ( 
.A(n_1441),
.Y(n_1496)
);

OR2x2_ASAP7_75t_L g1497 ( 
.A(n_1466),
.B(n_1415),
.Y(n_1497)
);

INVx2_ASAP7_75t_L g1498 ( 
.A(n_1441),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1449),
.Y(n_1499)
);

OR2x2_ASAP7_75t_L g1500 ( 
.A(n_1467),
.B(n_1436),
.Y(n_1500)
);

OR2x2_ASAP7_75t_L g1501 ( 
.A(n_1467),
.B(n_1419),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_L g1502 ( 
.A(n_1455),
.B(n_1445),
.Y(n_1502)
);

AND2x2_ASAP7_75t_L g1503 ( 
.A(n_1472),
.B(n_1430),
.Y(n_1503)
);

AND2x2_ASAP7_75t_L g1504 ( 
.A(n_1472),
.B(n_1465),
.Y(n_1504)
);

AND2x2_ASAP7_75t_L g1505 ( 
.A(n_1465),
.B(n_1430),
.Y(n_1505)
);

NOR2xp67_ASAP7_75t_L g1506 ( 
.A(n_1462),
.B(n_1430),
.Y(n_1506)
);

NAND2xp5_ASAP7_75t_L g1507 ( 
.A(n_1445),
.B(n_1440),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_SL g1508 ( 
.A(n_1446),
.B(n_1433),
.Y(n_1508)
);

INVx4_ASAP7_75t_L g1509 ( 
.A(n_1444),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_L g1510 ( 
.A(n_1458),
.B(n_1433),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_L g1511 ( 
.A(n_1507),
.B(n_1419),
.Y(n_1511)
);

OR2x2_ASAP7_75t_L g1512 ( 
.A(n_1493),
.B(n_1414),
.Y(n_1512)
);

NAND2xp5_ASAP7_75t_L g1513 ( 
.A(n_1502),
.B(n_1433),
.Y(n_1513)
);

OR2x2_ASAP7_75t_L g1514 ( 
.A(n_1474),
.B(n_1414),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1500),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1500),
.Y(n_1516)
);

HB1xp67_ASAP7_75t_L g1517 ( 
.A(n_1477),
.Y(n_1517)
);

OR2x2_ASAP7_75t_L g1518 ( 
.A(n_1474),
.B(n_1414),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1477),
.Y(n_1519)
);

AND2x2_ASAP7_75t_L g1520 ( 
.A(n_1481),
.B(n_1465),
.Y(n_1520)
);

CKINVDCx16_ASAP7_75t_R g1521 ( 
.A(n_1495),
.Y(n_1521)
);

OR2x2_ASAP7_75t_L g1522 ( 
.A(n_1483),
.B(n_1424),
.Y(n_1522)
);

OAI21xp33_ASAP7_75t_L g1523 ( 
.A1(n_1508),
.A2(n_1443),
.B(n_1446),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1478),
.Y(n_1524)
);

INVx2_ASAP7_75t_L g1525 ( 
.A(n_1487),
.Y(n_1525)
);

AND2x2_ASAP7_75t_L g1526 ( 
.A(n_1481),
.B(n_1462),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1478),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1479),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1479),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1480),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_L g1531 ( 
.A(n_1483),
.B(n_1458),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1480),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1489),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1489),
.Y(n_1534)
);

NOR2x1_ASAP7_75t_L g1535 ( 
.A(n_1509),
.B(n_1476),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1490),
.Y(n_1536)
);

AND2x4_ASAP7_75t_L g1537 ( 
.A(n_1509),
.B(n_1481),
.Y(n_1537)
);

OAI22xp5_ASAP7_75t_L g1538 ( 
.A1(n_1486),
.A2(n_1443),
.B1(n_1454),
.B2(n_1463),
.Y(n_1538)
);

INVx3_ASAP7_75t_L g1539 ( 
.A(n_1482),
.Y(n_1539)
);

NOR2x1_ASAP7_75t_L g1540 ( 
.A(n_1509),
.B(n_1352),
.Y(n_1540)
);

OAI22xp5_ASAP7_75t_L g1541 ( 
.A1(n_1497),
.A2(n_1454),
.B1(n_1463),
.B2(n_1471),
.Y(n_1541)
);

INVxp67_ASAP7_75t_L g1542 ( 
.A(n_1475),
.Y(n_1542)
);

AND2x4_ASAP7_75t_L g1543 ( 
.A(n_1509),
.B(n_1457),
.Y(n_1543)
);

NAND2xp5_ASAP7_75t_L g1544 ( 
.A(n_1492),
.B(n_1470),
.Y(n_1544)
);

OR2x2_ASAP7_75t_L g1545 ( 
.A(n_1497),
.B(n_1459),
.Y(n_1545)
);

NAND2xp5_ASAP7_75t_L g1546 ( 
.A(n_1492),
.B(n_1470),
.Y(n_1546)
);

OR2x2_ASAP7_75t_L g1547 ( 
.A(n_1491),
.B(n_1424),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1490),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1499),
.Y(n_1549)
);

OR2x2_ASAP7_75t_L g1550 ( 
.A(n_1491),
.B(n_1424),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1499),
.Y(n_1551)
);

AND2x2_ASAP7_75t_L g1552 ( 
.A(n_1481),
.B(n_1457),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1517),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1517),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1520),
.B(n_1504),
.Y(n_1555)
);

AND2x2_ASAP7_75t_L g1556 ( 
.A(n_1520),
.B(n_1504),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1519),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_L g1558 ( 
.A(n_1513),
.B(n_1494),
.Y(n_1558)
);

INVx2_ASAP7_75t_L g1559 ( 
.A(n_1525),
.Y(n_1559)
);

INVx2_ASAP7_75t_L g1560 ( 
.A(n_1525),
.Y(n_1560)
);

INVxp67_ASAP7_75t_SL g1561 ( 
.A(n_1542),
.Y(n_1561)
);

AND2x2_ASAP7_75t_L g1562 ( 
.A(n_1552),
.B(n_1475),
.Y(n_1562)
);

BUFx2_ASAP7_75t_L g1563 ( 
.A(n_1542),
.Y(n_1563)
);

OR2x2_ASAP7_75t_L g1564 ( 
.A(n_1512),
.B(n_1514),
.Y(n_1564)
);

INVx1_ASAP7_75t_SL g1565 ( 
.A(n_1521),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1552),
.B(n_1526),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1526),
.B(n_1506),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1535),
.B(n_1506),
.Y(n_1568)
);

HB1xp67_ASAP7_75t_L g1569 ( 
.A(n_1524),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1527),
.Y(n_1570)
);

OR2x2_ASAP7_75t_L g1571 ( 
.A(n_1518),
.B(n_1488),
.Y(n_1571)
);

AND2x2_ASAP7_75t_L g1572 ( 
.A(n_1543),
.B(n_1485),
.Y(n_1572)
);

AND2x2_ASAP7_75t_L g1573 ( 
.A(n_1543),
.B(n_1485),
.Y(n_1573)
);

AOI32xp33_ASAP7_75t_L g1574 ( 
.A1(n_1523),
.A2(n_1453),
.A3(n_1494),
.B1(n_1503),
.B2(n_1484),
.Y(n_1574)
);

OR2x2_ASAP7_75t_L g1575 ( 
.A(n_1511),
.B(n_1488),
.Y(n_1575)
);

AOI211x1_ASAP7_75t_SL g1576 ( 
.A1(n_1538),
.A2(n_1488),
.B(n_1510),
.C(n_1463),
.Y(n_1576)
);

INVx1_ASAP7_75t_SL g1577 ( 
.A(n_1540),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_L g1578 ( 
.A(n_1515),
.B(n_1503),
.Y(n_1578)
);

AND2x2_ASAP7_75t_L g1579 ( 
.A(n_1543),
.B(n_1505),
.Y(n_1579)
);

AND3x2_ASAP7_75t_L g1580 ( 
.A(n_1537),
.B(n_1464),
.C(n_1460),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_L g1581 ( 
.A(n_1516),
.B(n_1501),
.Y(n_1581)
);

NOR2xp33_ASAP7_75t_L g1582 ( 
.A(n_1537),
.B(n_1452),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_L g1583 ( 
.A(n_1528),
.B(n_1501),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1529),
.Y(n_1584)
);

INVx4_ASAP7_75t_L g1585 ( 
.A(n_1537),
.Y(n_1585)
);

INVx2_ASAP7_75t_L g1586 ( 
.A(n_1545),
.Y(n_1586)
);

INVx2_ASAP7_75t_L g1587 ( 
.A(n_1545),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1569),
.Y(n_1588)
);

OAI22xp33_ASAP7_75t_L g1589 ( 
.A1(n_1575),
.A2(n_1453),
.B1(n_1541),
.B2(n_1550),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1569),
.Y(n_1590)
);

OAI21xp33_ASAP7_75t_SL g1591 ( 
.A1(n_1574),
.A2(n_1539),
.B(n_1505),
.Y(n_1591)
);

NOR2x1_ASAP7_75t_L g1592 ( 
.A(n_1565),
.B(n_1563),
.Y(n_1592)
);

INVx2_ASAP7_75t_L g1593 ( 
.A(n_1555),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_L g1594 ( 
.A(n_1561),
.B(n_1531),
.Y(n_1594)
);

NOR2x1_ASAP7_75t_L g1595 ( 
.A(n_1565),
.B(n_1356),
.Y(n_1595)
);

AOI22xp5_ASAP7_75t_L g1596 ( 
.A1(n_1582),
.A2(n_1452),
.B1(n_1437),
.B2(n_1367),
.Y(n_1596)
);

AOI22xp33_ASAP7_75t_L g1597 ( 
.A1(n_1580),
.A2(n_1464),
.B1(n_1437),
.B2(n_1367),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_SL g1598 ( 
.A(n_1574),
.B(n_1463),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1553),
.Y(n_1599)
);

AOI22xp5_ASAP7_75t_L g1600 ( 
.A1(n_1582),
.A2(n_1367),
.B1(n_1498),
.B2(n_1496),
.Y(n_1600)
);

AOI211xp5_ASAP7_75t_L g1601 ( 
.A1(n_1575),
.A2(n_1532),
.B(n_1530),
.C(n_1539),
.Y(n_1601)
);

AOI22xp33_ASAP7_75t_SL g1602 ( 
.A1(n_1575),
.A2(n_1463),
.B1(n_1539),
.B2(n_1399),
.Y(n_1602)
);

AND2x2_ASAP7_75t_L g1603 ( 
.A(n_1566),
.B(n_1544),
.Y(n_1603)
);

AOI21xp5_ASAP7_75t_L g1604 ( 
.A1(n_1561),
.A2(n_1551),
.B(n_1534),
.Y(n_1604)
);

AOI22xp5_ASAP7_75t_L g1605 ( 
.A1(n_1580),
.A2(n_1587),
.B1(n_1586),
.B2(n_1559),
.Y(n_1605)
);

NOR2xp33_ASAP7_75t_L g1606 ( 
.A(n_1585),
.B(n_1577),
.Y(n_1606)
);

OR2x6_ASAP7_75t_L g1607 ( 
.A(n_1563),
.B(n_1356),
.Y(n_1607)
);

NOR2xp33_ASAP7_75t_L g1608 ( 
.A(n_1585),
.B(n_1522),
.Y(n_1608)
);

INVx1_ASAP7_75t_SL g1609 ( 
.A(n_1563),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_L g1610 ( 
.A(n_1564),
.B(n_1546),
.Y(n_1610)
);

OAI31xp33_ASAP7_75t_L g1611 ( 
.A1(n_1571),
.A2(n_1420),
.A3(n_1548),
.B(n_1536),
.Y(n_1611)
);

AOI21xp5_ASAP7_75t_L g1612 ( 
.A1(n_1568),
.A2(n_1549),
.B(n_1533),
.Y(n_1612)
);

NOR3xp33_ASAP7_75t_L g1613 ( 
.A(n_1592),
.B(n_1577),
.C(n_1554),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1609),
.Y(n_1614)
);

INVx1_ASAP7_75t_SL g1615 ( 
.A(n_1595),
.Y(n_1615)
);

O2A1O1Ixp33_ASAP7_75t_SL g1616 ( 
.A1(n_1598),
.A2(n_1571),
.B(n_1554),
.C(n_1553),
.Y(n_1616)
);

AOI22xp5_ASAP7_75t_L g1617 ( 
.A1(n_1605),
.A2(n_1587),
.B1(n_1586),
.B2(n_1559),
.Y(n_1617)
);

INVx2_ASAP7_75t_L g1618 ( 
.A(n_1609),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1593),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_1603),
.B(n_1566),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_SL g1621 ( 
.A(n_1589),
.B(n_1568),
.Y(n_1621)
);

OAI22xp5_ASAP7_75t_L g1622 ( 
.A1(n_1596),
.A2(n_1564),
.B1(n_1571),
.B2(n_1558),
.Y(n_1622)
);

INVx2_ASAP7_75t_L g1623 ( 
.A(n_1607),
.Y(n_1623)
);

INVxp67_ASAP7_75t_L g1624 ( 
.A(n_1606),
.Y(n_1624)
);

AOI221xp5_ASAP7_75t_SL g1625 ( 
.A1(n_1591),
.A2(n_1568),
.B1(n_1562),
.B2(n_1576),
.C(n_1581),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1588),
.Y(n_1626)
);

OAI31xp33_ASAP7_75t_L g1627 ( 
.A1(n_1611),
.A2(n_1587),
.A3(n_1586),
.B(n_1576),
.Y(n_1627)
);

AOI22xp5_ASAP7_75t_L g1628 ( 
.A1(n_1600),
.A2(n_1560),
.B1(n_1559),
.B2(n_1558),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_L g1629 ( 
.A(n_1610),
.B(n_1555),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1607),
.B(n_1566),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1607),
.B(n_1562),
.Y(n_1631)
);

A2O1A1Ixp33_ASAP7_75t_L g1632 ( 
.A1(n_1627),
.A2(n_1601),
.B(n_1597),
.C(n_1604),
.Y(n_1632)
);

AOI22xp5_ASAP7_75t_L g1633 ( 
.A1(n_1621),
.A2(n_1608),
.B1(n_1594),
.B2(n_1560),
.Y(n_1633)
);

NAND2xp5_ASAP7_75t_L g1634 ( 
.A(n_1620),
.B(n_1590),
.Y(n_1634)
);

OAI211xp5_ASAP7_75t_L g1635 ( 
.A1(n_1613),
.A2(n_1599),
.B(n_1602),
.C(n_1612),
.Y(n_1635)
);

INVx2_ASAP7_75t_L g1636 ( 
.A(n_1620),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_L g1637 ( 
.A(n_1629),
.B(n_1555),
.Y(n_1637)
);

AOI31xp33_ASAP7_75t_L g1638 ( 
.A1(n_1624),
.A2(n_1562),
.A3(n_1564),
.B(n_1557),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1618),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1618),
.Y(n_1640)
);

O2A1O1Ixp33_ASAP7_75t_L g1641 ( 
.A1(n_1616),
.A2(n_1557),
.B(n_1584),
.C(n_1570),
.Y(n_1641)
);

AOI21xp33_ASAP7_75t_L g1642 ( 
.A1(n_1615),
.A2(n_1560),
.B(n_1570),
.Y(n_1642)
);

NOR2xp33_ASAP7_75t_L g1643 ( 
.A(n_1638),
.B(n_1631),
.Y(n_1643)
);

BUFx2_ASAP7_75t_L g1644 ( 
.A(n_1636),
.Y(n_1644)
);

NAND4xp25_ASAP7_75t_L g1645 ( 
.A(n_1632),
.B(n_1633),
.C(n_1625),
.D(n_1634),
.Y(n_1645)
);

AOI22x1_ASAP7_75t_L g1646 ( 
.A1(n_1639),
.A2(n_1631),
.B1(n_1630),
.B2(n_1614),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_L g1647 ( 
.A(n_1637),
.B(n_1630),
.Y(n_1647)
);

AND2x2_ASAP7_75t_L g1648 ( 
.A(n_1640),
.B(n_1556),
.Y(n_1648)
);

NOR3x1_ASAP7_75t_L g1649 ( 
.A(n_1635),
.B(n_1619),
.C(n_1614),
.Y(n_1649)
);

OA211x2_ASAP7_75t_L g1650 ( 
.A1(n_1635),
.A2(n_1581),
.B(n_1583),
.C(n_1578),
.Y(n_1650)
);

AOI21xp5_ASAP7_75t_L g1651 ( 
.A1(n_1641),
.A2(n_1626),
.B(n_1617),
.Y(n_1651)
);

NAND3xp33_ASAP7_75t_L g1652 ( 
.A(n_1642),
.B(n_1623),
.C(n_1619),
.Y(n_1652)
);

AOI22xp33_ASAP7_75t_L g1653 ( 
.A1(n_1645),
.A2(n_1622),
.B1(n_1628),
.B2(n_1623),
.Y(n_1653)
);

NOR3xp33_ASAP7_75t_L g1654 ( 
.A(n_1652),
.B(n_1626),
.C(n_1585),
.Y(n_1654)
);

AOI322xp5_ASAP7_75t_L g1655 ( 
.A1(n_1643),
.A2(n_1583),
.A3(n_1584),
.B1(n_1578),
.B2(n_1556),
.C1(n_1567),
.C2(n_1572),
.Y(n_1655)
);

AOI211xp5_ASAP7_75t_L g1656 ( 
.A1(n_1651),
.A2(n_1573),
.B(n_1572),
.C(n_1567),
.Y(n_1656)
);

NAND4xp25_ASAP7_75t_L g1657 ( 
.A(n_1649),
.B(n_1585),
.C(n_1573),
.D(n_1572),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1644),
.Y(n_1658)
);

NAND5xp2_ASAP7_75t_SL g1659 ( 
.A(n_1653),
.B(n_1648),
.C(n_1650),
.D(n_1646),
.E(n_1647),
.Y(n_1659)
);

NAND5xp2_ASAP7_75t_SL g1660 ( 
.A(n_1654),
.B(n_1573),
.C(n_1579),
.D(n_1567),
.E(n_1585),
.Y(n_1660)
);

INVx2_ASAP7_75t_SL g1661 ( 
.A(n_1658),
.Y(n_1661)
);

AOI221xp5_ASAP7_75t_L g1662 ( 
.A1(n_1657),
.A2(n_1556),
.B1(n_1579),
.B2(n_1420),
.C(n_1487),
.Y(n_1662)
);

OAI311xp33_ASAP7_75t_L g1663 ( 
.A1(n_1655),
.A2(n_1384),
.A3(n_1579),
.B1(n_1547),
.C1(n_1337),
.Y(n_1663)
);

AND2x2_ASAP7_75t_L g1664 ( 
.A(n_1656),
.B(n_1482),
.Y(n_1664)
);

XOR2xp5_ASAP7_75t_L g1665 ( 
.A(n_1659),
.B(n_1337),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1661),
.Y(n_1666)
);

NOR2xp67_ASAP7_75t_L g1667 ( 
.A(n_1664),
.B(n_1482),
.Y(n_1667)
);

OR2x2_ASAP7_75t_L g1668 ( 
.A(n_1660),
.B(n_1418),
.Y(n_1668)
);

NAND2x1p5_ASAP7_75t_SL g1669 ( 
.A(n_1663),
.B(n_1337),
.Y(n_1669)
);

OR2x2_ASAP7_75t_L g1670 ( 
.A(n_1666),
.B(n_1662),
.Y(n_1670)
);

AO22x1_ASAP7_75t_L g1671 ( 
.A1(n_1665),
.A2(n_1669),
.B1(n_1667),
.B2(n_1668),
.Y(n_1671)
);

OAI21xp33_ASAP7_75t_SL g1672 ( 
.A1(n_1666),
.A2(n_1444),
.B(n_1450),
.Y(n_1672)
);

AOI21xp5_ASAP7_75t_L g1673 ( 
.A1(n_1671),
.A2(n_1392),
.B(n_1410),
.Y(n_1673)
);

AOI22xp5_ASAP7_75t_L g1674 ( 
.A1(n_1673),
.A2(n_1670),
.B1(n_1672),
.B2(n_1487),
.Y(n_1674)
);

OAI21xp33_ASAP7_75t_L g1675 ( 
.A1(n_1674),
.A2(n_1310),
.B(n_1463),
.Y(n_1675)
);

NOR2x1_ASAP7_75t_L g1676 ( 
.A(n_1674),
.B(n_1444),
.Y(n_1676)
);

OAI22x1_ASAP7_75t_L g1677 ( 
.A1(n_1676),
.A2(n_1450),
.B1(n_1444),
.B2(n_1471),
.Y(n_1677)
);

OAI21x1_ASAP7_75t_L g1678 ( 
.A1(n_1675),
.A2(n_1498),
.B(n_1496),
.Y(n_1678)
);

OAI22xp5_ASAP7_75t_SL g1679 ( 
.A1(n_1677),
.A2(n_1360),
.B1(n_1471),
.B2(n_1450),
.Y(n_1679)
);

AOI22xp5_ASAP7_75t_L g1680 ( 
.A1(n_1678),
.A2(n_1450),
.B1(n_1471),
.B2(n_1461),
.Y(n_1680)
);

NAND2x1p5_ASAP7_75t_L g1681 ( 
.A(n_1680),
.B(n_1360),
.Y(n_1681)
);

OAI21xp5_ASAP7_75t_SL g1682 ( 
.A1(n_1681),
.A2(n_1679),
.B(n_1351),
.Y(n_1682)
);

AOI22x1_ASAP7_75t_L g1683 ( 
.A1(n_1682),
.A2(n_1351),
.B1(n_1331),
.B2(n_1309),
.Y(n_1683)
);

OAI221xp5_ASAP7_75t_R g1684 ( 
.A1(n_1683),
.A2(n_1377),
.B1(n_1381),
.B2(n_1391),
.C(n_1459),
.Y(n_1684)
);

AOI211xp5_ASAP7_75t_L g1685 ( 
.A1(n_1684),
.A2(n_1351),
.B(n_1378),
.C(n_1349),
.Y(n_1685)
);


endmodule