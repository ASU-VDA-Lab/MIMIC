module fake_ariane_849_n_219 (n_8, n_24, n_7, n_22, n_1, n_6, n_13, n_20, n_27, n_29, n_17, n_4, n_2, n_18, n_32, n_28, n_9, n_11, n_34, n_26, n_3, n_14, n_0, n_33, n_19, n_30, n_31, n_16, n_5, n_12, n_15, n_21, n_23, n_10, n_25, n_219);

input n_8;
input n_24;
input n_7;
input n_22;
input n_1;
input n_6;
input n_13;
input n_20;
input n_27;
input n_29;
input n_17;
input n_4;
input n_2;
input n_18;
input n_32;
input n_28;
input n_9;
input n_11;
input n_34;
input n_26;
input n_3;
input n_14;
input n_0;
input n_33;
input n_19;
input n_30;
input n_31;
input n_16;
input n_5;
input n_12;
input n_15;
input n_21;
input n_23;
input n_10;
input n_25;

output n_219;

wire n_83;
wire n_56;
wire n_60;
wire n_190;
wire n_170;
wire n_160;
wire n_64;
wire n_179;
wire n_180;
wire n_124;
wire n_119;
wire n_167;
wire n_90;
wire n_195;
wire n_38;
wire n_213;
wire n_47;
wire n_110;
wire n_153;
wire n_197;
wire n_86;
wire n_75;
wire n_89;
wire n_67;
wire n_176;
wire n_149;
wire n_158;
wire n_172;
wire n_69;
wire n_95;
wire n_175;
wire n_92;
wire n_143;
wire n_183;
wire n_203;
wire n_150;
wire n_98;
wire n_74;
wire n_113;
wire n_114;
wire n_40;
wire n_181;
wire n_152;
wire n_120;
wire n_169;
wire n_106;
wire n_53;
wire n_173;
wire n_111;
wire n_115;
wire n_133;
wire n_66;
wire n_205;
wire n_71;
wire n_109;
wire n_208;
wire n_96;
wire n_156;
wire n_209;
wire n_49;
wire n_174;
wire n_100;
wire n_50;
wire n_187;
wire n_132;
wire n_62;
wire n_210;
wire n_147;
wire n_204;
wire n_200;
wire n_51;
wire n_166;
wire n_76;
wire n_218;
wire n_103;
wire n_79;
wire n_46;
wire n_84;
wire n_36;
wire n_199;
wire n_91;
wire n_159;
wire n_107;
wire n_189;
wire n_72;
wire n_105;
wire n_128;
wire n_217;
wire n_44;
wire n_82;
wire n_178;
wire n_42;
wire n_57;
wire n_131;
wire n_201;
wire n_70;
wire n_117;
wire n_139;
wire n_165;
wire n_85;
wire n_130;
wire n_144;
wire n_214;
wire n_48;
wire n_101;
wire n_94;
wire n_134;
wire n_188;
wire n_185;
wire n_58;
wire n_37;
wire n_65;
wire n_123;
wire n_212;
wire n_138;
wire n_112;
wire n_45;
wire n_162;
wire n_129;
wire n_126;
wire n_137;
wire n_122;
wire n_198;
wire n_148;
wire n_164;
wire n_52;
wire n_157;
wire n_184;
wire n_177;
wire n_135;
wire n_73;
wire n_77;
wire n_171;
wire n_121;
wire n_93;
wire n_118;
wire n_61;
wire n_108;
wire n_102;
wire n_182;
wire n_196;
wire n_125;
wire n_168;
wire n_43;
wire n_81;
wire n_87;
wire n_206;
wire n_207;
wire n_41;
wire n_140;
wire n_55;
wire n_191;
wire n_151;
wire n_136;
wire n_192;
wire n_80;
wire n_146;
wire n_211;
wire n_194;
wire n_97;
wire n_154;
wire n_215;
wire n_142;
wire n_161;
wire n_163;
wire n_88;
wire n_186;
wire n_141;
wire n_68;
wire n_116;
wire n_104;
wire n_202;
wire n_145;
wire n_78;
wire n_193;
wire n_39;
wire n_59;
wire n_63;
wire n_99;
wire n_216;
wire n_155;
wire n_127;
wire n_35;
wire n_54;

CKINVDCx5p33_ASAP7_75t_R g35 ( 
.A(n_34),
.Y(n_35)
);

INVxp33_ASAP7_75t_SL g36 ( 
.A(n_22),
.Y(n_36)
);

INVxp67_ASAP7_75t_SL g37 ( 
.A(n_25),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

INVxp33_ASAP7_75t_SL g39 ( 
.A(n_33),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

INVxp67_ASAP7_75t_SL g41 ( 
.A(n_26),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_4),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_0),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_11),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_8),
.Y(n_49)
);

CKINVDCx5p33_ASAP7_75t_R g50 ( 
.A(n_13),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_5),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_7),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_29),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_31),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_1),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_15),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_30),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_2),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_14),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_2),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_3),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_16),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_23),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

CKINVDCx5p33_ASAP7_75t_R g65 ( 
.A(n_35),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_52),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_58),
.Y(n_68)
);

CKINVDCx5p33_ASAP7_75t_R g69 ( 
.A(n_35),
.Y(n_69)
);

CKINVDCx5p33_ASAP7_75t_R g70 ( 
.A(n_60),
.Y(n_70)
);

CKINVDCx5p33_ASAP7_75t_R g71 ( 
.A(n_50),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_61),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_51),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

CKINVDCx5p33_ASAP7_75t_R g75 ( 
.A(n_50),
.Y(n_75)
);

BUFx2_ASAP7_75t_L g76 ( 
.A(n_51),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_38),
.B(n_0),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_49),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_R g79 ( 
.A(n_48),
.B(n_9),
.Y(n_79)
);

CKINVDCx5p33_ASAP7_75t_R g80 ( 
.A(n_36),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_38),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_49),
.Y(n_82)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_42),
.Y(n_83)
);

OAI21x1_ASAP7_75t_L g84 ( 
.A1(n_42),
.A2(n_24),
.B(n_21),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_R g85 ( 
.A(n_40),
.B(n_18),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_45),
.B(n_1),
.Y(n_86)
);

CKINVDCx5p33_ASAP7_75t_R g87 ( 
.A(n_36),
.Y(n_87)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_57),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_46),
.Y(n_89)
);

INVx3_ASAP7_75t_R g90 ( 
.A(n_76),
.Y(n_90)
);

NAND3xp33_ASAP7_75t_L g91 ( 
.A(n_65),
.B(n_57),
.C(n_62),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_64),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_78),
.A2(n_39),
.B1(n_59),
.B2(n_56),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_66),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_81),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_81),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_71),
.B(n_75),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_74),
.B(n_63),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_67),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_74),
.B(n_54),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_81),
.Y(n_101)
);

AND2x4_ASAP7_75t_L g102 ( 
.A(n_89),
.B(n_47),
.Y(n_102)
);

AND2x4_ASAP7_75t_L g103 ( 
.A(n_82),
.B(n_53),
.Y(n_103)
);

AND2x4_ASAP7_75t_L g104 ( 
.A(n_82),
.B(n_41),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_73),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_80),
.A2(n_55),
.B1(n_39),
.B2(n_37),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_65),
.B(n_55),
.Y(n_107)
);

AND2x4_ASAP7_75t_L g108 ( 
.A(n_83),
.B(n_88),
.Y(n_108)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_81),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_69),
.B(n_3),
.Y(n_110)
);

NOR2x1p5_ASAP7_75t_L g111 ( 
.A(n_70),
.B(n_4),
.Y(n_111)
);

NAND2x1p5_ASAP7_75t_L g112 ( 
.A(n_77),
.B(n_12),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_68),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_98),
.A2(n_86),
.B(n_84),
.Y(n_114)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_96),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_R g116 ( 
.A(n_97),
.B(n_80),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_92),
.Y(n_117)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_95),
.Y(n_118)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_95),
.Y(n_119)
);

CKINVDCx5p33_ASAP7_75t_R g120 ( 
.A(n_105),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_101),
.Y(n_121)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_104),
.Y(n_122)
);

HB1xp67_ASAP7_75t_L g123 ( 
.A(n_107),
.Y(n_123)
);

A2O1A1Ixp33_ASAP7_75t_L g124 ( 
.A1(n_93),
.A2(n_84),
.B(n_72),
.C(n_87),
.Y(n_124)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_109),
.Y(n_125)
);

BUFx2_ASAP7_75t_L g126 ( 
.A(n_105),
.Y(n_126)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_109),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_L g128 ( 
.A1(n_93),
.A2(n_88),
.B1(n_83),
.B2(n_81),
.Y(n_128)
);

AND2x4_ASAP7_75t_L g129 ( 
.A(n_102),
.B(n_83),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_104),
.B(n_69),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_94),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_100),
.B(n_87),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_101),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_104),
.B(n_88),
.Y(n_134)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_121),
.Y(n_135)
);

AND2x6_ASAP7_75t_L g136 ( 
.A(n_129),
.B(n_103),
.Y(n_136)
);

CKINVDCx6p67_ASAP7_75t_R g137 ( 
.A(n_126),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_132),
.B(n_106),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_114),
.A2(n_113),
.B(n_99),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_122),
.A2(n_110),
.B1(n_91),
.B2(n_102),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_117),
.Y(n_141)
);

AND2x2_ASAP7_75t_SL g142 ( 
.A(n_122),
.B(n_110),
.Y(n_142)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_121),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_L g144 ( 
.A1(n_122),
.A2(n_103),
.B1(n_102),
.B2(n_112),
.Y(n_144)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_118),
.Y(n_145)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_118),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_123),
.B(n_100),
.Y(n_147)
);

OAI22xp33_ASAP7_75t_L g148 ( 
.A1(n_130),
.A2(n_131),
.B1(n_112),
.B2(n_134),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_129),
.B(n_103),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_115),
.A2(n_96),
.B(n_108),
.Y(n_150)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_121),
.Y(n_151)
);

BUFx2_ASAP7_75t_SL g152 ( 
.A(n_129),
.Y(n_152)
);

NAND2x1p5_ASAP7_75t_L g153 ( 
.A(n_121),
.B(n_108),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_115),
.A2(n_124),
.B(n_127),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_116),
.A2(n_73),
.B1(n_79),
.B2(n_85),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_115),
.A2(n_96),
.B(n_108),
.Y(n_156)
);

AND2x4_ASAP7_75t_L g157 ( 
.A(n_128),
.B(n_111),
.Y(n_157)
);

CKINVDCx8_ASAP7_75t_R g158 ( 
.A(n_152),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_138),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_142),
.B(n_120),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_142),
.A2(n_124),
.B1(n_120),
.B2(n_125),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_144),
.A2(n_127),
.B1(n_125),
.B2(n_119),
.Y(n_162)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_145),
.Y(n_163)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_145),
.Y(n_164)
);

BUFx2_ASAP7_75t_L g165 ( 
.A(n_137),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_L g166 ( 
.A1(n_157),
.A2(n_116),
.B1(n_119),
.B2(n_133),
.Y(n_166)
);

OAI22xp33_ASAP7_75t_L g167 ( 
.A1(n_140),
.A2(n_133),
.B1(n_96),
.B2(n_7),
.Y(n_167)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_146),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_136),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_136),
.A2(n_133),
.B1(n_90),
.B2(n_6),
.Y(n_170)
);

BUFx10_ASAP7_75t_L g171 ( 
.A(n_157),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_136),
.B(n_133),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_146),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_157),
.A2(n_5),
.B1(n_6),
.B2(n_20),
.Y(n_174)
);

AND2x4_ASAP7_75t_L g175 ( 
.A(n_136),
.B(n_147),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_141),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_149),
.Y(n_177)
);

BUFx2_ASAP7_75t_L g178 ( 
.A(n_137),
.Y(n_178)
);

OR2x2_ASAP7_75t_L g179 ( 
.A(n_155),
.B(n_153),
.Y(n_179)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_153),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_163),
.Y(n_181)
);

HB1xp67_ASAP7_75t_L g182 ( 
.A(n_175),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_175),
.B(n_148),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_171),
.B(n_136),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_L g185 ( 
.A1(n_159),
.A2(n_144),
.B1(n_148),
.B2(n_143),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_L g186 ( 
.A1(n_160),
.A2(n_143),
.B1(n_135),
.B2(n_151),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_177),
.B(n_135),
.Y(n_187)
);

INVx2_ASAP7_75t_SL g188 ( 
.A(n_171),
.Y(n_188)
);

OAI22xp33_ASAP7_75t_L g189 ( 
.A1(n_167),
.A2(n_135),
.B1(n_151),
.B2(n_154),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_164),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_168),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_190),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_185),
.A2(n_169),
.B1(n_179),
.B2(n_167),
.Y(n_193)
);

OAI321xp33_ASAP7_75t_L g194 ( 
.A1(n_183),
.A2(n_161),
.A3(n_170),
.B1(n_166),
.B2(n_174),
.C(n_169),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g195 ( 
.A(n_182),
.B(n_165),
.Y(n_195)
);

OAI221xp5_ASAP7_75t_L g196 ( 
.A1(n_186),
.A2(n_174),
.B1(n_161),
.B2(n_176),
.C(n_158),
.Y(n_196)
);

AND2x4_ASAP7_75t_L g197 ( 
.A(n_184),
.B(n_178),
.Y(n_197)
);

OAI221xp5_ASAP7_75t_L g198 ( 
.A1(n_188),
.A2(n_187),
.B1(n_139),
.B2(n_172),
.C(n_180),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_188),
.B(n_173),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_192),
.B(n_191),
.Y(n_200)
);

INVxp67_ASAP7_75t_SL g201 ( 
.A(n_199),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_193),
.B(n_191),
.Y(n_202)
);

HB1xp67_ASAP7_75t_L g203 ( 
.A(n_195),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_198),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g205 ( 
.A(n_203),
.B(n_197),
.Y(n_205)
);

INVx1_ASAP7_75t_SL g206 ( 
.A(n_200),
.Y(n_206)
);

AOI221xp5_ASAP7_75t_L g207 ( 
.A1(n_206),
.A2(n_204),
.B1(n_196),
.B2(n_194),
.C(n_201),
.Y(n_207)
);

NOR2x1_ASAP7_75t_L g208 ( 
.A(n_205),
.B(n_204),
.Y(n_208)
);

O2A1O1Ixp5_ASAP7_75t_L g209 ( 
.A1(n_208),
.A2(n_205),
.B(n_197),
.C(n_202),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_207),
.A2(n_194),
.B(n_189),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_209),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_211),
.Y(n_212)
);

OAI211xp5_ASAP7_75t_L g213 ( 
.A1(n_212),
.A2(n_210),
.B(n_202),
.C(n_200),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_213),
.A2(n_184),
.B1(n_190),
.B2(n_181),
.Y(n_214)
);

NOR3xp33_ASAP7_75t_L g215 ( 
.A(n_214),
.B(n_150),
.C(n_156),
.Y(n_215)
);

BUFx4f_ASAP7_75t_SL g216 ( 
.A(n_215),
.Y(n_216)
);

INVxp67_ASAP7_75t_SL g217 ( 
.A(n_216),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_217),
.A2(n_181),
.B1(n_172),
.B2(n_151),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_218),
.A2(n_162),
.B(n_217),
.Y(n_219)
);


endmodule