module fake_jpeg_16060_n_343 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_343);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_343;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx10_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx16f_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_13),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_10),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_14),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_16),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_20),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_36),
.B(n_39),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_18),
.B(n_9),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_37),
.B(n_46),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_35),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_20),
.Y(n_39)
);

INVx13_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_45),
.B(n_17),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_20),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_27),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_47),
.B(n_33),
.Y(n_70)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_48),
.Y(n_87)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_51),
.Y(n_94)
);

OAI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_36),
.A2(n_34),
.B1(n_21),
.B2(n_22),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_53),
.A2(n_47),
.B1(n_46),
.B2(n_39),
.Y(n_72)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_54),
.Y(n_76)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_55),
.B(n_57),
.Y(n_80)
);

BUFx2_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_56),
.Y(n_81)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_58),
.B(n_62),
.Y(n_92)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_61),
.Y(n_75)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_64),
.B(n_66),
.Y(n_99)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_65),
.Y(n_82)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_67),
.B(n_70),
.Y(n_96)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_71),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_72),
.A2(n_26),
.B1(n_27),
.B2(n_33),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_59),
.B(n_44),
.C(n_37),
.Y(n_73)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_73),
.B(n_49),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_68),
.B(n_37),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_74),
.B(n_77),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_68),
.B(n_44),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_68),
.B(n_46),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_78),
.B(n_79),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_57),
.B(n_46),
.Y(n_79)
);

INVx1_ASAP7_75t_SL g83 ( 
.A(n_52),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_83),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_71),
.A2(n_31),
.B(n_28),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_84),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_56),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_85),
.B(n_45),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_58),
.B(n_47),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_86),
.B(n_90),
.Y(n_114)
);

INVx2_ASAP7_75t_SL g88 ( 
.A(n_50),
.Y(n_88)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_88),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_62),
.B(n_47),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_66),
.B(n_60),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_91),
.B(n_39),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_60),
.B(n_39),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_93),
.B(n_36),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_63),
.B(n_21),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_95),
.B(n_21),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_50),
.A2(n_64),
.B1(n_55),
.B2(n_54),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_97),
.A2(n_98),
.B1(n_36),
.B2(n_33),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_63),
.A2(n_18),
.B1(n_28),
.B2(n_25),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_77),
.A2(n_18),
.B1(n_25),
.B2(n_28),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_100),
.A2(n_102),
.B1(n_108),
.B2(n_83),
.Y(n_133)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_101),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_74),
.A2(n_25),
.B1(n_45),
.B2(n_34),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_103),
.B(n_126),
.Y(n_148)
);

OR2x4_ASAP7_75t_L g104 ( 
.A(n_78),
.B(n_21),
.Y(n_104)
);

MAJx2_ASAP7_75t_L g130 ( 
.A(n_104),
.B(n_113),
.C(n_84),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_107),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_95),
.A2(n_45),
.B1(n_34),
.B2(n_41),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_96),
.B(n_22),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_112),
.B(n_119),
.Y(n_134)
);

MAJx2_ASAP7_75t_L g113 ( 
.A(n_73),
.B(n_45),
.C(n_31),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_96),
.B(n_0),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_115),
.B(n_116),
.Y(n_143)
);

A2O1A1Ixp33_ASAP7_75t_L g117 ( 
.A1(n_79),
.A2(n_86),
.B(n_90),
.C(n_72),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_117),
.B(n_121),
.Y(n_156)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_91),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_118),
.Y(n_154)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_92),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_81),
.B(n_85),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_120),
.B(n_128),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_95),
.B(n_0),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g147 ( 
.A1(n_122),
.A2(n_125),
.B1(n_30),
.B2(n_29),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_95),
.B(n_97),
.Y(n_123)
);

AND2x2_ASAP7_75t_SL g138 ( 
.A(n_123),
.B(n_98),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_124),
.B(n_92),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_93),
.B(n_69),
.Y(n_126)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_75),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_127),
.B(n_76),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_76),
.Y(n_128)
);

INVx6_ASAP7_75t_L g129 ( 
.A(n_76),
.Y(n_129)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_129),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_130),
.A2(n_138),
.B(n_141),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_105),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_132),
.B(n_142),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_L g168 ( 
.A1(n_133),
.A2(n_147),
.B1(n_94),
.B2(n_87),
.Y(n_168)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_129),
.Y(n_135)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_135),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_109),
.A2(n_118),
.B1(n_114),
.B2(n_111),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_136),
.A2(n_157),
.B1(n_158),
.B2(n_100),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_139),
.B(n_110),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_124),
.B(n_99),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_140),
.B(n_31),
.C(n_17),
.Y(n_186)
);

OA21x2_ASAP7_75t_L g141 ( 
.A1(n_126),
.A2(n_99),
.B(n_80),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_105),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_119),
.B(n_80),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_145),
.B(n_155),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g149 ( 
.A(n_104),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_149),
.B(n_153),
.Y(n_183)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_150),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_127),
.B(n_81),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_151),
.B(n_152),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_116),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_128),
.B(n_88),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_114),
.B(n_89),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_109),
.A2(n_89),
.B1(n_88),
.B2(n_83),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_111),
.A2(n_38),
.B1(n_41),
.B2(n_82),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_154),
.A2(n_123),
.B1(n_102),
.B2(n_117),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_159),
.A2(n_149),
.B1(n_143),
.B2(n_141),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_160),
.B(n_32),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_156),
.A2(n_123),
.B(n_110),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_161),
.A2(n_174),
.B(n_177),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_131),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_163),
.B(n_167),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_138),
.A2(n_113),
.B1(n_107),
.B2(n_121),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_164),
.A2(n_166),
.B1(n_169),
.B2(n_172),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_165),
.B(n_168),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_152),
.A2(n_108),
.B1(n_122),
.B2(n_106),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_144),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_138),
.A2(n_107),
.B1(n_121),
.B2(n_115),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_154),
.A2(n_75),
.B1(n_82),
.B2(n_87),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_155),
.B(n_115),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_148),
.B(n_38),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_176),
.B(n_185),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_156),
.A2(n_27),
.B(n_26),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_139),
.B(n_49),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_178),
.B(n_179),
.C(n_186),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_140),
.B(n_31),
.Y(n_179)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_137),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_180),
.B(n_188),
.Y(n_201)
);

AND2x4_ASAP7_75t_L g181 ( 
.A(n_141),
.B(n_48),
.Y(n_181)
);

XNOR2x1_ASAP7_75t_L g199 ( 
.A(n_181),
.B(n_141),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_130),
.A2(n_94),
.B1(n_65),
.B2(n_61),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_182),
.A2(n_187),
.B1(n_41),
.B2(n_38),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_148),
.B(n_136),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_138),
.A2(n_51),
.B1(n_38),
.B2(n_41),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_144),
.Y(n_188)
);

XOR2x2_ASAP7_75t_L g189 ( 
.A(n_175),
.B(n_130),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_SL g237 ( 
.A(n_189),
.B(n_208),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_192),
.A2(n_199),
.B1(n_200),
.B2(n_204),
.Y(n_244)
);

OR2x2_ASAP7_75t_L g193 ( 
.A(n_181),
.B(n_137),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_193),
.B(n_215),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_178),
.B(n_143),
.C(n_158),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_194),
.B(n_207),
.C(n_209),
.Y(n_219)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_170),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_197),
.B(n_206),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_175),
.A2(n_145),
.B(n_142),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_180),
.B(n_134),
.Y(n_202)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_202),
.Y(n_223)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_171),
.Y(n_203)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_203),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_181),
.A2(n_146),
.B1(n_132),
.B2(n_133),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_181),
.A2(n_157),
.B1(n_134),
.B2(n_135),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_205),
.A2(n_183),
.B1(n_177),
.B2(n_169),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_182),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_160),
.B(n_31),
.Y(n_207)
);

MAJx2_ASAP7_75t_L g208 ( 
.A(n_179),
.B(n_31),
.C(n_32),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_164),
.B(n_17),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_173),
.B(n_131),
.Y(n_211)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_211),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g212 ( 
.A(n_184),
.Y(n_212)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_212),
.Y(n_234)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_213),
.Y(n_238)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_162),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_214),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_173),
.B(n_17),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_162),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_216),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_217),
.B(n_165),
.C(n_187),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_191),
.B(n_186),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_218),
.B(n_224),
.C(n_228),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_189),
.B(n_161),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_220),
.B(n_32),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_191),
.B(n_185),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_211),
.B(n_176),
.Y(n_226)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_226),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_229),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_210),
.B(n_174),
.Y(n_231)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_231),
.Y(n_261)
);

OA21x2_ASAP7_75t_SL g232 ( 
.A1(n_199),
.A2(n_174),
.B(n_166),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_SL g264 ( 
.A1(n_232),
.A2(n_19),
.B(n_30),
.Y(n_264)
);

HB1xp67_ASAP7_75t_L g233 ( 
.A(n_198),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_233),
.B(n_236),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_200),
.B(n_172),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_235),
.B(n_239),
.C(n_194),
.Y(n_252)
);

HB1xp67_ASAP7_75t_L g236 ( 
.A(n_215),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_217),
.B(n_163),
.C(n_41),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_206),
.A2(n_26),
.B1(n_69),
.B2(n_52),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_240),
.A2(n_241),
.B1(n_29),
.B2(n_23),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_195),
.A2(n_210),
.B1(n_196),
.B2(n_204),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_201),
.B(n_19),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_243),
.B(n_19),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g245 ( 
.A1(n_221),
.A2(n_193),
.B(n_205),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_SL g276 ( 
.A(n_245),
.B(n_264),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_222),
.A2(n_190),
.B(n_192),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g273 ( 
.A1(n_248),
.A2(n_266),
.B(n_222),
.Y(n_273)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_223),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_249),
.B(n_260),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_252),
.B(n_239),
.Y(n_274)
);

OAI22x1_ASAP7_75t_L g253 ( 
.A1(n_244),
.A2(n_213),
.B1(n_196),
.B2(n_190),
.Y(n_253)
);

XNOR2x1_ASAP7_75t_L g283 ( 
.A(n_253),
.B(n_256),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_254),
.B(n_255),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_227),
.B(n_209),
.Y(n_255)
);

XNOR2x1_ASAP7_75t_L g256 ( 
.A(n_220),
.B(n_207),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_218),
.B(n_208),
.C(n_38),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_257),
.B(n_259),
.C(n_228),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_238),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_258),
.B(n_240),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_224),
.B(n_17),
.C(n_35),
.Y(n_259)
);

HB1xp67_ASAP7_75t_L g260 ( 
.A(n_234),
.Y(n_260)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_225),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_262),
.B(n_230),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_263),
.B(n_265),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_219),
.B(n_32),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_SL g266 ( 
.A1(n_242),
.A2(n_30),
.B1(n_29),
.B2(n_23),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_267),
.B(n_23),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_265),
.B(n_219),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_270),
.B(n_275),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_267),
.B(n_241),
.Y(n_271)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_271),
.Y(n_290)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_272),
.Y(n_292)
);

OR2x2_ASAP7_75t_L g297 ( 
.A(n_273),
.B(n_258),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_274),
.B(n_277),
.C(n_278),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_250),
.B(n_237),
.C(n_235),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_250),
.B(n_237),
.C(n_231),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_279),
.B(n_281),
.C(n_257),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_247),
.B(n_229),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_280),
.B(n_282),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_252),
.B(n_226),
.C(n_35),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_259),
.B(n_10),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_285),
.B(n_245),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_283),
.A2(n_253),
.B1(n_248),
.B2(n_261),
.Y(n_286)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_286),
.Y(n_306)
);

AND2x2_ASAP7_75t_L g289 ( 
.A(n_283),
.B(n_246),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_289),
.B(n_295),
.Y(n_311)
);

HB1xp67_ASAP7_75t_L g291 ( 
.A(n_281),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_291),
.B(n_296),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_L g293 ( 
.A1(n_279),
.A2(n_277),
.B(n_278),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_293),
.A2(n_274),
.B(n_284),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g295 ( 
.A(n_268),
.Y(n_295)
);

HB1xp67_ASAP7_75t_L g296 ( 
.A(n_269),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_297),
.B(n_299),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_284),
.B(n_251),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_298),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_300),
.B(n_263),
.C(n_276),
.Y(n_302)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_301),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_302),
.B(n_311),
.C(n_304),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_294),
.B(n_276),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_303),
.B(n_307),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_294),
.B(n_256),
.C(n_10),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_305),
.B(n_309),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_290),
.A2(n_16),
.B1(n_15),
.B2(n_14),
.Y(n_307)
);

HB1xp67_ASAP7_75t_L g308 ( 
.A(n_287),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_308),
.B(n_313),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_300),
.B(n_16),
.C(n_13),
.Y(n_309)
);

A2O1A1Ixp33_ASAP7_75t_SL g312 ( 
.A1(n_297),
.A2(n_1),
.B(n_2),
.C(n_3),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_L g324 ( 
.A1(n_312),
.A2(n_1),
.B(n_2),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_295),
.B(n_13),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_310),
.A2(n_292),
.B1(n_289),
.B2(n_288),
.Y(n_317)
);

OR2x2_ASAP7_75t_L g329 ( 
.A(n_317),
.B(n_320),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_304),
.B(n_12),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_321),
.B(n_322),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_SL g322 ( 
.A(n_314),
.B(n_11),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_311),
.A2(n_11),
.B(n_2),
.Y(n_323)
);

OAI321xp33_ASAP7_75t_L g331 ( 
.A1(n_323),
.A2(n_324),
.A3(n_4),
.B1(n_5),
.B2(n_6),
.C(n_7),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_316),
.A2(n_306),
.B1(n_312),
.B2(n_5),
.Y(n_325)
);

INVxp67_ASAP7_75t_L g333 ( 
.A(n_325),
.Y(n_333)
);

AOI21x1_ASAP7_75t_L g326 ( 
.A1(n_319),
.A2(n_312),
.B(n_4),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_L g337 ( 
.A1(n_326),
.A2(n_327),
.B(n_5),
.Y(n_337)
);

AOI21x1_ASAP7_75t_L g327 ( 
.A1(n_315),
.A2(n_3),
.B(n_4),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_320),
.B(n_3),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_328),
.B(n_331),
.Y(n_335)
);

OAI21x1_ASAP7_75t_L g332 ( 
.A1(n_316),
.A2(n_4),
.B(n_5),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_SL g336 ( 
.A(n_332),
.B(n_7),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_329),
.B(n_318),
.C(n_6),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_334),
.B(n_336),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_SL g339 ( 
.A1(n_337),
.A2(n_330),
.B(n_6),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_SL g340 ( 
.A1(n_339),
.A2(n_335),
.B(n_338),
.Y(n_340)
);

AOI21xp5_ASAP7_75t_SL g341 ( 
.A1(n_340),
.A2(n_333),
.B(n_7),
.Y(n_341)
);

AND2x2_ASAP7_75t_L g342 ( 
.A(n_341),
.B(n_7),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_342),
.Y(n_343)
);


endmodule