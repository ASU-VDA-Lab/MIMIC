module fake_jpeg_2149_n_86 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_86);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_86;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

INVx6_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_19),
.Y(n_27)
);

INVx11_ASAP7_75t_SL g28 ( 
.A(n_3),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_21),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_20),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_18),
.B(n_10),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_15),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_34),
.B(n_36),
.Y(n_39)
);

BUFx10_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_35),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_31),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_37),
.B(n_32),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_L g40 ( 
.A1(n_33),
.A2(n_26),
.B1(n_29),
.B2(n_32),
.Y(n_40)
);

OR2x2_ASAP7_75t_L g50 ( 
.A(n_40),
.B(n_43),
.Y(n_50)
);

AO22x1_ASAP7_75t_SL g41 ( 
.A1(n_35),
.A2(n_30),
.B1(n_27),
.B2(n_29),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_41),
.B(n_42),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_36),
.B(n_30),
.Y(n_42)
);

INVx13_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

HB1xp67_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_42),
.B(n_27),
.C(n_35),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_47),
.B(n_52),
.Y(n_58)
);

OAI21xp5_ASAP7_75t_L g48 ( 
.A1(n_43),
.A2(n_34),
.B(n_35),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_L g57 ( 
.A1(n_48),
.A2(n_49),
.B(n_0),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_41),
.B(n_0),
.Y(n_49)
);

AND2x6_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_24),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_SL g55 ( 
.A1(n_51),
.A2(n_39),
.B(n_44),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_SL g64 ( 
.A1(n_55),
.A2(n_56),
.B(n_57),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_49),
.A2(n_44),
.B1(n_38),
.B2(n_11),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_47),
.B(n_1),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_59),
.B(n_61),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g60 ( 
.A1(n_45),
.A2(n_1),
.B(n_2),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_SL g68 ( 
.A1(n_60),
.A2(n_4),
.B(n_5),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_50),
.B(n_2),
.Y(n_61)
);

O2A1O1Ixp33_ASAP7_75t_L g62 ( 
.A1(n_54),
.A2(n_52),
.B(n_50),
.C(n_46),
.Y(n_62)
);

AOI221xp5_ASAP7_75t_L g73 ( 
.A1(n_62),
.A2(n_14),
.B1(n_22),
.B2(n_17),
.C(n_16),
.Y(n_73)
);

XNOR2xp5_ASAP7_75t_L g63 ( 
.A(n_58),
.B(n_12),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_63),
.B(n_68),
.C(n_69),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_54),
.B(n_3),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_65),
.B(n_67),
.Y(n_76)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_53),
.Y(n_66)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_66),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_56),
.B(n_4),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_59),
.B(n_5),
.Y(n_69)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_73),
.Y(n_78)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_62),
.Y(n_74)
);

XNOR2xp5_ASAP7_75t_L g79 ( 
.A(n_74),
.B(n_75),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_63),
.B(n_13),
.C(n_23),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_71),
.A2(n_64),
.B1(n_70),
.B2(n_9),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_77),
.A2(n_72),
.B1(n_76),
.B2(n_73),
.Y(n_80)
);

HB1xp67_ASAP7_75t_L g81 ( 
.A(n_80),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_81),
.B(n_79),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_SL g83 ( 
.A1(n_82),
.A2(n_77),
.B(n_78),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_83),
.A2(n_6),
.B(n_8),
.Y(n_84)
);

OAI21xp33_ASAP7_75t_L g85 ( 
.A1(n_84),
.A2(n_6),
.B(n_8),
.Y(n_85)
);

XOR2xp5_ASAP7_75t_L g86 ( 
.A(n_85),
.B(n_9),
.Y(n_86)
);


endmodule