module fake_jpeg_110_n_132 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_132);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_132;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_26),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_27),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_16),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_8),
.Y(n_41)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

BUFx16f_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_10),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_6),
.B(n_21),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_5),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_49),
.Y(n_58)
);

BUFx4f_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_50),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_51),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_42),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_52)
);

AOI21xp5_ASAP7_75t_L g65 ( 
.A1(n_52),
.A2(n_46),
.B(n_41),
.Y(n_65)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_53),
.Y(n_61)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_54),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_55),
.B(n_40),
.Y(n_56)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_49),
.B(n_48),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_57),
.B(n_63),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_51),
.B(n_46),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_53),
.B(n_48),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_64),
.B(n_55),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_65),
.A2(n_50),
.B1(n_41),
.B2(n_36),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_65),
.A2(n_54),
.B1(n_35),
.B2(n_47),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_66),
.A2(n_72),
.B1(n_60),
.B2(n_62),
.Y(n_90)
);

INVx13_ASAP7_75t_L g67 ( 
.A(n_59),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_67),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_63),
.B(n_37),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_69),
.B(n_73),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_70),
.B(n_76),
.Y(n_82)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_59),
.Y(n_71)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_71),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_58),
.A2(n_47),
.B1(n_36),
.B2(n_44),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_58),
.B(n_46),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_61),
.B(n_44),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_75),
.B(n_77),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_61),
.B(n_39),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_L g78 ( 
.A1(n_68),
.A2(n_45),
.B(n_39),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_78),
.B(n_4),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_74),
.B(n_38),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_79),
.B(n_86),
.Y(n_93)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_71),
.Y(n_80)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_80),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_73),
.B(n_76),
.C(n_66),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_83),
.B(n_89),
.C(n_18),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_72),
.B(n_0),
.Y(n_86)
);

AND2x2_ASAP7_75t_SL g88 ( 
.A(n_67),
.B(n_55),
.Y(n_88)
);

CKINVDCx14_ASAP7_75t_R g94 ( 
.A(n_88),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_68),
.B(n_60),
.C(n_50),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_90),
.B(n_3),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_81),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_91),
.B(n_96),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_82),
.A2(n_55),
.B(n_62),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_92),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_82),
.A2(n_60),
.B(n_2),
.Y(n_95)
);

INVx1_ASAP7_75t_SL g109 ( 
.A(n_95),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_84),
.B(n_1),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_81),
.A2(n_3),
.B(n_4),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_97),
.A2(n_103),
.B1(n_85),
.B2(n_87),
.Y(n_105)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_87),
.Y(n_99)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_99),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g100 ( 
.A(n_89),
.B(n_19),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_100),
.B(n_101),
.C(n_15),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_88),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_102),
.B(n_104),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_105),
.A2(n_7),
.B(n_9),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_95),
.A2(n_94),
.B1(n_101),
.B2(n_92),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_110),
.A2(n_114),
.B1(n_97),
.B2(n_9),
.Y(n_119)
);

AOI322xp5_ASAP7_75t_L g111 ( 
.A1(n_100),
.A2(n_22),
.A3(n_33),
.B1(n_32),
.B2(n_31),
.C1(n_30),
.C2(n_29),
.Y(n_111)
);

A2O1A1O1Ixp25_ASAP7_75t_L g120 ( 
.A1(n_111),
.A2(n_116),
.B(n_106),
.C(n_23),
.D(n_34),
.Y(n_120)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_98),
.Y(n_112)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_112),
.Y(n_122)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_99),
.Y(n_113)
);

HB1xp67_ASAP7_75t_L g117 ( 
.A(n_113),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_93),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_115),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_118),
.B(n_119),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_120),
.A2(n_121),
.B(n_116),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_122),
.A2(n_109),
.B1(n_107),
.B2(n_108),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_124),
.B(n_125),
.Y(n_126)
);

AOI31xp67_ASAP7_75t_L g127 ( 
.A1(n_124),
.A2(n_109),
.A3(n_107),
.B(n_117),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_127),
.A2(n_123),
.B1(n_117),
.B2(n_12),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_128),
.B(n_126),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_129),
.A2(n_14),
.B1(n_20),
.B2(n_24),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_130),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_131),
.B(n_11),
.Y(n_132)
);


endmodule