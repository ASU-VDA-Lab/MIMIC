module real_aes_8231_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_551;
wire n_320;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_363;
wire n_182;
wire n_754;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_527;
wire n_434;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_617;
wire n_552;
wire n_602;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_756;
wire n_147;
wire n_288;
wire n_404;
wire n_713;
wire n_598;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_217;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_765;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g105 ( .A(n_0), .Y(n_105) );
INVx1_ASAP7_75t_L g481 ( .A(n_1), .Y(n_481) );
INVx1_ASAP7_75t_L g194 ( .A(n_2), .Y(n_194) );
AOI22xp33_ASAP7_75t_L g526 ( .A1(n_3), .A2(n_38), .B1(n_155), .B2(n_511), .Y(n_526) );
AOI21xp33_ASAP7_75t_L g162 ( .A1(n_4), .A2(n_136), .B(n_163), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_5), .B(n_129), .Y(n_494) );
AND2x6_ASAP7_75t_L g141 ( .A(n_6), .B(n_142), .Y(n_141) );
AOI21xp5_ASAP7_75t_L g243 ( .A1(n_7), .A2(n_244), .B(n_245), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g110 ( .A(n_8), .B(n_111), .Y(n_110) );
NOR2xp33_ASAP7_75t_L g450 ( .A(n_8), .B(n_39), .Y(n_450) );
INVx1_ASAP7_75t_L g169 ( .A(n_9), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_10), .B(n_236), .Y(n_235) );
INVx1_ASAP7_75t_L g134 ( .A(n_11), .Y(n_134) );
INVx1_ASAP7_75t_L g475 ( .A(n_12), .Y(n_475) );
INVx1_ASAP7_75t_L g250 ( .A(n_13), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_14), .B(n_177), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_15), .B(n_130), .Y(n_552) );
AO32x2_ASAP7_75t_L g524 ( .A1(n_16), .A2(n_129), .A3(n_174), .B1(n_503), .B2(n_525), .Y(n_524) );
OAI22xp5_ASAP7_75t_L g118 ( .A1(n_17), .A2(n_119), .B1(n_120), .B2(n_445), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_17), .Y(n_119) );
NAND2xp5_ASAP7_75t_SL g521 ( .A(n_18), .B(n_155), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_19), .B(n_150), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_20), .B(n_130), .Y(n_484) );
AOI22xp33_ASAP7_75t_L g527 ( .A1(n_21), .A2(n_50), .B1(n_155), .B2(n_511), .Y(n_527) );
NAND2xp5_ASAP7_75t_SL g206 ( .A(n_22), .B(n_136), .Y(n_206) );
AOI22xp33_ASAP7_75t_SL g512 ( .A1(n_23), .A2(n_75), .B1(n_155), .B2(n_177), .Y(n_512) );
NAND2xp5_ASAP7_75t_SL g539 ( .A(n_24), .B(n_155), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_25), .B(n_158), .Y(n_157) );
A2O1A1Ixp33_ASAP7_75t_L g247 ( .A1(n_26), .A2(n_248), .B(n_249), .C(n_251), .Y(n_247) );
CKINVDCx20_ASAP7_75t_R g453 ( .A(n_27), .Y(n_453) );
BUFx6f_ASAP7_75t_L g140 ( .A(n_28), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_29), .B(n_171), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_30), .B(n_167), .Y(n_196) );
INVx1_ASAP7_75t_L g183 ( .A(n_31), .Y(n_183) );
AOI22xp33_ASAP7_75t_L g99 ( .A1(n_32), .A2(n_100), .B1(n_112), .B2(n_767), .Y(n_99) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_33), .B(n_171), .Y(n_541) );
INVx2_ASAP7_75t_L g139 ( .A(n_34), .Y(n_139) );
NAND2xp5_ASAP7_75t_SL g498 ( .A(n_35), .B(n_155), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_36), .B(n_171), .Y(n_523) );
A2O1A1Ixp33_ASAP7_75t_L g207 ( .A1(n_37), .A2(n_141), .B(n_145), .C(n_208), .Y(n_207) );
INVx1_ASAP7_75t_L g111 ( .A(n_39), .Y(n_111) );
INVx1_ASAP7_75t_L g181 ( .A(n_40), .Y(n_181) );
NAND2xp5_ASAP7_75t_SL g222 ( .A(n_41), .B(n_167), .Y(n_222) );
NAND2xp5_ASAP7_75t_SL g489 ( .A(n_42), .B(n_155), .Y(n_489) );
AOI22xp33_ASAP7_75t_L g510 ( .A1(n_43), .A2(n_85), .B1(n_213), .B2(n_511), .Y(n_510) );
NAND2xp5_ASAP7_75t_SL g492 ( .A(n_44), .B(n_155), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_45), .B(n_155), .Y(n_476) );
CKINVDCx16_ASAP7_75t_R g184 ( .A(n_46), .Y(n_184) );
OAI222xp33_ASAP7_75t_L g455 ( .A1(n_47), .A2(n_456), .B1(n_754), .B2(n_755), .C1(n_760), .C2(n_764), .Y(n_455) );
CKINVDCx16_ASAP7_75t_R g754 ( .A(n_47), .Y(n_754) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_48), .B(n_480), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_49), .B(n_136), .Y(n_238) );
AOI22xp33_ASAP7_75t_SL g550 ( .A1(n_51), .A2(n_60), .B1(n_155), .B2(n_177), .Y(n_550) );
AOI22xp5_ASAP7_75t_L g176 ( .A1(n_52), .A2(n_145), .B1(n_177), .B2(n_179), .Y(n_176) );
CKINVDCx20_ASAP7_75t_R g216 ( .A(n_53), .Y(n_216) );
NAND2xp5_ASAP7_75t_SL g502 ( .A(n_54), .B(n_155), .Y(n_502) );
CKINVDCx16_ASAP7_75t_R g191 ( .A(n_55), .Y(n_191) );
NAND2xp5_ASAP7_75t_SL g517 ( .A(n_56), .B(n_155), .Y(n_517) );
A2O1A1Ixp33_ASAP7_75t_L g165 ( .A1(n_57), .A2(n_154), .B(n_166), .C(n_168), .Y(n_165) );
CKINVDCx20_ASAP7_75t_R g226 ( .A(n_58), .Y(n_226) );
INVx1_ASAP7_75t_L g164 ( .A(n_59), .Y(n_164) );
INVx1_ASAP7_75t_L g142 ( .A(n_61), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_62), .B(n_155), .Y(n_482) );
INVx1_ASAP7_75t_L g133 ( .A(n_63), .Y(n_133) );
CKINVDCx20_ASAP7_75t_R g116 ( .A(n_64), .Y(n_116) );
AO32x2_ASAP7_75t_L g508 ( .A1(n_65), .A2(n_129), .A3(n_230), .B1(n_503), .B2(n_509), .Y(n_508) );
INVx1_ASAP7_75t_L g501 ( .A(n_66), .Y(n_501) );
INVx1_ASAP7_75t_L g536 ( .A(n_67), .Y(n_536) );
CKINVDCx20_ASAP7_75t_R g764 ( .A(n_68), .Y(n_764) );
A2O1A1Ixp33_ASAP7_75t_SL g149 ( .A1(n_69), .A2(n_150), .B(n_151), .C(n_154), .Y(n_149) );
INVxp67_ASAP7_75t_L g152 ( .A(n_70), .Y(n_152) );
NAND2xp5_ASAP7_75t_SL g537 ( .A(n_71), .B(n_177), .Y(n_537) );
INVx1_ASAP7_75t_L g108 ( .A(n_72), .Y(n_108) );
CKINVDCx20_ASAP7_75t_R g187 ( .A(n_73), .Y(n_187) );
INVx1_ASAP7_75t_L g219 ( .A(n_74), .Y(n_219) );
A2O1A1Ixp33_ASAP7_75t_L g220 ( .A1(n_76), .A2(n_141), .B(n_145), .C(n_221), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_77), .B(n_511), .Y(n_522) );
NAND2xp5_ASAP7_75t_SL g540 ( .A(n_78), .B(n_177), .Y(n_540) );
NAND2xp5_ASAP7_75t_SL g209 ( .A(n_79), .B(n_195), .Y(n_209) );
INVx2_ASAP7_75t_L g131 ( .A(n_80), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_81), .B(n_150), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_82), .B(n_177), .Y(n_490) );
A2O1A1Ixp33_ASAP7_75t_L g192 ( .A1(n_83), .A2(n_141), .B(n_145), .C(n_193), .Y(n_192) );
NAND3xp33_ASAP7_75t_SL g104 ( .A(n_84), .B(n_105), .C(n_106), .Y(n_104) );
OR2x2_ASAP7_75t_L g447 ( .A(n_84), .B(n_448), .Y(n_447) );
OR2x2_ASAP7_75t_L g458 ( .A(n_84), .B(n_449), .Y(n_458) );
INVx2_ASAP7_75t_L g462 ( .A(n_84), .Y(n_462) );
AOI22xp33_ASAP7_75t_L g549 ( .A1(n_86), .A2(n_98), .B1(n_177), .B2(n_178), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_87), .B(n_171), .Y(n_170) );
CKINVDCx20_ASAP7_75t_R g199 ( .A(n_88), .Y(n_199) );
A2O1A1Ixp33_ASAP7_75t_L g232 ( .A1(n_89), .A2(n_141), .B(n_145), .C(n_233), .Y(n_232) );
CKINVDCx20_ASAP7_75t_R g240 ( .A(n_90), .Y(n_240) );
INVx1_ASAP7_75t_L g148 ( .A(n_91), .Y(n_148) );
CKINVDCx16_ASAP7_75t_R g246 ( .A(n_92), .Y(n_246) );
NAND2xp5_ASAP7_75t_SL g234 ( .A(n_93), .B(n_195), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_94), .B(n_177), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_95), .B(n_129), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g107 ( .A(n_96), .B(n_108), .Y(n_107) );
AOI21xp5_ASAP7_75t_L g135 ( .A1(n_97), .A2(n_136), .B(n_143), .Y(n_135) );
INVx1_ASAP7_75t_L g100 ( .A(n_101), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
INVx2_ASAP7_75t_SL g769 ( .A(n_102), .Y(n_769) );
AND2x2_ASAP7_75t_SL g102 ( .A(n_103), .B(n_109), .Y(n_102) );
CKINVDCx16_ASAP7_75t_R g103 ( .A(n_104), .Y(n_103) );
AND2x2_ASAP7_75t_L g449 ( .A(n_105), .B(n_450), .Y(n_449) );
INVx1_ASAP7_75t_SL g106 ( .A(n_107), .Y(n_106) );
INVxp67_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
OAI21xp5_ASAP7_75t_L g112 ( .A1(n_113), .A2(n_117), .B(n_454), .Y(n_112) );
BUFx2_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
BUFx2_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
INVx2_ASAP7_75t_SL g766 ( .A(n_115), .Y(n_766) );
INVx2_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
AOI21xp5_ASAP7_75t_L g117 ( .A1(n_118), .A2(n_446), .B(n_451), .Y(n_117) );
INVx2_ASAP7_75t_L g445 ( .A(n_120), .Y(n_445) );
INVx1_ASAP7_75t_SL g459 ( .A(n_120), .Y(n_459) );
AOI22xp5_ASAP7_75t_L g755 ( .A1(n_120), .A2(n_756), .B1(n_758), .B2(n_759), .Y(n_755) );
INVx3_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
AND4x1_ASAP7_75t_L g121 ( .A(n_122), .B(n_363), .C(n_410), .D(n_430), .Y(n_121) );
NOR3xp33_ASAP7_75t_SL g122 ( .A(n_123), .B(n_293), .C(n_318), .Y(n_122) );
OAI211xp5_ASAP7_75t_SL g123 ( .A1(n_124), .A2(n_201), .B(n_253), .C(n_283), .Y(n_123) );
INVxp67_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
NOR2xp33_ASAP7_75t_L g125 ( .A(n_126), .B(n_172), .Y(n_125) );
INVx3_ASAP7_75t_SL g335 ( .A(n_126), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_126), .B(n_266), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_126), .B(n_188), .Y(n_416) );
AND2x2_ASAP7_75t_L g439 ( .A(n_126), .B(n_305), .Y(n_439) );
AND2x4_ASAP7_75t_L g126 ( .A(n_127), .B(n_160), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
AND2x2_ASAP7_75t_L g257 ( .A(n_128), .B(n_161), .Y(n_257) );
INVx3_ASAP7_75t_L g270 ( .A(n_128), .Y(n_270) );
AND2x2_ASAP7_75t_L g275 ( .A(n_128), .B(n_160), .Y(n_275) );
OR2x2_ASAP7_75t_L g326 ( .A(n_128), .B(n_267), .Y(n_326) );
BUFx2_ASAP7_75t_L g346 ( .A(n_128), .Y(n_346) );
AND2x2_ASAP7_75t_L g356 ( .A(n_128), .B(n_267), .Y(n_356) );
AND2x2_ASAP7_75t_L g362 ( .A(n_128), .B(n_173), .Y(n_362) );
OA21x2_ASAP7_75t_L g128 ( .A1(n_129), .A2(n_135), .B(n_157), .Y(n_128) );
INVx4_ASAP7_75t_L g159 ( .A(n_129), .Y(n_159) );
OA21x2_ASAP7_75t_L g486 ( .A1(n_129), .A2(n_487), .B(n_494), .Y(n_486) );
BUFx6f_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
INVx1_ASAP7_75t_L g174 ( .A(n_130), .Y(n_174) );
AND2x2_ASAP7_75t_L g130 ( .A(n_131), .B(n_132), .Y(n_130) );
AND2x2_ASAP7_75t_SL g171 ( .A(n_131), .B(n_132), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g132 ( .A(n_133), .B(n_134), .Y(n_132) );
BUFx2_ASAP7_75t_L g244 ( .A(n_136), .Y(n_244) );
AND2x4_ASAP7_75t_L g136 ( .A(n_137), .B(n_141), .Y(n_136) );
NAND2x1p5_ASAP7_75t_L g185 ( .A(n_137), .B(n_141), .Y(n_185) );
AND2x2_ASAP7_75t_L g137 ( .A(n_138), .B(n_140), .Y(n_137) );
INVx1_ASAP7_75t_L g480 ( .A(n_138), .Y(n_480) );
INVx1_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
INVx2_ASAP7_75t_L g146 ( .A(n_139), .Y(n_146) );
INVx1_ASAP7_75t_L g178 ( .A(n_139), .Y(n_178) );
INVx1_ASAP7_75t_L g147 ( .A(n_140), .Y(n_147) );
INVx1_ASAP7_75t_L g150 ( .A(n_140), .Y(n_150) );
INVx3_ASAP7_75t_L g153 ( .A(n_140), .Y(n_153) );
BUFx6f_ASAP7_75t_L g167 ( .A(n_140), .Y(n_167) );
BUFx6f_ASAP7_75t_L g180 ( .A(n_140), .Y(n_180) );
INVx4_ASAP7_75t_SL g156 ( .A(n_141), .Y(n_156) );
OAI21xp5_ASAP7_75t_L g473 ( .A1(n_141), .A2(n_474), .B(n_478), .Y(n_473) );
OAI21xp5_ASAP7_75t_L g487 ( .A1(n_141), .A2(n_488), .B(n_491), .Y(n_487) );
BUFx3_ASAP7_75t_L g503 ( .A(n_141), .Y(n_503) );
OAI21xp5_ASAP7_75t_L g515 ( .A1(n_141), .A2(n_516), .B(n_520), .Y(n_515) );
OAI21xp5_ASAP7_75t_L g534 ( .A1(n_141), .A2(n_535), .B(n_538), .Y(n_534) );
O2A1O1Ixp33_ASAP7_75t_L g143 ( .A1(n_144), .A2(n_148), .B(n_149), .C(n_156), .Y(n_143) );
O2A1O1Ixp33_ASAP7_75t_L g163 ( .A1(n_144), .A2(n_156), .B(n_164), .C(n_165), .Y(n_163) );
O2A1O1Ixp33_ASAP7_75t_L g245 ( .A1(n_144), .A2(n_156), .B(n_246), .C(n_247), .Y(n_245) );
INVx5_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
AND2x6_ASAP7_75t_L g145 ( .A(n_146), .B(n_147), .Y(n_145) );
BUFx6f_ASAP7_75t_L g155 ( .A(n_146), .Y(n_155) );
BUFx3_ASAP7_75t_L g213 ( .A(n_146), .Y(n_213) );
INVx1_ASAP7_75t_L g511 ( .A(n_146), .Y(n_511) );
INVx1_ASAP7_75t_L g519 ( .A(n_150), .Y(n_519) );
NOR2xp33_ASAP7_75t_L g151 ( .A(n_152), .B(n_153), .Y(n_151) );
NOR2xp33_ASAP7_75t_L g168 ( .A(n_153), .B(n_169), .Y(n_168) );
INVx5_ASAP7_75t_L g195 ( .A(n_153), .Y(n_195) );
OAI22xp5_ASAP7_75t_SL g509 ( .A1(n_153), .A2(n_167), .B1(n_510), .B2(n_512), .Y(n_509) );
O2A1O1Ixp5_ASAP7_75t_SL g535 ( .A1(n_154), .A2(n_195), .B(n_536), .C(n_537), .Y(n_535) );
INVx3_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
HB1xp67_ASAP7_75t_L g237 ( .A(n_155), .Y(n_237) );
OAI22xp33_ASAP7_75t_L g175 ( .A1(n_156), .A2(n_176), .B1(n_184), .B2(n_185), .Y(n_175) );
OA21x2_ASAP7_75t_L g161 ( .A1(n_158), .A2(n_162), .B(n_170), .Y(n_161) );
INVx3_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
NOR2xp33_ASAP7_75t_SL g215 ( .A(n_159), .B(n_216), .Y(n_215) );
AO21x1_ASAP7_75t_L g547 ( .A1(n_159), .A2(n_548), .B(n_551), .Y(n_547) );
NAND3xp33_ASAP7_75t_L g566 ( .A(n_159), .B(n_503), .C(n_548), .Y(n_566) );
INVx1_ASAP7_75t_SL g160 ( .A(n_161), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_161), .B(n_267), .Y(n_281) );
INVx2_ASAP7_75t_L g291 ( .A(n_161), .Y(n_291) );
AND2x2_ASAP7_75t_L g304 ( .A(n_161), .B(n_270), .Y(n_304) );
OR2x2_ASAP7_75t_L g315 ( .A(n_161), .B(n_267), .Y(n_315) );
AND2x2_ASAP7_75t_SL g361 ( .A(n_161), .B(n_362), .Y(n_361) );
BUFx2_ASAP7_75t_L g373 ( .A(n_161), .Y(n_373) );
AND2x2_ASAP7_75t_L g419 ( .A(n_161), .B(n_173), .Y(n_419) );
O2A1O1Ixp5_ASAP7_75t_L g500 ( .A1(n_166), .A2(n_479), .B(n_501), .C(n_502), .Y(n_500) );
AOI21xp5_ASAP7_75t_L g520 ( .A1(n_166), .A2(n_521), .B(n_522), .Y(n_520) );
INVx2_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
INVx4_ASAP7_75t_L g236 ( .A(n_167), .Y(n_236) );
OAI22xp5_ASAP7_75t_L g525 ( .A1(n_167), .A2(n_483), .B1(n_526), .B2(n_527), .Y(n_525) );
OAI22xp5_ASAP7_75t_L g548 ( .A1(n_167), .A2(n_483), .B1(n_549), .B2(n_550), .Y(n_548) );
INVx1_ASAP7_75t_L g200 ( .A(n_171), .Y(n_200) );
INVx2_ASAP7_75t_L g230 ( .A(n_171), .Y(n_230) );
OA21x2_ASAP7_75t_L g242 ( .A1(n_171), .A2(n_243), .B(n_252), .Y(n_242) );
OA21x2_ASAP7_75t_L g514 ( .A1(n_171), .A2(n_515), .B(n_523), .Y(n_514) );
OA21x2_ASAP7_75t_L g533 ( .A1(n_171), .A2(n_534), .B(n_541), .Y(n_533) );
INVx3_ASAP7_75t_SL g292 ( .A(n_172), .Y(n_292) );
OR2x2_ASAP7_75t_L g345 ( .A(n_172), .B(n_346), .Y(n_345) );
OR2x2_ASAP7_75t_L g172 ( .A(n_173), .B(n_188), .Y(n_172) );
INVx3_ASAP7_75t_L g267 ( .A(n_173), .Y(n_267) );
AND2x2_ASAP7_75t_L g334 ( .A(n_173), .B(n_189), .Y(n_334) );
HB1xp67_ASAP7_75t_L g402 ( .A(n_173), .Y(n_402) );
AOI33xp33_ASAP7_75t_L g406 ( .A1(n_173), .A2(n_335), .A3(n_342), .B1(n_351), .B2(n_407), .B3(n_408), .Y(n_406) );
AO21x2_ASAP7_75t_L g173 ( .A1(n_174), .A2(n_175), .B(n_186), .Y(n_173) );
NOR2xp33_ASAP7_75t_L g186 ( .A(n_174), .B(n_187), .Y(n_186) );
AO21x2_ASAP7_75t_L g189 ( .A1(n_174), .A2(n_190), .B(n_198), .Y(n_189) );
INVx2_ASAP7_75t_L g214 ( .A(n_174), .Y(n_214) );
INVx2_ASAP7_75t_L g197 ( .A(n_177), .Y(n_197) );
INVx3_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
OAI22xp5_ASAP7_75t_SL g179 ( .A1(n_180), .A2(n_181), .B1(n_182), .B2(n_183), .Y(n_179) );
INVx2_ASAP7_75t_L g182 ( .A(n_180), .Y(n_182) );
INVx4_ASAP7_75t_L g248 ( .A(n_180), .Y(n_248) );
OAI21xp5_ASAP7_75t_L g190 ( .A1(n_185), .A2(n_191), .B(n_192), .Y(n_190) );
OAI21xp5_ASAP7_75t_L g218 ( .A1(n_185), .A2(n_219), .B(n_220), .Y(n_218) );
INVx1_ASAP7_75t_L g255 ( .A(n_188), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_188), .B(n_270), .Y(n_269) );
NOR3xp33_ASAP7_75t_L g329 ( .A(n_188), .B(n_330), .C(n_332), .Y(n_329) );
AND2x2_ASAP7_75t_L g355 ( .A(n_188), .B(n_356), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_188), .B(n_362), .Y(n_365) );
AND2x2_ASAP7_75t_L g418 ( .A(n_188), .B(n_419), .Y(n_418) );
INVx3_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
INVx3_ASAP7_75t_L g274 ( .A(n_189), .Y(n_274) );
OR2x2_ASAP7_75t_L g368 ( .A(n_189), .B(n_267), .Y(n_368) );
O2A1O1Ixp33_ASAP7_75t_L g193 ( .A1(n_194), .A2(n_195), .B(n_196), .C(n_197), .Y(n_193) );
INVx2_ASAP7_75t_L g483 ( .A(n_195), .Y(n_483) );
AOI21xp5_ASAP7_75t_L g488 ( .A1(n_195), .A2(n_489), .B(n_490), .Y(n_488) );
AOI21xp5_ASAP7_75t_L g497 ( .A1(n_195), .A2(n_498), .B(n_499), .Y(n_497) );
O2A1O1Ixp33_ASAP7_75t_L g474 ( .A1(n_197), .A2(n_475), .B(n_476), .C(n_477), .Y(n_474) );
NOR2xp33_ASAP7_75t_L g198 ( .A(n_199), .B(n_200), .Y(n_198) );
NOR2xp33_ASAP7_75t_L g225 ( .A(n_200), .B(n_226), .Y(n_225) );
NOR2xp33_ASAP7_75t_L g239 ( .A(n_200), .B(n_240), .Y(n_239) );
OR2x2_ASAP7_75t_L g201 ( .A(n_202), .B(n_227), .Y(n_201) );
AOI32xp33_ASAP7_75t_L g319 ( .A1(n_202), .A2(n_320), .A3(n_322), .B1(n_324), .B2(n_327), .Y(n_319) );
NOR2xp67_ASAP7_75t_L g392 ( .A(n_202), .B(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g422 ( .A(n_202), .Y(n_422) );
INVx4_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
AND2x2_ASAP7_75t_L g354 ( .A(n_203), .B(n_338), .Y(n_354) );
AND2x2_ASAP7_75t_L g374 ( .A(n_203), .B(n_300), .Y(n_374) );
AND2x2_ASAP7_75t_L g442 ( .A(n_203), .B(n_360), .Y(n_442) );
AND2x2_ASAP7_75t_L g203 ( .A(n_204), .B(n_217), .Y(n_203) );
INVx3_ASAP7_75t_L g263 ( .A(n_204), .Y(n_263) );
AND2x2_ASAP7_75t_L g277 ( .A(n_204), .B(n_261), .Y(n_277) );
OR2x2_ASAP7_75t_L g282 ( .A(n_204), .B(n_260), .Y(n_282) );
INVx1_ASAP7_75t_L g289 ( .A(n_204), .Y(n_289) );
AND2x2_ASAP7_75t_L g297 ( .A(n_204), .B(n_271), .Y(n_297) );
AND2x2_ASAP7_75t_L g299 ( .A(n_204), .B(n_300), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_204), .B(n_338), .Y(n_337) );
INVx2_ASAP7_75t_L g352 ( .A(n_204), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_204), .B(n_437), .Y(n_436) );
OR2x6_ASAP7_75t_L g204 ( .A(n_205), .B(n_215), .Y(n_204) );
AOI21xp5_ASAP7_75t_SL g205 ( .A1(n_206), .A2(n_207), .B(n_214), .Y(n_205) );
AOI21xp5_ASAP7_75t_L g208 ( .A1(n_209), .A2(n_210), .B(n_211), .Y(n_208) );
AOI21xp5_ASAP7_75t_L g221 ( .A1(n_211), .A2(n_222), .B(n_223), .Y(n_221) );
INVx2_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
INVx2_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
INVx1_ASAP7_75t_L g251 ( .A(n_213), .Y(n_251) );
INVx1_ASAP7_75t_L g224 ( .A(n_214), .Y(n_224) );
OA21x2_ASAP7_75t_L g472 ( .A1(n_214), .A2(n_473), .B(n_484), .Y(n_472) );
OA21x2_ASAP7_75t_L g495 ( .A1(n_214), .A2(n_496), .B(n_504), .Y(n_495) );
INVx2_ASAP7_75t_L g261 ( .A(n_217), .Y(n_261) );
AND2x2_ASAP7_75t_L g307 ( .A(n_217), .B(n_228), .Y(n_307) );
AND2x2_ASAP7_75t_L g317 ( .A(n_217), .B(n_242), .Y(n_317) );
AO21x2_ASAP7_75t_L g217 ( .A1(n_218), .A2(n_224), .B(n_225), .Y(n_217) );
INVx2_ASAP7_75t_L g437 ( .A(n_227), .Y(n_437) );
OR2x2_ASAP7_75t_L g227 ( .A(n_228), .B(n_241), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_228), .B(n_261), .Y(n_260) );
INVx1_ASAP7_75t_L g278 ( .A(n_228), .Y(n_278) );
AND2x2_ASAP7_75t_L g322 ( .A(n_228), .B(n_323), .Y(n_322) );
AND2x2_ASAP7_75t_L g338 ( .A(n_228), .B(n_301), .Y(n_338) );
INVx2_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
INVx1_ASAP7_75t_L g286 ( .A(n_229), .Y(n_286) );
AND2x2_ASAP7_75t_L g300 ( .A(n_229), .B(n_301), .Y(n_300) );
AND2x2_ASAP7_75t_L g351 ( .A(n_229), .B(n_352), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_229), .B(n_261), .Y(n_383) );
AO21x2_ASAP7_75t_L g229 ( .A1(n_230), .A2(n_231), .B(n_239), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_232), .B(n_238), .Y(n_231) );
AOI21xp5_ASAP7_75t_L g233 ( .A1(n_234), .A2(n_235), .B(n_237), .Y(n_233) );
AND2x2_ASAP7_75t_L g262 ( .A(n_241), .B(n_263), .Y(n_262) );
INVx2_ASAP7_75t_L g323 ( .A(n_241), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_241), .B(n_331), .Y(n_330) );
INVx1_ASAP7_75t_L g360 ( .A(n_241), .Y(n_360) );
INVx1_ASAP7_75t_L g393 ( .A(n_241), .Y(n_393) );
INVx2_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
AND2x2_ASAP7_75t_L g271 ( .A(n_242), .B(n_261), .Y(n_271) );
INVx1_ASAP7_75t_L g301 ( .A(n_242), .Y(n_301) );
NOR2xp33_ASAP7_75t_L g249 ( .A(n_248), .B(n_250), .Y(n_249) );
INVx1_ASAP7_75t_L g477 ( .A(n_248), .Y(n_477) );
AOI21xp5_ASAP7_75t_L g538 ( .A1(n_248), .A2(n_539), .B(n_540), .Y(n_538) );
AOI221xp5_ASAP7_75t_L g253 ( .A1(n_254), .A2(n_258), .B1(n_264), .B2(n_271), .C(n_272), .Y(n_253) );
NOR2xp33_ASAP7_75t_L g254 ( .A(n_255), .B(n_256), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_255), .B(n_275), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_255), .B(n_338), .Y(n_415) );
INVx1_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_257), .B(n_305), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_257), .B(n_266), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_257), .B(n_280), .Y(n_409) );
AND2x2_ASAP7_75t_L g258 ( .A(n_259), .B(n_262), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
INVx2_ASAP7_75t_L g331 ( .A(n_261), .Y(n_331) );
AND2x2_ASAP7_75t_L g306 ( .A(n_262), .B(n_307), .Y(n_306) );
INVx1_ASAP7_75t_L g384 ( .A(n_262), .Y(n_384) );
AND2x2_ASAP7_75t_L g316 ( .A(n_263), .B(n_317), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_263), .B(n_286), .Y(n_332) );
AND2x2_ASAP7_75t_L g396 ( .A(n_263), .B(n_322), .Y(n_396) );
INVx1_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_266), .B(n_268), .Y(n_265) );
BUFx2_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
AND2x2_ASAP7_75t_L g305 ( .A(n_267), .B(n_274), .Y(n_305) );
AND2x2_ASAP7_75t_L g401 ( .A(n_268), .B(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_270), .B(n_314), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_271), .B(n_289), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_271), .B(n_278), .Y(n_366) );
AND2x2_ASAP7_75t_L g386 ( .A(n_271), .B(n_286), .Y(n_386) );
AND2x2_ASAP7_75t_L g407 ( .A(n_271), .B(n_351), .Y(n_407) );
OAI32xp33_ASAP7_75t_L g272 ( .A1(n_273), .A2(n_276), .A3(n_278), .B1(n_279), .B2(n_282), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_274), .B(n_275), .Y(n_273) );
INVx1_ASAP7_75t_SL g280 ( .A(n_274), .Y(n_280) );
NAND2x1_ASAP7_75t_L g321 ( .A(n_274), .B(n_304), .Y(n_321) );
OR2x2_ASAP7_75t_L g325 ( .A(n_274), .B(n_326), .Y(n_325) );
NOR2xp33_ASAP7_75t_L g426 ( .A(n_274), .B(n_373), .Y(n_426) );
INVx1_ASAP7_75t_L g294 ( .A(n_275), .Y(n_294) );
OAI221xp5_ASAP7_75t_SL g412 ( .A1(n_276), .A2(n_367), .B1(n_413), .B2(n_416), .C(n_417), .Y(n_412) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
AND2x2_ASAP7_75t_L g284 ( .A(n_277), .B(n_285), .Y(n_284) );
AND2x2_ASAP7_75t_L g327 ( .A(n_277), .B(n_300), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_277), .B(n_359), .Y(n_358) );
AND2x2_ASAP7_75t_L g405 ( .A(n_277), .B(n_338), .Y(n_405) );
INVxp67_ASAP7_75t_L g341 ( .A(n_278), .Y(n_341) );
OR2x2_ASAP7_75t_L g279 ( .A(n_280), .B(n_281), .Y(n_279) );
AND2x2_ASAP7_75t_L g411 ( .A(n_280), .B(n_398), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_280), .B(n_361), .Y(n_434) );
INVx1_ASAP7_75t_L g309 ( .A(n_282), .Y(n_309) );
NAND2xp5_ASAP7_75t_SL g390 ( .A(n_282), .B(n_391), .Y(n_390) );
OR2x2_ASAP7_75t_L g427 ( .A(n_282), .B(n_428), .Y(n_427) );
OAI21xp5_ASAP7_75t_SL g283 ( .A1(n_284), .A2(n_287), .B(n_290), .Y(n_283) );
AND2x2_ASAP7_75t_L g296 ( .A(n_285), .B(n_297), .Y(n_296) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
AND2x2_ASAP7_75t_L g380 ( .A(n_289), .B(n_300), .Y(n_380) );
AND2x2_ASAP7_75t_L g290 ( .A(n_291), .B(n_292), .Y(n_290) );
AND2x2_ASAP7_75t_L g398 ( .A(n_291), .B(n_356), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_291), .B(n_355), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_292), .B(n_304), .Y(n_378) );
OAI211xp5_ASAP7_75t_L g293 ( .A1(n_294), .A2(n_295), .B(n_298), .C(n_308), .Y(n_293) );
AOI221xp5_ASAP7_75t_L g328 ( .A1(n_294), .A2(n_329), .B1(n_333), .B2(n_336), .C(n_339), .Y(n_328) );
AOI31xp33_ASAP7_75t_L g423 ( .A1(n_294), .A2(n_424), .A3(n_425), .B(n_427), .Y(n_423) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
AOI22xp5_ASAP7_75t_L g298 ( .A1(n_299), .A2(n_302), .B1(n_304), .B2(n_306), .Y(n_298) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_304), .B(n_305), .Y(n_303) );
INVx1_ASAP7_75t_L g424 ( .A(n_304), .Y(n_424) );
INVx1_ASAP7_75t_L g387 ( .A(n_305), .Y(n_387) );
O2A1O1Ixp33_ASAP7_75t_L g430 ( .A1(n_307), .A2(n_431), .B(n_433), .C(n_435), .Y(n_430) );
AOI22xp33_ASAP7_75t_L g308 ( .A1(n_309), .A2(n_310), .B1(n_312), .B2(n_316), .Y(n_308) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_313), .B(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
OAI221xp5_ASAP7_75t_SL g403 ( .A1(n_315), .A2(n_349), .B1(n_368), .B2(n_404), .C(n_406), .Y(n_403) );
INVx1_ASAP7_75t_L g399 ( .A(n_316), .Y(n_399) );
INVx1_ASAP7_75t_L g353 ( .A(n_317), .Y(n_353) );
NAND3xp33_ASAP7_75t_SL g318 ( .A(n_319), .B(n_328), .C(n_343), .Y(n_318) );
OAI21xp33_ASAP7_75t_L g369 ( .A1(n_320), .A2(n_370), .B(n_374), .Y(n_369) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_322), .B(n_422), .Y(n_421) );
INVxp67_ASAP7_75t_L g429 ( .A(n_323), .Y(n_429) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
OR2x2_ASAP7_75t_L g367 ( .A(n_330), .B(n_350), .Y(n_367) );
INVx1_ASAP7_75t_L g342 ( .A(n_331), .Y(n_342) );
AND2x2_ASAP7_75t_L g333 ( .A(n_334), .B(n_335), .Y(n_333) );
INVx1_ASAP7_75t_L g340 ( .A(n_334), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_334), .B(n_372), .Y(n_371) );
NOR4xp25_ASAP7_75t_L g339 ( .A(n_335), .B(n_340), .C(n_341), .D(n_342), .Y(n_339) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
AOI222xp33_ASAP7_75t_L g343 ( .A1(n_344), .A2(n_348), .B1(n_354), .B2(n_355), .C1(n_357), .C2(n_361), .Y(n_343) );
NAND2xp5_ASAP7_75t_SL g344 ( .A(n_345), .B(n_347), .Y(n_344) );
INVx1_ASAP7_75t_L g441 ( .A(n_345), .Y(n_441) );
INVx1_ASAP7_75t_SL g348 ( .A(n_349), .Y(n_348) );
OR2x2_ASAP7_75t_L g349 ( .A(n_350), .B(n_353), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_357), .B(n_444), .Y(n_443) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
OAI21xp5_ASAP7_75t_SL g417 ( .A1(n_362), .A2(n_418), .B(n_420), .Y(n_417) );
NOR4xp25_ASAP7_75t_L g363 ( .A(n_364), .B(n_375), .C(n_388), .D(n_403), .Y(n_363) );
OAI221xp5_ASAP7_75t_SL g364 ( .A1(n_365), .A2(n_366), .B1(n_367), .B2(n_368), .C(n_369), .Y(n_364) );
INVx1_ASAP7_75t_L g444 ( .A(n_365), .Y(n_444) );
INVx1_ASAP7_75t_SL g370 ( .A(n_371), .Y(n_370) );
NOR2xp33_ASAP7_75t_L g414 ( .A(n_372), .B(n_415), .Y(n_414) );
INVx1_ASAP7_75t_SL g372 ( .A(n_373), .Y(n_372) );
OAI222xp33_ASAP7_75t_L g375 ( .A1(n_376), .A2(n_379), .B1(n_381), .B2(n_382), .C1(n_385), .C2(n_387), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
AOI211xp5_ASAP7_75t_L g410 ( .A1(n_380), .A2(n_411), .B(n_412), .C(n_423), .Y(n_410) );
OR2x2_ASAP7_75t_L g382 ( .A(n_383), .B(n_384), .Y(n_382) );
INVx1_ASAP7_75t_SL g385 ( .A(n_386), .Y(n_385) );
OAI222xp33_ASAP7_75t_L g388 ( .A1(n_389), .A2(n_394), .B1(n_395), .B2(n_397), .C1(n_399), .C2(n_400), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVxp67_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
AOI22xp5_ASAP7_75t_L g440 ( .A1(n_405), .A2(n_408), .B1(n_441), .B2(n_442), .Y(n_440) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
HB1xp67_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
OAI211xp5_ASAP7_75t_SL g435 ( .A1(n_436), .A2(n_438), .B(n_440), .C(n_443), .Y(n_435) );
INVx2_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
BUFx2_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
HB1xp67_ASAP7_75t_L g452 ( .A(n_447), .Y(n_452) );
NOR2x2_ASAP7_75t_L g763 ( .A(n_448), .B(n_462), .Y(n_763) );
INVx2_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
OR2x2_ASAP7_75t_L g461 ( .A(n_449), .B(n_462), .Y(n_461) );
OAI21xp5_ASAP7_75t_SL g454 ( .A1(n_451), .A2(n_455), .B(n_765), .Y(n_454) );
NOR2xp33_ASAP7_75t_SL g451 ( .A(n_452), .B(n_453), .Y(n_451) );
AOI22xp5_ASAP7_75t_L g456 ( .A1(n_457), .A2(n_459), .B1(n_460), .B2(n_463), .Y(n_456) );
INVx2_ASAP7_75t_L g757 ( .A(n_457), .Y(n_757) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx6_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVx1_ASAP7_75t_L g758 ( .A(n_461), .Y(n_758) );
INVx1_ASAP7_75t_L g759 ( .A(n_463), .Y(n_759) );
AND2x2_ASAP7_75t_SL g463 ( .A(n_464), .B(n_720), .Y(n_463) );
NOR3xp33_ASAP7_75t_L g464 ( .A(n_465), .B(n_624), .C(n_708), .Y(n_464) );
NAND4xp25_ASAP7_75t_L g465 ( .A(n_466), .B(n_567), .C(n_589), .D(n_605), .Y(n_465) );
AOI221xp5_ASAP7_75t_L g466 ( .A1(n_467), .A2(n_505), .B1(n_528), .B2(n_546), .C(n_553), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_469), .B(n_485), .Y(n_468) );
NAND2xp5_ASAP7_75t_SL g579 ( .A(n_469), .B(n_546), .Y(n_579) );
NAND4xp25_ASAP7_75t_L g619 ( .A(n_469), .B(n_607), .C(n_620), .D(n_622), .Y(n_619) );
INVxp67_ASAP7_75t_L g736 ( .A(n_469), .Y(n_736) );
INVx3_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
OR2x2_ASAP7_75t_L g618 ( .A(n_470), .B(n_556), .Y(n_618) );
AND2x2_ASAP7_75t_L g642 ( .A(n_470), .B(n_485), .Y(n_642) );
INVx2_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
AND2x2_ASAP7_75t_L g609 ( .A(n_471), .B(n_545), .Y(n_609) );
AND2x2_ASAP7_75t_L g649 ( .A(n_471), .B(n_630), .Y(n_649) );
AND2x2_ASAP7_75t_L g666 ( .A(n_471), .B(n_667), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_471), .B(n_486), .Y(n_690) );
INVx2_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
AND2x2_ASAP7_75t_L g544 ( .A(n_472), .B(n_545), .Y(n_544) );
AND2x2_ASAP7_75t_L g561 ( .A(n_472), .B(n_562), .Y(n_561) );
AND2x2_ASAP7_75t_L g573 ( .A(n_472), .B(n_486), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_472), .B(n_495), .Y(n_595) );
O2A1O1Ixp33_ASAP7_75t_L g478 ( .A1(n_479), .A2(n_481), .B(n_482), .C(n_483), .Y(n_478) );
INVx2_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
AOI21xp5_ASAP7_75t_L g491 ( .A1(n_483), .A2(n_492), .B(n_493), .Y(n_491) );
AND2x2_ASAP7_75t_L g576 ( .A(n_485), .B(n_577), .Y(n_576) );
AOI221xp5_ASAP7_75t_L g625 ( .A1(n_485), .A2(n_626), .B1(n_629), .B2(n_631), .C(n_635), .Y(n_625) );
AND2x2_ASAP7_75t_L g684 ( .A(n_485), .B(n_649), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_485), .B(n_666), .Y(n_718) );
AND2x2_ASAP7_75t_L g485 ( .A(n_486), .B(n_495), .Y(n_485) );
INVx3_ASAP7_75t_L g545 ( .A(n_486), .Y(n_545) );
AND2x2_ASAP7_75t_L g593 ( .A(n_486), .B(n_594), .Y(n_593) );
AND2x2_ASAP7_75t_L g647 ( .A(n_486), .B(n_562), .Y(n_647) );
AND2x2_ASAP7_75t_L g705 ( .A(n_486), .B(n_706), .Y(n_705) );
AND2x2_ASAP7_75t_L g546 ( .A(n_495), .B(n_547), .Y(n_546) );
INVx2_ASAP7_75t_L g562 ( .A(n_495), .Y(n_562) );
INVx1_ASAP7_75t_L g617 ( .A(n_495), .Y(n_617) );
HB1xp67_ASAP7_75t_L g623 ( .A(n_495), .Y(n_623) );
AND2x2_ASAP7_75t_L g668 ( .A(n_495), .B(n_545), .Y(n_668) );
OR2x2_ASAP7_75t_L g707 ( .A(n_495), .B(n_547), .Y(n_707) );
OAI21xp5_ASAP7_75t_L g496 ( .A1(n_497), .A2(n_500), .B(n_503), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_505), .B(n_587), .Y(n_586) );
AND2x2_ASAP7_75t_L g505 ( .A(n_506), .B(n_513), .Y(n_505) );
AND2x2_ASAP7_75t_L g703 ( .A(n_506), .B(n_700), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g735 ( .A(n_506), .B(n_685), .Y(n_735) );
BUFx2_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
AND2x2_ASAP7_75t_L g634 ( .A(n_507), .B(n_558), .Y(n_634) );
AND2x2_ASAP7_75t_L g683 ( .A(n_507), .B(n_531), .Y(n_683) );
INVx1_ASAP7_75t_L g729 ( .A(n_507), .Y(n_729) );
INVx1_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
BUFx6f_ASAP7_75t_L g543 ( .A(n_508), .Y(n_543) );
AND2x2_ASAP7_75t_L g584 ( .A(n_508), .B(n_558), .Y(n_584) );
INVx1_ASAP7_75t_L g601 ( .A(n_508), .Y(n_601) );
AND2x2_ASAP7_75t_L g607 ( .A(n_508), .B(n_524), .Y(n_607) );
AND2x2_ASAP7_75t_L g675 ( .A(n_513), .B(n_583), .Y(n_675) );
INVx2_ASAP7_75t_L g740 ( .A(n_513), .Y(n_740) );
AND2x2_ASAP7_75t_L g513 ( .A(n_514), .B(n_524), .Y(n_513) );
AND2x2_ASAP7_75t_L g557 ( .A(n_514), .B(n_558), .Y(n_557) );
OR2x2_ASAP7_75t_L g570 ( .A(n_514), .B(n_532), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_514), .B(n_531), .Y(n_598) );
INVx1_ASAP7_75t_L g604 ( .A(n_514), .Y(n_604) );
INVx1_ASAP7_75t_L g621 ( .A(n_514), .Y(n_621) );
HB1xp67_ASAP7_75t_L g633 ( .A(n_514), .Y(n_633) );
INVx2_ASAP7_75t_L g701 ( .A(n_514), .Y(n_701) );
AOI21xp5_ASAP7_75t_L g516 ( .A1(n_517), .A2(n_518), .B(n_519), .Y(n_516) );
INVx2_ASAP7_75t_L g558 ( .A(n_524), .Y(n_558) );
BUFx2_ASAP7_75t_L g655 ( .A(n_524), .Y(n_655) );
AND2x2_ASAP7_75t_L g700 ( .A(n_524), .B(n_701), .Y(n_700) );
INVx1_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_530), .B(n_542), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_530), .B(n_637), .Y(n_636) );
AOI21xp5_ASAP7_75t_L g723 ( .A1(n_530), .A2(n_699), .B(n_713), .Y(n_723) );
AND2x2_ASAP7_75t_L g748 ( .A(n_530), .B(n_634), .Y(n_748) );
BUFx2_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
INVx2_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
INVx1_ASAP7_75t_L g670 ( .A(n_532), .Y(n_670) );
AND2x2_ASAP7_75t_L g699 ( .A(n_532), .B(n_700), .Y(n_699) );
INVx2_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
HB1xp67_ASAP7_75t_L g583 ( .A(n_533), .Y(n_583) );
INVx2_ASAP7_75t_L g602 ( .A(n_533), .Y(n_602) );
OR2x2_ASAP7_75t_L g603 ( .A(n_533), .B(n_604), .Y(n_603) );
AND2x2_ASAP7_75t_L g542 ( .A(n_543), .B(n_544), .Y(n_542) );
INVx2_ASAP7_75t_L g556 ( .A(n_543), .Y(n_556) );
OR2x2_ASAP7_75t_L g569 ( .A(n_543), .B(n_570), .Y(n_569) );
AND2x2_ASAP7_75t_L g637 ( .A(n_543), .B(n_633), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_543), .B(n_733), .Y(n_732) );
OR2x2_ASAP7_75t_L g738 ( .A(n_543), .B(n_739), .Y(n_738) );
NAND2xp5_ASAP7_75t_L g750 ( .A(n_543), .B(n_675), .Y(n_750) );
AND2x2_ASAP7_75t_L g629 ( .A(n_544), .B(n_630), .Y(n_629) );
AND2x2_ASAP7_75t_L g652 ( .A(n_544), .B(n_546), .Y(n_652) );
INVx2_ASAP7_75t_L g564 ( .A(n_545), .Y(n_564) );
AND2x2_ASAP7_75t_L g592 ( .A(n_545), .B(n_565), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_545), .B(n_617), .Y(n_673) );
AND2x2_ASAP7_75t_L g587 ( .A(n_546), .B(n_588), .Y(n_587) );
INVx1_ASAP7_75t_L g734 ( .A(n_546), .Y(n_734) );
AND2x2_ASAP7_75t_L g746 ( .A(n_546), .B(n_609), .Y(n_746) );
AND2x2_ASAP7_75t_L g572 ( .A(n_547), .B(n_562), .Y(n_572) );
INVx1_ASAP7_75t_L g667 ( .A(n_547), .Y(n_667) );
INVx1_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
AND2x4_ASAP7_75t_L g565 ( .A(n_552), .B(n_566), .Y(n_565) );
INVxp67_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_555), .B(n_559), .Y(n_554) );
AND2x2_ASAP7_75t_L g555 ( .A(n_556), .B(n_557), .Y(n_555) );
NOR2xp33_ASAP7_75t_L g612 ( .A(n_556), .B(n_603), .Y(n_612) );
OR2x2_ASAP7_75t_L g744 ( .A(n_556), .B(n_745), .Y(n_744) );
AND2x2_ASAP7_75t_L g661 ( .A(n_557), .B(n_602), .Y(n_661) );
AND2x2_ASAP7_75t_L g669 ( .A(n_557), .B(n_670), .Y(n_669) );
AND2x2_ASAP7_75t_L g728 ( .A(n_557), .B(n_729), .Y(n_728) );
AND2x2_ASAP7_75t_L g752 ( .A(n_557), .B(n_599), .Y(n_752) );
NOR2xp67_ASAP7_75t_L g710 ( .A(n_558), .B(n_711), .Y(n_710) );
OR2x2_ASAP7_75t_L g739 ( .A(n_558), .B(n_602), .Y(n_739) );
INVx1_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
NAND2x1p5_ASAP7_75t_L g560 ( .A(n_561), .B(n_563), .Y(n_560) );
AND2x2_ASAP7_75t_L g591 ( .A(n_561), .B(n_592), .Y(n_591) );
INVxp67_ASAP7_75t_L g753 ( .A(n_561), .Y(n_753) );
NOR2x1_ASAP7_75t_L g563 ( .A(n_564), .B(n_565), .Y(n_563) );
INVx1_ASAP7_75t_L g588 ( .A(n_564), .Y(n_588) );
AND2x2_ASAP7_75t_L g639 ( .A(n_564), .B(n_572), .Y(n_639) );
NOR2xp33_ASAP7_75t_L g733 ( .A(n_564), .B(n_707), .Y(n_733) );
INVx2_ASAP7_75t_L g578 ( .A(n_565), .Y(n_578) );
INVx3_ASAP7_75t_L g630 ( .A(n_565), .Y(n_630) );
OR2x2_ASAP7_75t_L g658 ( .A(n_565), .B(n_659), .Y(n_658) );
AOI311xp33_ASAP7_75t_L g567 ( .A1(n_568), .A2(n_571), .A3(n_573), .B(n_574), .C(n_585), .Y(n_567) );
O2A1O1Ixp33_ASAP7_75t_L g605 ( .A1(n_568), .A2(n_606), .B(n_608), .C(n_610), .Y(n_605) );
INVx2_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
INVx2_ASAP7_75t_SL g590 ( .A(n_570), .Y(n_590) );
INVx2_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
AND2x2_ASAP7_75t_L g608 ( .A(n_572), .B(n_609), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_572), .B(n_588), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g741 ( .A(n_572), .B(n_573), .Y(n_741) );
AND2x2_ASAP7_75t_L g663 ( .A(n_573), .B(n_577), .Y(n_663) );
AOI21xp33_ASAP7_75t_L g574 ( .A1(n_575), .A2(n_579), .B(n_580), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
AND2x2_ASAP7_75t_L g721 ( .A(n_577), .B(n_609), .Y(n_721) );
INVx2_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
NOR2xp33_ASAP7_75t_L g594 ( .A(n_578), .B(n_595), .Y(n_594) );
INVx1_ASAP7_75t_L g615 ( .A(n_578), .Y(n_615) );
INVx1_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
AND2x2_ASAP7_75t_L g581 ( .A(n_582), .B(n_584), .Y(n_581) );
AND2x2_ASAP7_75t_L g606 ( .A(n_582), .B(n_607), .Y(n_606) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
INVx1_ASAP7_75t_L g651 ( .A(n_584), .Y(n_651) );
AND2x4_ASAP7_75t_L g713 ( .A(n_584), .B(n_682), .Y(n_713) );
INVx1_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
AOI222xp33_ASAP7_75t_L g664 ( .A1(n_587), .A2(n_653), .B1(n_665), .B2(n_669), .C1(n_671), .C2(n_675), .Y(n_664) );
A2O1A1Ixp33_ASAP7_75t_L g589 ( .A1(n_590), .A2(n_591), .B(n_593), .C(n_596), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_590), .B(n_634), .Y(n_657) );
INVx1_ASAP7_75t_L g679 ( .A(n_592), .Y(n_679) );
INVx1_ASAP7_75t_L g613 ( .A(n_594), .Y(n_613) );
OR2x2_ASAP7_75t_L g678 ( .A(n_595), .B(n_679), .Y(n_678) );
OAI21xp33_ASAP7_75t_SL g596 ( .A1(n_597), .A2(n_599), .B(n_603), .Y(n_596) );
NAND3xp33_ASAP7_75t_L g614 ( .A(n_597), .B(n_615), .C(n_616), .Y(n_614) );
AOI21xp5_ASAP7_75t_L g712 ( .A1(n_597), .A2(n_634), .B(n_713), .Y(n_712) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
INVx1_ASAP7_75t_SL g599 ( .A(n_600), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_601), .B(n_602), .Y(n_600) );
HB1xp67_ASAP7_75t_L g654 ( .A(n_601), .Y(n_654) );
AND2x2_ASAP7_75t_SL g620 ( .A(n_602), .B(n_621), .Y(n_620) );
INVx1_ASAP7_75t_L g711 ( .A(n_602), .Y(n_711) );
HB1xp67_ASAP7_75t_L g727 ( .A(n_602), .Y(n_727) );
INVx2_ASAP7_75t_L g685 ( .A(n_603), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_607), .B(n_628), .Y(n_627) );
INVx2_ASAP7_75t_L g659 ( .A(n_609), .Y(n_659) );
OAI221xp5_ASAP7_75t_L g610 ( .A1(n_611), .A2(n_613), .B1(n_614), .B2(n_618), .C(n_619), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
NAND2xp5_ASAP7_75t_SL g692 ( .A(n_613), .B(n_693), .Y(n_692) );
INVx1_ASAP7_75t_SL g747 ( .A(n_613), .Y(n_747) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
INVx2_ASAP7_75t_L g628 ( .A(n_620), .Y(n_628) );
NOR2xp33_ASAP7_75t_L g650 ( .A(n_620), .B(n_651), .Y(n_650) );
AND2x2_ASAP7_75t_L g686 ( .A(n_620), .B(n_634), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_620), .B(n_696), .Y(n_695) );
AND2x2_ASAP7_75t_L g719 ( .A(n_620), .B(n_654), .Y(n_719) );
BUFx3_ASAP7_75t_L g682 ( .A(n_621), .Y(n_682) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
NAND5xp2_ASAP7_75t_L g624 ( .A(n_625), .B(n_643), .C(n_664), .D(n_676), .E(n_691), .Y(n_624) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
AOI32xp33_ASAP7_75t_L g716 ( .A1(n_628), .A2(n_655), .A3(n_671), .B1(n_717), .B2(n_719), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_630), .B(n_689), .Y(n_688) );
AND2x2_ASAP7_75t_L g631 ( .A(n_632), .B(n_634), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
INVx1_ASAP7_75t_SL g640 ( .A(n_634), .Y(n_640) );
OAI22xp5_ASAP7_75t_L g635 ( .A1(n_636), .A2(n_638), .B1(n_640), .B2(n_641), .Y(n_635) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
INVx1_ASAP7_75t_SL g641 ( .A(n_642), .Y(n_641) );
AOI221xp5_ASAP7_75t_L g643 ( .A1(n_644), .A2(n_650), .B1(n_652), .B2(n_653), .C(n_656), .Y(n_643) );
INVx2_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
OR2x2_ASAP7_75t_L g645 ( .A(n_646), .B(n_648), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
AND2x2_ASAP7_75t_L g715 ( .A(n_647), .B(n_666), .Y(n_715) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
AOI221xp5_ASAP7_75t_L g730 ( .A1(n_652), .A2(n_713), .B1(n_731), .B2(n_736), .C(n_737), .Y(n_730) );
AND2x2_ASAP7_75t_L g653 ( .A(n_654), .B(n_655), .Y(n_653) );
INVx2_ASAP7_75t_L g696 ( .A(n_655), .Y(n_696) );
OAI22xp5_ASAP7_75t_L g656 ( .A1(n_657), .A2(n_658), .B1(n_660), .B2(n_662), .Y(n_656) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
INVx1_ASAP7_75t_SL g662 ( .A(n_663), .Y(n_662) );
AND2x2_ASAP7_75t_L g665 ( .A(n_666), .B(n_668), .Y(n_665) );
INVx1_ASAP7_75t_L g674 ( .A(n_666), .Y(n_674) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
OR2x2_ASAP7_75t_L g672 ( .A(n_673), .B(n_674), .Y(n_672) );
AOI222xp33_ASAP7_75t_L g676 ( .A1(n_677), .A2(n_680), .B1(n_684), .B2(n_685), .C1(n_686), .C2(n_687), .Y(n_676) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
AND2x2_ASAP7_75t_L g680 ( .A(n_681), .B(n_683), .Y(n_680) );
INVxp67_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
OAI22xp33_ASAP7_75t_L g731 ( .A1(n_685), .A2(n_732), .B1(n_734), .B2(n_735), .Y(n_731) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
INVx1_ASAP7_75t_SL g689 ( .A(n_690), .Y(n_689) );
AOI21xp5_ASAP7_75t_L g691 ( .A1(n_692), .A2(n_694), .B(n_697), .Y(n_691) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
AOI21xp33_ASAP7_75t_L g697 ( .A1(n_698), .A2(n_702), .B(n_704), .Y(n_697) );
INVx2_ASAP7_75t_SL g698 ( .A(n_699), .Y(n_698) );
INVx1_ASAP7_75t_L g745 ( .A(n_700), .Y(n_745) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
INVx1_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
INVx1_ASAP7_75t_SL g706 ( .A(n_707), .Y(n_706) );
A2O1A1Ixp33_ASAP7_75t_L g708 ( .A1(n_709), .A2(n_712), .B(n_714), .C(n_716), .Y(n_708) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
INVx1_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
AOI211xp5_ASAP7_75t_L g720 ( .A1(n_721), .A2(n_722), .B(n_724), .C(n_749), .Y(n_720) );
CKINVDCx16_ASAP7_75t_R g725 ( .A(n_721), .Y(n_725) );
INVxp67_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
OAI211xp5_ASAP7_75t_L g724 ( .A1(n_725), .A2(n_726), .B(n_730), .C(n_742), .Y(n_724) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_727), .B(n_728), .Y(n_726) );
AOI21xp33_ASAP7_75t_L g737 ( .A1(n_738), .A2(n_740), .B(n_741), .Y(n_737) );
AOI22xp5_ASAP7_75t_L g742 ( .A1(n_743), .A2(n_746), .B1(n_747), .B2(n_748), .Y(n_742) );
INVx1_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
AOI21xp33_ASAP7_75t_L g749 ( .A1(n_750), .A2(n_751), .B(n_753), .Y(n_749) );
INVx1_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
INVx1_ASAP7_75t_SL g756 ( .A(n_757), .Y(n_756) );
INVx1_ASAP7_75t_SL g760 ( .A(n_761), .Y(n_760) );
INVx1_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
INVx2_ASAP7_75t_L g762 ( .A(n_763), .Y(n_762) );
INVx2_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
INVx1_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
INVx1_ASAP7_75t_SL g768 ( .A(n_769), .Y(n_768) );
endmodule