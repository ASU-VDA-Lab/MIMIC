module fake_jpeg_27363_n_337 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_337);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_337;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_11),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_14),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_15),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_7),
.B(n_0),
.Y(n_28)
);

INVx11_ASAP7_75t_SL g29 ( 
.A(n_6),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

INVx13_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_35),
.Y(n_37)
);

INVx1_ASAP7_75t_SL g55 ( 
.A(n_37),
.Y(n_55)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_34),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_38),
.B(n_39),
.Y(n_58)
);

INVx2_ASAP7_75t_SL g39 ( 
.A(n_29),
.Y(n_39)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_44),
.B(n_45),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx2_ASAP7_75t_SL g69 ( 
.A(n_46),
.Y(n_69)
);

BUFx16f_ASAP7_75t_L g47 ( 
.A(n_26),
.Y(n_47)
);

CKINVDCx14_ASAP7_75t_R g51 ( 
.A(n_47),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_41),
.B(n_28),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_48),
.B(n_54),
.Y(n_72)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_52),
.Y(n_85)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_53),
.B(n_63),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_41),
.B(n_28),
.Y(n_54)
);

BUFx12_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_37),
.A2(n_19),
.B1(n_23),
.B2(n_34),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_57),
.A2(n_59),
.B1(n_46),
.B2(n_42),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_37),
.A2(n_19),
.B1(n_23),
.B2(n_34),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_42),
.A2(n_19),
.B1(n_23),
.B2(n_30),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_62),
.A2(n_46),
.B1(n_33),
.B2(n_25),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_43),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_64),
.B(n_43),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_44),
.B(n_28),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_65),
.B(n_68),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_44),
.B(n_28),
.Y(n_68)
);

OR2x2_ASAP7_75t_SL g70 ( 
.A(n_48),
.B(n_17),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_70),
.B(n_73),
.Y(n_111)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_67),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_67),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_74),
.B(n_78),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_54),
.B(n_36),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_75),
.B(n_88),
.C(n_91),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_65),
.B(n_33),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_77),
.B(n_81),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_58),
.B(n_17),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_58),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_79),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_62),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_80),
.B(n_84),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_68),
.B(n_36),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_66),
.Y(n_82)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_82),
.Y(n_108)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_66),
.Y(n_83)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_83),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_57),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_59),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_86),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_63),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_87),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_55),
.B(n_25),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_53),
.B(n_18),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_89),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_90),
.A2(n_40),
.B1(n_52),
.B2(n_30),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_55),
.B(n_25),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_69),
.Y(n_92)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_92),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_55),
.A2(n_32),
.B1(n_18),
.B2(n_20),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_93),
.A2(n_24),
.B1(n_27),
.B2(n_26),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_52),
.Y(n_94)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_94),
.Y(n_132)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_69),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_95),
.A2(n_100),
.B1(n_104),
.B2(n_105),
.Y(n_112)
);

OR2x2_ASAP7_75t_L g130 ( 
.A(n_97),
.B(n_98),
.Y(n_130)
);

NAND3xp33_ASAP7_75t_L g98 ( 
.A(n_50),
.B(n_11),
.C(n_15),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_56),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_99),
.Y(n_123)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_69),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_64),
.B(n_36),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_101),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_51),
.B(n_20),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_102),
.Y(n_129)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_60),
.Y(n_103)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_103),
.Y(n_127)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_69),
.Y(n_104)
);

BUFx4f_ASAP7_75t_SL g106 ( 
.A(n_56),
.Y(n_106)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_106),
.Y(n_131)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_106),
.Y(n_109)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_109),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_84),
.A2(n_49),
.B1(n_61),
.B2(n_38),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_110),
.A2(n_116),
.B1(n_117),
.B2(n_126),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_80),
.A2(n_50),
.B1(n_49),
.B2(n_61),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_113),
.Y(n_139)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_106),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_114),
.B(n_71),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_90),
.A2(n_49),
.B1(n_61),
.B2(n_50),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_81),
.A2(n_40),
.B1(n_51),
.B2(n_33),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_118),
.A2(n_93),
.B1(n_91),
.B2(n_88),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_75),
.A2(n_32),
.B1(n_35),
.B2(n_43),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_119),
.A2(n_135),
.B1(n_134),
.B2(n_133),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_75),
.A2(n_27),
.B1(n_24),
.B2(n_31),
.Y(n_135)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_110),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_137),
.B(n_145),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_124),
.B(n_76),
.C(n_72),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_138),
.B(n_146),
.C(n_149),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_136),
.A2(n_77),
.B(n_79),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_140),
.A2(n_164),
.B(n_168),
.Y(n_180)
);

CKINVDCx14_ASAP7_75t_R g186 ( 
.A(n_141),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_107),
.B(n_72),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_142),
.B(n_153),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_136),
.A2(n_73),
.B1(n_74),
.B2(n_87),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_144),
.A2(n_167),
.B1(n_132),
.B2(n_135),
.Y(n_172)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_116),
.Y(n_145)
);

MAJx2_ASAP7_75t_L g146 ( 
.A(n_124),
.B(n_76),
.C(n_70),
.Y(n_146)
);

BUFx24_ASAP7_75t_SL g147 ( 
.A(n_129),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_147),
.B(n_154),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_115),
.B(n_96),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_148),
.B(n_162),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_107),
.B(n_101),
.C(n_96),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_150),
.A2(n_157),
.B1(n_166),
.B2(n_117),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_112),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_151),
.B(n_152),
.Y(n_195)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_115),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_120),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_129),
.B(n_121),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_122),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_155),
.B(n_160),
.Y(n_194)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_120),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_156),
.B(n_163),
.Y(n_182)
);

MAJx2_ASAP7_75t_L g159 ( 
.A(n_111),
.B(n_97),
.C(n_26),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_159),
.B(n_131),
.C(n_31),
.Y(n_197)
);

BUFx5_ASAP7_75t_L g160 ( 
.A(n_109),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_121),
.B(n_82),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_161),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_122),
.B(n_83),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_128),
.B(n_104),
.Y(n_163)
);

OAI21x1_ASAP7_75t_L g164 ( 
.A1(n_126),
.A2(n_45),
.B(n_47),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_128),
.B(n_92),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_165),
.B(n_127),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_119),
.A2(n_100),
.B1(n_95),
.B2(n_103),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_114),
.A2(n_85),
.B1(n_106),
.B2(n_56),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_130),
.A2(n_111),
.B(n_134),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_169),
.B(n_187),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_172),
.A2(n_198),
.B(n_159),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_145),
.A2(n_132),
.B1(n_125),
.B2(n_108),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_173),
.A2(n_179),
.B1(n_189),
.B2(n_60),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_138),
.B(n_130),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_174),
.B(n_202),
.C(n_31),
.Y(n_213)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_158),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_175),
.B(n_191),
.Y(n_219)
);

HB1xp67_ASAP7_75t_L g176 ( 
.A(n_163),
.Y(n_176)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_176),
.Y(n_231)
);

HB1xp67_ASAP7_75t_L g177 ( 
.A(n_165),
.Y(n_177)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_177),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_137),
.A2(n_108),
.B1(n_125),
.B2(n_130),
.Y(n_179)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_166),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_183),
.B(n_190),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_150),
.A2(n_127),
.B1(n_123),
.B2(n_94),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_184),
.A2(n_47),
.B1(n_60),
.B2(n_22),
.Y(n_215)
);

INVx13_ASAP7_75t_L g187 ( 
.A(n_160),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_188),
.B(n_199),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_151),
.A2(n_85),
.B1(n_131),
.B2(n_123),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_168),
.B(n_21),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_152),
.B(n_21),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_153),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_192),
.B(n_196),
.Y(n_229)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_156),
.Y(n_196)
);

XNOR2x1_ASAP7_75t_L g214 ( 
.A(n_197),
.B(n_47),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_139),
.A2(n_0),
.B(n_1),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_142),
.B(n_45),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_144),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_200),
.B(n_201),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_149),
.B(n_31),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_146),
.B(n_56),
.C(n_85),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_170),
.A2(n_183),
.B1(n_169),
.B2(n_200),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_203),
.A2(n_220),
.B1(n_227),
.B2(n_199),
.Y(n_233)
);

OAI32xp33_ASAP7_75t_L g204 ( 
.A1(n_182),
.A2(n_140),
.A3(n_157),
.B1(n_164),
.B2(n_143),
.Y(n_204)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_204),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_195),
.A2(n_139),
.B(n_143),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g240 ( 
.A1(n_205),
.A2(n_211),
.B(n_217),
.Y(n_240)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_188),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_207),
.B(n_212),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_185),
.B(n_158),
.Y(n_209)
);

CKINVDCx14_ASAP7_75t_R g251 ( 
.A(n_209),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_194),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_210),
.Y(n_232)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_182),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_213),
.B(n_225),
.C(n_197),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_214),
.B(n_202),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_215),
.B(n_216),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_185),
.B(n_71),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_180),
.A2(n_0),
.B(n_1),
.Y(n_217)
);

OAI32xp33_ASAP7_75t_L g221 ( 
.A1(n_179),
.A2(n_22),
.A3(n_21),
.B1(n_8),
.B2(n_10),
.Y(n_221)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_221),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_180),
.A2(n_1),
.B(n_2),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_222),
.Y(n_247)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_173),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_223),
.B(n_220),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_191),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_224),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_193),
.B(n_22),
.C(n_14),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_184),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_178),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_230),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_233),
.A2(n_203),
.B1(n_223),
.B2(n_208),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_213),
.B(n_193),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_SL g256 ( 
.A(n_234),
.B(n_241),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_237),
.B(n_214),
.Y(n_265)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_229),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_242),
.B(n_243),
.Y(n_269)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_229),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_224),
.B(n_186),
.Y(n_244)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_244),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_225),
.B(n_201),
.C(n_174),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_245),
.B(n_250),
.C(n_211),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_210),
.B(n_187),
.Y(n_246)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_246),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_219),
.B(n_175),
.Y(n_248)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_248),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_226),
.B(n_178),
.C(n_172),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_252),
.B(n_254),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_219),
.Y(n_253)
);

A2O1A1Ixp33_ASAP7_75t_SL g272 ( 
.A1(n_253),
.A2(n_228),
.B(n_190),
.C(n_222),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_230),
.B(n_181),
.Y(n_254)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_253),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_257),
.B(n_261),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_258),
.A2(n_252),
.B1(n_254),
.B2(n_255),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_232),
.B(n_171),
.Y(n_260)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_260),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_232),
.B(n_226),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_235),
.A2(n_227),
.B1(n_215),
.B2(n_189),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_263),
.B(n_233),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_236),
.A2(n_205),
.B1(n_228),
.B2(n_181),
.Y(n_264)
);

AOI322xp5_ASAP7_75t_L g276 ( 
.A1(n_264),
.A2(n_240),
.A3(n_238),
.B1(n_249),
.B2(n_255),
.C1(n_221),
.C2(n_236),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_265),
.B(n_270),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_266),
.B(n_275),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_251),
.B(n_231),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_267),
.B(n_239),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_234),
.B(n_204),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_272),
.A2(n_247),
.B(n_240),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_245),
.B(n_207),
.C(n_218),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_273),
.B(n_237),
.C(n_250),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_235),
.A2(n_231),
.B1(n_206),
.B2(n_212),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_274),
.A2(n_238),
.B(n_243),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_SL g275 ( 
.A(n_241),
.B(n_218),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_276),
.B(n_272),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_277),
.A2(n_283),
.B(n_272),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_278),
.B(n_285),
.C(n_289),
.Y(n_295)
);

CKINVDCx14_ASAP7_75t_R g300 ( 
.A(n_279),
.Y(n_300)
);

OA21x2_ASAP7_75t_L g298 ( 
.A1(n_280),
.A2(n_270),
.B(n_272),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_281),
.A2(n_291),
.B1(n_292),
.B2(n_268),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_269),
.A2(n_247),
.B(n_242),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_256),
.B(n_239),
.C(n_206),
.Y(n_285)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_286),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_256),
.B(n_196),
.C(n_192),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_266),
.B(n_217),
.C(n_198),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_290),
.B(n_275),
.C(n_9),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_274),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_273),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_288),
.B(n_262),
.Y(n_293)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_293),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_283),
.Y(n_294)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_294),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_296),
.B(n_302),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_280),
.A2(n_271),
.B(n_259),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_SL g311 ( 
.A1(n_297),
.A2(n_290),
.B(n_292),
.Y(n_311)
);

OA21x2_ASAP7_75t_L g317 ( 
.A1(n_298),
.A2(n_299),
.B(n_9),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g302 ( 
.A(n_277),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_287),
.B(n_10),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_303),
.B(n_304),
.Y(n_315)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_281),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_305),
.B(n_284),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_306),
.B(n_291),
.C(n_284),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_295),
.B(n_278),
.C(n_289),
.Y(n_309)
);

OR2x2_ASAP7_75t_L g325 ( 
.A(n_309),
.B(n_310),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_295),
.B(n_285),
.C(n_282),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g319 ( 
.A1(n_311),
.A2(n_317),
.B(n_294),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_299),
.B(n_282),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_312),
.B(n_316),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_SL g323 ( 
.A(n_314),
.B(n_306),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_308),
.B(n_301),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g326 ( 
.A1(n_318),
.A2(n_321),
.B(n_322),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_L g329 ( 
.A1(n_319),
.A2(n_320),
.B(n_14),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_L g320 ( 
.A1(n_313),
.A2(n_302),
.B(n_298),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_SL g321 ( 
.A1(n_315),
.A2(n_307),
.B(n_317),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_SL g322 ( 
.A1(n_317),
.A2(n_300),
.B(n_296),
.Y(n_322)
);

AND2x2_ASAP7_75t_L g330 ( 
.A(n_323),
.B(n_324),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_325),
.B(n_309),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g331 ( 
.A1(n_327),
.A2(n_328),
.B(n_329),
.Y(n_331)
);

A2O1A1Ixp33_ASAP7_75t_L g328 ( 
.A1(n_318),
.A2(n_310),
.B(n_298),
.C(n_312),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_330),
.B(n_12),
.C(n_11),
.Y(n_332)
);

AOI321xp33_ASAP7_75t_L g333 ( 
.A1(n_332),
.A2(n_326),
.A3(n_12),
.B1(n_10),
.B2(n_6),
.C(n_3),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_333),
.B(n_331),
.C(n_12),
.Y(n_334)
);

AOI21xp5_ASAP7_75t_L g335 ( 
.A1(n_334),
.A2(n_4),
.B(n_5),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_335),
.B(n_5),
.Y(n_336)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_336),
.B(n_7),
.Y(n_337)
);


endmodule