module fake_jpeg_18023_n_85 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_8, n_15, n_7, n_85);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_8;
input n_15;
input n_7;

output n_85;

wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_30),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_23),
.B(n_24),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_27),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

CKINVDCx14_ASAP7_75t_R g41 ( 
.A(n_31),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

BUFx2_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_36),
.B(n_0),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_44),
.B(n_47),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_46),
.B(n_51),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_36),
.B(n_1),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_50),
.Y(n_54)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

BUFx12f_ASAP7_75t_SL g52 ( 
.A(n_51),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_52),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_44),
.B(n_34),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_53),
.B(n_3),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_44),
.B(n_41),
.Y(n_59)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_59),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_49),
.A2(n_43),
.B1(n_39),
.B2(n_32),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_60),
.A2(n_7),
.B1(n_8),
.B2(n_10),
.Y(n_67)
);

AND2x2_ASAP7_75t_SL g70 ( 
.A(n_62),
.B(n_64),
.Y(n_70)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_61),
.Y(n_63)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_63),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_55),
.Y(n_65)
);

O2A1O1Ixp33_ASAP7_75t_L g71 ( 
.A1(n_65),
.A2(n_66),
.B(n_67),
.C(n_57),
.Y(n_71)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_58),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_71),
.B(n_62),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_70),
.A2(n_56),
.B1(n_68),
.B2(n_69),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_72),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_73),
.B(n_74),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_71),
.B(n_54),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_L g77 ( 
.A1(n_75),
.A2(n_11),
.B(n_13),
.Y(n_77)
);

XOR2xp5_ASAP7_75t_L g78 ( 
.A(n_77),
.B(n_14),
.Y(n_78)
);

A2O1A1Ixp33_ASAP7_75t_SL g79 ( 
.A1(n_78),
.A2(n_15),
.B(n_16),
.C(n_17),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_79),
.B(n_18),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_80),
.B(n_21),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_81),
.B(n_22),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_82),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_83),
.A2(n_76),
.B1(n_26),
.B2(n_29),
.Y(n_84)
);

XOR2xp5_ASAP7_75t_L g85 ( 
.A(n_84),
.B(n_25),
.Y(n_85)
);


endmodule