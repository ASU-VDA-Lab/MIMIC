module real_jpeg_15938_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_646, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_646;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_598;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_630;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_643;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_640;
wire n_160;
wire n_211;
wire n_574;
wire n_627;
wire n_595;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_578;
wire n_456;
wire n_620;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_623;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_216;
wire n_202;
wire n_605;
wire n_483;
wire n_367;
wire n_639;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_621;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_601;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_393;
wire n_221;
wire n_489;
wire n_611;
wire n_104;
wire n_153;
wire n_634;
wire n_443;
wire n_599;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_607;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_98;
wire n_469;
wire n_378;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_214;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_631;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_470;
wire n_219;
wire n_372;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_593;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_590;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_612;
wire n_110;
wire n_195;
wire n_592;
wire n_533;
wire n_289;
wire n_117;
wire n_614;
wire n_193;
wire n_382;
wire n_411;
wire n_278;
wire n_314;
wire n_103;
wire n_559;
wire n_232;
wire n_582;
wire n_448;
wire n_615;
wire n_212;
wire n_579;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_583;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_589;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_644;
wire n_515;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_632;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_638;
wire n_497;
wire n_633;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_596;
wire n_617;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_594;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_604;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_586;
wire n_572;
wire n_548;
wire n_319;
wire n_487;
wire n_93;
wire n_242;
wire n_493;
wire n_637;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_613;
wire n_231;
wire n_44;
wire n_635;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_642;
wire n_172;
wire n_285;
wire n_531;
wire n_546;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_616;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_600;
wire n_392;
wire n_575;
wire n_375;
wire n_196;
wire n_298;
wire n_330;
wire n_450;
wire n_333;
wire n_492;
wire n_152;
wire n_584;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_622;
wire n_183;
wire n_248;
wire n_192;
wire n_624;
wire n_318;
wire n_537;
wire n_603;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_628;
wire n_413;
wire n_585;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_581;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_534;
wire n_181;
wire n_358;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_587;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_608;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_602;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_610;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_636;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_606;
wire n_245;
wire n_451;
wire n_626;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_597;
wire n_618;
wire n_609;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_619;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_588;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_568;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_130;
wire n_641;
wire n_225;
wire n_43;
wire n_438;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_629;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_591;
wire n_625;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

AND2x2_ASAP7_75t_L g22 ( 
.A(n_0),
.B(n_23),
.Y(n_22)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_1),
.A2(n_189),
.B1(n_191),
.B2(n_193),
.Y(n_188)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_1),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_1),
.A2(n_193),
.B1(n_382),
.B2(n_383),
.Y(n_381)
);

AOI22xp33_ASAP7_75t_L g592 ( 
.A1(n_1),
.A2(n_193),
.B1(n_593),
.B2(n_595),
.Y(n_592)
);

AOI22xp33_ASAP7_75t_SL g627 ( 
.A1(n_1),
.A2(n_193),
.B1(n_628),
.B2(n_631),
.Y(n_627)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_2),
.Y(n_112)
);

BUFx5_ASAP7_75t_L g133 ( 
.A(n_2),
.Y(n_133)
);

BUFx5_ASAP7_75t_L g344 ( 
.A(n_2),
.Y(n_344)
);

BUFx3_ASAP7_75t_L g449 ( 
.A(n_2),
.Y(n_449)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_3),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_3),
.B(n_174),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_3),
.B(n_285),
.Y(n_459)
);

OAI22xp5_ASAP7_75t_SL g490 ( 
.A1(n_3),
.A2(n_109),
.B1(n_491),
.B2(n_497),
.Y(n_490)
);

OAI32xp33_ASAP7_75t_L g508 ( 
.A1(n_3),
.A2(n_53),
.A3(n_432),
.B1(n_509),
.B2(n_513),
.Y(n_508)
);

AOI22xp33_ASAP7_75t_SL g522 ( 
.A1(n_3),
.A2(n_85),
.B1(n_523),
.B2(n_527),
.Y(n_522)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_4),
.Y(n_93)
);

INVx6_ASAP7_75t_L g155 ( 
.A(n_4),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_4),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_5),
.A2(n_86),
.B1(n_144),
.B2(n_145),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_5),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g315 ( 
.A1(n_5),
.A2(n_144),
.B1(n_316),
.B2(n_320),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g434 ( 
.A1(n_5),
.A2(n_144),
.B1(n_435),
.B2(n_438),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_SL g491 ( 
.A1(n_5),
.A2(n_144),
.B1(n_492),
.B2(n_496),
.Y(n_491)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_6),
.A2(n_21),
.B(n_22),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_7),
.A2(n_119),
.B1(n_123),
.B2(n_124),
.Y(n_118)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_7),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_7),
.A2(n_123),
.B1(n_229),
.B2(n_233),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_SL g356 ( 
.A1(n_7),
.A2(n_123),
.B1(n_357),
.B2(n_362),
.Y(n_356)
);

AOI22xp33_ASAP7_75t_SL g573 ( 
.A1(n_7),
.A2(n_123),
.B1(n_574),
.B2(n_575),
.Y(n_573)
);

AOI22xp33_ASAP7_75t_L g179 ( 
.A1(n_8),
.A2(n_125),
.B1(n_180),
.B2(n_183),
.Y(n_179)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_8),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g333 ( 
.A1(n_8),
.A2(n_183),
.B1(n_334),
.B2(n_336),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g579 ( 
.A1(n_8),
.A2(n_99),
.B1(n_183),
.B2(n_580),
.Y(n_579)
);

AOI22xp33_ASAP7_75t_SL g617 ( 
.A1(n_8),
.A2(n_183),
.B1(n_618),
.B2(n_619),
.Y(n_617)
);

BUFx5_ASAP7_75t_L g199 ( 
.A(n_9),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_9),
.Y(n_203)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_9),
.Y(n_220)
);

BUFx5_ASAP7_75t_L g418 ( 
.A(n_9),
.Y(n_418)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_10),
.Y(n_116)
);

BUFx12f_ASAP7_75t_L g122 ( 
.A(n_10),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_10),
.Y(n_130)
);

BUFx4f_ASAP7_75t_L g428 ( 
.A(n_10),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_11),
.A2(n_167),
.B1(n_170),
.B2(n_171),
.Y(n_166)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_11),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_11),
.A2(n_94),
.B1(n_170),
.B2(n_283),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g462 ( 
.A1(n_11),
.A2(n_170),
.B1(n_210),
.B2(n_463),
.Y(n_462)
);

AOI22xp33_ASAP7_75t_SL g469 ( 
.A1(n_11),
.A2(n_170),
.B1(n_470),
.B2(n_473),
.Y(n_469)
);

OAI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_12),
.A2(n_34),
.B1(n_39),
.B2(n_40),
.Y(n_33)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_12),
.A2(n_39),
.B1(n_257),
.B2(n_260),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g442 ( 
.A1(n_12),
.A2(n_39),
.B1(n_443),
.B2(n_445),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_L g531 ( 
.A1(n_12),
.A2(n_39),
.B1(n_532),
.B2(n_534),
.Y(n_531)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_13),
.Y(n_50)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_13),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_14),
.A2(n_135),
.B1(n_139),
.B2(n_141),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_14),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_L g205 ( 
.A1(n_14),
.A2(n_141),
.B1(n_206),
.B2(n_210),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_14),
.A2(n_74),
.B1(n_141),
.B2(n_376),
.Y(n_375)
);

OAI22xp33_ASAP7_75t_SL g601 ( 
.A1(n_14),
.A2(n_141),
.B1(n_148),
.B2(n_289),
.Y(n_601)
);

AOI22xp33_ASAP7_75t_L g239 ( 
.A1(n_15),
.A2(n_240),
.B1(n_244),
.B2(n_245),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_15),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_15),
.A2(n_244),
.B1(n_266),
.B2(n_270),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_15),
.A2(n_244),
.B1(n_305),
.B2(n_308),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_15),
.A2(n_244),
.B1(n_394),
.B2(n_396),
.Y(n_393)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_16),
.Y(n_64)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_16),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g209 ( 
.A(n_16),
.Y(n_209)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_16),
.Y(n_214)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_16),
.Y(n_232)
);

BUFx3_ASAP7_75t_L g243 ( 
.A(n_16),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g295 ( 
.A(n_16),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_17),
.A2(n_73),
.B1(n_78),
.B2(n_79),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_17),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_17),
.A2(n_78),
.B1(n_292),
.B2(n_293),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_17),
.A2(n_78),
.B1(n_350),
.B2(n_352),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_SL g451 ( 
.A1(n_17),
.A2(n_78),
.B1(n_452),
.B2(n_454),
.Y(n_451)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g88 ( 
.A(n_19),
.Y(n_88)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_19),
.Y(n_107)
);

BUFx5_ASAP7_75t_L g150 ( 
.A(n_19),
.Y(n_150)
);

BUFx3_ASAP7_75t_L g169 ( 
.A(n_19),
.Y(n_169)
);

BUFx8_ASAP7_75t_L g351 ( 
.A(n_19),
.Y(n_351)
);

AOI21xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_639),
.B(n_643),
.Y(n_23)
);

AO21x1_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_564),
.B(n_632),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_401),
.B(n_559),
.Y(n_25)
);

NAND3xp33_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_326),
.C(n_367),
.Y(n_26)
);

AOI21xp33_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_273),
.B(n_297),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g560 ( 
.A(n_28),
.B(n_273),
.C(n_561),
.Y(n_560)
);

XNOR2xp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_175),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_29),
.B(n_176),
.C(n_235),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_82),
.C(n_142),
.Y(n_29)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_31),
.B(n_142),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_32),
.A2(n_44),
.B1(n_72),
.B2(n_80),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_33),
.A2(n_281),
.B1(n_282),
.B2(n_285),
.Y(n_280)
);

HB1xp67_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_37),
.Y(n_272)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_37),
.Y(n_378)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_38),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g269 ( 
.A(n_38),
.Y(n_269)
);

BUFx5_ASAP7_75t_L g526 ( 
.A(n_38),
.Y(n_526)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_42),
.Y(n_319)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_43),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_43),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g321 ( 
.A(n_43),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_44),
.A2(n_72),
.B1(n_80),
.B2(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_44),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g355 ( 
.A1(n_44),
.A2(n_80),
.B1(n_265),
.B2(n_356),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_SL g521 ( 
.A1(n_44),
.A2(n_80),
.B1(n_315),
.B2(n_522),
.Y(n_521)
);

OAI22x1_ASAP7_75t_L g578 ( 
.A1(n_44),
.A2(n_80),
.B1(n_375),
.B2(n_579),
.Y(n_578)
);

OAI22xp5_ASAP7_75t_L g591 ( 
.A1(n_44),
.A2(n_80),
.B1(n_579),
.B2(n_592),
.Y(n_591)
);

AO21x2_ASAP7_75t_L g44 ( 
.A1(n_45),
.A2(n_53),
.B(n_61),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_51),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_50),
.Y(n_67)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_58),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_58),
.Y(n_594)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_60),
.Y(n_98)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_61),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_62),
.A2(n_65),
.B1(n_68),
.B2(n_71),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx4_ASAP7_75t_L g385 ( 
.A(n_63),
.Y(n_385)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_64),
.Y(n_222)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g537 ( 
.A(n_69),
.Y(n_537)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_70),
.Y(n_247)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_70),
.Y(n_423)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

HB1xp67_ASAP7_75t_L g79 ( 
.A(n_74),
.Y(n_79)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx6_ASAP7_75t_L g163 ( 
.A(n_77),
.Y(n_163)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_80),
.Y(n_285)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_82),
.B(n_276),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_83),
.B(n_108),
.Y(n_82)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_83),
.B(n_108),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_89),
.B1(n_99),
.B2(n_103),
.Y(n_83)
);

OAI21xp33_ASAP7_75t_SL g287 ( 
.A1(n_84),
.A2(n_85),
.B(n_288),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_86),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_85),
.B(n_420),
.Y(n_419)
);

OAI21xp33_ASAP7_75t_SL g431 ( 
.A1(n_85),
.A2(n_419),
.B(n_432),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_SL g486 ( 
.A(n_85),
.B(n_487),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_85),
.B(n_197),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_85),
.B(n_234),
.Y(n_513)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g354 ( 
.A(n_88),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_94),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_92),
.B(n_105),
.Y(n_104)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_95),
.Y(n_580)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g512 ( 
.A(n_102),
.Y(n_512)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

OA21x2_ASAP7_75t_L g151 ( 
.A1(n_104),
.A2(n_152),
.B(n_158),
.Y(n_151)
);

INVx6_ASAP7_75t_L g397 ( 
.A(n_105),
.Y(n_397)
);

BUFx2_ASAP7_75t_L g631 ( 
.A(n_105),
.Y(n_631)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx4_ASAP7_75t_L g259 ( 
.A(n_106),
.Y(n_259)
);

INVx5_ASAP7_75t_L g262 ( 
.A(n_106),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g630 ( 
.A(n_106),
.Y(n_630)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_107),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_109),
.A2(n_117),
.B1(n_131),
.B2(n_134),
.Y(n_108)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_109),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_109),
.A2(n_134),
.B1(n_179),
.B2(n_249),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_SL g341 ( 
.A1(n_109),
.A2(n_188),
.B(n_342),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_L g441 ( 
.A1(n_109),
.A2(n_442),
.B1(n_447),
.B2(n_450),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_SL g499 ( 
.A1(n_109),
.A2(n_131),
.B1(n_469),
.B2(n_491),
.Y(n_499)
);

OR2x2_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_113),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g489 ( 
.A(n_110),
.Y(n_489)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_110),
.Y(n_497)
);

INVx4_ASAP7_75t_SL g516 ( 
.A(n_110),
.Y(n_516)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_111),
.Y(n_252)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_112),
.Y(n_186)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g414 ( 
.A(n_116),
.Y(n_414)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_118),
.A2(n_184),
.B1(n_304),
.B2(n_311),
.Y(n_303)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

BUFx2_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx3_ASAP7_75t_L g444 ( 
.A(n_121),
.Y(n_444)
);

INVx3_ASAP7_75t_L g453 ( 
.A(n_121),
.Y(n_453)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_122),
.Y(n_140)
);

INVx5_ASAP7_75t_L g182 ( 
.A(n_122),
.Y(n_182)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_122),
.Y(n_192)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_122),
.Y(n_310)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_129),
.Y(n_457)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_129),
.Y(n_495)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g138 ( 
.A(n_130),
.Y(n_138)
);

INVx6_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

BUFx12f_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_138),
.Y(n_474)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx3_ASAP7_75t_L g307 ( 
.A(n_140),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_143),
.A2(n_151),
.B1(n_165),
.B2(n_174),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_143),
.A2(n_151),
.B1(n_174),
.B2(n_287),
.Y(n_286)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx2_ASAP7_75t_SL g255 ( 
.A(n_151),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g599 ( 
.A1(n_151),
.A2(n_174),
.B1(n_600),
.B2(n_601),
.Y(n_599)
);

OAI21xp5_ASAP7_75t_SL g640 ( 
.A1(n_151),
.A2(n_174),
.B(n_641),
.Y(n_640)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_156),
.Y(n_152)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx3_ASAP7_75t_SL g154 ( 
.A(n_155),
.Y(n_154)
);

INVx3_ASAP7_75t_L g618 ( 
.A(n_156),
.Y(n_618)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx6_ASAP7_75t_L g395 ( 
.A(n_157),
.Y(n_395)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_158),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g348 ( 
.A1(n_158),
.A2(n_255),
.B1(n_256),
.B2(n_349),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_SL g392 ( 
.A1(n_158),
.A2(n_255),
.B1(n_349),
.B2(n_393),
.Y(n_392)
);

AOI22x1_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_161),
.B1(n_163),
.B2(n_164),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_160),
.Y(n_164)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_162),
.Y(n_284)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_162),
.Y(n_596)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_166),
.A2(n_255),
.B1(n_256),
.B2(n_263),
.Y(n_254)
);

INVx3_ASAP7_75t_L g619 ( 
.A(n_167),
.Y(n_619)
);

INVx5_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

BUFx12f_ASAP7_75t_L g173 ( 
.A(n_169),
.Y(n_173)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx5_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_SL g263 ( 
.A(n_174),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_235),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_194),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g363 ( 
.A1(n_177),
.A2(n_195),
.B(n_215),
.Y(n_363)
);

AOI22x1_ASAP7_75t_SL g177 ( 
.A1(n_178),
.A2(n_184),
.B1(n_185),
.B2(n_187),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_181),
.A2(n_192),
.B1(n_199),
.B2(n_200),
.Y(n_198)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_181),
.Y(n_446)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_182),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g467 ( 
.A1(n_184),
.A2(n_468),
.B1(n_475),
.B2(n_476),
.Y(n_467)
);

AOI22xp5_ASAP7_75t_L g514 ( 
.A1(n_184),
.A2(n_304),
.B1(n_451),
.B2(n_515),
.Y(n_514)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx6_ASAP7_75t_L g312 ( 
.A(n_186),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_215),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_196),
.B(n_204),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_196),
.A2(n_216),
.B1(n_291),
.B2(n_296),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_SL g379 ( 
.A1(n_196),
.A2(n_216),
.B1(n_380),
.B2(n_381),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g430 ( 
.A1(n_196),
.A2(n_216),
.B1(n_431),
.B2(n_434),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_SL g461 ( 
.A1(n_196),
.A2(n_216),
.B1(n_434),
.B2(n_462),
.Y(n_461)
);

AOI22xp5_ASAP7_75t_L g530 ( 
.A1(n_196),
.A2(n_216),
.B1(n_462),
.B2(n_531),
.Y(n_530)
);

OA21x2_ASAP7_75t_L g581 ( 
.A1(n_196),
.A2(n_216),
.B(n_381),
.Y(n_581)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_197),
.A2(n_228),
.B1(n_238),
.B2(n_239),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_197),
.A2(n_205),
.B1(n_238),
.B2(n_333),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g547 ( 
.A1(n_197),
.A2(n_238),
.B1(n_548),
.B2(n_549),
.Y(n_547)
);

BUFx2_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

AND2x2_ASAP7_75t_SL g216 ( 
.A(n_198),
.B(n_217),
.Y(n_216)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx6_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

HB1xp67_ASAP7_75t_L g224 ( 
.A(n_203),
.Y(n_224)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

BUFx2_ASAP7_75t_L g234 ( 
.A(n_208),
.Y(n_234)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_209),
.Y(n_437)
);

BUFx6f_ASAP7_75t_L g439 ( 
.A(n_209),
.Y(n_439)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx4_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_213),
.Y(n_339)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_214),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_216),
.B(n_227),
.Y(n_215)
);

INVx1_ASAP7_75t_SL g238 ( 
.A(n_216),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_218),
.A2(n_221),
.B1(n_223),
.B2(n_225),
.Y(n_217)
);

BUFx2_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx4_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx6_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g433 ( 
.A(n_226),
.Y(n_433)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

BUFx3_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_SL g233 ( 
.A(n_234),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_253),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g329 ( 
.A(n_236),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_237),
.B(n_248),
.Y(n_236)
);

XOR2x2_ASAP7_75t_L g277 ( 
.A(n_237),
.B(n_248),
.Y(n_277)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_239),
.Y(n_296)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_242),
.Y(n_410)
);

INVx3_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_245),
.Y(n_463)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

BUFx2_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_264),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_254),
.B(n_264),
.C(n_329),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g572 ( 
.A1(n_255),
.A2(n_263),
.B1(n_393),
.B2(n_573),
.Y(n_572)
);

OAI22xp5_ASAP7_75t_SL g615 ( 
.A1(n_255),
.A2(n_263),
.B1(n_616),
.B2(n_617),
.Y(n_615)
);

OAI22xp5_ASAP7_75t_SL g626 ( 
.A1(n_255),
.A2(n_263),
.B1(n_617),
.B2(n_627),
.Y(n_626)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

BUFx6f_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx4_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx6_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx4_ASAP7_75t_L g289 ( 
.A(n_262),
.Y(n_289)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_269),
.Y(n_361)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx3_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

BUFx3_ASAP7_75t_L g362 ( 
.A(n_272),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_277),
.C(n_278),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_274),
.A2(n_275),
.B1(n_324),
.B2(n_325),
.Y(n_323)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_277),
.B(n_279),
.Y(n_324)
);

HB1xp67_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_286),
.C(n_290),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_280),
.B(n_290),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_281),
.A2(n_282),
.B1(n_285),
.B2(n_314),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_281),
.A2(n_285),
.B1(n_373),
.B2(n_374),
.Y(n_372)
);

OAI21xp33_ASAP7_75t_R g613 ( 
.A1(n_281),
.A2(n_285),
.B(n_614),
.Y(n_613)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_286),
.B(n_300),
.Y(n_299)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g549 ( 
.A(n_291),
.Y(n_549)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

BUFx12f_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx4_ASAP7_75t_L g335 ( 
.A(n_295),
.Y(n_335)
);

BUFx6f_ASAP7_75t_L g533 ( 
.A(n_295),
.Y(n_533)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_323),
.Y(n_297)
);

OR2x2_ASAP7_75t_L g561 ( 
.A(n_298),
.B(n_323),
.Y(n_561)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_301),
.C(n_302),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g555 ( 
.A(n_299),
.B(n_556),
.Y(n_555)
);

XNOR2xp5_ASAP7_75t_L g556 ( 
.A(n_301),
.B(n_302),
.Y(n_556)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_313),
.C(n_322),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g543 ( 
.A(n_303),
.B(n_322),
.Y(n_543)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx6_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g542 ( 
.A(n_313),
.B(n_543),
.Y(n_542)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

INVx6_ASAP7_75t_L g528 ( 
.A(n_321),
.Y(n_528)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_324),
.Y(n_325)
);

A2O1A1O1Ixp25_ASAP7_75t_L g559 ( 
.A1(n_326),
.A2(n_367),
.B(n_560),
.C(n_562),
.D(n_563),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_327),
.B(n_366),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g562 ( 
.A(n_327),
.B(n_366),
.Y(n_562)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_330),
.Y(n_327)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_328),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_331),
.A2(n_346),
.B1(n_364),
.B2(n_365),
.Y(n_330)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_331),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_331),
.B(n_365),
.C(n_400),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_332),
.A2(n_340),
.B1(n_341),
.B2(n_345),
.Y(n_331)
);

INVxp67_ASAP7_75t_L g345 ( 
.A(n_332),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_332),
.B(n_341),
.Y(n_388)
);

INVxp67_ASAP7_75t_L g380 ( 
.A(n_333),
.Y(n_380)
);

HB1xp67_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_335),
.Y(n_382)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_340),
.A2(n_341),
.B1(n_391),
.B2(n_392),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_SL g584 ( 
.A1(n_340),
.A2(n_398),
.B1(n_585),
.B2(n_646),
.Y(n_584)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

BUFx3_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_346),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_347),
.B(n_363),
.Y(n_346)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_348),
.B(n_355),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_348),
.B(n_355),
.C(n_363),
.Y(n_369)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_351),
.Y(n_576)
);

INVx1_ASAP7_75t_SL g352 ( 
.A(n_353),
.Y(n_352)
);

INVx3_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

INVxp67_ASAP7_75t_L g373 ( 
.A(n_356),
.Y(n_373)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

INVx3_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_SL g367 ( 
.A(n_368),
.B(n_399),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g563 ( 
.A(n_368),
.B(n_399),
.Y(n_563)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_369),
.B(n_370),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g604 ( 
.A(n_369),
.B(n_605),
.C(n_606),
.Y(n_604)
);

XNOR2xp5_ASAP7_75t_L g370 ( 
.A(n_371),
.B(n_387),
.Y(n_370)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_371),
.Y(n_606)
);

OAI21xp5_ASAP7_75t_SL g371 ( 
.A1(n_372),
.A2(n_379),
.B(n_386),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_372),
.B(n_379),
.Y(n_386)
);

INVxp67_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

BUFx6f_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_386),
.Y(n_583)
);

AOI22xp5_ASAP7_75t_L g608 ( 
.A1(n_386),
.A2(n_570),
.B1(n_583),
.B2(n_609),
.Y(n_608)
);

INVxp67_ASAP7_75t_L g605 ( 
.A(n_387),
.Y(n_605)
);

OAI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_388),
.A2(n_389),
.B1(n_390),
.B2(n_398),
.Y(n_387)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_388),
.Y(n_398)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

HB1xp67_ASAP7_75t_L g585 ( 
.A(n_392),
.Y(n_585)
);

INVx3_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_396),
.Y(n_574)
);

INVx3_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

AOI21x1_ASAP7_75t_L g401 ( 
.A1(n_402),
.A2(n_554),
.B(n_558),
.Y(n_401)
);

OAI21x1_ASAP7_75t_L g402 ( 
.A1(n_403),
.A2(n_539),
.B(n_553),
.Y(n_402)
);

AOI21x1_ASAP7_75t_SL g403 ( 
.A1(n_404),
.A2(n_504),
.B(n_538),
.Y(n_403)
);

OAI21x1_ASAP7_75t_L g404 ( 
.A1(n_405),
.A2(n_465),
.B(n_503),
.Y(n_404)
);

AND2x2_ASAP7_75t_L g405 ( 
.A(n_406),
.B(n_440),
.Y(n_405)
);

OR2x2_ASAP7_75t_L g503 ( 
.A(n_406),
.B(n_440),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_407),
.B(n_429),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_L g477 ( 
.A1(n_407),
.A2(n_429),
.B1(n_430),
.B2(n_478),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_407),
.Y(n_478)
);

OAI32xp33_ASAP7_75t_L g407 ( 
.A1(n_408),
.A2(n_411),
.A3(n_415),
.B1(n_419),
.B2(n_424),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

BUFx3_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

INVx3_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_414),
.Y(n_472)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_416),
.B(n_425),
.Y(n_424)
);

BUFx2_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

HB1xp67_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

INVx5_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_427),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

INVx5_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

BUFx2_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_441),
.B(n_458),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_441),
.B(n_460),
.C(n_464),
.Y(n_505)
);

INVxp67_ASAP7_75t_L g476 ( 
.A(n_442),
.Y(n_476)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_446),
.Y(n_445)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_447),
.Y(n_475)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

BUFx3_ASAP7_75t_L g448 ( 
.A(n_449),
.Y(n_448)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_451),
.Y(n_450)
);

BUFx2_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_455),
.Y(n_454)
);

BUFx2_ASAP7_75t_L g455 ( 
.A(n_456),
.Y(n_455)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_456),
.Y(n_485)
);

BUFx6f_ASAP7_75t_L g456 ( 
.A(n_457),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_L g458 ( 
.A1(n_459),
.A2(n_460),
.B1(n_461),
.B2(n_464),
.Y(n_458)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_459),
.Y(n_464)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_461),
.Y(n_460)
);

AOI21xp5_ASAP7_75t_L g465 ( 
.A1(n_466),
.A2(n_479),
.B(n_502),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_467),
.B(n_477),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_467),
.B(n_477),
.Y(n_502)
);

INVxp67_ASAP7_75t_L g468 ( 
.A(n_469),
.Y(n_468)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_470),
.Y(n_496)
);

BUFx2_ASAP7_75t_L g470 ( 
.A(n_471),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_472),
.Y(n_471)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_474),
.Y(n_473)
);

OAI21xp5_ASAP7_75t_L g479 ( 
.A1(n_480),
.A2(n_498),
.B(n_501),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_481),
.B(n_490),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_482),
.B(n_486),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_483),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_484),
.Y(n_483)
);

HB1xp67_ASAP7_75t_L g484 ( 
.A(n_485),
.Y(n_484)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_488),
.Y(n_487)
);

BUFx3_ASAP7_75t_L g488 ( 
.A(n_489),
.Y(n_488)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_493),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_494),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_495),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_499),
.B(n_500),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_499),
.B(n_500),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_505),
.B(n_506),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_505),
.B(n_506),
.Y(n_538)
);

XOR2xp5_ASAP7_75t_L g506 ( 
.A(n_507),
.B(n_519),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g552 ( 
.A(n_507),
.B(n_520),
.C(n_530),
.Y(n_552)
);

AOI22xp5_ASAP7_75t_L g507 ( 
.A1(n_508),
.A2(n_514),
.B1(n_517),
.B2(n_518),
.Y(n_507)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_508),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_508),
.B(n_518),
.Y(n_546)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_510),
.Y(n_509)
);

INVx3_ASAP7_75t_L g510 ( 
.A(n_511),
.Y(n_510)
);

BUFx6f_ASAP7_75t_L g511 ( 
.A(n_512),
.Y(n_511)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_514),
.Y(n_518)
);

INVx4_ASAP7_75t_L g515 ( 
.A(n_516),
.Y(n_515)
);

OAI22xp5_ASAP7_75t_SL g519 ( 
.A1(n_520),
.A2(n_521),
.B1(n_529),
.B2(n_530),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_521),
.Y(n_520)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_524),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_525),
.Y(n_524)
);

INVx2_ASAP7_75t_SL g525 ( 
.A(n_526),
.Y(n_525)
);

INVx6_ASAP7_75t_L g527 ( 
.A(n_528),
.Y(n_527)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_530),
.Y(n_529)
);

INVxp67_ASAP7_75t_L g548 ( 
.A(n_531),
.Y(n_548)
);

HB1xp67_ASAP7_75t_L g532 ( 
.A(n_533),
.Y(n_532)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_535),
.Y(n_534)
);

INVx3_ASAP7_75t_L g535 ( 
.A(n_536),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_537),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_L g539 ( 
.A(n_540),
.B(n_552),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_540),
.B(n_552),
.Y(n_553)
);

OAI22xp5_ASAP7_75t_SL g540 ( 
.A1(n_541),
.A2(n_542),
.B1(n_544),
.B2(n_545),
.Y(n_540)
);

MAJIxp5_ASAP7_75t_L g557 ( 
.A(n_541),
.B(n_547),
.C(n_550),
.Y(n_557)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_542),
.Y(n_541)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_545),
.Y(n_544)
);

OAI22xp5_ASAP7_75t_SL g545 ( 
.A1(n_546),
.A2(n_547),
.B1(n_550),
.B2(n_551),
.Y(n_545)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_546),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_547),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_SL g554 ( 
.A(n_555),
.B(n_557),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_555),
.B(n_557),
.Y(n_558)
);

NOR3xp33_ASAP7_75t_L g564 ( 
.A(n_565),
.B(n_610),
.C(n_624),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_566),
.B(n_603),
.Y(n_565)
);

INVxp67_ASAP7_75t_SL g566 ( 
.A(n_567),
.Y(n_566)
);

OAI21xp5_ASAP7_75t_L g634 ( 
.A1(n_567),
.A2(n_635),
.B(n_636),
.Y(n_634)
);

NOR2xp67_ASAP7_75t_L g567 ( 
.A(n_568),
.B(n_586),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_568),
.B(n_586),
.Y(n_636)
);

MAJIxp5_ASAP7_75t_L g568 ( 
.A(n_569),
.B(n_583),
.C(n_584),
.Y(n_568)
);

HB1xp67_ASAP7_75t_L g569 ( 
.A(n_570),
.Y(n_569)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_570),
.Y(n_609)
);

AOI22xp5_ASAP7_75t_L g570 ( 
.A1(n_571),
.A2(n_572),
.B1(n_577),
.B2(n_582),
.Y(n_570)
);

MAJIxp5_ASAP7_75t_L g587 ( 
.A(n_571),
.B(n_578),
.C(n_581),
.Y(n_587)
);

OAI22xp5_ASAP7_75t_L g588 ( 
.A1(n_571),
.A2(n_572),
.B1(n_589),
.B2(n_602),
.Y(n_588)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_572),
.Y(n_571)
);

MAJIxp5_ASAP7_75t_L g621 ( 
.A(n_572),
.B(n_622),
.C(n_623),
.Y(n_621)
);

INVxp67_ASAP7_75t_L g600 ( 
.A(n_573),
.Y(n_600)
);

INVx3_ASAP7_75t_L g575 ( 
.A(n_576),
.Y(n_575)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_577),
.Y(n_582)
);

XNOR2xp5_ASAP7_75t_L g577 ( 
.A(n_578),
.B(n_581),
.Y(n_577)
);

OAI22xp5_ASAP7_75t_L g590 ( 
.A1(n_581),
.A2(n_591),
.B1(n_597),
.B2(n_598),
.Y(n_590)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_581),
.Y(n_598)
);

MAJIxp5_ASAP7_75t_L g620 ( 
.A(n_581),
.B(n_597),
.C(n_599),
.Y(n_620)
);

XOR2xp5_ASAP7_75t_L g607 ( 
.A(n_584),
.B(n_608),
.Y(n_607)
);

XNOR2xp5_ASAP7_75t_L g586 ( 
.A(n_587),
.B(n_588),
.Y(n_586)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_587),
.Y(n_623)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_589),
.Y(n_602)
);

HB1xp67_ASAP7_75t_L g622 ( 
.A(n_589),
.Y(n_622)
);

XNOR2x1_ASAP7_75t_L g589 ( 
.A(n_590),
.B(n_599),
.Y(n_589)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_591),
.Y(n_597)
);

INVxp67_ASAP7_75t_L g614 ( 
.A(n_592),
.Y(n_614)
);

BUFx2_ASAP7_75t_L g593 ( 
.A(n_594),
.Y(n_593)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_596),
.Y(n_595)
);

INVxp67_ASAP7_75t_L g616 ( 
.A(n_601),
.Y(n_616)
);

OR2x2_ASAP7_75t_L g603 ( 
.A(n_604),
.B(n_607),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_604),
.B(n_607),
.Y(n_635)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_611),
.Y(n_610)
);

A2O1A1O1Ixp25_ASAP7_75t_L g633 ( 
.A1(n_611),
.A2(n_625),
.B(n_634),
.C(n_637),
.D(n_638),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_612),
.B(n_621),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_612),
.B(n_626),
.Y(n_625)
);

NOR2xp33_ASAP7_75t_L g637 ( 
.A(n_612),
.B(n_621),
.Y(n_637)
);

NOR2xp33_ASAP7_75t_L g638 ( 
.A(n_612),
.B(n_626),
.Y(n_638)
);

FAx1_ASAP7_75t_SL g612 ( 
.A(n_613),
.B(n_615),
.CI(n_620),
.CON(n_612),
.SN(n_612)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_625),
.Y(n_624)
);

OR2x2_ASAP7_75t_L g639 ( 
.A(n_626),
.B(n_640),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_626),
.B(n_640),
.Y(n_644)
);

HB1xp67_ASAP7_75t_L g642 ( 
.A(n_627),
.Y(n_642)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_629),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_630),
.Y(n_629)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_633),
.Y(n_632)
);

CKINVDCx16_ASAP7_75t_R g641 ( 
.A(n_642),
.Y(n_641)
);

CKINVDCx16_ASAP7_75t_R g643 ( 
.A(n_644),
.Y(n_643)
);


endmodule