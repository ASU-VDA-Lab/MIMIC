module fake_jpeg_21315_n_325 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_325);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_325;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_13;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_11;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_145;
wire n_20;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_12;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_7),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g13 ( 
.A(n_9),
.B(n_10),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_1),
.Y(n_14)
);

BUFx10_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_10),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx10_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_24),
.B(n_25),
.Y(n_39)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_22),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_12),
.Y(n_28)
);

OR2x2_ASAP7_75t_L g35 ( 
.A(n_28),
.B(n_32),
.Y(n_35)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_22),
.Y(n_32)
);

BUFx10_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_28),
.A2(n_23),
.B1(n_14),
.B2(n_19),
.Y(n_37)
);

OA22x2_ASAP7_75t_L g51 ( 
.A1(n_37),
.A2(n_35),
.B1(n_29),
.B2(n_30),
.Y(n_51)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_45),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_45),
.Y(n_48)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

INVx13_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_49),
.Y(n_77)
);

OR2x2_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_28),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_50),
.B(n_51),
.Y(n_72)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_52),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_35),
.B(n_13),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_53),
.B(n_57),
.Y(n_66)
);

OAI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_38),
.A2(n_27),
.B1(n_32),
.B2(n_23),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_54),
.A2(n_41),
.B1(n_43),
.B2(n_44),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_35),
.B(n_29),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_55),
.B(n_56),
.Y(n_63)
);

OR2x2_ASAP7_75t_L g56 ( 
.A(n_37),
.B(n_32),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_38),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_58),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_59),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_35),
.B(n_30),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_60),
.B(n_40),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_38),
.B(n_13),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_61),
.B(n_18),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_56),
.B(n_31),
.C(n_39),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_64),
.B(n_78),
.C(n_51),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_68),
.B(n_54),
.Y(n_93)
);

OAI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_56),
.A2(n_40),
.B1(n_41),
.B2(n_27),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_69),
.A2(n_75),
.B1(n_79),
.B2(n_44),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_70),
.B(n_73),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_57),
.A2(n_40),
.B1(n_23),
.B2(n_42),
.Y(n_71)
);

AO21x1_ASAP7_75t_L g90 ( 
.A1(n_71),
.A2(n_26),
.B(n_42),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_60),
.B(n_45),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_61),
.B(n_18),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_74),
.B(n_51),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_56),
.A2(n_39),
.B1(n_43),
.B2(n_41),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_L g78 ( 
.A(n_53),
.B(n_39),
.Y(n_78)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_76),
.Y(n_81)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_81),
.Y(n_128)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_69),
.Y(n_82)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_82),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_66),
.B(n_50),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_83),
.B(n_85),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_66),
.B(n_50),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_73),
.A2(n_50),
.B1(n_51),
.B2(n_55),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_86),
.A2(n_88),
.B1(n_72),
.B2(n_63),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_68),
.B(n_51),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_87),
.B(n_97),
.Y(n_112)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_65),
.Y(n_89)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_89),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g102 ( 
.A1(n_90),
.A2(n_79),
.B(n_43),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_77),
.A2(n_52),
.B1(n_44),
.B2(n_42),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_91),
.A2(n_77),
.B1(n_62),
.B2(n_52),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_65),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_92),
.B(n_96),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_93),
.B(n_80),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_94),
.B(n_64),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_95),
.B(n_33),
.Y(n_124)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_67),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_72),
.B(n_51),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_70),
.B(n_31),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_98),
.B(n_31),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_76),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_99),
.Y(n_103)
);

NOR2x1_ASAP7_75t_L g100 ( 
.A(n_72),
.B(n_26),
.Y(n_100)
);

OAI21x1_ASAP7_75t_L g114 ( 
.A1(n_100),
.A2(n_26),
.B(n_24),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_97),
.A2(n_72),
.B(n_75),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_101),
.A2(n_102),
.B(n_114),
.Y(n_148)
);

BUFx24_ASAP7_75t_SL g104 ( 
.A(n_83),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_104),
.B(n_49),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_107),
.A2(n_110),
.B1(n_116),
.B2(n_34),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_108),
.B(n_25),
.C(n_24),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_82),
.A2(n_64),
.B1(n_63),
.B2(n_71),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_109),
.B(n_115),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_88),
.A2(n_78),
.B1(n_74),
.B2(n_58),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g161 ( 
.A1(n_111),
.A2(n_121),
.B1(n_21),
.B2(n_46),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_87),
.A2(n_18),
.B(n_17),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_113),
.A2(n_17),
.B(n_92),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_86),
.A2(n_58),
.B1(n_80),
.B2(n_67),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_89),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_118),
.B(n_120),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_95),
.A2(n_48),
.B1(n_47),
.B2(n_14),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_119),
.A2(n_129),
.B1(n_76),
.B2(n_46),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_85),
.Y(n_120)
);

OAI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_93),
.A2(n_17),
.B1(n_14),
.B2(n_36),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_91),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_122),
.B(n_124),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_123),
.B(n_125),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_94),
.A2(n_84),
.B1(n_98),
.B2(n_100),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_84),
.B(n_48),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_126),
.B(n_99),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_90),
.A2(n_48),
.B1(n_47),
.B2(n_36),
.Y(n_129)
);

CKINVDCx14_ASAP7_75t_R g170 ( 
.A(n_130),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_106),
.A2(n_90),
.B(n_100),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_131),
.A2(n_148),
.B(n_134),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_132),
.B(n_143),
.Y(n_168)
);

NAND3xp33_ASAP7_75t_L g133 ( 
.A(n_106),
.B(n_36),
.C(n_8),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_133),
.A2(n_134),
.B(n_142),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_115),
.B(n_31),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g135 ( 
.A(n_128),
.Y(n_135)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_135),
.Y(n_174)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_127),
.Y(n_136)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_136),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_110),
.B(n_81),
.Y(n_139)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_139),
.Y(n_182)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_127),
.Y(n_141)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_141),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_105),
.B(n_31),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_120),
.B(n_96),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_118),
.B(n_96),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_144),
.B(n_145),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_117),
.B(n_49),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_126),
.B(n_47),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_146),
.B(n_149),
.Y(n_186)
);

INVxp33_ASAP7_75t_L g147 ( 
.A(n_116),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_147),
.B(n_157),
.Y(n_169)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_117),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_128),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_150),
.B(n_155),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_151),
.B(n_33),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_152),
.A2(n_165),
.B1(n_46),
.B2(n_34),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_108),
.B(n_125),
.C(n_101),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_153),
.B(n_16),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_107),
.B(n_99),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_156),
.Y(n_171)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_128),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_119),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_158),
.A2(n_162),
.B(n_164),
.Y(n_166)
);

OR2x2_ASAP7_75t_L g159 ( 
.A(n_112),
.B(n_26),
.Y(n_159)
);

A2O1A1Ixp33_ASAP7_75t_SL g173 ( 
.A1(n_159),
.A2(n_114),
.B(n_129),
.C(n_124),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_109),
.B(n_59),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_160),
.Y(n_194)
);

OAI21xp33_ASAP7_75t_SL g176 ( 
.A1(n_161),
.A2(n_123),
.B(n_111),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_112),
.B(n_59),
.Y(n_162)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_103),
.Y(n_163)
);

BUFx4f_ASAP7_75t_SL g183 ( 
.A(n_163),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_105),
.B(n_59),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_137),
.A2(n_113),
.B(n_102),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_167),
.A2(n_177),
.B(n_179),
.Y(n_216)
);

AO22x1_ASAP7_75t_L g219 ( 
.A1(n_173),
.A2(n_164),
.B1(n_157),
.B2(n_150),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_176),
.A2(n_187),
.B1(n_188),
.B2(n_142),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_148),
.A2(n_108),
.B(n_21),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_180),
.A2(n_191),
.B1(n_155),
.B2(n_154),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_138),
.A2(n_46),
.B1(n_34),
.B2(n_21),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_181),
.A2(n_136),
.B1(n_141),
.B2(n_134),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_158),
.A2(n_21),
.B1(n_11),
.B2(n_16),
.Y(n_184)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_184),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_131),
.A2(n_21),
.B(n_26),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_140),
.A2(n_21),
.B(n_26),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_189),
.B(n_190),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_153),
.B(n_16),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_165),
.A2(n_152),
.B1(n_138),
.B2(n_154),
.Y(n_191)
);

OAI21xp33_ASAP7_75t_L g192 ( 
.A1(n_140),
.A2(n_10),
.B(n_9),
.Y(n_192)
);

A2O1A1Ixp33_ASAP7_75t_SL g215 ( 
.A1(n_192),
.A2(n_6),
.B(n_9),
.C(n_8),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_195),
.B(n_151),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_178),
.B(n_146),
.Y(n_196)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_196),
.Y(n_231)
);

CKINVDCx14_ASAP7_75t_R g243 ( 
.A(n_197),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_199),
.B(n_191),
.Y(n_222)
);

OR2x2_ASAP7_75t_L g200 ( 
.A(n_169),
.B(n_137),
.Y(n_200)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_200),
.Y(n_234)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_186),
.Y(n_202)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_202),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_203),
.A2(n_173),
.B1(n_172),
.B2(n_183),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_190),
.B(n_195),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_204),
.B(n_219),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_205),
.A2(n_209),
.B1(n_194),
.B2(n_180),
.Y(n_224)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_193),
.Y(n_206)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_206),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_175),
.B(n_143),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_207),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_179),
.B(n_159),
.C(n_162),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_208),
.B(n_210),
.C(n_177),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_171),
.A2(n_144),
.B1(n_149),
.B2(n_142),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_189),
.B(n_159),
.C(n_145),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_185),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_211),
.B(n_212),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_168),
.B(n_130),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_174),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_213),
.B(n_214),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_170),
.B(n_163),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_215),
.A2(n_8),
.B1(n_7),
.B2(n_6),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_182),
.B(n_135),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_217),
.B(n_218),
.Y(n_233)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_183),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_166),
.Y(n_220)
);

AOI21xp33_ASAP7_75t_L g242 ( 
.A1(n_220),
.A2(n_6),
.B(n_5),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_221),
.B(n_205),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_222),
.B(n_226),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_224),
.A2(n_228),
.B1(n_0),
.B2(n_1),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_198),
.B(n_187),
.Y(n_226)
);

XNOR2x1_ASAP7_75t_L g227 ( 
.A(n_216),
.B(n_173),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_227),
.B(n_237),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_203),
.A2(n_194),
.B1(n_171),
.B2(n_173),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_198),
.B(n_181),
.C(n_188),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_229),
.B(n_235),
.C(n_238),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_230),
.B(n_197),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_199),
.B(n_183),
.C(n_192),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_216),
.B(n_204),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_210),
.B(n_219),
.C(n_208),
.Y(n_238)
);

AND2x2_ASAP7_75t_L g246 ( 
.A(n_239),
.B(n_200),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_242),
.A2(n_5),
.B1(n_6),
.B2(n_2),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_244),
.B(n_247),
.Y(n_264)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_233),
.Y(n_245)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_245),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_246),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_223),
.B(n_207),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_232),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_248),
.B(n_250),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_249),
.A2(n_259),
.B1(n_238),
.B2(n_229),
.Y(n_265)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_234),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_231),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_251),
.B(n_253),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_240),
.B(n_196),
.Y(n_253)
);

NAND3xp33_ASAP7_75t_L g254 ( 
.A(n_243),
.B(n_201),
.C(n_215),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g272 ( 
.A1(n_254),
.A2(n_5),
.B(n_1),
.Y(n_272)
);

AO22x1_ASAP7_75t_L g255 ( 
.A1(n_227),
.A2(n_209),
.B1(n_215),
.B2(n_59),
.Y(n_255)
);

AO21x1_ASAP7_75t_L g269 ( 
.A1(n_255),
.A2(n_258),
.B(n_235),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_228),
.B(n_215),
.Y(n_256)
);

BUFx2_ASAP7_75t_L g274 ( 
.A(n_256),
.Y(n_274)
);

NAND2xp33_ASAP7_75t_L g263 ( 
.A(n_257),
.B(n_230),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_225),
.B(n_59),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_241),
.A2(n_11),
.B1(n_5),
.B2(n_20),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_260),
.A2(n_246),
.B1(n_224),
.B2(n_255),
.Y(n_267)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_263),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_265),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_267),
.A2(n_262),
.B1(n_261),
.B2(n_11),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_252),
.B(n_222),
.C(n_221),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_268),
.B(n_271),
.C(n_277),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_269),
.A2(n_270),
.B(n_272),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_259),
.A2(n_236),
.B(n_237),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_252),
.B(n_236),
.C(n_226),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_244),
.B(n_22),
.C(n_15),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_273),
.A2(n_262),
.B(n_254),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_279),
.B(n_280),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_L g281 ( 
.A1(n_269),
.A2(n_261),
.B(n_1),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_281),
.B(n_282),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_264),
.A2(n_266),
.B(n_276),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_274),
.B(n_20),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_283),
.B(n_285),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_274),
.B(n_20),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_268),
.B(n_22),
.C(n_15),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_286),
.B(n_271),
.C(n_277),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_275),
.B(n_15),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_287),
.B(n_289),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_267),
.B(n_22),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_290),
.B(n_0),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_265),
.B(n_24),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_291),
.B(n_24),
.Y(n_299)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_293),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_284),
.B(n_270),
.C(n_272),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_294),
.B(n_295),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_284),
.B(n_24),
.C(n_25),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_288),
.B(n_24),
.C(n_25),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_296),
.B(n_298),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_299),
.A2(n_25),
.B1(n_33),
.B2(n_4),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_288),
.B(n_24),
.C(n_25),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_302),
.B(n_280),
.C(n_281),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_290),
.B(n_0),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g312 ( 
.A(n_303),
.B(n_3),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_304),
.B(n_305),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_300),
.B(n_286),
.C(n_278),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_L g306 ( 
.A1(n_301),
.A2(n_2),
.B(n_3),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_306),
.B(n_307),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_297),
.A2(n_2),
.B(n_3),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_310),
.A2(n_299),
.B(n_4),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_312),
.B(n_292),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_313),
.B(n_315),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_314),
.B(n_311),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_318),
.B(n_308),
.C(n_309),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_319),
.B(n_317),
.Y(n_320)
);

NAND3xp33_ASAP7_75t_L g321 ( 
.A(n_320),
.B(n_316),
.C(n_309),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_321),
.A2(n_25),
.B1(n_33),
.B2(n_3),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_322),
.B(n_25),
.C(n_33),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_323),
.B(n_33),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_324),
.A2(n_4),
.B1(n_33),
.B2(n_41),
.Y(n_325)
);


endmodule