module fake_aes_880_n_48 (n_11, n_1, n_2, n_13, n_12, n_6, n_4, n_3, n_9, n_5, n_14, n_7, n_10, n_8, n_0, n_48);
input n_11;
input n_1;
input n_2;
input n_13;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_14;
input n_7;
input n_10;
input n_8;
input n_0;
output n_48;
wire n_45;
wire n_20;
wire n_38;
wire n_44;
wire n_36;
wire n_47;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_46;
wire n_25;
wire n_16;
wire n_26;
wire n_33;
wire n_30;
wire n_18;
wire n_32;
wire n_41;
wire n_35;
wire n_17;
wire n_15;
wire n_42;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_43;
wire n_40;
wire n_27;
wire n_39;
CKINVDCx16_ASAP7_75t_R g15 ( .A(n_3), .Y(n_15) );
OAI22xp5_ASAP7_75t_L g16 ( .A1(n_1), .A2(n_10), .B1(n_6), .B2(n_14), .Y(n_16) );
CKINVDCx5p33_ASAP7_75t_R g17 ( .A(n_4), .Y(n_17) );
INVx5_ASAP7_75t_L g18 ( .A(n_13), .Y(n_18) );
CKINVDCx5p33_ASAP7_75t_R g19 ( .A(n_7), .Y(n_19) );
CKINVDCx5p33_ASAP7_75t_R g20 ( .A(n_2), .Y(n_20) );
BUFx2_ASAP7_75t_L g21 ( .A(n_1), .Y(n_21) );
INVx2_ASAP7_75t_L g22 ( .A(n_12), .Y(n_22) );
INVx1_ASAP7_75t_L g23 ( .A(n_0), .Y(n_23) );
AND3x1_ASAP7_75t_L g24 ( .A(n_23), .B(n_0), .C(n_2), .Y(n_24) );
CKINVDCx5p33_ASAP7_75t_R g25 ( .A(n_15), .Y(n_25) );
INVx3_ASAP7_75t_L g26 ( .A(n_22), .Y(n_26) );
NAND2xp5_ASAP7_75t_L g27 ( .A(n_21), .B(n_3), .Y(n_27) );
INVx1_ASAP7_75t_L g28 ( .A(n_22), .Y(n_28) );
AOI22xp33_ASAP7_75t_SL g29 ( .A1(n_27), .A2(n_16), .B1(n_20), .B2(n_17), .Y(n_29) );
INVx2_ASAP7_75t_L g30 ( .A(n_26), .Y(n_30) );
INVx3_ASAP7_75t_SL g31 ( .A(n_25), .Y(n_31) );
AND2x2_ASAP7_75t_L g32 ( .A(n_31), .B(n_27), .Y(n_32) );
AND2x2_ASAP7_75t_L g33 ( .A(n_29), .B(n_24), .Y(n_33) );
AND2x2_ASAP7_75t_L g34 ( .A(n_32), .B(n_29), .Y(n_34) );
NAND2xp5_ASAP7_75t_L g35 ( .A(n_33), .B(n_30), .Y(n_35) );
AOI22xp33_ASAP7_75t_SL g36 ( .A1(n_34), .A2(n_24), .B1(n_26), .B2(n_28), .Y(n_36) );
NOR2x1_ASAP7_75t_SL g37 ( .A(n_35), .B(n_28), .Y(n_37) );
NAND2xp5_ASAP7_75t_L g38 ( .A(n_34), .B(n_26), .Y(n_38) );
INVx1_ASAP7_75t_L g39 ( .A(n_38), .Y(n_39) );
AOI22xp5_ASAP7_75t_L g40 ( .A1(n_36), .A2(n_26), .B1(n_19), .B2(n_18), .Y(n_40) );
OAI221xp5_ASAP7_75t_L g41 ( .A1(n_37), .A2(n_18), .B1(n_4), .B2(n_8), .C(n_9), .Y(n_41) );
INVx1_ASAP7_75t_L g42 ( .A(n_39), .Y(n_42) );
INVx1_ASAP7_75t_L g43 ( .A(n_41), .Y(n_43) );
AND2x2_ASAP7_75t_L g44 ( .A(n_40), .B(n_18), .Y(n_44) );
OR2x2_ASAP7_75t_L g45 ( .A(n_42), .B(n_18), .Y(n_45) );
INVx1_ASAP7_75t_L g46 ( .A(n_43), .Y(n_46) );
AOI22xp5_ASAP7_75t_L g47 ( .A1(n_46), .A2(n_44), .B1(n_5), .B2(n_11), .Y(n_47) );
NAND2xp5_ASAP7_75t_L g48 ( .A(n_47), .B(n_45), .Y(n_48) );
endmodule