module fake_jpeg_15604_n_140 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_140);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_140;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_138;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx1_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_0),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_9),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

AND2x2_ASAP7_75t_L g16 ( 
.A(n_11),
.B(n_9),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_4),
.B(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_7),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_21),
.B(n_0),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_26),
.B(n_28),
.Y(n_33)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_29),
.B(n_32),
.Y(n_37)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

BUFx4f_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_21),
.B(n_1),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_31),
.Y(n_34)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_26),
.B(n_21),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_36),
.B(n_40),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_26),
.B(n_22),
.Y(n_40)
);

OA22x2_ASAP7_75t_SL g41 ( 
.A1(n_32),
.A2(n_16),
.B1(n_20),
.B2(n_19),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_41),
.B(n_32),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_22),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_45),
.B(n_53),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

HB1xp67_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

INVx13_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_49),
.B(n_51),
.Y(n_77)
);

AND2x4_ASAP7_75t_L g50 ( 
.A(n_38),
.B(n_29),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_SL g67 ( 
.A1(n_50),
.A2(n_28),
.B(n_25),
.Y(n_67)
);

INVx13_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_52),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_33),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_54),
.B(n_56),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_55),
.A2(n_58),
.B1(n_16),
.B2(n_27),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_37),
.A2(n_27),
.B1(n_29),
.B2(n_25),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_37),
.B(n_13),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_57),
.B(n_14),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_42),
.A2(n_25),
.B1(n_29),
.B2(n_27),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_41),
.B(n_30),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_59),
.B(n_41),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_61),
.A2(n_17),
.B1(n_12),
.B2(n_23),
.Y(n_88)
);

INVx2_ASAP7_75t_SL g65 ( 
.A(n_46),
.Y(n_65)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_65),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_66),
.B(n_71),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_67),
.A2(n_46),
.B(n_43),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_69),
.B(n_70),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_59),
.B(n_41),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_55),
.B(n_30),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_55),
.B(n_30),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_73),
.B(n_74),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_44),
.B(n_28),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_48),
.Y(n_75)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_75),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_56),
.B(n_12),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_76),
.B(n_16),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_64),
.A2(n_50),
.B1(n_35),
.B2(n_52),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_78),
.A2(n_79),
.B1(n_75),
.B2(n_72),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_69),
.A2(n_50),
.B1(n_35),
.B2(n_51),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_L g81 ( 
.A(n_70),
.B(n_50),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_81),
.B(n_83),
.C(n_90),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_61),
.A2(n_67),
.B1(n_76),
.B2(n_71),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_82),
.A2(n_84),
.B(n_60),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g83 ( 
.A(n_73),
.B(n_16),
.Y(n_83)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_63),
.Y(n_86)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_86),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_87),
.B(n_74),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_88),
.B(n_77),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g90 ( 
.A(n_62),
.B(n_30),
.Y(n_90)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_63),
.Y(n_93)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_93),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_94),
.A2(n_103),
.B(n_85),
.Y(n_108)
);

OAI22x1_ASAP7_75t_L g95 ( 
.A1(n_84),
.A2(n_47),
.B1(n_53),
.B2(n_68),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_95),
.A2(n_99),
.B1(n_101),
.B2(n_104),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_97),
.A2(n_105),
.B1(n_91),
.B2(n_89),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_92),
.A2(n_72),
.B1(n_49),
.B2(n_43),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_81),
.B(n_60),
.C(n_46),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_102),
.B(n_31),
.C(n_17),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_82),
.A2(n_65),
.B1(n_47),
.B2(n_23),
.Y(n_104)
);

AOI22x1_ASAP7_75t_L g105 ( 
.A1(n_78),
.A2(n_53),
.B1(n_65),
.B2(n_31),
.Y(n_105)
);

OAI21xp33_ASAP7_75t_SL g119 ( 
.A1(n_106),
.A2(n_114),
.B(n_24),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_108),
.A2(n_110),
.B(n_98),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_96),
.B(n_90),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_109),
.B(n_113),
.C(n_13),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_103),
.A2(n_80),
.B(n_79),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_105),
.A2(n_95),
.B1(n_101),
.B2(n_99),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_111),
.A2(n_112),
.B1(n_24),
.B2(n_20),
.Y(n_118)
);

A2O1A1O1Ixp25_ASAP7_75t_L g112 ( 
.A1(n_96),
.A2(n_83),
.B(n_88),
.C(n_31),
.D(n_23),
.Y(n_112)
);

NAND2xp33_ASAP7_75t_SL g114 ( 
.A(n_104),
.B(n_102),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_106),
.B(n_100),
.Y(n_115)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_115),
.Y(n_123)
);

CKINVDCx14_ASAP7_75t_R g116 ( 
.A(n_107),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_116),
.B(n_120),
.Y(n_127)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_117),
.Y(n_124)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_118),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_119),
.B(n_121),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_109),
.B(n_19),
.C(n_14),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_121),
.B(n_113),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_125),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_124),
.A2(n_119),
.B(n_114),
.Y(n_128)
);

AOI322xp5_ASAP7_75t_L g134 ( 
.A1(n_128),
.A2(n_131),
.A3(n_1),
.B1(n_2),
.B2(n_3),
.C1(n_4),
.C2(n_5),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_123),
.B(n_10),
.Y(n_130)
);

BUFx24_ASAP7_75t_SL g133 ( 
.A(n_130),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_126),
.A2(n_122),
.B1(n_127),
.B2(n_112),
.Y(n_131)
);

OR2x2_ASAP7_75t_L g132 ( 
.A(n_125),
.B(n_1),
.Y(n_132)
);

AOI311xp33_ASAP7_75t_L g136 ( 
.A1(n_132),
.A2(n_3),
.A3(n_6),
.B(n_8),
.C(n_22),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_134),
.Y(n_138)
);

AOI322xp5_ASAP7_75t_L g135 ( 
.A1(n_129),
.A2(n_2),
.A3(n_3),
.B1(n_4),
.B2(n_5),
.C1(n_6),
.C2(n_7),
.Y(n_135)
);

HB1xp67_ASAP7_75t_L g137 ( 
.A(n_135),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_138),
.A2(n_136),
.B(n_133),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_139),
.B(n_137),
.Y(n_140)
);


endmodule