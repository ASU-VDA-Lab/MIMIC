module fake_jpeg_11010_n_174 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_174);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_174;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g46 ( 
.A(n_21),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_42),
.Y(n_47)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_20),
.Y(n_49)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

BUFx4f_ASAP7_75t_SL g51 ( 
.A(n_34),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_27),
.Y(n_53)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_5),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_29),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_30),
.Y(n_58)
);

BUFx12_ASAP7_75t_L g59 ( 
.A(n_0),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_32),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_13),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_2),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_39),
.B(n_26),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

BUFx10_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_8),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_1),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_19),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_24),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_43),
.Y(n_70)
);

INVx11_ASAP7_75t_L g71 ( 
.A(n_28),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_4),
.Y(n_72)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_61),
.Y(n_73)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_73),
.Y(n_88)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_62),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_74),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_56),
.B(n_0),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_75),
.B(n_67),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_63),
.B(n_61),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_76),
.B(n_77),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_71),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_78),
.Y(n_97)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_46),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_79),
.Y(n_95)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_65),
.Y(n_80)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_80),
.Y(n_86)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_66),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_81),
.B(n_70),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_51),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g92 ( 
.A(n_82),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_75),
.B(n_67),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_85),
.B(n_68),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_87),
.B(n_90),
.Y(n_114)
);

NOR2x1_ASAP7_75t_L g89 ( 
.A(n_76),
.B(n_72),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_89),
.B(n_93),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_78),
.Y(n_90)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_91),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_82),
.B(n_47),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_75),
.B(n_47),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_94),
.B(n_96),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_75),
.B(n_49),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_97),
.Y(n_98)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_98),
.Y(n_122)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_97),
.Y(n_99)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_99),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g100 ( 
.A(n_83),
.B(n_89),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_SL g140 ( 
.A(n_100),
.B(n_111),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_95),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_103),
.B(n_104),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_95),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_88),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_105),
.B(n_106),
.Y(n_130)
);

OAI32xp33_ASAP7_75t_L g106 ( 
.A1(n_84),
.A2(n_65),
.A3(n_57),
.B1(n_64),
.B2(n_59),
.Y(n_106)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_92),
.Y(n_107)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_107),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_109),
.B(n_115),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_84),
.B(n_68),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_110),
.B(n_112),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_86),
.B(n_49),
.C(n_50),
.Y(n_111)
);

AO22x1_ASAP7_75t_L g112 ( 
.A1(n_92),
.A2(n_59),
.B1(n_60),
.B2(n_69),
.Y(n_112)
);

HB1xp67_ASAP7_75t_L g113 ( 
.A(n_92),
.Y(n_113)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_113),
.Y(n_136)
);

AND2x6_ASAP7_75t_L g115 ( 
.A(n_83),
.B(n_25),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_97),
.A2(n_55),
.B1(n_52),
.B2(n_53),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_116),
.A2(n_6),
.B(n_7),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_83),
.B(n_58),
.C(n_54),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_117),
.B(n_11),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_83),
.A2(n_1),
.B(n_2),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_118),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_85),
.B(n_3),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_119),
.B(n_3),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_113),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_120),
.B(n_126),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_101),
.A2(n_48),
.B1(n_4),
.B2(n_5),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_124),
.A2(n_133),
.B1(n_132),
.B2(n_137),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_127),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_105),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_128),
.B(n_139),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_114),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_129),
.A2(n_130),
.B1(n_131),
.B2(n_138),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_101),
.B(n_9),
.Y(n_132)
);

OAI21xp33_ASAP7_75t_L g148 ( 
.A1(n_132),
.A2(n_133),
.B(n_134),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_102),
.B(n_9),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_102),
.B(n_10),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_138),
.B(n_141),
.Y(n_147)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_108),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_110),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_125),
.B(n_12),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_142),
.B(n_151),
.Y(n_159)
);

INVx13_ASAP7_75t_L g143 ( 
.A(n_121),
.Y(n_143)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_143),
.Y(n_158)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_136),
.Y(n_145)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_145),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_146),
.A2(n_154),
.B(n_156),
.Y(n_161)
);

NOR3xp33_ASAP7_75t_L g162 ( 
.A(n_150),
.B(n_153),
.C(n_155),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_140),
.B(n_15),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_130),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_134),
.Y(n_154)
);

AO21x2_ASAP7_75t_L g155 ( 
.A1(n_123),
.A2(n_22),
.B(n_23),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_135),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_152),
.A2(n_122),
.B(n_33),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_157),
.A2(n_163),
.B(n_147),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_151),
.A2(n_31),
.B(n_36),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_164),
.B(n_165),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_161),
.B(n_149),
.C(n_142),
.Y(n_165)
);

XNOR2x1_ASAP7_75t_SL g166 ( 
.A(n_159),
.B(n_148),
.Y(n_166)
);

AOI321xp33_ASAP7_75t_L g167 ( 
.A1(n_166),
.A2(n_158),
.A3(n_144),
.B1(n_162),
.B2(n_160),
.C(n_155),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_167),
.B(n_155),
.C(n_162),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_169),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_170),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_171),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_172),
.B(n_168),
.Y(n_173)
);

XNOR2x2_ASAP7_75t_SL g174 ( 
.A(n_173),
.B(n_37),
.Y(n_174)
);


endmodule