module real_jpeg_14330_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_357, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_357;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_216;
wire n_202;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_0),
.Y(n_54)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

BUFx4f_ASAP7_75t_L g52 ( 
.A(n_2),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_3),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_3),
.B(n_31),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_3),
.B(n_68),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_3),
.B(n_52),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_3),
.B(n_63),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_3),
.B(n_46),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_4),
.B(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_4),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_4),
.B(n_63),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_4),
.B(n_68),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_4),
.B(n_31),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_4),
.B(n_27),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_4),
.B(n_54),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_5),
.B(n_35),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_5),
.B(n_52),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_5),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_5),
.B(n_54),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_5),
.B(n_63),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_5),
.B(n_31),
.Y(n_287)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_7),
.B(n_63),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_7),
.B(n_46),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_7),
.B(n_27),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_7),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_7),
.B(n_31),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_8),
.B(n_27),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_8),
.B(n_52),
.Y(n_81)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_8),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_8),
.B(n_46),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_8),
.B(n_68),
.Y(n_304)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_9),
.Y(n_47)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_10),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_11),
.B(n_27),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_11),
.B(n_63),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_11),
.B(n_68),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_11),
.B(n_52),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_11),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_11),
.B(n_46),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_11),
.B(n_31),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_11),
.B(n_35),
.Y(n_302)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_13),
.B(n_31),
.Y(n_30)
);

AND2x2_ASAP7_75t_SL g53 ( 
.A(n_13),
.B(n_54),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_13),
.B(n_68),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_13),
.B(n_46),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_13),
.B(n_52),
.Y(n_103)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_13),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_13),
.B(n_27),
.Y(n_141)
);

AND2x2_ASAP7_75t_SL g288 ( 
.A(n_13),
.B(n_63),
.Y(n_288)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_14),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_15),
.B(n_27),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_15),
.B(n_63),
.Y(n_73)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_15),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_15),
.B(n_31),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_15),
.B(n_54),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_15),
.B(n_68),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_148),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_147),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_121),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_20),
.B(n_121),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_83),
.C(n_107),
.Y(n_20)
);

XOR2xp5_ASAP7_75t_L g346 ( 
.A(n_21),
.B(n_347),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_65),
.C(n_77),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_22),
.A2(n_23),
.B1(n_341),
.B2(n_342),
.Y(n_340)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_40),
.B2(n_41),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_24),
.B(n_42),
.C(n_59),
.Y(n_109)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

XOR2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_29),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_26),
.B(n_30),
.C(n_33),
.Y(n_106)
);

INVx5_ASAP7_75t_SL g174 ( 
.A(n_27),
.Y(n_174)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g29 ( 
.A1(n_30),
.A2(n_32),
.B1(n_33),
.B2(n_39),
.Y(n_29)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_38),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_34),
.B(n_118),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_34),
.B(n_50),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_34),
.B(n_205),
.Y(n_276)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx13_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_38),
.B(n_164),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_38),
.B(n_174),
.Y(n_226)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_42),
.A2(n_43),
.B1(n_58),
.B2(n_59),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_45),
.B1(n_48),
.B2(n_57),
.Y(n_43)
);

CKINVDCx16_ASAP7_75t_R g44 ( 
.A(n_45),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_45),
.B(n_53),
.C(n_55),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_46),
.Y(n_90)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_48),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_49),
.A2(n_53),
.B1(n_55),
.B2(n_56),
.Y(n_48)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_49),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_49),
.A2(n_55),
.B1(n_141),
.B2(n_142),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_50),
.B(n_51),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_51),
.B(n_205),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_51),
.B(n_91),
.Y(n_294)
);

INVx13_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_53),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_53),
.B(n_67),
.C(n_71),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_53),
.A2(n_56),
.B1(n_67),
.B2(n_80),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_53),
.A2(n_56),
.B1(n_166),
.B2(n_167),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_53),
.B(n_166),
.Y(n_182)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_54),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_55),
.B(n_141),
.C(n_276),
.Y(n_297)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_61),
.C(n_62),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_60),
.A2(n_62),
.B1(n_138),
.B2(n_316),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_60),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_61),
.B(n_315),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_62),
.A2(n_138),
.B1(n_139),
.B2(n_140),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_62),
.Y(n_138)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_64),
.B(n_93),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g342 ( 
.A(n_65),
.B(n_77),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_72),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_66),
.B(n_73),
.C(n_75),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_67),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_67),
.A2(n_80),
.B1(n_233),
.B2(n_234),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_67),
.B(n_233),
.Y(n_265)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_69),
.B(n_162),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_69),
.B(n_205),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

XOR2xp5_ASAP7_75t_L g78 ( 
.A(n_71),
.B(n_79),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_73),
.A2(n_74),
.B1(n_75),
.B2(n_76),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_73),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_74),
.A2(n_75),
.B1(n_102),
.B2(n_103),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_74),
.A2(n_75),
.B1(n_116),
.B2(n_117),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_74),
.B(n_117),
.C(n_119),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_74),
.B(n_99),
.C(n_103),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_74),
.A2(n_75),
.B1(n_186),
.B2(n_187),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_75),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_75),
.B(n_186),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_81),
.C(n_82),
.Y(n_77)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_78),
.B(n_325),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_L g325 ( 
.A1(n_81),
.A2(n_82),
.B1(n_326),
.B2(n_327),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_81),
.Y(n_327)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_82),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_83),
.B(n_107),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_85),
.B1(n_95),
.B2(n_96),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_84),
.B(n_97),
.C(n_106),
.Y(n_123)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_87),
.B1(n_88),
.B2(n_94),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_86),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_86),
.B(n_89),
.C(n_92),
.Y(n_144)
);

CKINVDCx14_ASAP7_75t_R g87 ( 
.A(n_88),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_92),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_91),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_90),
.B(n_162),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_93),
.B(n_164),
.Y(n_272)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_97),
.A2(n_98),
.B1(n_105),
.B2(n_106),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_99),
.A2(n_100),
.B1(n_101),
.B2(n_104),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_99),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_99),
.A2(n_104),
.B1(n_285),
.B2(n_286),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_99),
.B(n_288),
.C(n_289),
.Y(n_318)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_102),
.A2(n_103),
.B1(n_141),
.B2(n_142),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_102),
.A2(n_103),
.B1(n_228),
.B2(n_229),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_103),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_103),
.B(n_226),
.C(n_228),
.Y(n_266)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_109),
.B1(n_110),
.B2(n_111),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_108),
.B(n_112),
.C(n_120),
.Y(n_146)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_120),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_113),
.A2(n_114),
.B1(n_115),
.B2(n_119),
.Y(n_112)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_113),
.Y(n_119)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_146),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_124),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_136),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_126),
.A2(n_127),
.B1(n_128),
.B2(n_129),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_130),
.A2(n_131),
.B1(n_132),
.B2(n_135),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_131),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_132),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_SL g132 ( 
.A(n_133),
.B(n_134),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_SL g136 ( 
.A(n_137),
.B(n_143),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_141),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_145),
.Y(n_143)
);

AOI321xp33_ASAP7_75t_L g148 ( 
.A1(n_149),
.A2(n_334),
.A3(n_344),
.B1(n_348),
.B2(n_353),
.C(n_357),
.Y(n_148)
);

NOR3xp33_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_279),
.C(n_329),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_250),
.B(n_278),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_152),
.A2(n_220),
.B(n_249),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_153),
.A2(n_189),
.B(n_219),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_168),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_154),
.B(n_168),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_159),
.C(n_165),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_155),
.A2(n_171),
.B1(n_172),
.B2(n_180),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_155),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_155),
.B(n_216),
.Y(n_215)
);

FAx1_ASAP7_75t_SL g155 ( 
.A(n_156),
.B(n_157),
.CI(n_158),
.CON(n_155),
.SN(n_155)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_159),
.A2(n_160),
.B1(n_165),
.B2(n_217),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_160),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_163),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_SL g198 ( 
.A(n_161),
.B(n_163),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_162),
.B(n_174),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_164),
.B(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_165),
.Y(n_217)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_169),
.A2(n_170),
.B1(n_181),
.B2(n_188),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_171),
.B(n_180),
.C(n_188),
.Y(n_221)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_172),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_175),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_173),
.B(n_176),
.C(n_179),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_176),
.A2(n_177),
.B1(n_178),
.B2(n_179),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_178),
.Y(n_179)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_181),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_SL g181 ( 
.A(n_182),
.B(n_183),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_182),
.B(n_184),
.C(n_185),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_185),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_186),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_186),
.A2(n_187),
.B1(n_304),
.B2(n_305),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_186),
.B(n_302),
.C(n_305),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_190),
.A2(n_213),
.B(n_218),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_191),
.A2(n_202),
.B(n_212),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_197),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_192),
.B(n_197),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_193),
.B(n_195),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_193),
.A2(n_194),
.B1(n_195),
.B2(n_196),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_194),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_196),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_199),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_198),
.B(n_200),
.C(n_201),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_201),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_203),
.A2(n_207),
.B(n_211),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_206),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_204),
.B(n_206),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_208),
.B(n_210),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_215),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_214),
.B(n_215),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_222),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_221),
.B(n_222),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_223),
.A2(n_224),
.B1(n_235),
.B2(n_236),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_223),
.B(n_237),
.C(n_248),
.Y(n_251)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_230),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_225),
.B(n_231),
.C(n_232),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_SL g225 ( 
.A(n_226),
.B(n_227),
.Y(n_225)
);

CKINVDCx14_ASAP7_75t_R g228 ( 
.A(n_229),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_232),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_237),
.A2(n_238),
.B1(n_247),
.B2(n_248),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_239),
.A2(n_240),
.B1(n_241),
.B2(n_246),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_239),
.B(n_243),
.C(n_245),
.Y(n_269)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_241),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_242),
.A2(n_243),
.B1(n_244),
.B2(n_245),
.Y(n_241)
);

CKINVDCx14_ASAP7_75t_R g245 ( 
.A(n_242),
.Y(n_245)
);

CKINVDCx14_ASAP7_75t_R g243 ( 
.A(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_252),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g278 ( 
.A(n_251),
.B(n_252),
.Y(n_278)
);

AOI22xp33_ASAP7_75t_SL g252 ( 
.A1(n_253),
.A2(n_254),
.B1(n_268),
.B2(n_277),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_255),
.A2(n_256),
.B1(n_257),
.B2(n_267),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_255),
.B(n_267),
.C(n_277),
.Y(n_330)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_257),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_258),
.A2(n_259),
.B1(n_263),
.B2(n_264),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_258),
.B(n_265),
.C(n_266),
.Y(n_298)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

BUFx24_ASAP7_75t_SL g354 ( 
.A(n_259),
.Y(n_354)
);

FAx1_ASAP7_75t_SL g259 ( 
.A(n_260),
.B(n_261),
.CI(n_262),
.CON(n_259),
.SN(n_259)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_260),
.B(n_261),
.C(n_262),
.Y(n_307)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_SL g264 ( 
.A(n_265),
.B(n_266),
.Y(n_264)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_268),
.Y(n_277)
);

BUFx24_ASAP7_75t_SL g356 ( 
.A(n_268),
.Y(n_356)
);

FAx1_ASAP7_75t_SL g268 ( 
.A(n_269),
.B(n_270),
.CI(n_274),
.CON(n_268),
.SN(n_268)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_269),
.B(n_270),
.C(n_274),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_271),
.A2(n_272),
.B(n_273),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_271),
.B(n_272),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_273),
.A2(n_307),
.B1(n_308),
.B2(n_309),
.Y(n_306)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_273),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_SL g274 ( 
.A(n_275),
.B(n_276),
.Y(n_274)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

AOI21xp33_ASAP7_75t_L g349 ( 
.A1(n_280),
.A2(n_350),
.B(n_351),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_311),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_281),
.B(n_311),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_299),
.C(n_310),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_282),
.B(n_332),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_SL g282 ( 
.A(n_283),
.B(n_298),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_291),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_284),
.B(n_291),
.C(n_298),
.Y(n_328)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_287),
.A2(n_288),
.B1(n_289),
.B2(n_290),
.Y(n_286)
);

CKINVDCx16_ASAP7_75t_R g289 ( 
.A(n_287),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_288),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_297),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_293),
.A2(n_294),
.B1(n_295),
.B2(n_296),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_294),
.B(n_295),
.C(n_297),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_296),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g332 ( 
.A1(n_299),
.A2(n_300),
.B1(n_310),
.B2(n_333),
.Y(n_332)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_SL g300 ( 
.A(n_301),
.B(n_306),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_301),
.B(n_307),
.C(n_309),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_SL g301 ( 
.A(n_302),
.B(n_303),
.Y(n_301)
);

CKINVDCx14_ASAP7_75t_R g305 ( 
.A(n_304),
.Y(n_305)
);

CKINVDCx14_ASAP7_75t_R g308 ( 
.A(n_307),
.Y(n_308)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_310),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_328),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_320),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_313),
.B(n_320),
.C(n_328),
.Y(n_336)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_317),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_314),
.B(n_318),
.C(n_319),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_319),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_SL g320 ( 
.A(n_321),
.B(n_322),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_321),
.B(n_323),
.C(n_324),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_324),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_331),
.Y(n_329)
);

AND2x2_ASAP7_75t_L g350 ( 
.A(n_330),
.B(n_331),
.Y(n_350)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_SL g348 ( 
.A1(n_335),
.A2(n_349),
.B(n_352),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_336),
.B(n_337),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_336),
.B(n_337),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_343),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_339),
.B(n_340),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_339),
.B(n_340),
.C(n_343),
.Y(n_345)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_345),
.B(n_346),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_345),
.B(n_346),
.Y(n_353)
);


endmodule