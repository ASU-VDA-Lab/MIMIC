module real_aes_2221_n_105 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_104, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_105);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_104;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_105;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_485;
wire n_822;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_357;
wire n_287;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_571;
wire n_376;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_556;
wire n_341;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_504;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_505;
wire n_527;
wire n_434;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_617;
wire n_552;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_146;
wire n_807;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_831;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_575;
wire n_210;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_639;
wire n_587;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_601;
wire n_307;
wire n_661;
wire n_463;
wire n_804;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_237;
wire n_797;
wire n_668;
NAND2xp5_ASAP7_75t_L g534 ( .A(n_0), .B(n_231), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g116 ( .A(n_1), .B(n_117), .Y(n_116) );
INVx1_ASAP7_75t_L g165 ( .A(n_2), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_3), .B(n_537), .Y(n_556) );
NAND2xp33_ASAP7_75t_SL g527 ( .A(n_4), .B(n_186), .Y(n_527) );
NAND2xp5_ASAP7_75t_SL g222 ( .A(n_5), .B(n_199), .Y(n_222) );
INVx1_ASAP7_75t_L g519 ( .A(n_6), .Y(n_519) );
INVx1_ASAP7_75t_L g256 ( .A(n_7), .Y(n_256) );
CKINVDCx16_ASAP7_75t_R g117 ( .A(n_8), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g273 ( .A(n_9), .Y(n_273) );
AND2x2_ASAP7_75t_L g554 ( .A(n_10), .B(n_155), .Y(n_554) );
INVx2_ASAP7_75t_L g156 ( .A(n_11), .Y(n_156) );
AND3x1_ASAP7_75t_L g114 ( .A(n_12), .B(n_34), .C(n_115), .Y(n_114) );
CKINVDCx16_ASAP7_75t_R g128 ( .A(n_12), .Y(n_128) );
INVx1_ASAP7_75t_L g232 ( .A(n_13), .Y(n_232) );
AOI221x1_ASAP7_75t_L g522 ( .A1(n_14), .A2(n_188), .B1(n_523), .B2(n_525), .C(n_526), .Y(n_522) );
OAI22xp5_ASAP7_75t_SL g808 ( .A1(n_14), .A2(n_59), .B1(n_809), .B2(n_810), .Y(n_808) );
INVxp67_ASAP7_75t_L g810 ( .A(n_14), .Y(n_810) );
NAND2xp5_ASAP7_75t_SL g590 ( .A(n_15), .B(n_537), .Y(n_590) );
NOR2xp33_ASAP7_75t_SL g111 ( .A(n_16), .B(n_112), .Y(n_111) );
INVx1_ASAP7_75t_L g131 ( .A(n_16), .Y(n_131) );
INVx1_ASAP7_75t_L g229 ( .A(n_17), .Y(n_229) );
INVx1_ASAP7_75t_SL g177 ( .A(n_18), .Y(n_177) );
NAND2xp5_ASAP7_75t_SL g202 ( .A(n_19), .B(n_180), .Y(n_202) );
AOI33xp33_ASAP7_75t_L g247 ( .A1(n_20), .A2(n_49), .A3(n_162), .B1(n_173), .B2(n_248), .B3(n_249), .Y(n_247) );
AOI21xp5_ASAP7_75t_L g557 ( .A1(n_21), .A2(n_525), .B(n_558), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_22), .B(n_231), .Y(n_559) );
AOI221xp5_ASAP7_75t_SL g599 ( .A1(n_23), .A2(n_39), .B1(n_525), .B2(n_537), .C(n_600), .Y(n_599) );
INVx1_ASAP7_75t_L g266 ( .A(n_24), .Y(n_266) );
OR2x2_ASAP7_75t_L g157 ( .A(n_25), .B(n_93), .Y(n_157) );
OA21x2_ASAP7_75t_L g190 ( .A1(n_25), .A2(n_93), .B(n_156), .Y(n_190) );
INVxp67_ASAP7_75t_L g521 ( .A(n_26), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_27), .B(n_234), .Y(n_594) );
AND2x2_ASAP7_75t_L g548 ( .A(n_28), .B(n_154), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_29), .B(n_160), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g125 ( .A(n_30), .B(n_126), .Y(n_125) );
AOI21xp5_ASAP7_75t_L g532 ( .A1(n_31), .A2(n_525), .B(n_533), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_32), .B(n_234), .Y(n_601) );
AND2x2_ASAP7_75t_L g167 ( .A(n_33), .B(n_168), .Y(n_167) );
INVx1_ASAP7_75t_L g172 ( .A(n_33), .Y(n_172) );
AND2x2_ASAP7_75t_L g186 ( .A(n_33), .B(n_165), .Y(n_186) );
OR2x6_ASAP7_75t_L g129 ( .A(n_34), .B(n_130), .Y(n_129) );
CKINVDCx20_ASAP7_75t_R g268 ( .A(n_35), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_36), .B(n_160), .Y(n_293) );
AOI22xp5_ASAP7_75t_L g194 ( .A1(n_37), .A2(n_189), .B1(n_195), .B2(n_199), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_38), .B(n_204), .Y(n_203) );
AOI22xp5_ASAP7_75t_L g566 ( .A1(n_40), .A2(n_85), .B1(n_170), .B2(n_525), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_41), .B(n_180), .Y(n_179) );
AOI22xp33_ASAP7_75t_L g105 ( .A1(n_42), .A2(n_106), .B1(n_118), .B2(n_831), .Y(n_105) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_43), .B(n_231), .Y(n_546) );
NAND2xp5_ASAP7_75t_SL g258 ( .A(n_44), .B(n_206), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_45), .B(n_180), .Y(n_257) );
CKINVDCx5p33_ASAP7_75t_R g198 ( .A(n_46), .Y(n_198) );
AND2x2_ASAP7_75t_L g538 ( .A(n_47), .B(n_154), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_48), .B(n_154), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_50), .B(n_180), .Y(n_297) );
CKINVDCx20_ASAP7_75t_R g445 ( .A(n_51), .Y(n_445) );
OAI22xp5_ASAP7_75t_L g820 ( .A1(n_51), .A2(n_64), .B1(n_445), .B2(n_821), .Y(n_820) );
NAND2xp5_ASAP7_75t_L g828 ( .A(n_52), .B(n_829), .Y(n_828) );
INVx1_ASAP7_75t_L g163 ( .A(n_53), .Y(n_163) );
INVx1_ASAP7_75t_L g182 ( .A(n_53), .Y(n_182) );
AOI22x1_ASAP7_75t_L g135 ( .A1(n_54), .A2(n_136), .B1(n_137), .B2(n_138), .Y(n_135) );
CKINVDCx20_ASAP7_75t_R g136 ( .A(n_54), .Y(n_136) );
AND2x2_ASAP7_75t_L g298 ( .A(n_55), .B(n_154), .Y(n_298) );
AOI221xp5_ASAP7_75t_L g254 ( .A1(n_56), .A2(n_78), .B1(n_160), .B2(n_170), .C(n_255), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_57), .B(n_160), .Y(n_215) );
NAND2xp5_ASAP7_75t_SL g547 ( .A(n_58), .B(n_537), .Y(n_547) );
INVx1_ASAP7_75t_L g809 ( .A(n_59), .Y(n_809) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_60), .B(n_189), .Y(n_275) );
AOI21xp5_ASAP7_75t_SL g211 ( .A1(n_61), .A2(n_170), .B(n_212), .Y(n_211) );
AND2x2_ASAP7_75t_L g575 ( .A(n_62), .B(n_154), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_63), .B(n_234), .Y(n_535) );
CKINVDCx20_ASAP7_75t_R g821 ( .A(n_64), .Y(n_821) );
INVx1_ASAP7_75t_L g225 ( .A(n_65), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_66), .B(n_231), .Y(n_573) );
AND2x2_ASAP7_75t_SL g595 ( .A(n_67), .B(n_155), .Y(n_595) );
AOI21xp5_ASAP7_75t_L g543 ( .A1(n_68), .A2(n_525), .B(n_544), .Y(n_543) );
INVx1_ASAP7_75t_L g296 ( .A(n_69), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_70), .B(n_234), .Y(n_560) );
AND2x2_ASAP7_75t_SL g567 ( .A(n_71), .B(n_206), .Y(n_567) );
XOR2xp5_ASAP7_75t_L g134 ( .A(n_72), .B(n_135), .Y(n_134) );
OAI22xp5_ASAP7_75t_L g138 ( .A1(n_73), .A2(n_104), .B1(n_139), .B2(n_140), .Y(n_138) );
CKINVDCx20_ASAP7_75t_R g139 ( .A(n_73), .Y(n_139) );
AOI21xp5_ASAP7_75t_L g294 ( .A1(n_74), .A2(n_170), .B(n_295), .Y(n_294) );
OAI22xp5_ASAP7_75t_L g818 ( .A1(n_75), .A2(n_819), .B1(n_820), .B2(n_822), .Y(n_818) );
CKINVDCx20_ASAP7_75t_R g819 ( .A(n_75), .Y(n_819) );
INVx1_ASAP7_75t_L g168 ( .A(n_76), .Y(n_168) );
INVx1_ASAP7_75t_L g184 ( .A(n_76), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_77), .B(n_160), .Y(n_250) );
AND2x2_ASAP7_75t_L g187 ( .A(n_79), .B(n_188), .Y(n_187) );
INVx1_ASAP7_75t_L g226 ( .A(n_80), .Y(n_226) );
AOI21xp5_ASAP7_75t_L g169 ( .A1(n_81), .A2(n_170), .B(n_176), .Y(n_169) );
A2O1A1Ixp33_ASAP7_75t_L g200 ( .A1(n_82), .A2(n_170), .B(n_201), .C(n_205), .Y(n_200) );
AOI22xp5_ASAP7_75t_L g565 ( .A1(n_83), .A2(n_88), .B1(n_160), .B2(n_537), .Y(n_565) );
NAND2xp5_ASAP7_75t_SL g574 ( .A(n_84), .B(n_537), .Y(n_574) );
INVx1_ASAP7_75t_L g112 ( .A(n_86), .Y(n_112) );
AND2x2_ASAP7_75t_SL g209 ( .A(n_87), .B(n_188), .Y(n_209) );
AOI22xp5_ASAP7_75t_L g244 ( .A1(n_89), .A2(n_170), .B1(n_245), .B2(n_246), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_90), .B(n_231), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_91), .B(n_231), .Y(n_602) );
AOI21xp5_ASAP7_75t_L g570 ( .A1(n_92), .A2(n_525), .B(n_571), .Y(n_570) );
INVx1_ASAP7_75t_L g213 ( .A(n_94), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_95), .B(n_234), .Y(n_572) );
AND2x2_ASAP7_75t_L g251 ( .A(n_96), .B(n_188), .Y(n_251) );
A2O1A1Ixp33_ASAP7_75t_L g263 ( .A1(n_97), .A2(n_264), .B(n_265), .C(n_267), .Y(n_263) );
INVxp67_ASAP7_75t_L g524 ( .A(n_98), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_99), .B(n_537), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_100), .B(n_234), .Y(n_545) );
AOI21xp5_ASAP7_75t_L g591 ( .A1(n_101), .A2(n_525), .B(n_592), .Y(n_591) );
BUFx2_ASAP7_75t_L g123 ( .A(n_102), .Y(n_123) );
INVx1_ASAP7_75t_SL g806 ( .A(n_102), .Y(n_806) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_103), .B(n_180), .Y(n_214) );
CKINVDCx20_ASAP7_75t_R g140 ( .A(n_104), .Y(n_140) );
INVx1_ASAP7_75t_SL g106 ( .A(n_107), .Y(n_106) );
CKINVDCx20_ASAP7_75t_R g107 ( .A(n_108), .Y(n_107) );
INVx1_ASAP7_75t_SL g108 ( .A(n_109), .Y(n_108) );
INVx1_ASAP7_75t_SL g832 ( .A(n_109), .Y(n_832) );
OR2x2_ASAP7_75t_L g109 ( .A(n_110), .B(n_113), .Y(n_109) );
CKINVDCx16_ASAP7_75t_R g110 ( .A(n_111), .Y(n_110) );
NAND2xp5_ASAP7_75t_L g130 ( .A(n_112), .B(n_131), .Y(n_130) );
INVx1_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
INVx2_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
AO21x2_ASAP7_75t_L g118 ( .A1(n_119), .A2(n_124), .B(n_804), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx2_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
HB1xp67_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
HB1xp67_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
NAND2xp5_ASAP7_75t_L g124 ( .A(n_125), .B(n_132), .Y(n_124) );
INVx3_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
OR2x2_ASAP7_75t_L g127 ( .A(n_128), .B(n_129), .Y(n_127) );
AND2x6_ASAP7_75t_SL g509 ( .A(n_128), .B(n_129), .Y(n_509) );
OR2x6_ASAP7_75t_SL g800 ( .A(n_128), .B(n_801), .Y(n_800) );
NAND2xp5_ASAP7_75t_L g827 ( .A(n_128), .B(n_801), .Y(n_827) );
CKINVDCx5p33_ASAP7_75t_R g801 ( .A(n_129), .Y(n_801) );
AOI22xp33_ASAP7_75t_L g132 ( .A1(n_133), .A2(n_134), .B1(n_141), .B2(n_802), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
INVx1_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
OAI22x1_ASAP7_75t_L g141 ( .A1(n_142), .A2(n_508), .B1(n_510), .B2(n_798), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
OAI22xp5_ASAP7_75t_L g802 ( .A1(n_143), .A2(n_508), .B1(n_511), .B2(n_803), .Y(n_802) );
AND3x1_ASAP7_75t_L g143 ( .A(n_144), .B(n_502), .C(n_505), .Y(n_143) );
NAND5xp2_ASAP7_75t_L g144 ( .A(n_145), .B(n_402), .C(n_432), .D(n_446), .E(n_472), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
OAI21xp33_ASAP7_75t_L g502 ( .A1(n_146), .A2(n_445), .B(n_503), .Y(n_502) );
INVx1_ASAP7_75t_L g815 ( .A(n_146), .Y(n_815) );
NAND2xp5_ASAP7_75t_L g146 ( .A(n_147), .B(n_351), .Y(n_146) );
NOR3xp33_ASAP7_75t_SL g147 ( .A(n_148), .B(n_299), .C(n_333), .Y(n_147) );
A2O1A1Ixp33_ASAP7_75t_L g148 ( .A1(n_149), .A2(n_216), .B(n_238), .C(n_277), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g149 ( .A(n_150), .B(n_191), .Y(n_149) );
BUFx2_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_151), .B(n_289), .Y(n_354) );
AND2x2_ASAP7_75t_L g441 ( .A(n_151), .B(n_219), .Y(n_441) );
HB1xp67_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
OR2x2_ASAP7_75t_L g237 ( .A(n_152), .B(n_208), .Y(n_237) );
INVx1_ASAP7_75t_L g279 ( .A(n_152), .Y(n_279) );
INVx2_ASAP7_75t_L g284 ( .A(n_152), .Y(n_284) );
HB1xp67_ASAP7_75t_L g312 ( .A(n_152), .Y(n_312) );
INVx1_ASAP7_75t_L g326 ( .A(n_152), .Y(n_326) );
AND2x2_ASAP7_75t_L g330 ( .A(n_152), .B(n_221), .Y(n_330) );
AND2x2_ASAP7_75t_L g411 ( .A(n_152), .B(n_220), .Y(n_411) );
AO21x2_ASAP7_75t_L g152 ( .A1(n_153), .A2(n_158), .B(n_187), .Y(n_152) );
AO21x2_ASAP7_75t_L g541 ( .A1(n_153), .A2(n_542), .B(n_548), .Y(n_541) );
AO21x2_ASAP7_75t_L g568 ( .A1(n_153), .A2(n_569), .B(n_575), .Y(n_568) );
AO21x2_ASAP7_75t_L g606 ( .A1(n_153), .A2(n_542), .B(n_548), .Y(n_606) );
CKINVDCx5p33_ASAP7_75t_R g153 ( .A(n_154), .Y(n_153) );
OA21x2_ASAP7_75t_L g598 ( .A1(n_154), .A2(n_599), .B(n_603), .Y(n_598) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
AND2x2_ASAP7_75t_SL g155 ( .A(n_156), .B(n_157), .Y(n_155) );
AND2x4_ASAP7_75t_L g199 ( .A(n_156), .B(n_157), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_159), .B(n_169), .Y(n_158) );
INVx1_ASAP7_75t_L g276 ( .A(n_160), .Y(n_276) );
AOI22xp5_ASAP7_75t_L g517 ( .A1(n_160), .A2(n_170), .B1(n_518), .B2(n_520), .Y(n_517) );
AND2x4_ASAP7_75t_L g160 ( .A(n_161), .B(n_166), .Y(n_160) );
INVx1_ASAP7_75t_L g196 ( .A(n_161), .Y(n_196) );
AND2x2_ASAP7_75t_L g161 ( .A(n_162), .B(n_164), .Y(n_161) );
OR2x6_ASAP7_75t_L g178 ( .A(n_162), .B(n_174), .Y(n_178) );
INVxp33_ASAP7_75t_L g248 ( .A(n_162), .Y(n_248) );
INVx2_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
AND2x2_ASAP7_75t_L g175 ( .A(n_163), .B(n_165), .Y(n_175) );
AND2x4_ASAP7_75t_L g234 ( .A(n_163), .B(n_183), .Y(n_234) );
HB1xp67_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
INVx1_ASAP7_75t_L g197 ( .A(n_166), .Y(n_197) );
BUFx3_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
AND2x6_ASAP7_75t_L g525 ( .A(n_167), .B(n_175), .Y(n_525) );
INVx2_ASAP7_75t_L g174 ( .A(n_168), .Y(n_174) );
AND2x6_ASAP7_75t_L g231 ( .A(n_168), .B(n_181), .Y(n_231) );
INVxp67_ASAP7_75t_L g274 ( .A(n_170), .Y(n_274) );
AND2x4_ASAP7_75t_L g170 ( .A(n_171), .B(n_175), .Y(n_170) );
NOR2x1p5_ASAP7_75t_L g171 ( .A(n_172), .B(n_173), .Y(n_171) );
INVx1_ASAP7_75t_L g249 ( .A(n_173), .Y(n_249) );
INVx3_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
O2A1O1Ixp33_ASAP7_75t_SL g176 ( .A1(n_177), .A2(n_178), .B(n_179), .C(n_185), .Y(n_176) );
INVx2_ASAP7_75t_L g204 ( .A(n_178), .Y(n_204) );
O2A1O1Ixp33_ASAP7_75t_L g212 ( .A1(n_178), .A2(n_185), .B(n_213), .C(n_214), .Y(n_212) );
OAI22xp5_ASAP7_75t_L g224 ( .A1(n_178), .A2(n_225), .B1(n_226), .B2(n_227), .Y(n_224) );
O2A1O1Ixp33_ASAP7_75t_SL g255 ( .A1(n_178), .A2(n_185), .B(n_256), .C(n_257), .Y(n_255) );
INVxp67_ASAP7_75t_L g264 ( .A(n_178), .Y(n_264) );
O2A1O1Ixp33_ASAP7_75t_L g295 ( .A1(n_178), .A2(n_185), .B(n_296), .C(n_297), .Y(n_295) );
INVx1_ASAP7_75t_L g227 ( .A(n_180), .Y(n_227) );
AND2x4_ASAP7_75t_L g537 ( .A(n_180), .B(n_186), .Y(n_537) );
AND2x4_ASAP7_75t_L g180 ( .A(n_181), .B(n_183), .Y(n_180) );
INVx2_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
INVx2_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
AOI21xp5_ASAP7_75t_L g201 ( .A1(n_185), .A2(n_202), .B(n_203), .Y(n_201) );
NOR2xp33_ASAP7_75t_L g235 ( .A(n_185), .B(n_199), .Y(n_235) );
INVx1_ASAP7_75t_L g245 ( .A(n_185), .Y(n_245) );
AOI21xp5_ASAP7_75t_L g533 ( .A1(n_185), .A2(n_534), .B(n_535), .Y(n_533) );
AOI21xp5_ASAP7_75t_L g544 ( .A1(n_185), .A2(n_545), .B(n_546), .Y(n_544) );
AOI21xp5_ASAP7_75t_L g558 ( .A1(n_185), .A2(n_559), .B(n_560), .Y(n_558) );
AOI21xp5_ASAP7_75t_L g571 ( .A1(n_185), .A2(n_572), .B(n_573), .Y(n_571) );
AOI21xp5_ASAP7_75t_L g592 ( .A1(n_185), .A2(n_593), .B(n_594), .Y(n_592) );
AOI21xp5_ASAP7_75t_L g600 ( .A1(n_185), .A2(n_601), .B(n_602), .Y(n_600) );
INVx5_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
HB1xp67_ASAP7_75t_L g267 ( .A(n_186), .Y(n_267) );
OAI22xp5_ASAP7_75t_L g262 ( .A1(n_188), .A2(n_263), .B1(n_268), .B2(n_269), .Y(n_262) );
INVx3_ASAP7_75t_L g269 ( .A(n_188), .Y(n_269) );
INVx4_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_189), .B(n_272), .Y(n_271) );
AOI21x1_ASAP7_75t_L g530 ( .A1(n_189), .A2(n_531), .B(n_538), .Y(n_530) );
INVx3_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
BUFx4f_ASAP7_75t_L g206 ( .A(n_190), .Y(n_206) );
AND2x4_ASAP7_75t_SL g191 ( .A(n_192), .B(n_207), .Y(n_191) );
HB1xp67_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
INVx2_ASAP7_75t_L g236 ( .A(n_193), .Y(n_236) );
AND2x2_ASAP7_75t_L g280 ( .A(n_193), .B(n_221), .Y(n_280) );
AND2x2_ASAP7_75t_L g301 ( .A(n_193), .B(n_208), .Y(n_301) );
INVx1_ASAP7_75t_L g324 ( .A(n_193), .Y(n_324) );
AND2x4_ASAP7_75t_L g391 ( .A(n_193), .B(n_220), .Y(n_391) );
AND2x2_ASAP7_75t_L g193 ( .A(n_194), .B(n_200), .Y(n_193) );
NOR3xp33_ASAP7_75t_L g195 ( .A(n_196), .B(n_197), .C(n_198), .Y(n_195) );
AOI21xp5_ASAP7_75t_L g210 ( .A1(n_199), .A2(n_211), .B(n_215), .Y(n_210) );
NOR2xp33_ASAP7_75t_L g518 ( .A(n_199), .B(n_519), .Y(n_518) );
NOR2xp33_ASAP7_75t_L g520 ( .A(n_199), .B(n_521), .Y(n_520) );
NOR2xp33_ASAP7_75t_L g523 ( .A(n_199), .B(n_524), .Y(n_523) );
NOR3xp33_ASAP7_75t_L g526 ( .A(n_199), .B(n_227), .C(n_527), .Y(n_526) );
AOI21xp5_ASAP7_75t_L g555 ( .A1(n_199), .A2(n_556), .B(n_557), .Y(n_555) );
AO21x2_ASAP7_75t_L g242 ( .A1(n_205), .A2(n_243), .B(n_251), .Y(n_242) );
AO21x2_ASAP7_75t_L g306 ( .A1(n_205), .A2(n_243), .B(n_251), .Y(n_306) );
AOI21x1_ASAP7_75t_L g563 ( .A1(n_205), .A2(n_564), .B(n_567), .Y(n_563) );
INVx2_ASAP7_75t_SL g205 ( .A(n_206), .Y(n_205) );
OA21x2_ASAP7_75t_L g253 ( .A1(n_206), .A2(n_254), .B(n_258), .Y(n_253) );
AOI21xp5_ASAP7_75t_L g589 ( .A1(n_206), .A2(n_590), .B(n_591), .Y(n_589) );
AND2x4_ASAP7_75t_L g407 ( .A(n_207), .B(n_324), .Y(n_407) );
OR2x2_ASAP7_75t_L g448 ( .A(n_207), .B(n_449), .Y(n_448) );
NOR2xp67_ASAP7_75t_SL g467 ( .A(n_207), .B(n_340), .Y(n_467) );
NOR2x1_ASAP7_75t_L g485 ( .A(n_207), .B(n_399), .Y(n_485) );
INVx4_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
NOR2x1_ASAP7_75t_SL g285 ( .A(n_208), .B(n_221), .Y(n_285) );
AND2x4_ASAP7_75t_L g323 ( .A(n_208), .B(n_324), .Y(n_323) );
BUFx6f_ASAP7_75t_L g329 ( .A(n_208), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_208), .B(n_283), .Y(n_361) );
INVx2_ASAP7_75t_L g375 ( .A(n_208), .Y(n_375) );
NAND2xp5_ASAP7_75t_SL g397 ( .A(n_208), .B(n_327), .Y(n_397) );
AND2x2_ASAP7_75t_L g489 ( .A(n_208), .B(n_347), .Y(n_489) );
OR2x6_ASAP7_75t_L g208 ( .A(n_209), .B(n_210), .Y(n_208) );
INVx1_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
NOR2x1_ASAP7_75t_L g217 ( .A(n_218), .B(n_237), .Y(n_217) );
INVx2_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_219), .B(n_326), .Y(n_340) );
AND2x2_ASAP7_75t_SL g349 ( .A(n_219), .B(n_329), .Y(n_349) );
AND2x2_ASAP7_75t_L g219 ( .A(n_220), .B(n_236), .Y(n_219) );
INVx1_ASAP7_75t_L g327 ( .A(n_220), .Y(n_327) );
INVx3_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
INVx2_ASAP7_75t_L g347 ( .A(n_221), .Y(n_347) );
AND2x4_ASAP7_75t_L g221 ( .A(n_222), .B(n_223), .Y(n_221) );
OAI21xp5_ASAP7_75t_L g223 ( .A1(n_224), .A2(n_228), .B(n_235), .Y(n_223) );
NOR2xp33_ASAP7_75t_L g265 ( .A(n_227), .B(n_266), .Y(n_265) );
OAI22xp5_ASAP7_75t_L g228 ( .A1(n_229), .A2(n_230), .B1(n_232), .B2(n_233), .Y(n_228) );
INVxp67_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
INVxp67_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
INVx1_ASAP7_75t_L g380 ( .A(n_236), .Y(n_380) );
INVx2_ASAP7_75t_SL g425 ( .A(n_237), .Y(n_425) );
INVx1_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
AND2x2_ASAP7_75t_L g239 ( .A(n_240), .B(n_259), .Y(n_239) );
NAND2x1p5_ASAP7_75t_L g334 ( .A(n_240), .B(n_335), .Y(n_334) );
BUFx2_ASAP7_75t_L g371 ( .A(n_240), .Y(n_371) );
AND2x2_ASAP7_75t_L g495 ( .A(n_240), .B(n_320), .Y(n_495) );
AND2x2_ASAP7_75t_L g240 ( .A(n_241), .B(n_252), .Y(n_240) );
AND2x4_ASAP7_75t_L g308 ( .A(n_241), .B(n_290), .Y(n_308) );
INVx1_ASAP7_75t_L g319 ( .A(n_241), .Y(n_319) );
AND2x2_ASAP7_75t_L g350 ( .A(n_241), .B(n_305), .Y(n_350) );
INVx2_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_242), .B(n_253), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_242), .B(n_291), .Y(n_382) );
NAND2xp5_ASAP7_75t_SL g243 ( .A(n_244), .B(n_250), .Y(n_243) );
INVx1_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
INVxp67_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
INVx2_ASAP7_75t_L g288 ( .A(n_253), .Y(n_288) );
AND2x4_ASAP7_75t_L g356 ( .A(n_253), .B(n_357), .Y(n_356) );
INVx1_ASAP7_75t_L g368 ( .A(n_253), .Y(n_368) );
INVx1_ASAP7_75t_L g410 ( .A(n_253), .Y(n_410) );
HB1xp67_ASAP7_75t_L g422 ( .A(n_253), .Y(n_422) );
AND2x2_ASAP7_75t_L g438 ( .A(n_253), .B(n_261), .Y(n_438) );
BUFx2_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
AND2x2_ASAP7_75t_L g385 ( .A(n_260), .B(n_343), .Y(n_385) );
INVx1_ASAP7_75t_SL g387 ( .A(n_260), .Y(n_387) );
AND2x2_ASAP7_75t_L g408 ( .A(n_260), .B(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
AND2x4_ASAP7_75t_L g287 ( .A(n_261), .B(n_288), .Y(n_287) );
INVx1_ASAP7_75t_L g315 ( .A(n_261), .Y(n_315) );
INVx2_ASAP7_75t_L g321 ( .A(n_261), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_261), .B(n_291), .Y(n_336) );
OR2x2_ASAP7_75t_L g261 ( .A(n_262), .B(n_270), .Y(n_261) );
AO21x2_ASAP7_75t_L g291 ( .A1(n_269), .A2(n_292), .B(n_298), .Y(n_291) );
AO21x2_ASAP7_75t_L g305 ( .A1(n_269), .A2(n_292), .B(n_298), .Y(n_305) );
OAI22xp5_ASAP7_75t_L g270 ( .A1(n_271), .A2(n_274), .B1(n_275), .B2(n_276), .Y(n_270) );
INVx1_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
OAI21xp5_ASAP7_75t_L g277 ( .A1(n_278), .A2(n_281), .B(n_286), .Y(n_277) );
INVx1_ASAP7_75t_L g417 ( .A(n_278), .Y(n_417) );
AND2x2_ASAP7_75t_L g278 ( .A(n_279), .B(n_280), .Y(n_278) );
INVx2_ASAP7_75t_L g337 ( .A(n_280), .Y(n_337) );
AND2x2_ASAP7_75t_L g393 ( .A(n_280), .B(n_329), .Y(n_393) );
AND2x2_ASAP7_75t_L g281 ( .A(n_282), .B(n_285), .Y(n_281) );
INVx1_ASAP7_75t_L g307 ( .A(n_282), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_282), .B(n_323), .Y(n_369) );
NOR2xp33_ASAP7_75t_L g398 ( .A(n_282), .B(n_399), .Y(n_398) );
AND2x2_ASAP7_75t_L g414 ( .A(n_282), .B(n_407), .Y(n_414) );
AND2x2_ASAP7_75t_L g488 ( .A(n_282), .B(n_489), .Y(n_488) );
INVx3_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
HB1xp67_ASAP7_75t_L g476 ( .A(n_283), .Y(n_476) );
INVx2_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
HB1xp67_ASAP7_75t_L g396 ( .A(n_284), .Y(n_396) );
AND2x2_ASAP7_75t_L g309 ( .A(n_285), .B(n_310), .Y(n_309) );
OAI21xp33_ASAP7_75t_L g497 ( .A1(n_285), .A2(n_498), .B(n_500), .Y(n_497) );
AND2x2_ASAP7_75t_L g286 ( .A(n_287), .B(n_289), .Y(n_286) );
INVx3_ASAP7_75t_L g383 ( .A(n_287), .Y(n_383) );
NAND2x1_ASAP7_75t_SL g427 ( .A(n_287), .B(n_428), .Y(n_427) );
AND2x2_ASAP7_75t_L g430 ( .A(n_287), .B(n_308), .Y(n_430) );
AND2x2_ASAP7_75t_L g342 ( .A(n_289), .B(n_343), .Y(n_342) );
OR2x2_ASAP7_75t_L g479 ( .A(n_289), .B(n_480), .Y(n_479) );
AND2x2_ASAP7_75t_L g490 ( .A(n_289), .B(n_438), .Y(n_490) );
INVx3_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
NAND2x1p5_ASAP7_75t_L g366 ( .A(n_290), .B(n_367), .Y(n_366) );
INVx3_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
AND2x2_ASAP7_75t_L g421 ( .A(n_291), .B(n_422), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_293), .B(n_294), .Y(n_292) );
OAI21xp5_ASAP7_75t_SL g299 ( .A1(n_300), .A2(n_313), .B(n_316), .Y(n_299) );
AOI22xp5_ASAP7_75t_L g300 ( .A1(n_301), .A2(n_302), .B1(n_308), .B2(n_309), .Y(n_300) );
HB1xp67_ASAP7_75t_L g358 ( .A(n_301), .Y(n_358) );
AND2x2_ASAP7_75t_L g302 ( .A(n_303), .B(n_307), .Y(n_302) );
AND2x2_ASAP7_75t_L g331 ( .A(n_303), .B(n_332), .Y(n_331) );
AND2x2_ASAP7_75t_L g437 ( .A(n_303), .B(n_438), .Y(n_437) );
AOI22xp5_ASAP7_75t_L g455 ( .A1(n_303), .A2(n_456), .B1(n_457), .B2(n_458), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_303), .B(n_464), .Y(n_463) );
AND2x4_ASAP7_75t_L g303 ( .A(n_304), .B(n_306), .Y(n_303) );
INVx2_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
AND2x2_ASAP7_75t_L g320 ( .A(n_305), .B(n_321), .Y(n_320) );
NOR2xp67_ASAP7_75t_L g401 ( .A(n_305), .B(n_321), .Y(n_401) );
NOR2x1_ASAP7_75t_L g409 ( .A(n_305), .B(n_410), .Y(n_409) );
INVx2_ASAP7_75t_L g357 ( .A(n_306), .Y(n_357) );
AND2x2_ASAP7_75t_L g365 ( .A(n_306), .B(n_321), .Y(n_365) );
INVx1_ASAP7_75t_L g428 ( .A(n_306), .Y(n_428) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
NAND2x1_ASAP7_75t_L g346 ( .A(n_311), .B(n_347), .Y(n_346) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
AND2x2_ASAP7_75t_L g458 ( .A(n_314), .B(n_343), .Y(n_458) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
INVx2_ASAP7_75t_L g332 ( .A(n_315), .Y(n_332) );
AND2x2_ASAP7_75t_L g355 ( .A(n_315), .B(n_356), .Y(n_355) );
AND2x2_ASAP7_75t_L g443 ( .A(n_315), .B(n_350), .Y(n_443) );
AOI22xp5_ASAP7_75t_L g316 ( .A1(n_317), .A2(n_322), .B1(n_328), .B2(n_331), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
OR2x2_ASAP7_75t_L g451 ( .A(n_318), .B(n_452), .Y(n_451) );
NAND2x1p5_ASAP7_75t_L g318 ( .A(n_319), .B(n_320), .Y(n_318) );
AND2x2_ASAP7_75t_L g481 ( .A(n_321), .B(n_368), .Y(n_481) );
AND2x2_ASAP7_75t_SL g322 ( .A(n_323), .B(n_325), .Y(n_322) );
INVx2_ASAP7_75t_L g348 ( .A(n_323), .Y(n_348) );
OAI21xp33_ASAP7_75t_SL g494 ( .A1(n_323), .A2(n_495), .B(n_496), .Y(n_494) );
AND2x4_ASAP7_75t_SL g325 ( .A(n_326), .B(n_327), .Y(n_325) );
HB1xp67_ASAP7_75t_L g484 ( .A(n_326), .Y(n_484) );
AND2x2_ASAP7_75t_L g328 ( .A(n_329), .B(n_330), .Y(n_328) );
O2A1O1Ixp33_ASAP7_75t_SL g426 ( .A1(n_329), .A2(n_427), .B(n_429), .C(n_431), .Y(n_426) );
AND2x2_ASAP7_75t_SL g378 ( .A(n_330), .B(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g431 ( .A(n_330), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_330), .B(n_407), .Y(n_471) );
INVx1_ASAP7_75t_SL g338 ( .A(n_331), .Y(n_338) );
AND2x2_ASAP7_75t_L g419 ( .A(n_332), .B(n_356), .Y(n_419) );
INVx1_ASAP7_75t_L g464 ( .A(n_332), .Y(n_464) );
OAI221xp5_ASAP7_75t_L g333 ( .A1(n_334), .A2(n_337), .B1(n_338), .B2(n_339), .C(n_341), .Y(n_333) );
HB1xp67_ASAP7_75t_L g453 ( .A(n_334), .Y(n_453) );
INVx2_ASAP7_75t_SL g335 ( .A(n_336), .Y(n_335) );
OR2x2_ASAP7_75t_L g501 ( .A(n_336), .B(n_344), .Y(n_501) );
OR2x2_ASAP7_75t_L g360 ( .A(n_337), .B(n_361), .Y(n_360) );
NOR2x1_ASAP7_75t_L g373 ( .A(n_337), .B(n_374), .Y(n_373) );
NOR2xp33_ASAP7_75t_L g460 ( .A(n_337), .B(n_461), .Y(n_460) );
OR2x2_ASAP7_75t_L g499 ( .A(n_337), .B(n_396), .Y(n_499) );
BUFx2_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
AOI32xp33_ASAP7_75t_L g341 ( .A1(n_342), .A2(n_345), .A3(n_348), .B1(n_349), .B2(n_350), .Y(n_341) );
INVx1_ASAP7_75t_L g362 ( .A(n_343), .Y(n_362) );
INVx2_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
NOR2xp33_ASAP7_75t_L g405 ( .A(n_345), .B(n_406), .Y(n_405) );
INVx2_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
INVx1_ASAP7_75t_L g457 ( .A(n_346), .Y(n_457) );
OAI22xp33_ASAP7_75t_SL g439 ( .A1(n_348), .A2(n_440), .B1(n_442), .B2(n_444), .Y(n_439) );
INVx1_ASAP7_75t_L g470 ( .A(n_349), .Y(n_470) );
AOI211x1_ASAP7_75t_L g351 ( .A1(n_352), .A2(n_358), .B(n_359), .C(n_376), .Y(n_351) );
AND2x2_ASAP7_75t_L g352 ( .A(n_353), .B(n_355), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_353), .B(n_438), .Y(n_444) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
AND2x4_ASAP7_75t_L g400 ( .A(n_356), .B(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g466 ( .A(n_356), .Y(n_466) );
OAI222xp33_ASAP7_75t_L g359 ( .A1(n_360), .A2(n_362), .B1(n_363), .B2(n_369), .C1(n_370), .C2(n_372), .Y(n_359) );
INVxp67_ASAP7_75t_L g456 ( .A(n_360), .Y(n_456) );
OR2x2_ASAP7_75t_L g363 ( .A(n_364), .B(n_366), .Y(n_363) );
NOR2xp33_ASAP7_75t_L g496 ( .A(n_364), .B(n_449), .Y(n_496) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
AND2x2_ASAP7_75t_L g412 ( .A(n_365), .B(n_409), .Y(n_412) );
INVx3_ASAP7_75t_L g452 ( .A(n_367), .Y(n_452) );
BUFx3_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
AND2x2_ASAP7_75t_L g390 ( .A(n_375), .B(n_391), .Y(n_390) );
OAI221xp5_ASAP7_75t_L g376 ( .A1(n_377), .A2(n_381), .B1(n_384), .B2(n_389), .C(n_392), .Y(n_376) );
INVx1_ASAP7_75t_SL g377 ( .A(n_378), .Y(n_377) );
OAI21xp5_ASAP7_75t_L g434 ( .A1(n_378), .A2(n_435), .B(n_437), .Y(n_434) );
INVx2_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
OR2x2_ASAP7_75t_L g381 ( .A(n_382), .B(n_383), .Y(n_381) );
INVx1_ASAP7_75t_L g388 ( .A(n_382), .Y(n_388) );
OR2x2_ASAP7_75t_L g492 ( .A(n_383), .B(n_428), .Y(n_492) );
NOR2xp67_ASAP7_75t_L g384 ( .A(n_385), .B(n_386), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_386), .B(n_414), .Y(n_413) );
AND2x2_ASAP7_75t_L g386 ( .A(n_387), .B(n_388), .Y(n_386) );
OAI21xp5_ASAP7_75t_L g486 ( .A1(n_389), .A2(n_418), .B(n_487), .Y(n_486) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
OAI21xp5_ASAP7_75t_L g468 ( .A1(n_390), .A2(n_462), .B(n_469), .Y(n_468) );
INVx4_ASAP7_75t_L g399 ( .A(n_391), .Y(n_399) );
OAI31xp33_ASAP7_75t_SL g392 ( .A1(n_393), .A2(n_394), .A3(n_398), .B(n_400), .Y(n_392) );
INVx1_ASAP7_75t_L g450 ( .A(n_394), .Y(n_450) );
NOR2x1_ASAP7_75t_L g394 ( .A(n_395), .B(n_397), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx2_ASAP7_75t_L g424 ( .A(n_399), .Y(n_424) );
AND2x2_ASAP7_75t_L g402 ( .A(n_403), .B(n_415), .Y(n_402) );
NAND4xp25_ASAP7_75t_L g503 ( .A(n_403), .B(n_415), .C(n_434), .D(n_504), .Y(n_503) );
AND2x2_ASAP7_75t_L g403 ( .A(n_404), .B(n_413), .Y(n_403) );
AOI22xp5_ASAP7_75t_L g404 ( .A1(n_405), .A2(n_408), .B1(n_411), .B2(n_412), .Y(n_404) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
AND2x2_ASAP7_75t_L g475 ( .A(n_407), .B(n_476), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_408), .B(n_428), .Y(n_436) );
INVx1_ASAP7_75t_SL g449 ( .A(n_411), .Y(n_449) );
NOR2xp33_ASAP7_75t_L g415 ( .A(n_416), .B(n_426), .Y(n_415) );
OAI22xp5_ASAP7_75t_L g416 ( .A1(n_417), .A2(n_418), .B1(n_420), .B2(n_423), .Y(n_416) );
INVx3_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVxp67_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
NAND2x1_ASAP7_75t_L g423 ( .A(n_424), .B(n_425), .Y(n_423) );
AOI22xp5_ASAP7_75t_L g487 ( .A1(n_425), .A2(n_488), .B1(n_490), .B2(n_491), .Y(n_487) );
INVx2_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
NOR3xp33_ASAP7_75t_L g432 ( .A(n_433), .B(n_439), .C(n_445), .Y(n_432) );
INVxp67_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g504 ( .A(n_439), .Y(n_504) );
INVx2_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
OAI21xp33_ASAP7_75t_L g505 ( .A1(n_445), .A2(n_506), .B(n_507), .Y(n_505) );
INVxp33_ASAP7_75t_L g506 ( .A(n_446), .Y(n_506) );
AND2x2_ASAP7_75t_L g814 ( .A(n_446), .B(n_472), .Y(n_814) );
NOR2xp67_ASAP7_75t_L g446 ( .A(n_447), .B(n_454), .Y(n_446) );
AOI22xp33_ASAP7_75t_L g447 ( .A1(n_448), .A2(n_450), .B1(n_451), .B2(n_453), .Y(n_447) );
OAI21xp5_ASAP7_75t_L g473 ( .A1(n_451), .A2(n_474), .B(n_477), .Y(n_473) );
INVx2_ASAP7_75t_L g461 ( .A(n_452), .Y(n_461) );
NAND3xp33_ASAP7_75t_SL g454 ( .A(n_455), .B(n_459), .C(n_468), .Y(n_454) );
AOI22xp5_ASAP7_75t_L g459 ( .A1(n_460), .A2(n_462), .B1(n_465), .B2(n_467), .Y(n_459) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx1_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_470), .B(n_471), .Y(n_469) );
INVxp33_ASAP7_75t_SL g507 ( .A(n_472), .Y(n_507) );
NOR3x1_ASAP7_75t_L g472 ( .A(n_473), .B(n_486), .C(n_493), .Y(n_472) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_478), .B(n_482), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
INVx2_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
INVx1_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_484), .B(n_485), .Y(n_483) );
INVx1_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
NAND2xp5_ASAP7_75t_SL g493 ( .A(n_494), .B(n_497), .Y(n_493) );
INVx1_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
INVx1_ASAP7_75t_SL g500 ( .A(n_501), .Y(n_500) );
INVx1_ASAP7_75t_L g816 ( .A(n_503), .Y(n_816) );
CKINVDCx11_ASAP7_75t_R g508 ( .A(n_509), .Y(n_508) );
INVx3_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
AND2x4_ASAP7_75t_L g511 ( .A(n_512), .B(n_675), .Y(n_511) );
NOR4xp25_ASAP7_75t_L g512 ( .A(n_513), .B(n_618), .C(n_657), .D(n_664), .Y(n_512) );
OAI221xp5_ASAP7_75t_L g513 ( .A1(n_514), .A2(n_539), .B1(n_576), .B2(n_585), .C(n_604), .Y(n_513) );
OR2x2_ASAP7_75t_L g748 ( .A(n_514), .B(n_610), .Y(n_748) );
INVx1_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
AND2x2_ASAP7_75t_L g663 ( .A(n_515), .B(n_588), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_515), .B(n_683), .Y(n_682) );
AND2x2_ASAP7_75t_SL g728 ( .A(n_515), .B(n_729), .Y(n_728) );
AND2x4_ASAP7_75t_L g515 ( .A(n_516), .B(n_528), .Y(n_515) );
AND2x4_ASAP7_75t_SL g587 ( .A(n_516), .B(n_588), .Y(n_587) );
INVx3_ASAP7_75t_L g609 ( .A(n_516), .Y(n_609) );
AND2x2_ASAP7_75t_L g644 ( .A(n_516), .B(n_617), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_516), .B(n_529), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_516), .B(n_611), .Y(n_696) );
OR2x2_ASAP7_75t_L g774 ( .A(n_516), .B(n_588), .Y(n_774) );
AND2x4_ASAP7_75t_L g516 ( .A(n_517), .B(n_522), .Y(n_516) );
INVx2_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
AND2x2_ASAP7_75t_L g596 ( .A(n_529), .B(n_597), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_529), .B(n_617), .Y(n_616) );
INVx1_ASAP7_75t_L g622 ( .A(n_529), .Y(n_622) );
OR2x2_ASAP7_75t_L g627 ( .A(n_529), .B(n_611), .Y(n_627) );
AND2x2_ASAP7_75t_L g640 ( .A(n_529), .B(n_598), .Y(n_640) );
HB1xp67_ASAP7_75t_L g643 ( .A(n_529), .Y(n_643) );
INVx1_ASAP7_75t_L g655 ( .A(n_529), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_529), .B(n_609), .Y(n_720) );
INVx3_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_532), .B(n_536), .Y(n_531) );
NAND2xp5_ASAP7_75t_SL g539 ( .A(n_540), .B(n_549), .Y(n_539) );
HB1xp67_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
OR2x2_ASAP7_75t_L g584 ( .A(n_541), .B(n_568), .Y(n_584) );
AND2x4_ASAP7_75t_L g614 ( .A(n_541), .B(n_553), .Y(n_614) );
INVx2_ASAP7_75t_L g648 ( .A(n_541), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_541), .B(n_568), .Y(n_706) );
AND2x2_ASAP7_75t_L g753 ( .A(n_541), .B(n_582), .Y(n_753) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_543), .B(n_547), .Y(n_542) );
AOI222xp33_ASAP7_75t_L g741 ( .A1(n_549), .A2(n_613), .B1(n_656), .B2(n_716), .C1(n_742), .C2(n_744), .Y(n_741) );
INVx1_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_551), .B(n_561), .Y(n_550) );
AND2x2_ASAP7_75t_L g660 ( .A(n_551), .B(n_580), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_551), .B(n_711), .Y(n_710) );
AND2x2_ASAP7_75t_L g789 ( .A(n_551), .B(n_629), .Y(n_789) );
INVx2_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
AOI21xp5_ASAP7_75t_L g619 ( .A1(n_552), .A2(n_620), .B(n_624), .Y(n_619) );
AND2x2_ASAP7_75t_L g700 ( .A(n_552), .B(n_583), .Y(n_700) );
OR2x2_ASAP7_75t_L g725 ( .A(n_552), .B(n_584), .Y(n_725) );
INVx2_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
INVx5_ASAP7_75t_L g579 ( .A(n_553), .Y(n_579) );
AND2x2_ASAP7_75t_L g666 ( .A(n_553), .B(n_648), .Y(n_666) );
AND2x2_ASAP7_75t_L g692 ( .A(n_553), .B(n_568), .Y(n_692) );
OR2x2_ASAP7_75t_L g695 ( .A(n_553), .B(n_582), .Y(n_695) );
HB1xp67_ASAP7_75t_L g713 ( .A(n_553), .Y(n_713) );
AND2x4_ASAP7_75t_SL g770 ( .A(n_553), .B(n_647), .Y(n_770) );
OR2x2_ASAP7_75t_L g779 ( .A(n_553), .B(n_606), .Y(n_779) );
OR2x6_ASAP7_75t_L g553 ( .A(n_554), .B(n_555), .Y(n_553) );
INVx1_ASAP7_75t_L g612 ( .A(n_561), .Y(n_612) );
AOI221xp5_ASAP7_75t_SL g730 ( .A1(n_561), .A2(n_614), .B1(n_731), .B2(n_733), .C(n_734), .Y(n_730) );
AND2x2_ASAP7_75t_L g561 ( .A(n_562), .B(n_568), .Y(n_561) );
OR2x2_ASAP7_75t_L g669 ( .A(n_562), .B(n_639), .Y(n_669) );
OR2x2_ASAP7_75t_L g679 ( .A(n_562), .B(n_680), .Y(n_679) );
OR2x2_ASAP7_75t_L g705 ( .A(n_562), .B(n_706), .Y(n_705) );
AND2x4_ASAP7_75t_L g711 ( .A(n_562), .B(n_630), .Y(n_711) );
NOR2xp33_ASAP7_75t_L g723 ( .A(n_562), .B(n_694), .Y(n_723) );
INVx2_ASAP7_75t_L g736 ( .A(n_562), .Y(n_736) );
NAND2xp5_ASAP7_75t_SL g757 ( .A(n_562), .B(n_614), .Y(n_757) );
AND2x2_ASAP7_75t_L g761 ( .A(n_562), .B(n_583), .Y(n_761) );
AND2x2_ASAP7_75t_L g769 ( .A(n_562), .B(n_770), .Y(n_769) );
BUFx6f_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
INVx2_ASAP7_75t_L g582 ( .A(n_563), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_565), .B(n_566), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_568), .B(n_579), .Y(n_578) );
AND2x2_ASAP7_75t_L g613 ( .A(n_568), .B(n_582), .Y(n_613) );
INVx2_ASAP7_75t_L g630 ( .A(n_568), .Y(n_630) );
AND2x4_ASAP7_75t_L g647 ( .A(n_568), .B(n_648), .Y(n_647) );
HB1xp67_ASAP7_75t_L g752 ( .A(n_568), .Y(n_752) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_570), .B(n_574), .Y(n_569) );
NOR2xp33_ASAP7_75t_L g576 ( .A(n_577), .B(n_580), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
OR2x2_ASAP7_75t_L g759 ( .A(n_578), .B(n_581), .Y(n_759) );
AND2x4_ASAP7_75t_L g605 ( .A(n_579), .B(n_606), .Y(n_605) );
AND2x2_ASAP7_75t_L g646 ( .A(n_579), .B(n_647), .Y(n_646) );
AND2x2_ASAP7_75t_L g673 ( .A(n_579), .B(n_613), .Y(n_673) );
AND2x2_ASAP7_75t_L g580 ( .A(n_581), .B(n_583), .Y(n_580) );
AND2x2_ASAP7_75t_L g777 ( .A(n_581), .B(n_778), .Y(n_777) );
BUFx2_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
AND2x2_ASAP7_75t_L g629 ( .A(n_582), .B(n_630), .Y(n_629) );
OAI21xp5_ASAP7_75t_SL g649 ( .A1(n_583), .A2(n_650), .B(n_656), .Y(n_649) );
INVx2_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
INVx1_ASAP7_75t_SL g585 ( .A(n_586), .Y(n_585) );
AND2x2_ASAP7_75t_L g586 ( .A(n_587), .B(n_596), .Y(n_586) );
INVx1_ASAP7_75t_SL g703 ( .A(n_587), .Y(n_703) );
AND2x2_ASAP7_75t_L g733 ( .A(n_587), .B(n_643), .Y(n_733) );
AND2x4_ASAP7_75t_L g744 ( .A(n_587), .B(n_745), .Y(n_744) );
OR2x2_ASAP7_75t_L g610 ( .A(n_588), .B(n_611), .Y(n_610) );
INVx2_ASAP7_75t_L g617 ( .A(n_588), .Y(n_617) );
AND2x4_ASAP7_75t_L g623 ( .A(n_588), .B(n_609), .Y(n_623) );
INVx2_ASAP7_75t_L g634 ( .A(n_588), .Y(n_634) );
INVx1_ASAP7_75t_L g683 ( .A(n_588), .Y(n_683) );
OR2x2_ASAP7_75t_L g704 ( .A(n_588), .B(n_688), .Y(n_704) );
OR2x2_ASAP7_75t_L g718 ( .A(n_588), .B(n_598), .Y(n_718) );
HB1xp67_ASAP7_75t_L g784 ( .A(n_588), .Y(n_784) );
NAND2xp5_ASAP7_75t_L g790 ( .A(n_588), .B(n_640), .Y(n_790) );
OR2x6_ASAP7_75t_L g588 ( .A(n_589), .B(n_595), .Y(n_588) );
INVx1_ASAP7_75t_L g635 ( .A(n_596), .Y(n_635) );
AND2x2_ASAP7_75t_L g768 ( .A(n_596), .B(n_634), .Y(n_768) );
AND2x2_ASAP7_75t_L g793 ( .A(n_596), .B(n_623), .Y(n_793) );
INVx2_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
INVx2_ASAP7_75t_L g611 ( .A(n_598), .Y(n_611) );
BUFx3_ASAP7_75t_L g653 ( .A(n_598), .Y(n_653) );
HB1xp67_ASAP7_75t_L g680 ( .A(n_598), .Y(n_680) );
INVx1_ASAP7_75t_L g689 ( .A(n_598), .Y(n_689) );
AOI33xp33_ASAP7_75t_L g604 ( .A1(n_605), .A2(n_607), .A3(n_612), .B1(n_613), .B2(n_614), .B3(n_615), .Y(n_604) );
AOI21x1_ASAP7_75t_SL g707 ( .A1(n_605), .A2(n_629), .B(n_691), .Y(n_707) );
INVx2_ASAP7_75t_L g737 ( .A(n_605), .Y(n_737) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_605), .B(n_736), .Y(n_743) );
AND2x2_ASAP7_75t_L g691 ( .A(n_606), .B(n_692), .Y(n_691) );
INVx1_ASAP7_75t_SL g607 ( .A(n_608), .Y(n_607) );
OR2x2_ASAP7_75t_L g608 ( .A(n_609), .B(n_610), .Y(n_608) );
AND2x2_ASAP7_75t_L g654 ( .A(n_609), .B(n_655), .Y(n_654) );
INVx2_ASAP7_75t_L g755 ( .A(n_610), .Y(n_755) );
HB1xp67_ASAP7_75t_L g745 ( .A(n_611), .Y(n_745) );
OAI32xp33_ASAP7_75t_L g794 ( .A1(n_612), .A2(n_614), .A3(n_790), .B1(n_795), .B2(n_797), .Y(n_794) );
AND2x2_ASAP7_75t_L g712 ( .A(n_613), .B(n_713), .Y(n_712) );
INVx2_ASAP7_75t_SL g702 ( .A(n_614), .Y(n_702) );
AND2x2_ASAP7_75t_L g767 ( .A(n_614), .B(n_711), .Y(n_767) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
OAI221xp5_ASAP7_75t_L g618 ( .A1(n_619), .A2(n_628), .B1(n_631), .B2(n_645), .C(n_649), .Y(n_618) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_622), .B(n_623), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_622), .B(n_689), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_623), .B(n_626), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g738 ( .A(n_623), .B(n_739), .Y(n_738) );
NAND2xp5_ASAP7_75t_L g762 ( .A(n_623), .B(n_763), .Y(n_762) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
INVx1_ASAP7_75t_L g672 ( .A(n_627), .Y(n_672) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
NOR3xp33_ASAP7_75t_L g631 ( .A(n_632), .B(n_636), .C(n_641), .Y(n_631) );
INVx1_ASAP7_75t_SL g632 ( .A(n_633), .Y(n_632) );
OAI22xp33_ASAP7_75t_L g734 ( .A1(n_633), .A2(n_695), .B1(n_735), .B2(n_738), .Y(n_734) );
OR2x2_ASAP7_75t_L g633 ( .A(n_634), .B(n_635), .Y(n_633) );
INVx1_ASAP7_75t_L g638 ( .A(n_634), .Y(n_638) );
NOR2x1p5_ASAP7_75t_L g652 ( .A(n_634), .B(n_653), .Y(n_652) );
HB1xp67_ASAP7_75t_L g674 ( .A(n_634), .Y(n_674) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
OAI322xp33_ASAP7_75t_L g701 ( .A1(n_637), .A2(n_679), .A3(n_702), .B1(n_703), .B2(n_704), .C1(n_705), .C2(n_707), .Y(n_701) );
OR2x2_ASAP7_75t_L g637 ( .A(n_638), .B(n_639), .Y(n_637) );
A2O1A1Ixp33_ASAP7_75t_L g657 ( .A1(n_639), .A2(n_658), .B(n_659), .C(n_661), .Y(n_657) );
OR2x2_ASAP7_75t_L g749 ( .A(n_639), .B(n_703), .Y(n_749) );
INVx2_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
AND2x2_ASAP7_75t_L g656 ( .A(n_640), .B(n_644), .Y(n_656) );
INVx1_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_643), .B(n_644), .Y(n_642) );
INVx2_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
AND2x2_ASAP7_75t_L g662 ( .A(n_646), .B(n_663), .Y(n_662) );
INVx3_ASAP7_75t_SL g694 ( .A(n_647), .Y(n_694) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_651), .B(n_715), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_652), .B(n_654), .Y(n_651) );
INVx1_ASAP7_75t_SL g698 ( .A(n_654), .Y(n_698) );
HB1xp67_ASAP7_75t_L g740 ( .A(n_655), .Y(n_740) );
OR2x6_ASAP7_75t_SL g795 ( .A(n_658), .B(n_796), .Y(n_795) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
INVxp67_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
AOI211xp5_ASAP7_75t_L g785 ( .A1(n_663), .A2(n_786), .B(n_787), .C(n_794), .Y(n_785) );
O2A1O1Ixp33_ASAP7_75t_SL g664 ( .A1(n_665), .A2(n_667), .B(n_670), .C(n_674), .Y(n_664) );
OAI211xp5_ASAP7_75t_SL g676 ( .A1(n_665), .A2(n_677), .B(n_684), .C(n_708), .Y(n_676) );
INVx2_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
INVx3_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
INVxp67_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
AND2x2_ASAP7_75t_L g671 ( .A(n_672), .B(n_673), .Y(n_671) );
NOR3xp33_ASAP7_75t_L g675 ( .A(n_676), .B(n_721), .C(n_765), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_678), .B(n_681), .Y(n_677) );
INVx1_ASAP7_75t_SL g678 ( .A(n_679), .Y(n_678) );
HB1xp67_ASAP7_75t_L g772 ( .A(n_680), .Y(n_772) );
INVx1_ASAP7_75t_SL g681 ( .A(n_682), .Y(n_681) );
INVx1_ASAP7_75t_L g727 ( .A(n_683), .Y(n_727) );
NOR3xp33_ASAP7_75t_SL g684 ( .A(n_685), .B(n_697), .C(n_701), .Y(n_684) );
OAI22xp5_ASAP7_75t_L g685 ( .A1(n_686), .A2(n_690), .B1(n_693), .B2(n_696), .Y(n_685) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g729 ( .A(n_689), .Y(n_729) );
INVxp67_ASAP7_75t_SL g796 ( .A(n_689), .Y(n_796) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
OR2x2_ASAP7_75t_L g693 ( .A(n_694), .B(n_695), .Y(n_693) );
INVx1_ASAP7_75t_SL g782 ( .A(n_695), .Y(n_782) );
NOR2xp33_ASAP7_75t_L g697 ( .A(n_698), .B(n_699), .Y(n_697) );
OR2x2_ASAP7_75t_L g732 ( .A(n_698), .B(n_718), .Y(n_732) );
OR2x2_ASAP7_75t_L g783 ( .A(n_698), .B(n_784), .Y(n_783) );
INVx2_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
INVx1_ASAP7_75t_L g781 ( .A(n_706), .Y(n_781) );
OR2x2_ASAP7_75t_L g797 ( .A(n_706), .B(n_736), .Y(n_797) );
OAI21xp33_ASAP7_75t_L g708 ( .A1(n_709), .A2(n_712), .B(n_714), .Y(n_708) );
OAI31xp33_ASAP7_75t_L g722 ( .A1(n_709), .A2(n_723), .A3(n_724), .B(n_726), .Y(n_722) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
AND2x2_ASAP7_75t_L g716 ( .A(n_717), .B(n_719), .Y(n_716) );
INVx1_ASAP7_75t_SL g717 ( .A(n_718), .Y(n_717) );
AND2x4_ASAP7_75t_L g754 ( .A(n_719), .B(n_755), .Y(n_754) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
NAND4xp25_ASAP7_75t_SL g721 ( .A(n_722), .B(n_730), .C(n_741), .D(n_746), .Y(n_721) );
INVx1_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
AND2x2_ASAP7_75t_L g726 ( .A(n_727), .B(n_728), .Y(n_726) );
HB1xp67_ASAP7_75t_L g764 ( .A(n_729), .Y(n_764) );
INVx1_ASAP7_75t_SL g731 ( .A(n_732), .Y(n_731) );
OR2x2_ASAP7_75t_L g735 ( .A(n_736), .B(n_737), .Y(n_735) );
INVxp67_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
INVx1_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
AOI221xp5_ASAP7_75t_L g746 ( .A1(n_747), .A2(n_750), .B1(n_754), .B2(n_756), .C(n_758), .Y(n_746) );
NAND2xp33_ASAP7_75t_SL g747 ( .A(n_748), .B(n_749), .Y(n_747) );
INVx1_ASAP7_75t_L g791 ( .A(n_750), .Y(n_791) );
AND2x2_ASAP7_75t_SL g750 ( .A(n_751), .B(n_753), .Y(n_750) );
INVx1_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
INVx1_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
AOI21xp33_ASAP7_75t_L g758 ( .A1(n_759), .A2(n_760), .B(n_762), .Y(n_758) );
INVx1_ASAP7_75t_L g786 ( .A(n_760), .Y(n_786) );
INVx2_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
INVx1_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
NAND2xp5_ASAP7_75t_SL g765 ( .A(n_766), .B(n_785), .Y(n_765) );
AOI221xp5_ASAP7_75t_L g766 ( .A1(n_767), .A2(n_768), .B1(n_769), .B2(n_771), .C(n_775), .Y(n_766) );
AND2x2_ASAP7_75t_L g771 ( .A(n_772), .B(n_773), .Y(n_771) );
INVx1_ASAP7_75t_SL g773 ( .A(n_774), .Y(n_773) );
AOI21xp33_ASAP7_75t_L g775 ( .A1(n_776), .A2(n_780), .B(n_783), .Y(n_775) );
INVxp33_ASAP7_75t_L g776 ( .A(n_777), .Y(n_776) );
INVx1_ASAP7_75t_SL g778 ( .A(n_779), .Y(n_778) );
NAND2xp5_ASAP7_75t_L g780 ( .A(n_781), .B(n_782), .Y(n_780) );
OAI22xp5_ASAP7_75t_L g787 ( .A1(n_788), .A2(n_790), .B1(n_791), .B2(n_792), .Y(n_787) );
INVx1_ASAP7_75t_L g788 ( .A(n_789), .Y(n_788) );
INVx1_ASAP7_75t_L g792 ( .A(n_793), .Y(n_792) );
CKINVDCx5p33_ASAP7_75t_R g798 ( .A(n_799), .Y(n_798) );
CKINVDCx20_ASAP7_75t_R g803 ( .A(n_799), .Y(n_803) );
CKINVDCx11_ASAP7_75t_R g799 ( .A(n_800), .Y(n_799) );
OAI21xp5_ASAP7_75t_L g804 ( .A1(n_805), .A2(n_807), .B(n_828), .Y(n_804) );
INVx2_ASAP7_75t_SL g805 ( .A(n_806), .Y(n_805) );
OAI21xp5_ASAP7_75t_L g807 ( .A1(n_808), .A2(n_811), .B(n_823), .Y(n_807) );
AOI21xp5_ASAP7_75t_L g823 ( .A1(n_808), .A2(n_824), .B(n_825), .Y(n_823) );
INVxp67_ASAP7_75t_SL g811 ( .A(n_812), .Y(n_811) );
INVx1_ASAP7_75t_L g824 ( .A(n_812), .Y(n_824) );
XNOR2xp5_ASAP7_75t_L g812 ( .A(n_813), .B(n_817), .Y(n_812) );
NAND3x1_ASAP7_75t_L g813 ( .A(n_814), .B(n_815), .C(n_816), .Y(n_813) );
CKINVDCx5p33_ASAP7_75t_R g817 ( .A(n_818), .Y(n_817) );
INVx1_ASAP7_75t_L g822 ( .A(n_820), .Y(n_822) );
CKINVDCx11_ASAP7_75t_R g830 ( .A(n_825), .Y(n_830) );
CKINVDCx20_ASAP7_75t_R g825 ( .A(n_826), .Y(n_825) );
BUFx3_ASAP7_75t_L g826 ( .A(n_827), .Y(n_826) );
CKINVDCx20_ASAP7_75t_R g829 ( .A(n_830), .Y(n_829) );
CKINVDCx20_ASAP7_75t_R g831 ( .A(n_832), .Y(n_831) );
endmodule