module fake_jpeg_14317_n_459 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_459);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_459;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_260;
wire n_199;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

INVx6_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_13),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_10),
.Y(n_33)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_7),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_7),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_3),
.B(n_2),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_3),
.Y(n_43)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_15),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_7),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_7),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_42),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_48),
.B(n_54),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_18),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_49),
.Y(n_108)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_20),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g122 ( 
.A(n_50),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_18),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_51),
.Y(n_112)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_20),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g119 ( 
.A(n_52),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_42),
.B(n_15),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_53),
.B(n_55),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_19),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_19),
.B(n_14),
.Y(n_55)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

INVx11_ASAP7_75t_L g138 ( 
.A(n_56),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_18),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_57),
.Y(n_144)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_20),
.Y(n_58)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_58),
.Y(n_117)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_27),
.Y(n_59)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_59),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_18),
.Y(n_60)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_60),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_21),
.B(n_13),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_61),
.B(n_64),
.Y(n_147)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_62),
.Y(n_102)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_16),
.Y(n_63)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_63),
.Y(n_107)
);

INVx2_ASAP7_75t_R g64 ( 
.A(n_27),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_32),
.Y(n_65)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_65),
.Y(n_109)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

INVx5_ASAP7_75t_L g145 ( 
.A(n_66),
.Y(n_145)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_30),
.Y(n_67)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_67),
.Y(n_110)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_30),
.Y(n_68)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_68),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_32),
.Y(n_69)
);

INVx6_ASAP7_75t_L g129 ( 
.A(n_69),
.Y(n_129)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_70),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_16),
.B(n_1),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_71),
.B(n_77),
.Y(n_103)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_35),
.Y(n_72)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_72),
.Y(n_99)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_31),
.Y(n_73)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_73),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_40),
.Y(n_74)
);

INVx5_ASAP7_75t_L g146 ( 
.A(n_74),
.Y(n_146)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_31),
.Y(n_75)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_75),
.Y(n_104)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_24),
.Y(n_76)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_76),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_24),
.Y(n_77)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_35),
.Y(n_78)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_78),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_32),
.Y(n_79)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_79),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_32),
.Y(n_80)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_80),
.Y(n_141)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_40),
.Y(n_81)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_81),
.Y(n_116)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_35),
.Y(n_82)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_82),
.Y(n_124)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_40),
.Y(n_83)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_83),
.Y(n_118)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_25),
.Y(n_84)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_84),
.Y(n_133)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_40),
.Y(n_85)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_85),
.Y(n_121)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_40),
.Y(n_86)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_86),
.Y(n_139)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_23),
.Y(n_87)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_87),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_44),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_88),
.B(n_89),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_21),
.B(n_1),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_36),
.Y(n_90)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_90),
.Y(n_142)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_36),
.Y(n_91)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_91),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_22),
.B(n_3),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_92),
.B(n_95),
.Y(n_115)
);

BUFx12f_ASAP7_75t_L g93 ( 
.A(n_36),
.Y(n_93)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_93),
.Y(n_136)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_23),
.Y(n_94)
);

HB1xp67_ASAP7_75t_L g101 ( 
.A(n_94),
.Y(n_101)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_25),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_91),
.A2(n_29),
.B1(n_39),
.B2(n_44),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_97),
.A2(n_98),
.B1(n_100),
.B2(n_128),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_62),
.A2(n_23),
.B1(n_44),
.B2(n_17),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_50),
.A2(n_17),
.B1(n_31),
.B2(n_36),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_64),
.B(n_28),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_125),
.B(n_130),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_49),
.A2(n_29),
.B1(n_39),
.B2(n_17),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_126),
.A2(n_140),
.B1(n_69),
.B2(n_26),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_50),
.A2(n_29),
.B1(n_39),
.B2(n_41),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_56),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_73),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_131),
.B(n_93),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_L g132 ( 
.A1(n_51),
.A2(n_65),
.B1(n_90),
.B2(n_57),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_132),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_197)
);

INVx5_ASAP7_75t_SL g137 ( 
.A(n_66),
.Y(n_137)
);

INVx4_ASAP7_75t_SL g182 ( 
.A(n_137),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_60),
.A2(n_39),
.B1(n_45),
.B2(n_43),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_66),
.A2(n_46),
.B1(n_41),
.B2(n_47),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_149),
.A2(n_70),
.B1(n_37),
.B2(n_43),
.Y(n_154)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_72),
.Y(n_150)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_150),
.Y(n_167)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_133),
.Y(n_151)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_151),
.Y(n_199)
);

A2O1A1Ixp33_ASAP7_75t_L g152 ( 
.A1(n_147),
.A2(n_46),
.B(n_47),
.C(n_34),
.Y(n_152)
);

A2O1A1Ixp33_ASAP7_75t_L g207 ( 
.A1(n_152),
.A2(n_138),
.B(n_128),
.C(n_98),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_147),
.B(n_45),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_153),
.B(n_161),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_154),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_101),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_155),
.B(n_163),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_105),
.B(n_82),
.Y(n_156)
);

INVx1_ASAP7_75t_SL g221 ( 
.A(n_156),
.Y(n_221)
);

OA22x2_ASAP7_75t_SL g157 ( 
.A1(n_110),
.A2(n_75),
.B1(n_87),
.B2(n_52),
.Y(n_157)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_157),
.Y(n_224)
);

OA22x2_ASAP7_75t_L g158 ( 
.A1(n_132),
.A2(n_78),
.B1(n_80),
.B2(n_79),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_158),
.Y(n_223)
);

BUFx12f_ASAP7_75t_L g159 ( 
.A(n_122),
.Y(n_159)
);

INVx4_ASAP7_75t_L g225 ( 
.A(n_159),
.Y(n_225)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_107),
.Y(n_160)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_160),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_123),
.B(n_103),
.Y(n_161)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_134),
.Y(n_162)
);

INVx4_ASAP7_75t_L g226 ( 
.A(n_162),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_113),
.Y(n_163)
);

BUFx3_ASAP7_75t_L g164 ( 
.A(n_122),
.Y(n_164)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_164),
.Y(n_222)
);

BUFx2_ASAP7_75t_L g166 ( 
.A(n_137),
.Y(n_166)
);

INVx11_ASAP7_75t_L g202 ( 
.A(n_166),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_96),
.B(n_74),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_168),
.B(n_172),
.Y(n_205)
);

OAI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_169),
.A2(n_142),
.B1(n_119),
.B2(n_6),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_115),
.A2(n_22),
.B(n_37),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_170),
.A2(n_111),
.B(n_138),
.Y(n_204)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_148),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_171),
.B(n_184),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_143),
.B(n_33),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_114),
.B(n_33),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_173),
.B(n_176),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_116),
.B(n_28),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_174),
.B(n_175),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_118),
.B(n_26),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_121),
.B(n_70),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_139),
.B(n_149),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_177),
.B(n_198),
.Y(n_209)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_146),
.Y(n_178)
);

INVx6_ASAP7_75t_L g237 ( 
.A(n_178),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_99),
.B(n_93),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_179),
.B(n_181),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_180),
.B(n_186),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_120),
.B(n_94),
.Y(n_181)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_127),
.Y(n_184)
);

INVx1_ASAP7_75t_SL g185 ( 
.A(n_124),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g235 ( 
.A(n_185),
.B(n_188),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_102),
.B(n_58),
.Y(n_186)
);

INVx8_ASAP7_75t_L g187 ( 
.A(n_108),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g232 ( 
.A1(n_187),
.A2(n_191),
.B1(n_192),
.B2(n_194),
.Y(n_232)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_135),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_135),
.Y(n_189)
);

AND2x2_ASAP7_75t_L g236 ( 
.A(n_189),
.B(n_190),
.Y(n_236)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_141),
.Y(n_190)
);

INVx6_ASAP7_75t_L g191 ( 
.A(n_108),
.Y(n_191)
);

INVx5_ASAP7_75t_L g192 ( 
.A(n_134),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_102),
.B(n_4),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_193),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_112),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_112),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_195),
.A2(n_106),
.B1(n_109),
.B2(n_129),
.Y(n_208)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_117),
.B(n_4),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_196),
.B(n_100),
.C(n_136),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_197),
.A2(n_129),
.B1(n_109),
.B2(n_106),
.Y(n_215)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_141),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_204),
.B(n_207),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_208),
.Y(n_255)
);

AND2x2_ASAP7_75t_SL g210 ( 
.A(n_177),
.B(n_153),
.Y(n_210)
);

MAJx2_ASAP7_75t_L g268 ( 
.A(n_210),
.B(n_211),
.C(n_188),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_151),
.B(n_104),
.C(n_144),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_212),
.B(n_214),
.C(n_220),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_183),
.A2(n_117),
.B1(n_111),
.B2(n_145),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_213),
.A2(n_229),
.B(n_170),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_160),
.B(n_144),
.C(n_146),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_215),
.A2(n_233),
.B1(n_196),
.B2(n_166),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_217),
.A2(n_164),
.B1(n_156),
.B2(n_185),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_174),
.B(n_142),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_175),
.B(n_4),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_227),
.B(n_228),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_152),
.B(n_5),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_196),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_197),
.A2(n_157),
.B1(n_158),
.B2(n_169),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_231),
.B(n_223),
.Y(n_247)
);

OAI22x1_ASAP7_75t_SL g233 ( 
.A1(n_157),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_210),
.B(n_156),
.C(n_184),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_240),
.B(n_250),
.C(n_221),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_205),
.B(n_165),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_241),
.B(n_260),
.Y(n_300)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_199),
.Y(n_242)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_242),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_243),
.A2(n_265),
.B1(n_267),
.B2(n_231),
.Y(n_283)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_199),
.Y(n_244)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_244),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_236),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_245),
.B(n_252),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_247),
.A2(n_224),
.B1(n_233),
.B2(n_219),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_249),
.A2(n_213),
.B1(n_216),
.B2(n_204),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_210),
.B(n_167),
.C(n_171),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_230),
.Y(n_251)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_251),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_236),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_236),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_253),
.B(n_254),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_203),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_256),
.A2(n_235),
.B1(n_226),
.B2(n_222),
.Y(n_303)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_230),
.Y(n_257)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_257),
.Y(n_298)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_206),
.Y(n_258)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_258),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_201),
.B(n_161),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_259),
.B(n_262),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_201),
.B(n_167),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_200),
.B(n_182),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_261),
.B(n_263),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_220),
.B(n_227),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_200),
.B(n_182),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_206),
.Y(n_264)
);

INVx1_ASAP7_75t_SL g295 ( 
.A(n_264),
.Y(n_295)
);

AOI22xp33_ASAP7_75t_L g265 ( 
.A1(n_223),
.A2(n_158),
.B1(n_187),
.B2(n_162),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_209),
.B(n_198),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_266),
.B(n_269),
.Y(n_293)
);

AOI22xp33_ASAP7_75t_L g267 ( 
.A1(n_224),
.A2(n_158),
.B1(n_190),
.B2(n_189),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_268),
.B(n_235),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_209),
.B(n_178),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_206),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_270),
.B(n_235),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_234),
.B(n_192),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_271),
.B(n_273),
.Y(n_291)
);

AOI22xp33_ASAP7_75t_SL g272 ( 
.A1(n_216),
.A2(n_159),
.B1(n_191),
.B2(n_195),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_272),
.A2(n_232),
.B(n_208),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_234),
.B(n_159),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_239),
.B(n_218),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_274),
.B(n_280),
.C(n_282),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_SL g309 ( 
.A(n_275),
.B(n_288),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_276),
.A2(n_283),
.B1(n_290),
.B2(n_299),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_278),
.A2(n_303),
.B(n_305),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_268),
.B(n_211),
.C(n_221),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_268),
.B(n_214),
.C(n_212),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g314 ( 
.A1(n_285),
.A2(n_261),
.B1(n_263),
.B2(n_249),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_239),
.B(n_228),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_248),
.A2(n_219),
.B(n_207),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g307 ( 
.A(n_289),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_247),
.A2(n_267),
.B1(n_265),
.B2(n_243),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_271),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_292),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_273),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_297),
.B(n_302),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_266),
.A2(n_215),
.B1(n_238),
.B2(n_229),
.Y(n_299)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_301),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_269),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_304),
.B(n_240),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_248),
.A2(n_202),
.B(n_225),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_259),
.B(n_226),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_306),
.B(n_264),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_281),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_308),
.B(n_324),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_314),
.A2(n_334),
.B1(n_295),
.B2(n_299),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_283),
.A2(n_239),
.B1(n_255),
.B2(n_250),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_L g359 ( 
.A1(n_315),
.A2(n_329),
.B1(n_295),
.B2(n_285),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_316),
.B(n_319),
.C(n_331),
.Y(n_348)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_277),
.Y(n_318)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_318),
.Y(n_353)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_280),
.B(n_240),
.Y(n_319)
);

A2O1A1O1Ixp25_ASAP7_75t_L g320 ( 
.A1(n_289),
.A2(n_260),
.B(n_262),
.C(n_246),
.D(n_250),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_SL g343 ( 
.A1(n_320),
.A2(n_332),
.B(n_303),
.Y(n_343)
);

OA21x2_ASAP7_75t_SL g321 ( 
.A1(n_281),
.A2(n_246),
.B(n_254),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_SL g337 ( 
.A(n_321),
.B(n_323),
.Y(n_337)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_277),
.Y(n_322)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_322),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_300),
.B(n_241),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_284),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_284),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_325),
.B(n_326),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_279),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_296),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_327),
.B(n_328),
.Y(n_361)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_296),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_290),
.A2(n_245),
.B1(n_252),
.B2(n_253),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_274),
.B(n_258),
.Y(n_331)
);

AOI21xp5_ASAP7_75t_L g332 ( 
.A1(n_305),
.A2(n_272),
.B(n_256),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_333),
.B(n_336),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_302),
.A2(n_270),
.B1(n_257),
.B2(n_251),
.Y(n_334)
);

BUFx2_ASAP7_75t_L g335 ( 
.A(n_294),
.Y(n_335)
);

INVxp67_ASAP7_75t_L g341 ( 
.A(n_335),
.Y(n_341)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_298),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_319),
.B(n_282),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g368 ( 
.A(n_339),
.B(n_340),
.Y(n_368)
);

XOR2xp5_ASAP7_75t_L g340 ( 
.A(n_309),
.B(n_304),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_330),
.B(n_275),
.Y(n_342)
);

XOR2xp5_ASAP7_75t_L g371 ( 
.A(n_342),
.B(n_354),
.Y(n_371)
);

AOI21xp5_ASAP7_75t_L g372 ( 
.A1(n_343),
.A2(n_350),
.B(n_312),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_344),
.A2(n_345),
.B1(n_352),
.B2(n_294),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_307),
.A2(n_276),
.B1(n_292),
.B2(n_288),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_310),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g364 ( 
.A(n_346),
.B(n_356),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_330),
.B(n_309),
.C(n_316),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_349),
.B(n_355),
.C(n_291),
.Y(n_369)
);

OAI21xp5_ASAP7_75t_SL g350 ( 
.A1(n_312),
.A2(n_278),
.B(n_287),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_307),
.A2(n_293),
.B1(n_297),
.B2(n_279),
.Y(n_352)
);

XOR2xp5_ASAP7_75t_L g354 ( 
.A(n_331),
.B(n_286),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_315),
.B(n_286),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_310),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_311),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_SL g376 ( 
.A(n_357),
.B(n_359),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_333),
.B(n_293),
.Y(n_360)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_360),
.Y(n_363)
);

CKINVDCx16_ASAP7_75t_R g362 ( 
.A(n_329),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_362),
.B(n_313),
.Y(n_383)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_338),
.Y(n_365)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_365),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_351),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_SL g391 ( 
.A(n_366),
.B(n_374),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_L g367 ( 
.A(n_342),
.B(n_291),
.Y(n_367)
);

XOR2xp5_ASAP7_75t_L g392 ( 
.A(n_367),
.B(n_372),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_369),
.B(n_379),
.C(n_381),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_338),
.B(n_334),
.Y(n_370)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_370),
.Y(n_397)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_358),
.Y(n_373)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_373),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_337),
.B(n_287),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_361),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_375),
.B(n_378),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_360),
.B(n_306),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_377),
.Y(n_399)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_347),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_339),
.B(n_317),
.C(n_313),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_347),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_L g394 ( 
.A1(n_380),
.A2(n_378),
.B1(n_335),
.B2(n_353),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_348),
.B(n_355),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_352),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_382),
.B(n_383),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_SL g384 ( 
.A(n_349),
.B(n_317),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_384),
.B(n_343),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_385),
.A2(n_354),
.B1(n_344),
.B2(n_345),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_381),
.B(n_348),
.C(n_340),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_387),
.B(n_390),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_371),
.B(n_369),
.C(n_368),
.Y(n_390)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_393),
.Y(n_404)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_394),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_SL g413 ( 
.A(n_396),
.B(n_398),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_364),
.B(n_353),
.Y(n_398)
);

BUFx2_ASAP7_75t_L g400 ( 
.A(n_373),
.Y(n_400)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_400),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_SL g402 ( 
.A1(n_370),
.A2(n_365),
.B1(n_376),
.B2(n_363),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_402),
.A2(n_403),
.B1(n_385),
.B2(n_379),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_SL g403 ( 
.A1(n_363),
.A2(n_332),
.B1(n_350),
.B2(n_320),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_SL g424 ( 
.A1(n_405),
.A2(n_407),
.B1(n_408),
.B2(n_393),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_386),
.B(n_371),
.C(n_368),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_406),
.B(n_415),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_L g407 ( 
.A1(n_402),
.A2(n_377),
.B1(n_380),
.B2(n_375),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_397),
.A2(n_372),
.B1(n_341),
.B2(n_322),
.Y(n_408)
);

XOR2xp5_ASAP7_75t_L g410 ( 
.A(n_392),
.B(n_367),
.Y(n_410)
);

XOR2xp5_ASAP7_75t_L g418 ( 
.A(n_410),
.B(n_387),
.Y(n_418)
);

A2O1A1Ixp33_ASAP7_75t_SL g412 ( 
.A1(n_403),
.A2(n_336),
.B(n_318),
.C(n_341),
.Y(n_412)
);

NAND2x1p5_ASAP7_75t_R g421 ( 
.A(n_412),
.B(n_388),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_SL g414 ( 
.A(n_391),
.B(n_244),
.Y(n_414)
);

CKINVDCx14_ASAP7_75t_R g420 ( 
.A(n_414),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_386),
.B(n_301),
.C(n_298),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_SL g417 ( 
.A(n_401),
.B(n_242),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_417),
.B(n_401),
.Y(n_423)
);

AND2x2_ASAP7_75t_L g433 ( 
.A(n_418),
.B(n_412),
.Y(n_433)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_404),
.A2(n_397),
.B1(n_395),
.B2(n_399),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_SL g437 ( 
.A1(n_419),
.A2(n_427),
.B1(n_225),
.B2(n_194),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_421),
.B(n_423),
.Y(n_431)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_416),
.Y(n_422)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_422),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_424),
.B(n_428),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_SL g425 ( 
.A1(n_407),
.A2(n_389),
.B1(n_409),
.B2(n_395),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_SL g439 ( 
.A(n_425),
.B(n_426),
.Y(n_439)
);

OAI21xp5_ASAP7_75t_SL g426 ( 
.A1(n_408),
.A2(n_399),
.B(n_388),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_413),
.A2(n_400),
.B1(n_392),
.B2(n_415),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_SL g428 ( 
.A1(n_412),
.A2(n_390),
.B1(n_406),
.B2(n_411),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_410),
.B(n_222),
.C(n_202),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_430),
.B(n_237),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_SL g447 ( 
.A(n_433),
.B(n_437),
.Y(n_447)
);

AND2x2_ASAP7_75t_L g434 ( 
.A(n_418),
.B(n_412),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_434),
.B(n_435),
.Y(n_442)
);

AND2x2_ASAP7_75t_L g435 ( 
.A(n_429),
.B(n_237),
.Y(n_435)
);

INVxp67_ASAP7_75t_L g443 ( 
.A(n_436),
.Y(n_443)
);

OAI21xp5_ASAP7_75t_SL g440 ( 
.A1(n_427),
.A2(n_8),
.B(n_10),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_SL g446 ( 
.A(n_440),
.B(n_426),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_432),
.B(n_420),
.Y(n_441)
);

AOI21xp5_ASAP7_75t_L g448 ( 
.A1(n_441),
.A2(n_444),
.B(n_445),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_438),
.B(n_428),
.C(n_424),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_439),
.B(n_425),
.Y(n_445)
);

NOR3xp33_ASAP7_75t_L g450 ( 
.A(n_446),
.B(n_436),
.C(n_421),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_442),
.B(n_439),
.C(n_431),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_449),
.B(n_451),
.C(n_443),
.Y(n_452)
);

INVxp67_ASAP7_75t_L g453 ( 
.A(n_450),
.Y(n_453)
);

OAI21xp5_ASAP7_75t_SL g451 ( 
.A1(n_447),
.A2(n_419),
.B(n_430),
.Y(n_451)
);

XOR2xp5_ASAP7_75t_L g455 ( 
.A(n_452),
.B(n_454),
.Y(n_455)
);

OAI21xp5_ASAP7_75t_SL g454 ( 
.A1(n_448),
.A2(n_443),
.B(n_11),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_453),
.B(n_8),
.C(n_11),
.Y(n_456)
);

BUFx24_ASAP7_75t_SL g457 ( 
.A(n_456),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_L g458 ( 
.A1(n_457),
.A2(n_12),
.B1(n_455),
.B2(n_453),
.Y(n_458)
);

XOR2xp5_ASAP7_75t_L g459 ( 
.A(n_458),
.B(n_12),
.Y(n_459)
);


endmodule