module real_jpeg_20805_n_18 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_290, n_11, n_14, n_7, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_290;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_18;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_286;
wire n_288;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_194;
wire n_153;
wire n_104;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_281;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_237;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_285;
wire n_112;
wire n_42;
wire n_268;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_137;
wire n_31;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_258;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_277;
wire n_226;
wire n_185;
wire n_125;
wire n_240;
wire n_209;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_128;
wire n_167;
wire n_213;
wire n_179;
wire n_202;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_283;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_269;
wire n_96;
wire n_253;
wire n_273;
wire n_89;

AOI22xp33_ASAP7_75t_L g132 ( 
.A1(n_0),
.A2(n_28),
.B1(n_37),
.B2(n_133),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_0),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_0),
.A2(n_66),
.B1(n_67),
.B2(n_133),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_0),
.A2(n_45),
.B1(n_46),
.B2(n_133),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_0),
.A2(n_32),
.B1(n_33),
.B2(n_133),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_1),
.A2(n_66),
.B1(n_67),
.B2(n_91),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_1),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_1),
.A2(n_32),
.B1(n_33),
.B2(n_91),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_1),
.A2(n_28),
.B1(n_37),
.B2(n_91),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_L g211 ( 
.A1(n_1),
.A2(n_45),
.B1(n_46),
.B2(n_91),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_2),
.A2(n_32),
.B1(n_33),
.B2(n_50),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_2),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_2),
.A2(n_45),
.B1(n_46),
.B2(n_50),
.Y(n_85)
);

BUFx16f_ASAP7_75t_L g66 ( 
.A(n_3),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_4),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_4),
.B(n_72),
.Y(n_165)
);

AOI21xp33_ASAP7_75t_L g185 ( 
.A1(n_4),
.A2(n_16),
.B(n_45),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_4),
.A2(n_32),
.B1(n_33),
.B2(n_137),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_4),
.A2(n_81),
.B1(n_82),
.B2(n_194),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_4),
.B(n_59),
.Y(n_206)
);

AOI21xp33_ASAP7_75t_L g223 ( 
.A1(n_4),
.A2(n_37),
.B(n_224),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_5),
.A2(n_65),
.B1(n_66),
.B2(n_67),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_5),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_5),
.A2(n_28),
.B1(n_37),
.B2(n_65),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_5),
.A2(n_32),
.B1(n_33),
.B2(n_65),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_5),
.A2(n_45),
.B1(n_46),
.B2(n_65),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_6),
.A2(n_28),
.B1(n_37),
.B2(n_39),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_6),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_6),
.A2(n_32),
.B1(n_33),
.B2(n_39),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_6),
.A2(n_39),
.B1(n_45),
.B2(n_46),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_7),
.A2(n_32),
.B1(n_33),
.B2(n_48),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_7),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_7),
.A2(n_28),
.B1(n_37),
.B2(n_48),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_7),
.A2(n_45),
.B1(n_46),
.B2(n_48),
.Y(n_102)
);

BUFx10_ASAP7_75t_L g45 ( 
.A(n_8),
.Y(n_45)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_9),
.Y(n_82)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_9),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_10),
.A2(n_66),
.B1(n_67),
.B2(n_112),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_10),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_10),
.A2(n_28),
.B1(n_37),
.B2(n_112),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_10),
.A2(n_45),
.B1(n_46),
.B2(n_112),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_10),
.A2(n_32),
.B1(n_33),
.B2(n_112),
.Y(n_227)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_12),
.A2(n_66),
.B1(n_67),
.B2(n_139),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_12),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_12),
.A2(n_28),
.B1(n_37),
.B2(n_139),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_12),
.A2(n_32),
.B1(n_33),
.B2(n_139),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_12),
.A2(n_45),
.B1(n_46),
.B2(n_139),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_13),
.A2(n_28),
.B1(n_36),
.B2(n_37),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_13),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_13),
.A2(n_36),
.B1(n_66),
.B2(n_67),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_13),
.A2(n_32),
.B1(n_33),
.B2(n_36),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_13),
.A2(n_36),
.B1(n_45),
.B2(n_46),
.Y(n_153)
);

INVx13_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_14),
.A2(n_29),
.B1(n_32),
.B2(n_33),
.Y(n_31)
);

OAI32xp33_ASAP7_75t_L g218 ( 
.A1(n_14),
.A2(n_33),
.A3(n_37),
.B1(n_219),
.B2(n_220),
.Y(n_218)
);

INVx13_ASAP7_75t_L g70 ( 
.A(n_15),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_15),
.A2(n_28),
.B1(n_37),
.B2(n_70),
.Y(n_72)
);

OAI22xp33_ASAP7_75t_L g42 ( 
.A1(n_16),
.A2(n_32),
.B1(n_33),
.B2(n_43),
.Y(n_42)
);

INVx6_ASAP7_75t_SL g43 ( 
.A(n_16),
.Y(n_43)
);

OA22x2_ASAP7_75t_L g44 ( 
.A1(n_16),
.A2(n_43),
.B1(n_45),
.B2(n_46),
.Y(n_44)
);

BUFx3_ASAP7_75t_SL g33 ( 
.A(n_17),
.Y(n_33)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_115),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_113),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_92),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_21),
.B(n_92),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_77),
.B2(n_78),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_51),
.B2(n_52),
.Y(n_23)
);

CKINVDCx14_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_25),
.A2(n_26),
.B(n_40),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_40),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_27),
.A2(n_31),
.B1(n_34),
.B2(n_38),
.Y(n_26)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_27),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_27),
.A2(n_31),
.B1(n_132),
.B2(n_134),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_27),
.A2(n_31),
.B1(n_134),
.B2(n_147),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_27),
.A2(n_31),
.B1(n_163),
.B2(n_223),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_27),
.A2(n_31),
.B1(n_108),
.B2(n_147),
.Y(n_266)
);

A2O1A1Ixp33_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_29),
.B(n_30),
.C(n_31),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_28),
.B(n_29),
.Y(n_30)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_28),
.A2(n_71),
.B1(n_136),
.B2(n_151),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_28),
.B(n_137),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_29),
.B(n_32),
.Y(n_219)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_31),
.Y(n_59)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

A2O1A1Ixp33_ASAP7_75t_L g184 ( 
.A1(n_33),
.A2(n_43),
.B(n_137),
.C(n_185),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_35),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_35),
.A2(n_57),
.B1(n_59),
.B2(n_107),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_37),
.B(n_70),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_38),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_41),
.A2(n_44),
.B1(n_47),
.B2(n_49),
.Y(n_40)
);

AOI21xp5_ASAP7_75t_SL g61 ( 
.A1(n_41),
.A2(n_44),
.B(n_49),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_41),
.A2(n_44),
.B1(n_47),
.B2(n_87),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_41),
.A2(n_44),
.B1(n_87),
.B2(n_105),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_41),
.A2(n_44),
.B1(n_105),
.B2(n_125),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_41),
.A2(n_44),
.B1(n_125),
.B2(n_129),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_41),
.A2(n_44),
.B1(n_188),
.B2(n_189),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_41),
.A2(n_44),
.B1(n_189),
.B2(n_209),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_41),
.A2(n_44),
.B1(n_209),
.B2(n_227),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_41),
.A2(n_44),
.B1(n_129),
.B2(n_227),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_44),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_44),
.B(n_137),
.Y(n_192)
);

INVx13_ASAP7_75t_L g46 ( 
.A(n_45),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_45),
.B(n_82),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_46),
.B(n_197),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_52),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_53),
.A2(n_62),
.B1(n_75),
.B2(n_76),
.Y(n_52)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_53),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_54),
.A2(n_55),
.B1(n_60),
.B2(n_61),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_56),
.A2(n_57),
.B1(n_58),
.B2(n_59),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_57),
.A2(n_59),
.B1(n_162),
.B2(n_164),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_61),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_62),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_63),
.A2(n_68),
.B1(n_73),
.B2(n_74),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_64),
.A2(n_69),
.B1(n_72),
.B2(n_89),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_66),
.Y(n_67)
);

O2A1O1Ixp33_ASAP7_75t_L g69 ( 
.A1(n_66),
.A2(n_70),
.B(n_71),
.C(n_72),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_66),
.B(n_70),
.Y(n_71)
);

HAxp5_ASAP7_75t_SL g136 ( 
.A(n_66),
.B(n_137),
.CON(n_136),
.SN(n_136)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_68),
.A2(n_74),
.B1(n_90),
.B2(n_111),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_68),
.A2(n_74),
.B1(n_144),
.B2(n_145),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_68),
.A2(n_74),
.B1(n_111),
.B2(n_145),
.Y(n_265)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_69),
.A2(n_72),
.B1(n_136),
.B2(n_138),
.Y(n_135)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_72),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_78),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_79),
.A2(n_80),
.B1(n_88),
.B2(n_290),
.Y(n_78)
);

XOR2xp5_ASAP7_75t_L g93 ( 
.A(n_79),
.B(n_94),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_86),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_80),
.A2(n_88),
.B1(n_95),
.B2(n_96),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_80),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_80),
.A2(n_86),
.B1(n_96),
.B2(n_280),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_83),
.B(n_85),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_81),
.A2(n_85),
.B1(n_102),
.B2(n_103),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_81),
.A2(n_102),
.B1(n_103),
.B2(n_123),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_81),
.A2(n_103),
.B1(n_123),
.B2(n_153),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_81),
.A2(n_82),
.B1(n_153),
.B2(n_168),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_81),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_81),
.A2(n_82),
.B1(n_179),
.B2(n_194),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_81),
.A2(n_83),
.B1(n_181),
.B2(n_211),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_81),
.A2(n_82),
.B1(n_168),
.B2(n_211),
.Y(n_217)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_82),
.Y(n_84)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_84),
.A2(n_177),
.B1(n_178),
.B2(n_180),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_86),
.Y(n_280)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_88),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_90),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_97),
.C(n_98),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_93),
.B(n_97),
.Y(n_287)
);

AOI22xp33_ASAP7_75t_SL g285 ( 
.A1(n_98),
.A2(n_99),
.B1(n_286),
.B2(n_287),
.Y(n_285)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_99),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_106),
.C(n_109),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_100),
.B(n_276),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_104),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_101),
.B(n_104),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_103),
.B(n_137),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_106),
.A2(n_109),
.B1(n_110),
.B2(n_277),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_106),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_110),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_116),
.A2(n_283),
.B(n_288),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g116 ( 
.A1(n_117),
.A2(n_270),
.B(n_282),
.Y(n_116)
);

O2A1O1Ixp33_ASAP7_75t_SL g117 ( 
.A1(n_118),
.A2(n_169),
.B(n_252),
.C(n_269),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_154),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_119),
.B(n_154),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_140),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_126),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_121),
.B(n_126),
.C(n_140),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_124),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_122),
.B(n_124),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_130),
.C(n_135),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_127),
.A2(n_128),
.B1(n_130),
.B2(n_131),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_128),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_132),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_SL g155 ( 
.A(n_135),
.B(n_156),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_138),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_SL g140 ( 
.A(n_141),
.B(n_149),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_142),
.A2(n_143),
.B1(n_146),
.B2(n_148),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_142),
.B(n_148),
.C(n_149),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_143),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_146),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_152),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_150),
.B(n_152),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_157),
.C(n_159),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_155),
.B(n_249),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_157),
.A2(n_158),
.B1(n_159),
.B2(n_160),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_158),
.Y(n_157)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_165),
.C(n_166),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_161),
.B(n_237),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_165),
.A2(n_166),
.B1(n_167),
.B2(n_238),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_165),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_167),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_170),
.B(n_251),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_171),
.A2(n_246),
.B(n_250),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_172),
.A2(n_232),
.B(n_245),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_173),
.A2(n_213),
.B(n_231),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_174),
.A2(n_201),
.B(n_212),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_175),
.A2(n_190),
.B(n_200),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_182),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_176),
.B(n_182),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_181),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_183),
.A2(n_184),
.B1(n_186),
.B2(n_187),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_184),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_184),
.B(n_186),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_187),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_191),
.A2(n_195),
.B(n_199),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_193),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_192),
.B(n_193),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_198),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_203),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_202),
.B(n_203),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_210),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_205),
.A2(n_206),
.B1(n_207),
.B2(n_208),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_205),
.B(n_208),
.C(n_210),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_206),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_208),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_215),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_214),
.B(n_215),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_216),
.A2(n_221),
.B1(n_229),
.B2(n_230),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_216),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_218),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_217),
.B(n_218),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_220),
.Y(n_224)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_221),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_222),
.A2(n_225),
.B1(n_226),
.B2(n_228),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_222),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_225),
.B(n_228),
.C(n_229),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_226),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_234),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_233),
.B(n_234),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_235),
.A2(n_236),
.B1(n_239),
.B2(n_240),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_235),
.B(n_242),
.C(n_243),
.Y(n_247)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_241),
.A2(n_242),
.B1(n_243),
.B2(n_244),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_241),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_242),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_248),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_247),
.B(n_248),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_254),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_253),
.B(n_254),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_255),
.A2(n_256),
.B1(n_257),
.B2(n_268),
.Y(n_254)
);

CKINVDCx14_ASAP7_75t_R g268 ( 
.A(n_255),
.Y(n_268)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_258),
.A2(n_259),
.B1(n_260),
.B2(n_261),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_258),
.B(n_261),
.C(n_268),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_259),
.Y(n_258)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_263),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_262),
.B(n_264),
.C(n_267),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_264),
.A2(n_265),
.B1(n_266),
.B2(n_267),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_265),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_266),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_272),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_271),
.B(n_272),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_281),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_274),
.A2(n_275),
.B1(n_278),
.B2(n_279),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_274),
.B(n_279),
.C(n_281),
.Y(n_284)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

CKINVDCx16_ASAP7_75t_R g278 ( 
.A(n_279),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_285),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g288 ( 
.A(n_284),
.B(n_285),
.Y(n_288)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);


endmodule