module fake_jpeg_30319_n_510 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_510);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_510;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_14),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx2_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx8_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_15),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_1),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_12),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

BUFx16f_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

OR2x2_ASAP7_75t_L g36 ( 
.A(n_1),
.B(n_8),
.Y(n_36)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_2),
.Y(n_46)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_10),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_10),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_4),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_2),
.Y(n_50)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_16),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_36),
.B(n_16),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_52),
.B(n_55),
.Y(n_102)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

BUFx8_ASAP7_75t_L g145 ( 
.A(n_53),
.Y(n_145)
);

BUFx10_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

INVxp33_ASAP7_75t_L g129 ( 
.A(n_54),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_35),
.Y(n_55)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_32),
.Y(n_56)
);

INVx11_ASAP7_75t_L g110 ( 
.A(n_56),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_26),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_57),
.Y(n_108)
);

INVx4_ASAP7_75t_SL g58 ( 
.A(n_34),
.Y(n_58)
);

CKINVDCx14_ASAP7_75t_R g147 ( 
.A(n_58),
.Y(n_147)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_59),
.Y(n_112)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_60),
.Y(n_124)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_61),
.Y(n_114)
);

BUFx4f_ASAP7_75t_L g62 ( 
.A(n_34),
.Y(n_62)
);

HB1xp67_ASAP7_75t_L g118 ( 
.A(n_62),
.Y(n_118)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_63),
.Y(n_119)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_32),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_64),
.Y(n_141)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_65),
.Y(n_125)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_66),
.Y(n_107)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_21),
.Y(n_67)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_67),
.Y(n_139)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_26),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_68),
.Y(n_152)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_21),
.Y(n_69)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_69),
.Y(n_149)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_21),
.Y(n_70)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_70),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_26),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_71),
.Y(n_158)
);

BUFx8_ASAP7_75t_L g72 ( 
.A(n_35),
.Y(n_72)
);

CKINVDCx9p33_ASAP7_75t_R g132 ( 
.A(n_72),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_20),
.B(n_15),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_73),
.B(n_75),
.Y(n_111)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_26),
.Y(n_74)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_74),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_35),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_36),
.B(n_15),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_76),
.B(n_89),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_18),
.Y(n_77)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_77),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_18),
.Y(n_78)
);

INVx6_ASAP7_75t_L g144 ( 
.A(n_78),
.Y(n_144)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_51),
.Y(n_79)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_79),
.Y(n_157)
);

BUFx10_ASAP7_75t_L g80 ( 
.A(n_20),
.Y(n_80)
);

INVx1_ASAP7_75t_SL g136 ( 
.A(n_80),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_18),
.Y(n_81)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_81),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_27),
.Y(n_82)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_82),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_32),
.Y(n_83)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_83),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_27),
.Y(n_84)
);

INVx5_ASAP7_75t_L g143 ( 
.A(n_84),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_27),
.Y(n_85)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_85),
.Y(n_115)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_51),
.Y(n_86)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_86),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_37),
.Y(n_87)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_87),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_29),
.Y(n_88)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_88),
.Y(n_146)
);

INVx2_ASAP7_75t_SL g89 ( 
.A(n_36),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_37),
.Y(n_90)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_90),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_29),
.Y(n_91)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_91),
.Y(n_151)
);

INVx11_ASAP7_75t_L g92 ( 
.A(n_29),
.Y(n_92)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_92),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_30),
.Y(n_93)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_93),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_47),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_94),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_30),
.Y(n_95)
);

BUFx12f_ASAP7_75t_L g155 ( 
.A(n_95),
.Y(n_155)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_30),
.Y(n_96)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_96),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_17),
.B(n_13),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_97),
.B(n_23),
.Y(n_117)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_19),
.Y(n_98)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_98),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_19),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_99),
.B(n_20),
.Y(n_156)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_28),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_100),
.B(n_20),
.Y(n_122)
);

BUFx2_ASAP7_75t_R g104 ( 
.A(n_62),
.Y(n_104)
);

CKINVDCx14_ASAP7_75t_R g192 ( 
.A(n_104),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_96),
.A2(n_19),
.B1(n_40),
.B2(n_44),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g171 ( 
.A1(n_105),
.A2(n_95),
.B1(n_93),
.B2(n_88),
.Y(n_171)
);

AND2x6_ASAP7_75t_L g106 ( 
.A(n_89),
.B(n_23),
.Y(n_106)
);

AOI21xp33_ASAP7_75t_L g164 ( 
.A1(n_106),
.A2(n_80),
.B(n_46),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_117),
.B(n_142),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_122),
.B(n_156),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_53),
.B(n_17),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_123),
.B(n_126),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_73),
.B(n_31),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_53),
.B(n_31),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_127),
.B(n_135),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_77),
.A2(n_38),
.B1(n_44),
.B2(n_45),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_133),
.A2(n_68),
.B1(n_74),
.B2(n_91),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_56),
.A2(n_45),
.B1(n_48),
.B2(n_24),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_134),
.A2(n_48),
.B(n_25),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_58),
.B(n_22),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_80),
.B(n_22),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_72),
.B(n_24),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_150),
.B(n_43),
.Y(n_190)
);

INVx6_ASAP7_75t_SL g153 ( 
.A(n_54),
.Y(n_153)
);

INVx13_ASAP7_75t_L g174 ( 
.A(n_153),
.Y(n_174)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_124),
.Y(n_159)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_159),
.Y(n_220)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_120),
.Y(n_160)
);

INVx4_ASAP7_75t_L g235 ( 
.A(n_160),
.Y(n_235)
);

CKINVDCx16_ASAP7_75t_R g236 ( 
.A(n_162),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_163),
.A2(n_171),
.B1(n_185),
.B2(n_105),
.Y(n_244)
);

XNOR2x1_ASAP7_75t_SL g230 ( 
.A(n_164),
.B(n_20),
.Y(n_230)
);

INVx5_ASAP7_75t_L g165 ( 
.A(n_110),
.Y(n_165)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_165),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_147),
.A2(n_83),
.B1(n_90),
.B2(n_87),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_166),
.A2(n_196),
.B1(n_205),
.B2(n_206),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_102),
.B(n_25),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_167),
.B(n_168),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_113),
.B(n_41),
.Y(n_168)
);

HB1xp67_ASAP7_75t_L g169 ( 
.A(n_107),
.Y(n_169)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_169),
.Y(n_245)
);

HB1xp67_ASAP7_75t_L g170 ( 
.A(n_140),
.Y(n_170)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_170),
.Y(n_253)
);

AND2x4_ASAP7_75t_L g172 ( 
.A(n_106),
.B(n_54),
.Y(n_172)
);

AND2x2_ASAP7_75t_SL g237 ( 
.A(n_172),
.B(n_44),
.Y(n_237)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_112),
.Y(n_175)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_175),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_114),
.B(n_39),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_177),
.B(n_186),
.Y(n_228)
);

INVx5_ASAP7_75t_L g178 ( 
.A(n_110),
.Y(n_178)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_178),
.Y(n_222)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_120),
.Y(n_179)
);

INVx3_ASAP7_75t_L g238 ( 
.A(n_179),
.Y(n_238)
);

BUFx10_ASAP7_75t_L g181 ( 
.A(n_132),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_181),
.Y(n_242)
);

INVx6_ASAP7_75t_L g182 ( 
.A(n_108),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_182),
.Y(n_224)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_125),
.Y(n_183)
);

BUFx3_ASAP7_75t_L g232 ( 
.A(n_183),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_108),
.Y(n_184)
);

INVx8_ASAP7_75t_L g217 ( 
.A(n_184),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_111),
.A2(n_85),
.B1(n_84),
.B2(n_82),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_147),
.B(n_41),
.Y(n_186)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_139),
.Y(n_187)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_187),
.Y(n_223)
);

OA22x2_ASAP7_75t_SL g188 ( 
.A1(n_149),
.A2(n_81),
.B1(n_78),
.B2(n_71),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_188),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_158),
.Y(n_189)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_189),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_190),
.B(n_198),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_158),
.Y(n_191)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_191),
.Y(n_226)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_137),
.Y(n_193)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_193),
.Y(n_239)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_101),
.Y(n_194)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_194),
.Y(n_243)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_121),
.Y(n_195)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_195),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_128),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_157),
.B(n_39),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_197),
.B(n_199),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_129),
.B(n_43),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_154),
.B(n_50),
.Y(n_199)
);

BUFx12f_ASAP7_75t_L g200 ( 
.A(n_116),
.Y(n_200)
);

BUFx16f_ASAP7_75t_L g219 ( 
.A(n_200),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_129),
.B(n_118),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_201),
.B(n_203),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_131),
.B(n_50),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_202),
.B(n_208),
.Y(n_218)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_130),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_118),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_204),
.B(n_207),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_128),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_109),
.A2(n_64),
.B1(n_143),
.B2(n_19),
.Y(n_206)
);

INVx6_ASAP7_75t_L g207 ( 
.A(n_144),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_144),
.B(n_46),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_138),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_209),
.B(n_119),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_155),
.A2(n_138),
.B1(n_121),
.B2(n_115),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g247 ( 
.A1(n_210),
.A2(n_136),
.B1(n_155),
.B2(n_141),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_188),
.A2(n_103),
.B1(n_148),
.B2(n_151),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_215),
.A2(n_233),
.B1(n_248),
.B2(n_251),
.Y(n_270)
);

OR2x2_ASAP7_75t_L g221 ( 
.A(n_161),
.B(n_136),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_221),
.B(n_237),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_230),
.B(n_174),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_188),
.A2(n_103),
.B1(n_148),
.B2(n_146),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_172),
.B(n_152),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_240),
.B(n_241),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_172),
.B(n_152),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_244),
.A2(n_207),
.B1(n_182),
.B2(n_196),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_247),
.A2(n_210),
.B1(n_192),
.B2(n_206),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_L g248 ( 
.A1(n_171),
.A2(n_155),
.B1(n_119),
.B2(n_57),
.Y(n_248)
);

CKINVDCx16_ASAP7_75t_R g264 ( 
.A(n_249),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_180),
.B(n_176),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_250),
.B(n_173),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_172),
.A2(n_141),
.B1(n_38),
.B2(n_40),
.Y(n_251)
);

AO22x1_ASAP7_75t_L g252 ( 
.A1(n_166),
.A2(n_94),
.B1(n_145),
.B2(n_33),
.Y(n_252)
);

AO22x1_ASAP7_75t_SL g289 ( 
.A1(n_252),
.A2(n_145),
.B1(n_181),
.B2(n_33),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_254),
.A2(n_289),
.B1(n_243),
.B2(n_242),
.Y(n_316)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_217),
.Y(n_256)
);

BUFx2_ASAP7_75t_L g321 ( 
.A(n_256),
.Y(n_321)
);

INVx3_ASAP7_75t_L g257 ( 
.A(n_217),
.Y(n_257)
);

INVx3_ASAP7_75t_L g298 ( 
.A(n_257),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_258),
.B(n_267),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_212),
.A2(n_194),
.B1(n_160),
.B2(n_195),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_259),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_260),
.A2(n_226),
.B1(n_223),
.B2(n_245),
.Y(n_324)
);

AOI22xp33_ASAP7_75t_L g261 ( 
.A1(n_212),
.A2(n_205),
.B1(n_191),
.B2(n_189),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_L g323 ( 
.A1(n_261),
.A2(n_263),
.B1(n_226),
.B2(n_225),
.Y(n_323)
);

INVx13_ASAP7_75t_L g262 ( 
.A(n_219),
.Y(n_262)
);

INVxp33_ASAP7_75t_L g315 ( 
.A(n_262),
.Y(n_315)
);

AOI22xp33_ASAP7_75t_L g263 ( 
.A1(n_244),
.A2(n_184),
.B1(n_179),
.B2(n_165),
.Y(n_263)
);

INVx4_ASAP7_75t_L g265 ( 
.A(n_211),
.Y(n_265)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_265),
.Y(n_306)
);

OR2x2_ASAP7_75t_SL g266 ( 
.A(n_230),
.B(n_174),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_266),
.B(n_271),
.C(n_236),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_232),
.Y(n_267)
);

INVx3_ASAP7_75t_L g268 ( 
.A(n_224),
.Y(n_268)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_268),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_232),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_269),
.B(n_275),
.Y(n_313)
);

BUFx2_ASAP7_75t_L g272 ( 
.A(n_224),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_272),
.Y(n_293)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_213),
.Y(n_273)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_273),
.Y(n_314)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_220),
.Y(n_274)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_274),
.Y(n_317)
);

CKINVDCx16_ASAP7_75t_R g275 ( 
.A(n_243),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_228),
.B(n_200),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_276),
.B(n_279),
.Y(n_318)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_213),
.Y(n_277)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_277),
.Y(n_319)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_220),
.Y(n_278)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_278),
.Y(n_322)
);

INVx13_ASAP7_75t_L g279 ( 
.A(n_219),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_239),
.Y(n_280)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_280),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_215),
.A2(n_38),
.B1(n_40),
.B2(n_178),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_282),
.B(n_283),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_214),
.B(n_33),
.Y(n_283)
);

INVx1_ASAP7_75t_SL g284 ( 
.A(n_219),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_284),
.B(n_242),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_SL g285 ( 
.A1(n_240),
.A2(n_200),
.B(n_145),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_285),
.A2(n_252),
.B(n_234),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_227),
.B(n_33),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_286),
.B(n_288),
.Y(n_296)
);

BUFx6f_ASAP7_75t_L g287 ( 
.A(n_211),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_287),
.Y(n_303)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_239),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_229),
.B(n_33),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_290),
.B(n_181),
.Y(n_301)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_222),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_291),
.Y(n_307)
);

INVx3_ASAP7_75t_L g292 ( 
.A(n_222),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_292),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_281),
.A2(n_216),
.B(n_252),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_SL g339 ( 
.A1(n_295),
.A2(n_300),
.B(n_289),
.Y(n_339)
);

OR2x2_ASAP7_75t_L g297 ( 
.A(n_255),
.B(n_241),
.Y(n_297)
);

INVx1_ASAP7_75t_SL g340 ( 
.A(n_297),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_299),
.B(n_262),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_301),
.B(n_302),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_283),
.B(n_218),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_L g304 ( 
.A1(n_281),
.A2(n_221),
.B(n_214),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_L g331 ( 
.A1(n_304),
.A2(n_325),
.B(n_277),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_264),
.B(n_218),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_309),
.B(n_311),
.Y(n_360)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_310),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_SL g311 ( 
.A(n_271),
.B(n_231),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_266),
.B(n_237),
.C(n_251),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_312),
.B(n_270),
.C(n_282),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_316),
.A2(n_238),
.B1(n_235),
.B2(n_278),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_260),
.A2(n_233),
.B1(n_237),
.B2(n_225),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_320),
.A2(n_324),
.B1(n_265),
.B2(n_292),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_323),
.B(n_270),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_L g325 ( 
.A1(n_259),
.A2(n_246),
.B(n_253),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_273),
.B(n_223),
.Y(n_329)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_329),
.Y(n_353)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_299),
.B(n_285),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_330),
.B(n_342),
.C(n_350),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_L g390 ( 
.A1(n_331),
.A2(n_333),
.B1(n_354),
.B2(n_307),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_310),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_332),
.B(n_334),
.Y(n_373)
);

NOR3xp33_ASAP7_75t_L g334 ( 
.A(n_309),
.B(n_288),
.C(n_280),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_327),
.B(n_253),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_SL g384 ( 
.A(n_335),
.B(n_337),
.Y(n_384)
);

AND2x6_ASAP7_75t_L g336 ( 
.A(n_295),
.B(n_279),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_SL g387 ( 
.A1(n_336),
.A2(n_339),
.B(n_345),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_327),
.B(n_267),
.Y(n_337)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_314),
.Y(n_341)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_341),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_343),
.A2(n_305),
.B1(n_296),
.B2(n_328),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_313),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_344),
.B(n_351),
.Y(n_367)
);

OAI21xp5_ASAP7_75t_L g345 ( 
.A1(n_295),
.A2(n_289),
.B(n_284),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_314),
.Y(n_346)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_346),
.Y(n_366)
);

BUFx6f_ASAP7_75t_L g347 ( 
.A(n_298),
.Y(n_347)
);

BUFx2_ASAP7_75t_L g371 ( 
.A(n_347),
.Y(n_371)
);

OAI22xp33_ASAP7_75t_SL g349 ( 
.A1(n_294),
.A2(n_257),
.B1(n_256),
.B2(n_272),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_349),
.A2(n_355),
.B1(n_324),
.B2(n_328),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_311),
.B(n_246),
.C(n_235),
.Y(n_350)
);

OAI21xp5_ASAP7_75t_L g351 ( 
.A1(n_300),
.A2(n_245),
.B(n_238),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_329),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_352),
.B(n_358),
.Y(n_369)
);

AOI22xp33_ASAP7_75t_SL g354 ( 
.A1(n_321),
.A2(n_291),
.B1(n_287),
.B2(n_268),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_356),
.B(n_357),
.C(n_359),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_304),
.B(n_274),
.C(n_28),
.Y(n_357)
);

AND2x6_ASAP7_75t_L g358 ( 
.A(n_316),
.B(n_13),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_312),
.B(n_28),
.Y(n_359)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_321),
.Y(n_361)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_361),
.Y(n_372)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_319),
.Y(n_362)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_362),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_L g401 ( 
.A1(n_363),
.A2(n_385),
.B1(n_391),
.B2(n_351),
.Y(n_401)
);

AO22x1_ASAP7_75t_SL g370 ( 
.A1(n_348),
.A2(n_320),
.B1(n_305),
.B2(n_325),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_370),
.B(n_343),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_374),
.A2(n_382),
.B1(n_322),
.B2(n_317),
.Y(n_409)
);

XNOR2x2_ASAP7_75t_L g375 ( 
.A(n_340),
.B(n_297),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_SL g397 ( 
.A(n_375),
.B(n_331),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_330),
.B(n_356),
.C(n_359),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_376),
.B(n_383),
.C(n_393),
.Y(n_394)
);

OR2x2_ASAP7_75t_L g378 ( 
.A(n_340),
.B(n_297),
.Y(n_378)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_378),
.Y(n_399)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_341),
.Y(n_379)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_379),
.Y(n_419)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_346),
.Y(n_380)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_380),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_360),
.B(n_302),
.Y(n_381)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_381),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_345),
.A2(n_296),
.B1(n_326),
.B2(n_319),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_350),
.B(n_318),
.C(n_326),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_355),
.A2(n_307),
.B1(n_303),
.B2(n_293),
.Y(n_385)
);

OR2x2_ASAP7_75t_L g386 ( 
.A(n_353),
.B(n_303),
.Y(n_386)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_386),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_360),
.B(n_315),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_SL g416 ( 
.A(n_388),
.B(n_389),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_338),
.B(n_301),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_SL g408 ( 
.A1(n_390),
.A2(n_361),
.B1(n_322),
.B2(n_317),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_358),
.A2(n_293),
.B1(n_321),
.B2(n_306),
.Y(n_391)
);

CKINVDCx16_ASAP7_75t_R g392 ( 
.A(n_362),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_SL g417 ( 
.A(n_392),
.B(n_0),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_357),
.B(n_306),
.C(n_308),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_365),
.B(n_376),
.C(n_368),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_395),
.B(n_387),
.C(n_373),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_386),
.B(n_298),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_396),
.B(n_398),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_397),
.B(n_403),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_SL g398 ( 
.A(n_369),
.B(n_347),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_400),
.B(n_370),
.Y(n_430)
);

HB1xp67_ASAP7_75t_L g437 ( 
.A(n_401),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_L g403 ( 
.A(n_365),
.B(n_339),
.Y(n_403)
);

XOR2xp5_ASAP7_75t_L g404 ( 
.A(n_368),
.B(n_342),
.Y(n_404)
);

XOR2xp5_ASAP7_75t_L g425 ( 
.A(n_404),
.B(n_405),
.Y(n_425)
);

XOR2xp5_ASAP7_75t_L g405 ( 
.A(n_383),
.B(n_336),
.Y(n_405)
);

XOR2xp5_ASAP7_75t_L g406 ( 
.A(n_393),
.B(n_308),
.Y(n_406)
);

XOR2xp5_ASAP7_75t_L g428 ( 
.A(n_406),
.B(n_410),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_SL g426 ( 
.A1(n_408),
.A2(n_409),
.B1(n_411),
.B2(n_363),
.Y(n_426)
);

XOR2xp5_ASAP7_75t_L g410 ( 
.A(n_382),
.B(n_28),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_374),
.A2(n_12),
.B1(n_1),
.B2(n_2),
.Y(n_411)
);

OAI22xp33_ASAP7_75t_SL g412 ( 
.A1(n_375),
.A2(n_47),
.B1(n_3),
.B2(n_4),
.Y(n_412)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_412),
.Y(n_427)
);

XOR2xp5_ASAP7_75t_L g413 ( 
.A(n_367),
.B(n_28),
.Y(n_413)
);

XOR2xp5_ASAP7_75t_L g439 ( 
.A(n_413),
.B(n_379),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_384),
.B(n_0),
.Y(n_414)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_414),
.Y(n_433)
);

OAI21xp5_ASAP7_75t_L g415 ( 
.A1(n_378),
.A2(n_47),
.B(n_3),
.Y(n_415)
);

INVxp67_ASAP7_75t_L g422 ( 
.A(n_415),
.Y(n_422)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_417),
.Y(n_435)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_418),
.Y(n_420)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_420),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_423),
.B(n_431),
.C(n_432),
.Y(n_449)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_416),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_SL g454 ( 
.A(n_424),
.B(n_440),
.Y(n_454)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_426),
.A2(n_410),
.B1(n_413),
.B2(n_405),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_430),
.B(n_434),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_394),
.B(n_387),
.C(n_391),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_394),
.B(n_385),
.C(n_364),
.Y(n_432)
);

INVxp67_ASAP7_75t_L g434 ( 
.A(n_408),
.Y(n_434)
);

MAJx2_ASAP7_75t_L g436 ( 
.A(n_395),
.B(n_370),
.C(n_380),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_436),
.B(n_403),
.C(n_404),
.Y(n_451)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_399),
.Y(n_438)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_438),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_439),
.B(n_397),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_SL g440 ( 
.A(n_407),
.B(n_377),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_L g465 ( 
.A1(n_441),
.A2(n_429),
.B1(n_377),
.B2(n_366),
.Y(n_465)
);

MAJx2_ASAP7_75t_L g470 ( 
.A(n_443),
.B(n_451),
.C(n_455),
.Y(n_470)
);

BUFx2_ASAP7_75t_L g444 ( 
.A(n_427),
.Y(n_444)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_444),
.Y(n_464)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_421),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_445),
.B(n_446),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_432),
.B(n_414),
.Y(n_446)
);

AOI21x1_ASAP7_75t_L g447 ( 
.A1(n_423),
.A2(n_400),
.B(n_415),
.Y(n_447)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_447),
.Y(n_472)
);

BUFx12_ASAP7_75t_L g448 ( 
.A(n_436),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_448),
.B(n_450),
.Y(n_468)
);

CKINVDCx16_ASAP7_75t_R g450 ( 
.A(n_433),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_425),
.B(n_406),
.C(n_409),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_455),
.B(n_428),
.C(n_431),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_435),
.B(n_411),
.Y(n_456)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_456),
.Y(n_469)
);

AOI21xp5_ASAP7_75t_L g457 ( 
.A1(n_434),
.A2(n_419),
.B(n_402),
.Y(n_457)
);

OAI21xp5_ASAP7_75t_SL g459 ( 
.A1(n_457),
.A2(n_422),
.B(n_366),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_458),
.B(n_5),
.C(n_8),
.Y(n_484)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_459),
.Y(n_482)
);

AOI22xp5_ASAP7_75t_L g460 ( 
.A1(n_457),
.A2(n_437),
.B1(n_422),
.B2(n_439),
.Y(n_460)
);

OAI22xp5_ASAP7_75t_L g477 ( 
.A1(n_460),
.A2(n_466),
.B1(n_471),
.B2(n_452),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_449),
.B(n_425),
.C(n_428),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_461),
.B(n_442),
.C(n_448),
.Y(n_481)
);

XOR2xp5_ASAP7_75t_L g462 ( 
.A(n_451),
.B(n_429),
.Y(n_462)
);

XOR2xp5_ASAP7_75t_L g476 ( 
.A(n_462),
.B(n_465),
.Y(n_476)
);

AOI22xp5_ASAP7_75t_L g466 ( 
.A1(n_444),
.A2(n_364),
.B1(n_372),
.B2(n_371),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_L g467 ( 
.A1(n_454),
.A2(n_372),
.B1(n_371),
.B2(n_4),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_467),
.B(n_442),
.Y(n_480)
);

XOR2xp5_ASAP7_75t_L g483 ( 
.A(n_470),
.B(n_5),
.Y(n_483)
);

AOI22xp5_ASAP7_75t_L g471 ( 
.A1(n_447),
.A2(n_0),
.B1(n_3),
.B2(n_5),
.Y(n_471)
);

OAI21xp5_ASAP7_75t_SL g473 ( 
.A1(n_463),
.A2(n_449),
.B(n_453),
.Y(n_473)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_473),
.Y(n_487)
);

XOR2x1_ASAP7_75t_SL g474 ( 
.A(n_468),
.B(n_448),
.Y(n_474)
);

OAI21x1_ASAP7_75t_L g489 ( 
.A1(n_474),
.A2(n_475),
.B(n_485),
.Y(n_489)
);

AOI21xp5_ASAP7_75t_L g475 ( 
.A1(n_472),
.A2(n_453),
.B(n_441),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_477),
.B(n_478),
.Y(n_493)
);

INVxp67_ASAP7_75t_L g478 ( 
.A(n_459),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_SL g479 ( 
.A(n_463),
.B(n_452),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_479),
.B(n_480),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_481),
.B(n_483),
.C(n_484),
.Y(n_490)
);

AOI21xp5_ASAP7_75t_L g485 ( 
.A1(n_461),
.A2(n_8),
.B(n_9),
.Y(n_485)
);

XOR2xp5_ASAP7_75t_L g486 ( 
.A(n_481),
.B(n_460),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_486),
.B(n_476),
.C(n_466),
.Y(n_498)
);

MAJx2_ASAP7_75t_L g488 ( 
.A(n_474),
.B(n_458),
.C(n_462),
.Y(n_488)
);

XNOR2xp5_ASAP7_75t_L g499 ( 
.A(n_488),
.B(n_10),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_476),
.B(n_470),
.C(n_469),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g496 ( 
.A(n_491),
.B(n_492),
.Y(n_496)
);

OAI21xp5_ASAP7_75t_L g492 ( 
.A1(n_482),
.A2(n_464),
.B(n_471),
.Y(n_492)
);

NOR2xp67_ASAP7_75t_L g495 ( 
.A(n_489),
.B(n_478),
.Y(n_495)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_495),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_494),
.B(n_483),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_SL g502 ( 
.A(n_497),
.B(n_499),
.Y(n_502)
);

OAI21xp5_ASAP7_75t_L g503 ( 
.A1(n_498),
.A2(n_500),
.B(n_490),
.Y(n_503)
);

AND2x2_ASAP7_75t_L g500 ( 
.A(n_487),
.B(n_493),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_503),
.B(n_488),
.C(n_486),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_502),
.B(n_496),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_504),
.B(n_505),
.C(n_501),
.Y(n_506)
);

A2O1A1Ixp33_ASAP7_75t_L g507 ( 
.A1(n_506),
.A2(n_11),
.B(n_495),
.C(n_503),
.Y(n_507)
);

INVxp33_ASAP7_75t_L g508 ( 
.A(n_507),
.Y(n_508)
);

XOR2xp5_ASAP7_75t_L g509 ( 
.A(n_508),
.B(n_11),
.Y(n_509)
);

XOR2xp5_ASAP7_75t_L g510 ( 
.A(n_509),
.B(n_11),
.Y(n_510)
);


endmodule