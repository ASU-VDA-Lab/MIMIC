module real_aes_6828_n_100 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_100);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_100;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_364;
wire n_421;
wire n_319;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_455;
wire n_504;
wire n_310;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_502;
wire n_434;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_349;
wire n_336;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_753;
wire n_741;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_546;
wire n_151;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_175;
wire n_241;
wire n_168;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g173 ( .A1(n_0), .A2(n_174), .B(n_177), .C(n_181), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_1), .B(n_165), .Y(n_184) );
INVx1_ASAP7_75t_L g112 ( .A(n_2), .Y(n_112) );
NAND2xp5_ASAP7_75t_SL g209 ( .A(n_3), .B(n_175), .Y(n_209) );
A2O1A1Ixp33_ASAP7_75t_L g504 ( .A1(n_4), .A2(n_138), .B(n_141), .C(n_505), .Y(n_504) );
AOI21xp5_ASAP7_75t_L g529 ( .A1(n_5), .A2(n_133), .B(n_530), .Y(n_529) );
AOI21xp5_ASAP7_75t_L g229 ( .A1(n_6), .A2(n_133), .B(n_230), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_7), .B(n_165), .Y(n_536) );
AO21x2_ASAP7_75t_L g238 ( .A1(n_8), .A2(n_167), .B(n_239), .Y(n_238) );
AOI222xp33_ASAP7_75t_L g115 ( .A1(n_9), .A2(n_116), .B1(n_727), .B2(n_728), .C1(n_731), .C2(n_734), .Y(n_115) );
AND2x6_ASAP7_75t_L g138 ( .A(n_10), .B(n_139), .Y(n_138) );
A2O1A1Ixp33_ASAP7_75t_L g255 ( .A1(n_11), .A2(n_138), .B(n_141), .C(n_256), .Y(n_255) );
INVx1_ASAP7_75t_L g496 ( .A(n_12), .Y(n_496) );
NOR2xp33_ASAP7_75t_L g113 ( .A(n_13), .B(n_40), .Y(n_113) );
NAND2xp5_ASAP7_75t_SL g507 ( .A(n_14), .B(n_180), .Y(n_507) );
INVx1_ASAP7_75t_L g159 ( .A(n_15), .Y(n_159) );
NAND2xp5_ASAP7_75t_SL g245 ( .A(n_16), .B(n_175), .Y(n_245) );
NAND2xp5_ASAP7_75t_SL g750 ( .A(n_17), .B(n_751), .Y(n_750) );
A2O1A1Ixp33_ASAP7_75t_L g515 ( .A1(n_18), .A2(n_176), .B(n_516), .C(n_518), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_19), .B(n_165), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_20), .B(n_153), .Y(n_473) );
A2O1A1Ixp33_ASAP7_75t_L g140 ( .A1(n_21), .A2(n_141), .B(n_144), .C(n_152), .Y(n_140) );
A2O1A1Ixp33_ASAP7_75t_L g545 ( .A1(n_22), .A2(n_179), .B(n_247), .C(n_546), .Y(n_545) );
NAND2xp5_ASAP7_75t_SL g481 ( .A(n_23), .B(n_180), .Y(n_481) );
NAND2xp5_ASAP7_75t_SL g458 ( .A(n_24), .B(n_180), .Y(n_458) );
CKINVDCx16_ASAP7_75t_R g477 ( .A(n_25), .Y(n_477) );
INVx1_ASAP7_75t_L g457 ( .A(n_26), .Y(n_457) );
A2O1A1Ixp33_ASAP7_75t_L g241 ( .A1(n_27), .A2(n_141), .B(n_152), .C(n_242), .Y(n_241) );
BUFx6f_ASAP7_75t_L g137 ( .A(n_28), .Y(n_137) );
CKINVDCx20_ASAP7_75t_R g503 ( .A(n_29), .Y(n_503) );
INVx1_ASAP7_75t_L g471 ( .A(n_30), .Y(n_471) );
AOI21xp5_ASAP7_75t_L g169 ( .A1(n_31), .A2(n_133), .B(n_170), .Y(n_169) );
INVx2_ASAP7_75t_L g136 ( .A(n_32), .Y(n_136) );
A2O1A1Ixp33_ASAP7_75t_L g190 ( .A1(n_33), .A2(n_191), .B(n_192), .C(n_196), .Y(n_190) );
CKINVDCx20_ASAP7_75t_R g509 ( .A(n_34), .Y(n_509) );
A2O1A1Ixp33_ASAP7_75t_L g532 ( .A1(n_35), .A2(n_179), .B(n_533), .C(n_535), .Y(n_532) );
INVxp67_ASAP7_75t_L g472 ( .A(n_36), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_37), .B(n_244), .Y(n_243) );
A2O1A1Ixp33_ASAP7_75t_L g455 ( .A1(n_38), .A2(n_141), .B(n_152), .C(n_456), .Y(n_455) );
CKINVDCx14_ASAP7_75t_R g531 ( .A(n_39), .Y(n_531) );
A2O1A1Ixp33_ASAP7_75t_L g493 ( .A1(n_41), .A2(n_181), .B(n_494), .C(n_495), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g131 ( .A(n_42), .B(n_132), .Y(n_131) );
CKINVDCx20_ASAP7_75t_R g260 ( .A(n_43), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_44), .B(n_175), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_45), .B(n_133), .Y(n_240) );
CKINVDCx20_ASAP7_75t_R g460 ( .A(n_46), .Y(n_460) );
CKINVDCx20_ASAP7_75t_R g468 ( .A(n_47), .Y(n_468) );
A2O1A1Ixp33_ASAP7_75t_L g220 ( .A1(n_48), .A2(n_191), .B(n_196), .C(n_221), .Y(n_220) );
INVx1_ASAP7_75t_L g178 ( .A(n_49), .Y(n_178) );
INVx1_ASAP7_75t_L g222 ( .A(n_50), .Y(n_222) );
INVx1_ASAP7_75t_L g544 ( .A(n_51), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_52), .B(n_133), .Y(n_219) );
CKINVDCx20_ASAP7_75t_R g161 ( .A(n_53), .Y(n_161) );
CKINVDCx14_ASAP7_75t_R g492 ( .A(n_54), .Y(n_492) );
INVx1_ASAP7_75t_L g139 ( .A(n_55), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_56), .B(n_133), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_57), .B(n_165), .Y(n_235) );
A2O1A1Ixp33_ASAP7_75t_L g232 ( .A1(n_58), .A2(n_151), .B(n_207), .C(n_233), .Y(n_232) );
INVx1_ASAP7_75t_L g158 ( .A(n_59), .Y(n_158) );
INVx1_ASAP7_75t_SL g534 ( .A(n_60), .Y(n_534) );
CKINVDCx20_ASAP7_75t_R g106 ( .A(n_61), .Y(n_106) );
NAND2xp5_ASAP7_75t_SL g194 ( .A(n_62), .B(n_175), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_63), .B(n_165), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_64), .B(n_176), .Y(n_257) );
INVx1_ASAP7_75t_L g480 ( .A(n_65), .Y(n_480) );
CKINVDCx16_ASAP7_75t_R g171 ( .A(n_66), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g145 ( .A(n_67), .B(n_146), .Y(n_145) );
A2O1A1Ixp33_ASAP7_75t_L g204 ( .A1(n_68), .A2(n_141), .B(n_196), .C(n_205), .Y(n_204) );
CKINVDCx16_ASAP7_75t_R g231 ( .A(n_69), .Y(n_231) );
INVx1_ASAP7_75t_L g105 ( .A(n_70), .Y(n_105) );
AOI21xp5_ASAP7_75t_L g490 ( .A1(n_71), .A2(n_133), .B(n_491), .Y(n_490) );
AOI222xp33_ASAP7_75t_SL g100 ( .A1(n_72), .A2(n_101), .B1(n_114), .B2(n_737), .C1(n_742), .C2(n_753), .Y(n_100) );
AOI22xp5_ASAP7_75t_L g745 ( .A1(n_72), .A2(n_92), .B1(n_746), .B2(n_747), .Y(n_745) );
CKINVDCx20_ASAP7_75t_R g747 ( .A(n_72), .Y(n_747) );
CKINVDCx20_ASAP7_75t_R g484 ( .A(n_73), .Y(n_484) );
AOI21xp5_ASAP7_75t_L g512 ( .A1(n_74), .A2(n_133), .B(n_513), .Y(n_512) );
OAI22xp5_ASAP7_75t_L g728 ( .A1(n_75), .A2(n_99), .B1(n_729), .B2(n_730), .Y(n_728) );
CKINVDCx20_ASAP7_75t_R g730 ( .A(n_75), .Y(n_730) );
AOI21xp5_ASAP7_75t_L g466 ( .A1(n_76), .A2(n_132), .B(n_467), .Y(n_466) );
CKINVDCx16_ASAP7_75t_R g454 ( .A(n_77), .Y(n_454) );
INVx1_ASAP7_75t_L g514 ( .A(n_78), .Y(n_514) );
NAND2xp5_ASAP7_75t_SL g148 ( .A(n_79), .B(n_149), .Y(n_148) );
CKINVDCx20_ASAP7_75t_R g198 ( .A(n_80), .Y(n_198) );
AOI21xp5_ASAP7_75t_L g542 ( .A1(n_81), .A2(n_133), .B(n_543), .Y(n_542) );
INVx1_ASAP7_75t_L g517 ( .A(n_82), .Y(n_517) );
INVx2_ASAP7_75t_L g156 ( .A(n_83), .Y(n_156) );
INVx1_ASAP7_75t_L g506 ( .A(n_84), .Y(n_506) );
CKINVDCx20_ASAP7_75t_R g214 ( .A(n_85), .Y(n_214) );
NAND2xp5_ASAP7_75t_SL g258 ( .A(n_86), .B(n_180), .Y(n_258) );
OR2x2_ASAP7_75t_L g109 ( .A(n_87), .B(n_110), .Y(n_109) );
OR2x2_ASAP7_75t_L g119 ( .A(n_87), .B(n_111), .Y(n_119) );
INVx2_ASAP7_75t_L g446 ( .A(n_87), .Y(n_446) );
A2O1A1Ixp33_ASAP7_75t_L g478 ( .A1(n_88), .A2(n_141), .B(n_196), .C(n_479), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_89), .B(n_133), .Y(n_189) );
INVx1_ASAP7_75t_L g193 ( .A(n_90), .Y(n_193) );
INVxp67_ASAP7_75t_L g234 ( .A(n_91), .Y(n_234) );
CKINVDCx20_ASAP7_75t_R g746 ( .A(n_92), .Y(n_746) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_93), .B(n_167), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g104 ( .A(n_94), .B(n_105), .Y(n_104) );
INVx1_ASAP7_75t_L g206 ( .A(n_95), .Y(n_206) );
INVx1_ASAP7_75t_L g253 ( .A(n_96), .Y(n_253) );
INVx2_ASAP7_75t_L g547 ( .A(n_97), .Y(n_547) );
AND2x2_ASAP7_75t_L g224 ( .A(n_98), .B(n_155), .Y(n_224) );
CKINVDCx20_ASAP7_75t_R g729 ( .A(n_99), .Y(n_729) );
INVx1_ASAP7_75t_SL g101 ( .A(n_102), .Y(n_101) );
NAND2xp33_ASAP7_75t_L g102 ( .A(n_103), .B(n_107), .Y(n_102) );
NOR2xp33_ASAP7_75t_SL g103 ( .A(n_104), .B(n_106), .Y(n_103) );
INVx1_ASAP7_75t_SL g741 ( .A(n_104), .Y(n_741) );
INVx1_ASAP7_75t_L g740 ( .A(n_106), .Y(n_740) );
OA21x2_ASAP7_75t_L g754 ( .A1(n_106), .A2(n_741), .B(n_752), .Y(n_754) );
INVx1_ASAP7_75t_SL g107 ( .A(n_108), .Y(n_107) );
INVx1_ASAP7_75t_SL g108 ( .A(n_109), .Y(n_108) );
HB1xp67_ASAP7_75t_L g749 ( .A(n_109), .Y(n_749) );
BUFx2_ASAP7_75t_L g752 ( .A(n_109), .Y(n_752) );
NOR2x2_ASAP7_75t_L g733 ( .A(n_110), .B(n_446), .Y(n_733) );
INVx2_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
OR2x2_ASAP7_75t_L g445 ( .A(n_111), .B(n_446), .Y(n_445) );
AND2x2_ASAP7_75t_L g111 ( .A(n_112), .B(n_113), .Y(n_111) );
INVxp67_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
OAI22xp5_ASAP7_75t_L g116 ( .A1(n_117), .A2(n_120), .B1(n_443), .B2(n_447), .Y(n_116) );
OAI22xp5_ASAP7_75t_SL g734 ( .A1(n_117), .A2(n_121), .B1(n_735), .B2(n_736), .Y(n_734) );
INVx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
OAI22xp5_ASAP7_75t_L g743 ( .A1(n_120), .A2(n_121), .B1(n_744), .B2(n_745), .Y(n_743) );
INVx2_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
AND2x2_ASAP7_75t_SL g121 ( .A(n_122), .B(n_398), .Y(n_121) );
NOR2xp33_ASAP7_75t_L g122 ( .A(n_123), .B(n_333), .Y(n_122) );
NAND4xp25_ASAP7_75t_SL g123 ( .A(n_124), .B(n_278), .C(n_302), .D(n_325), .Y(n_123) );
AOI221xp5_ASAP7_75t_L g124 ( .A1(n_125), .A2(n_215), .B1(n_249), .B2(n_262), .C(n_265), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
NAND2xp5_ASAP7_75t_L g126 ( .A(n_127), .B(n_185), .Y(n_126) );
AOI22xp33_ASAP7_75t_L g268 ( .A1(n_127), .A2(n_163), .B1(n_216), .B2(n_269), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_127), .B(n_186), .Y(n_336) );
AND2x2_ASAP7_75t_L g355 ( .A(n_127), .B(n_356), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_127), .B(n_339), .Y(n_425) );
AND2x4_ASAP7_75t_L g127 ( .A(n_128), .B(n_163), .Y(n_127) );
AND2x2_ASAP7_75t_L g293 ( .A(n_128), .B(n_186), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_128), .B(n_308), .Y(n_307) );
OR2x2_ASAP7_75t_L g316 ( .A(n_128), .B(n_317), .Y(n_316) );
AND2x2_ASAP7_75t_L g321 ( .A(n_128), .B(n_164), .Y(n_321) );
INVx2_ASAP7_75t_L g353 ( .A(n_128), .Y(n_353) );
HB1xp67_ASAP7_75t_L g397 ( .A(n_128), .Y(n_397) );
AND2x2_ASAP7_75t_L g414 ( .A(n_128), .B(n_291), .Y(n_414) );
INVx5_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
AND2x2_ASAP7_75t_L g332 ( .A(n_129), .B(n_291), .Y(n_332) );
AND2x4_ASAP7_75t_L g346 ( .A(n_129), .B(n_163), .Y(n_346) );
HB1xp67_ASAP7_75t_L g350 ( .A(n_129), .Y(n_350) );
AND2x2_ASAP7_75t_L g370 ( .A(n_129), .B(n_285), .Y(n_370) );
AND2x2_ASAP7_75t_L g420 ( .A(n_129), .B(n_187), .Y(n_420) );
AND2x2_ASAP7_75t_L g430 ( .A(n_129), .B(n_164), .Y(n_430) );
OR2x6_ASAP7_75t_L g129 ( .A(n_130), .B(n_160), .Y(n_129) );
AOI21xp5_ASAP7_75t_SL g130 ( .A1(n_131), .A2(n_140), .B(n_153), .Y(n_130) );
BUFx2_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
AND2x4_ASAP7_75t_L g133 ( .A(n_134), .B(n_138), .Y(n_133) );
NAND2x1p5_ASAP7_75t_L g254 ( .A(n_134), .B(n_138), .Y(n_254) );
AND2x2_ASAP7_75t_L g134 ( .A(n_135), .B(n_137), .Y(n_134) );
INVx1_ASAP7_75t_L g151 ( .A(n_135), .Y(n_151) );
INVx1_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
INVx2_ASAP7_75t_L g142 ( .A(n_136), .Y(n_142) );
INVx1_ASAP7_75t_L g248 ( .A(n_136), .Y(n_248) );
INVx1_ASAP7_75t_L g143 ( .A(n_137), .Y(n_143) );
BUFx6f_ASAP7_75t_L g147 ( .A(n_137), .Y(n_147) );
INVx3_ASAP7_75t_L g176 ( .A(n_137), .Y(n_176) );
BUFx6f_ASAP7_75t_L g180 ( .A(n_137), .Y(n_180) );
INVx1_ASAP7_75t_L g244 ( .A(n_137), .Y(n_244) );
BUFx3_ASAP7_75t_L g152 ( .A(n_138), .Y(n_152) );
INVx4_ASAP7_75t_SL g183 ( .A(n_138), .Y(n_183) );
INVx5_ASAP7_75t_L g172 ( .A(n_141), .Y(n_172) );
AND2x6_ASAP7_75t_L g141 ( .A(n_142), .B(n_143), .Y(n_141) );
BUFx3_ASAP7_75t_L g182 ( .A(n_142), .Y(n_182) );
BUFx6f_ASAP7_75t_L g211 ( .A(n_142), .Y(n_211) );
AOI21xp5_ASAP7_75t_L g144 ( .A1(n_145), .A2(n_148), .B(n_150), .Y(n_144) );
INVx2_ASAP7_75t_L g149 ( .A(n_146), .Y(n_149) );
INVx2_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx4_ASAP7_75t_L g208 ( .A(n_147), .Y(n_208) );
O2A1O1Ixp33_ASAP7_75t_L g192 ( .A1(n_149), .A2(n_193), .B(n_194), .C(n_195), .Y(n_192) );
O2A1O1Ixp33_ASAP7_75t_L g221 ( .A1(n_149), .A2(n_195), .B(n_222), .C(n_223), .Y(n_221) );
O2A1O1Ixp33_ASAP7_75t_L g479 ( .A1(n_149), .A2(n_480), .B(n_481), .C(n_482), .Y(n_479) );
O2A1O1Ixp5_ASAP7_75t_L g505 ( .A1(n_149), .A2(n_482), .B(n_506), .C(n_507), .Y(n_505) );
O2A1O1Ixp33_ASAP7_75t_L g456 ( .A1(n_150), .A2(n_175), .B(n_457), .C(n_458), .Y(n_456) );
INVx2_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
NAND2xp5_ASAP7_75t_SL g469 ( .A(n_151), .B(n_470), .Y(n_469) );
INVx1_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
NOR2xp33_ASAP7_75t_L g483 ( .A(n_154), .B(n_484), .Y(n_483) );
INVx2_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx1_ASAP7_75t_L g162 ( .A(n_155), .Y(n_162) );
AOI21xp5_ASAP7_75t_L g188 ( .A1(n_155), .A2(n_189), .B(n_190), .Y(n_188) );
AOI21xp5_ASAP7_75t_L g218 ( .A1(n_155), .A2(n_219), .B(n_220), .Y(n_218) );
O2A1O1Ixp33_ASAP7_75t_L g453 ( .A1(n_155), .A2(n_254), .B(n_454), .C(n_455), .Y(n_453) );
OA21x2_ASAP7_75t_L g489 ( .A1(n_155), .A2(n_490), .B(n_497), .Y(n_489) );
AND2x2_ASAP7_75t_SL g155 ( .A(n_156), .B(n_157), .Y(n_155) );
AND2x2_ASAP7_75t_L g168 ( .A(n_156), .B(n_157), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_158), .B(n_159), .Y(n_157) );
NOR2xp33_ASAP7_75t_L g160 ( .A(n_161), .B(n_162), .Y(n_160) );
AO21x2_ASAP7_75t_L g501 ( .A1(n_162), .A2(n_502), .B(n_508), .Y(n_501) );
AND2x2_ASAP7_75t_L g286 ( .A(n_163), .B(n_186), .Y(n_286) );
HB1xp67_ASAP7_75t_L g301 ( .A(n_163), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_163), .B(n_328), .Y(n_327) );
INVx1_ASAP7_75t_L g376 ( .A(n_163), .Y(n_376) );
INVx2_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
AND2x2_ASAP7_75t_L g264 ( .A(n_164), .B(n_201), .Y(n_264) );
AND2x2_ASAP7_75t_L g291 ( .A(n_164), .B(n_202), .Y(n_291) );
OA21x2_ASAP7_75t_L g164 ( .A1(n_165), .A2(n_169), .B(n_184), .Y(n_164) );
INVx3_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
NOR2xp33_ASAP7_75t_L g197 ( .A(n_166), .B(n_198), .Y(n_197) );
AO21x2_ASAP7_75t_L g202 ( .A1(n_166), .A2(n_203), .B(n_213), .Y(n_202) );
NOR2xp33_ASAP7_75t_L g213 ( .A(n_166), .B(n_214), .Y(n_213) );
AO21x2_ASAP7_75t_L g251 ( .A1(n_166), .A2(n_252), .B(n_259), .Y(n_251) );
NOR2xp33_ASAP7_75t_L g459 ( .A(n_166), .B(n_460), .Y(n_459) );
AO21x2_ASAP7_75t_L g475 ( .A1(n_166), .A2(n_476), .B(n_483), .Y(n_475) );
NOR2xp33_ASAP7_75t_L g508 ( .A(n_166), .B(n_509), .Y(n_508) );
INVx4_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
HB1xp67_ASAP7_75t_L g228 ( .A(n_167), .Y(n_228) );
AOI21xp5_ASAP7_75t_L g239 ( .A1(n_167), .A2(n_240), .B(n_241), .Y(n_239) );
BUFx6f_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
INVx1_ASAP7_75t_L g261 ( .A(n_168), .Y(n_261) );
O2A1O1Ixp33_ASAP7_75t_SL g170 ( .A1(n_171), .A2(n_172), .B(n_173), .C(n_183), .Y(n_170) );
INVx2_ASAP7_75t_L g191 ( .A(n_172), .Y(n_191) );
O2A1O1Ixp33_ASAP7_75t_L g230 ( .A1(n_172), .A2(n_183), .B(n_231), .C(n_232), .Y(n_230) );
O2A1O1Ixp33_ASAP7_75t_SL g467 ( .A1(n_172), .A2(n_183), .B(n_468), .C(n_469), .Y(n_467) );
O2A1O1Ixp33_ASAP7_75t_SL g491 ( .A1(n_172), .A2(n_183), .B(n_492), .C(n_493), .Y(n_491) );
O2A1O1Ixp33_ASAP7_75t_SL g513 ( .A1(n_172), .A2(n_183), .B(n_514), .C(n_515), .Y(n_513) );
O2A1O1Ixp33_ASAP7_75t_L g530 ( .A1(n_172), .A2(n_183), .B(n_531), .C(n_532), .Y(n_530) );
O2A1O1Ixp33_ASAP7_75t_SL g543 ( .A1(n_172), .A2(n_183), .B(n_544), .C(n_545), .Y(n_543) );
INVx2_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
NOR2xp33_ASAP7_75t_L g233 ( .A(n_175), .B(n_234), .Y(n_233) );
OAI22xp33_ASAP7_75t_L g470 ( .A1(n_175), .A2(n_208), .B1(n_471), .B2(n_472), .Y(n_470) );
INVx5_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
NOR2xp33_ASAP7_75t_L g495 ( .A(n_176), .B(n_496), .Y(n_495) );
NOR2xp33_ASAP7_75t_L g177 ( .A(n_178), .B(n_179), .Y(n_177) );
NOR2xp33_ASAP7_75t_L g533 ( .A(n_179), .B(n_534), .Y(n_533) );
INVx4_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
INVx2_ASAP7_75t_L g494 ( .A(n_180), .Y(n_494) );
INVx2_ASAP7_75t_L g482 ( .A(n_181), .Y(n_482) );
INVx2_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
HB1xp67_ASAP7_75t_L g195 ( .A(n_182), .Y(n_195) );
INVx1_ASAP7_75t_L g518 ( .A(n_182), .Y(n_518) );
INVx1_ASAP7_75t_L g196 ( .A(n_183), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_185), .B(n_350), .Y(n_349) );
AND2x2_ASAP7_75t_L g185 ( .A(n_186), .B(n_199), .Y(n_185) );
OR2x2_ASAP7_75t_L g317 ( .A(n_186), .B(n_200), .Y(n_317) );
AND2x2_ASAP7_75t_L g354 ( .A(n_186), .B(n_264), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_186), .B(n_285), .Y(n_365) );
HB1xp67_ASAP7_75t_L g369 ( .A(n_186), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_186), .B(n_321), .Y(n_438) );
INVx5_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
BUFx2_ASAP7_75t_L g263 ( .A(n_187), .Y(n_263) );
AND2x2_ASAP7_75t_L g272 ( .A(n_187), .B(n_200), .Y(n_272) );
AND2x2_ASAP7_75t_L g388 ( .A(n_187), .B(n_283), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_187), .B(n_321), .Y(n_410) );
OR2x6_ASAP7_75t_L g187 ( .A(n_188), .B(n_197), .Y(n_187) );
INVx1_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
HB1xp67_ASAP7_75t_L g356 ( .A(n_200), .Y(n_356) );
INVx2_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
HB1xp67_ASAP7_75t_L g308 ( .A(n_201), .Y(n_308) );
INVx2_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
BUFx2_ASAP7_75t_L g285 ( .A(n_202), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_204), .B(n_212), .Y(n_203) );
O2A1O1Ixp33_ASAP7_75t_L g205 ( .A1(n_206), .A2(n_207), .B(n_209), .C(n_210), .Y(n_205) );
INVx1_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
NOR2xp33_ASAP7_75t_L g516 ( .A(n_208), .B(n_517), .Y(n_516) );
NOR2xp33_ASAP7_75t_L g546 ( .A(n_208), .B(n_547), .Y(n_546) );
HB1xp67_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
INVx3_ASAP7_75t_L g535 ( .A(n_211), .Y(n_535) );
NOR2xp33_ASAP7_75t_L g215 ( .A(n_216), .B(n_225), .Y(n_215) );
NOR2xp33_ASAP7_75t_L g417 ( .A(n_216), .B(n_298), .Y(n_417) );
HB1xp67_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
NOR2xp33_ASAP7_75t_L g249 ( .A(n_217), .B(n_250), .Y(n_249) );
AND2x2_ASAP7_75t_L g269 ( .A(n_217), .B(n_270), .Y(n_269) );
INVx5_ASAP7_75t_SL g277 ( .A(n_217), .Y(n_277) );
OR2x2_ASAP7_75t_L g300 ( .A(n_217), .B(n_270), .Y(n_300) );
OR2x2_ASAP7_75t_L g310 ( .A(n_217), .B(n_311), .Y(n_310) );
AND2x2_ASAP7_75t_L g373 ( .A(n_217), .B(n_227), .Y(n_373) );
AND2x2_ASAP7_75t_SL g411 ( .A(n_217), .B(n_226), .Y(n_411) );
NOR4xp25_ASAP7_75t_L g432 ( .A(n_217), .B(n_353), .C(n_433), .D(n_434), .Y(n_432) );
AND2x2_ASAP7_75t_L g442 ( .A(n_217), .B(n_274), .Y(n_442) );
OR2x6_ASAP7_75t_L g217 ( .A(n_218), .B(n_224), .Y(n_217) );
INVx2_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
AND2x2_ASAP7_75t_L g267 ( .A(n_226), .B(n_263), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_226), .B(n_269), .Y(n_436) );
AND2x2_ASAP7_75t_L g226 ( .A(n_227), .B(n_236), .Y(n_226) );
OR2x2_ASAP7_75t_L g276 ( .A(n_227), .B(n_277), .Y(n_276) );
INVx3_ASAP7_75t_L g283 ( .A(n_227), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_227), .B(n_251), .Y(n_295) );
INVxp67_ASAP7_75t_L g298 ( .A(n_227), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_227), .B(n_270), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_227), .B(n_237), .Y(n_364) );
AND2x2_ASAP7_75t_L g379 ( .A(n_227), .B(n_274), .Y(n_379) );
OR2x2_ASAP7_75t_L g408 ( .A(n_227), .B(n_237), .Y(n_408) );
OA21x2_ASAP7_75t_L g227 ( .A1(n_228), .A2(n_229), .B(n_235), .Y(n_227) );
OA21x2_ASAP7_75t_L g511 ( .A1(n_228), .A2(n_512), .B(n_519), .Y(n_511) );
OA21x2_ASAP7_75t_L g528 ( .A1(n_228), .A2(n_529), .B(n_536), .Y(n_528) );
OA21x2_ASAP7_75t_L g541 ( .A1(n_228), .A2(n_542), .B(n_548), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_236), .B(n_313), .Y(n_312) );
NOR2xp33_ASAP7_75t_L g416 ( .A(n_236), .B(n_277), .Y(n_416) );
OR2x2_ASAP7_75t_L g437 ( .A(n_236), .B(n_314), .Y(n_437) );
INVx1_ASAP7_75t_SL g236 ( .A(n_237), .Y(n_236) );
OR2x2_ASAP7_75t_L g250 ( .A(n_237), .B(n_251), .Y(n_250) );
AND2x2_ASAP7_75t_L g274 ( .A(n_237), .B(n_270), .Y(n_274) );
NAND2xp5_ASAP7_75t_SL g289 ( .A(n_237), .B(n_251), .Y(n_289) );
AND2x2_ASAP7_75t_L g359 ( .A(n_237), .B(n_283), .Y(n_359) );
AND2x2_ASAP7_75t_L g393 ( .A(n_237), .B(n_277), .Y(n_393) );
INVx2_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_238), .B(n_277), .Y(n_296) );
AND2x2_ASAP7_75t_L g324 ( .A(n_238), .B(n_251), .Y(n_324) );
AOI21xp5_ASAP7_75t_L g242 ( .A1(n_243), .A2(n_245), .B(n_246), .Y(n_242) );
AOI21xp5_ASAP7_75t_L g256 ( .A1(n_246), .A2(n_257), .B(n_258), .Y(n_256) );
INVx2_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
INVx3_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_249), .B(n_332), .Y(n_331) );
AOI221xp5_ASAP7_75t_L g391 ( .A1(n_250), .A2(n_339), .B1(n_375), .B2(n_392), .C(n_394), .Y(n_391) );
INVx5_ASAP7_75t_SL g270 ( .A(n_251), .Y(n_270) );
OAI21xp5_ASAP7_75t_L g252 ( .A1(n_253), .A2(n_254), .B(n_255), .Y(n_252) );
OAI21xp5_ASAP7_75t_L g476 ( .A1(n_254), .A2(n_477), .B(n_478), .Y(n_476) );
OAI21xp5_ASAP7_75t_L g502 ( .A1(n_254), .A2(n_503), .B(n_504), .Y(n_502) );
NOR2xp33_ASAP7_75t_L g259 ( .A(n_260), .B(n_261), .Y(n_259) );
INVx2_ASAP7_75t_L g465 ( .A(n_261), .Y(n_465) );
AND2x2_ASAP7_75t_L g262 ( .A(n_263), .B(n_264), .Y(n_262) );
OAI33xp33_ASAP7_75t_L g290 ( .A1(n_263), .A2(n_291), .A3(n_292), .B1(n_294), .B2(n_297), .B3(n_301), .Y(n_290) );
OR2x2_ASAP7_75t_L g306 ( .A(n_263), .B(n_307), .Y(n_306) );
AOI322xp5_ASAP7_75t_L g415 ( .A1(n_263), .A2(n_332), .A3(n_339), .B1(n_416), .B2(n_417), .C1(n_418), .C2(n_421), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_263), .B(n_291), .Y(n_433) );
A2O1A1Ixp33_ASAP7_75t_SL g439 ( .A1(n_263), .A2(n_291), .B(n_440), .C(n_442), .Y(n_439) );
AOI221xp5_ASAP7_75t_L g278 ( .A1(n_264), .A2(n_279), .B1(n_284), .B2(n_287), .C(n_290), .Y(n_278) );
INVx1_ASAP7_75t_L g371 ( .A(n_264), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_264), .B(n_420), .Y(n_419) );
OAI22xp33_ASAP7_75t_L g265 ( .A1(n_266), .A2(n_268), .B1(n_271), .B2(n_273), .Y(n_265) );
INVx1_ASAP7_75t_SL g266 ( .A(n_267), .Y(n_266) );
AND2x2_ASAP7_75t_L g348 ( .A(n_269), .B(n_283), .Y(n_348) );
AND2x2_ASAP7_75t_L g406 ( .A(n_269), .B(n_407), .Y(n_406) );
OR2x2_ASAP7_75t_L g314 ( .A(n_270), .B(n_277), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_270), .B(n_283), .Y(n_342) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_272), .B(n_345), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_272), .B(n_350), .Y(n_404) );
OAI321xp33_ASAP7_75t_L g423 ( .A1(n_272), .A2(n_345), .A3(n_424), .B1(n_425), .B2(n_426), .C(n_427), .Y(n_423) );
INVx1_ASAP7_75t_L g390 ( .A(n_273), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_274), .B(n_275), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_274), .B(n_281), .Y(n_280) );
AND2x2_ASAP7_75t_L g329 ( .A(n_274), .B(n_277), .Y(n_329) );
AOI321xp33_ASAP7_75t_L g387 ( .A1(n_274), .A2(n_291), .A3(n_388), .B1(n_389), .B2(n_390), .C(n_391), .Y(n_387) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
OR2x2_ASAP7_75t_L g304 ( .A(n_276), .B(n_289), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_277), .B(n_283), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_277), .B(n_359), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_277), .B(n_363), .Y(n_400) );
INVx1_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
AND2x4_ASAP7_75t_L g323 ( .A(n_281), .B(n_324), .Y(n_323) );
INVx2_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
OR2x2_ASAP7_75t_L g288 ( .A(n_282), .B(n_289), .Y(n_288) );
INVx1_ASAP7_75t_L g396 ( .A(n_283), .Y(n_396) );
AND2x2_ASAP7_75t_L g284 ( .A(n_285), .B(n_286), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_286), .B(n_339), .Y(n_338) );
INVx2_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
INVx1_ASAP7_75t_L g319 ( .A(n_291), .Y(n_319) );
INVx1_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
NOR2xp33_ASAP7_75t_L g377 ( .A(n_293), .B(n_328), .Y(n_377) );
OR2x2_ASAP7_75t_L g294 ( .A(n_295), .B(n_296), .Y(n_294) );
OR2x2_ASAP7_75t_L g341 ( .A(n_296), .B(n_342), .Y(n_341) );
INVx1_ASAP7_75t_SL g386 ( .A(n_296), .Y(n_386) );
OAI22xp5_ASAP7_75t_L g343 ( .A1(n_297), .A2(n_344), .B1(n_347), .B2(n_349), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_298), .B(n_299), .Y(n_297) );
INVx1_ASAP7_75t_SL g299 ( .A(n_300), .Y(n_299) );
OR2x2_ASAP7_75t_L g441 ( .A(n_300), .B(n_364), .Y(n_441) );
AOI221xp5_ASAP7_75t_L g302 ( .A1(n_303), .A2(n_305), .B1(n_309), .B2(n_315), .C(n_318), .Y(n_302) );
INVx1_ASAP7_75t_SL g303 ( .A(n_304), .Y(n_303) );
INVx2_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
BUFx2_ASAP7_75t_L g339 ( .A(n_308), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_310), .B(n_312), .Y(n_309) );
INVx1_ASAP7_75t_SL g385 ( .A(n_311), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_313), .B(n_363), .Y(n_362) );
AOI21xp5_ASAP7_75t_L g380 ( .A1(n_313), .A2(n_381), .B(n_383), .Y(n_380) );
INVx2_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
OR2x2_ASAP7_75t_L g426 ( .A(n_314), .B(n_408), .Y(n_426) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
INVx2_ASAP7_75t_SL g328 ( .A(n_317), .Y(n_328) );
AOI21xp33_ASAP7_75t_L g318 ( .A1(n_319), .A2(n_320), .B(n_322), .Y(n_318) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
INVx2_ASAP7_75t_SL g322 ( .A(n_323), .Y(n_322) );
AND2x2_ASAP7_75t_L g372 ( .A(n_324), .B(n_373), .Y(n_372) );
INVxp67_ASAP7_75t_L g434 ( .A(n_324), .Y(n_434) );
AOI21xp5_ASAP7_75t_L g325 ( .A1(n_326), .A2(n_329), .B(n_330), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_328), .B(n_346), .Y(n_382) );
INVxp67_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
INVx1_ASAP7_75t_L g403 ( .A(n_332), .Y(n_403) );
NAND5xp2_ASAP7_75t_L g333 ( .A(n_334), .B(n_351), .C(n_360), .D(n_380), .E(n_387), .Y(n_333) );
O2A1O1Ixp33_ASAP7_75t_L g334 ( .A1(n_335), .A2(n_337), .B(n_340), .C(n_343), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
INVx1_ASAP7_75t_L g375 ( .A(n_339), .Y(n_375) );
CKINVDCx16_ASAP7_75t_R g340 ( .A(n_341), .Y(n_340) );
INVx1_ASAP7_75t_SL g345 ( .A(n_346), .Y(n_345) );
NOR2xp33_ASAP7_75t_L g412 ( .A(n_347), .B(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVx1_ASAP7_75t_L g389 ( .A(n_349), .Y(n_389) );
OAI21xp5_ASAP7_75t_SL g351 ( .A1(n_352), .A2(n_355), .B(n_357), .Y(n_351) );
AOI221xp5_ASAP7_75t_L g405 ( .A1(n_352), .A2(n_406), .B1(n_409), .B2(n_411), .C(n_412), .Y(n_405) );
AND2x2_ASAP7_75t_L g352 ( .A(n_353), .B(n_354), .Y(n_352) );
AOI321xp33_ASAP7_75t_L g360 ( .A1(n_353), .A2(n_361), .A3(n_365), .B1(n_366), .B2(n_372), .C(n_374), .Y(n_360) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx1_ASAP7_75t_SL g363 ( .A(n_364), .Y(n_363) );
INVx1_ASAP7_75t_L g431 ( .A(n_365), .Y(n_431) );
NAND2xp5_ASAP7_75t_SL g366 ( .A(n_367), .B(n_371), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
AND2x2_ASAP7_75t_L g383 ( .A(n_368), .B(n_384), .Y(n_383) );
AND2x2_ASAP7_75t_L g368 ( .A(n_369), .B(n_370), .Y(n_368) );
NOR2xp67_ASAP7_75t_SL g395 ( .A(n_369), .B(n_376), .Y(n_395) );
AOI321xp33_ASAP7_75t_SL g427 ( .A1(n_372), .A2(n_428), .A3(n_429), .B1(n_430), .B2(n_431), .C(n_432), .Y(n_427) );
O2A1O1Ixp33_ASAP7_75t_L g374 ( .A1(n_375), .A2(n_376), .B(n_377), .C(n_378), .Y(n_374) );
INVx1_ASAP7_75t_SL g378 ( .A(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
AND2x2_ASAP7_75t_L g384 ( .A(n_385), .B(n_386), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_385), .B(n_393), .Y(n_422) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
NAND3xp33_ASAP7_75t_L g394 ( .A(n_395), .B(n_396), .C(n_397), .Y(n_394) );
NOR3xp33_ASAP7_75t_L g398 ( .A(n_399), .B(n_423), .C(n_435), .Y(n_398) );
OAI211xp5_ASAP7_75t_SL g399 ( .A1(n_400), .A2(n_401), .B(n_405), .C(n_415), .Y(n_399) );
INVxp67_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
NAND2xp5_ASAP7_75t_SL g402 ( .A(n_403), .B(n_404), .Y(n_402) );
OAI221xp5_ASAP7_75t_L g435 ( .A1(n_404), .A2(n_436), .B1(n_437), .B2(n_438), .C(n_439), .Y(n_435) );
INVx1_ASAP7_75t_L g424 ( .A(n_406), .Y(n_424) );
INVx1_ASAP7_75t_SL g407 ( .A(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_SL g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx1_ASAP7_75t_SL g428 ( .A(n_426), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
CKINVDCx14_ASAP7_75t_R g440 ( .A(n_441), .Y(n_440) );
INVx2_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx2_ASAP7_75t_L g736 ( .A(n_444), .Y(n_736) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx2_ASAP7_75t_L g735 ( .A(n_447), .Y(n_735) );
OR4x2_ASAP7_75t_L g447 ( .A(n_448), .B(n_617), .C(n_664), .D(n_704), .Y(n_447) );
NAND3xp33_ASAP7_75t_SL g448 ( .A(n_449), .B(n_563), .C(n_592), .Y(n_448) );
AOI211xp5_ASAP7_75t_L g449 ( .A1(n_450), .A2(n_485), .B(n_520), .C(n_556), .Y(n_449) );
O2A1O1Ixp33_ASAP7_75t_L g592 ( .A1(n_450), .A2(n_576), .B(n_593), .C(n_597), .Y(n_592) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_452), .B(n_461), .Y(n_451) );
NAND2xp5_ASAP7_75t_SL g554 ( .A(n_452), .B(n_555), .Y(n_554) );
INVx3_ASAP7_75t_SL g559 ( .A(n_452), .Y(n_559) );
HB1xp67_ASAP7_75t_L g571 ( .A(n_452), .Y(n_571) );
AND2x4_ASAP7_75t_L g575 ( .A(n_452), .B(n_527), .Y(n_575) );
AND2x2_ASAP7_75t_L g586 ( .A(n_452), .B(n_475), .Y(n_586) );
OR2x2_ASAP7_75t_L g610 ( .A(n_452), .B(n_523), .Y(n_610) );
AND2x2_ASAP7_75t_L g623 ( .A(n_452), .B(n_528), .Y(n_623) );
AND2x2_ASAP7_75t_L g663 ( .A(n_452), .B(n_649), .Y(n_663) );
AND2x2_ASAP7_75t_L g670 ( .A(n_452), .B(n_633), .Y(n_670) );
AND2x2_ASAP7_75t_L g700 ( .A(n_452), .B(n_462), .Y(n_700) );
OR2x6_ASAP7_75t_L g452 ( .A(n_453), .B(n_459), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_461), .B(n_627), .Y(n_639) );
AND2x2_ASAP7_75t_L g461 ( .A(n_462), .B(n_474), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_462), .B(n_570), .Y(n_569) );
OR2x2_ASAP7_75t_L g577 ( .A(n_462), .B(n_474), .Y(n_577) );
BUFx3_ASAP7_75t_L g585 ( .A(n_462), .Y(n_585) );
OR2x2_ASAP7_75t_L g606 ( .A(n_462), .B(n_488), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_462), .B(n_627), .Y(n_717) );
OA21x2_ASAP7_75t_L g462 ( .A1(n_463), .A2(n_466), .B(n_473), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
AO21x2_ASAP7_75t_L g523 ( .A1(n_464), .A2(n_524), .B(n_525), .Y(n_523) );
INVx1_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
INVx1_ASAP7_75t_L g524 ( .A(n_466), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_473), .Y(n_525) );
AND2x2_ASAP7_75t_L g526 ( .A(n_474), .B(n_527), .Y(n_526) );
INVx1_ASAP7_75t_L g570 ( .A(n_474), .Y(n_570) );
AND2x2_ASAP7_75t_L g633 ( .A(n_474), .B(n_528), .Y(n_633) );
AOI221xp5_ASAP7_75t_L g635 ( .A1(n_474), .A2(n_636), .B1(n_638), .B2(n_640), .C(n_641), .Y(n_635) );
AND2x2_ASAP7_75t_L g649 ( .A(n_474), .B(n_523), .Y(n_649) );
AND2x2_ASAP7_75t_L g675 ( .A(n_474), .B(n_559), .Y(n_675) );
INVx2_ASAP7_75t_SL g474 ( .A(n_475), .Y(n_474) );
AND2x2_ASAP7_75t_L g555 ( .A(n_475), .B(n_528), .Y(n_555) );
BUFx2_ASAP7_75t_L g689 ( .A(n_475), .Y(n_689) );
INVx1_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
OAI32xp33_ASAP7_75t_L g655 ( .A1(n_486), .A2(n_616), .A3(n_630), .B1(n_656), .B2(n_657), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_487), .B(n_498), .Y(n_486) );
AND2x2_ASAP7_75t_L g596 ( .A(n_487), .B(n_540), .Y(n_596) );
INVx1_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
OR2x2_ASAP7_75t_L g578 ( .A(n_488), .B(n_579), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_488), .B(n_589), .Y(n_588) );
AND2x2_ASAP7_75t_L g650 ( .A(n_488), .B(n_540), .Y(n_650) );
AND2x2_ASAP7_75t_L g661 ( .A(n_488), .B(n_553), .Y(n_661) );
BUFx3_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
OR2x2_ASAP7_75t_L g562 ( .A(n_489), .B(n_541), .Y(n_562) );
AND2x2_ASAP7_75t_L g566 ( .A(n_489), .B(n_541), .Y(n_566) );
AND2x2_ASAP7_75t_L g601 ( .A(n_489), .B(n_552), .Y(n_601) );
AND2x2_ASAP7_75t_L g608 ( .A(n_489), .B(n_510), .Y(n_608) );
OAI211xp5_ASAP7_75t_L g613 ( .A1(n_489), .A2(n_559), .B(n_570), .C(n_614), .Y(n_613) );
INVx2_ASAP7_75t_L g667 ( .A(n_489), .Y(n_667) );
NOR2xp33_ASAP7_75t_L g678 ( .A(n_489), .B(n_500), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_498), .B(n_550), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_498), .B(n_566), .Y(n_656) );
INVx1_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
OR2x2_ASAP7_75t_L g561 ( .A(n_499), .B(n_562), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_500), .B(n_510), .Y(n_499) );
AND2x2_ASAP7_75t_L g553 ( .A(n_500), .B(n_511), .Y(n_553) );
OR2x2_ASAP7_75t_L g568 ( .A(n_500), .B(n_511), .Y(n_568) );
AND2x2_ASAP7_75t_L g591 ( .A(n_500), .B(n_552), .Y(n_591) );
INVx1_ASAP7_75t_L g595 ( .A(n_500), .Y(n_595) );
AND2x2_ASAP7_75t_L g614 ( .A(n_500), .B(n_551), .Y(n_614) );
OAI22xp33_ASAP7_75t_L g624 ( .A1(n_500), .A2(n_579), .B1(n_625), .B2(n_626), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_500), .B(n_667), .Y(n_691) );
AND2x2_ASAP7_75t_L g706 ( .A(n_500), .B(n_566), .Y(n_706) );
INVx4_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
BUFx3_ASAP7_75t_L g538 ( .A(n_501), .Y(n_538) );
AND2x2_ASAP7_75t_L g580 ( .A(n_501), .B(n_511), .Y(n_580) );
AND2x2_ASAP7_75t_L g582 ( .A(n_501), .B(n_540), .Y(n_582) );
AND3x2_ASAP7_75t_L g644 ( .A(n_501), .B(n_608), .C(n_645), .Y(n_644) );
AND2x2_ASAP7_75t_L g679 ( .A(n_510), .B(n_551), .Y(n_679) );
INVx1_ASAP7_75t_SL g510 ( .A(n_511), .Y(n_510) );
AND2x2_ASAP7_75t_L g540 ( .A(n_511), .B(n_541), .Y(n_540) );
HB1xp67_ASAP7_75t_L g589 ( .A(n_511), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_511), .B(n_550), .Y(n_612) );
NAND3xp33_ASAP7_75t_L g719 ( .A(n_511), .B(n_591), .C(n_667), .Y(n_719) );
OAI22xp5_ASAP7_75t_L g520 ( .A1(n_521), .A2(n_537), .B1(n_549), .B2(n_554), .Y(n_520) );
INVx1_ASAP7_75t_SL g521 ( .A(n_522), .Y(n_521) );
AND2x2_ASAP7_75t_L g522 ( .A(n_523), .B(n_526), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_523), .B(n_616), .Y(n_615) );
INVx1_ASAP7_75t_SL g631 ( .A(n_523), .Y(n_631) );
OAI31xp33_ASAP7_75t_L g647 ( .A1(n_526), .A2(n_648), .A3(n_649), .B(n_650), .Y(n_647) );
AND2x2_ASAP7_75t_L g672 ( .A(n_526), .B(n_559), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_526), .B(n_585), .Y(n_718) );
AND2x2_ASAP7_75t_L g627 ( .A(n_527), .B(n_559), .Y(n_627) );
AND2x2_ASAP7_75t_L g688 ( .A(n_527), .B(n_689), .Y(n_688) );
INVx2_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
AND2x2_ASAP7_75t_L g558 ( .A(n_528), .B(n_559), .Y(n_558) );
INVx1_ASAP7_75t_L g616 ( .A(n_528), .Y(n_616) );
OR2x2_ASAP7_75t_L g537 ( .A(n_538), .B(n_539), .Y(n_537) );
CKINVDCx16_ASAP7_75t_R g637 ( .A(n_538), .Y(n_637) );
NOR2xp33_ASAP7_75t_L g690 ( .A(n_539), .B(n_691), .Y(n_690) );
INVx1_ASAP7_75t_SL g539 ( .A(n_540), .Y(n_539) );
AOI221x1_ASAP7_75t_SL g604 ( .A1(n_540), .A2(n_605), .B1(n_607), .B2(n_609), .C(n_611), .Y(n_604) );
INVx2_ASAP7_75t_L g552 ( .A(n_541), .Y(n_552) );
HB1xp67_ASAP7_75t_L g646 ( .A(n_541), .Y(n_646) );
INVx1_ASAP7_75t_L g634 ( .A(n_549), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_550), .B(n_553), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_550), .B(n_567), .Y(n_659) );
INVx1_ASAP7_75t_SL g722 ( .A(n_550), .Y(n_722) );
INVx2_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
INVx2_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
AND2x2_ASAP7_75t_L g640 ( .A(n_553), .B(n_566), .Y(n_640) );
INVx1_ASAP7_75t_L g708 ( .A(n_554), .Y(n_708) );
NOR2xp33_ASAP7_75t_L g721 ( .A(n_554), .B(n_637), .Y(n_721) );
INVx2_ASAP7_75t_SL g560 ( .A(n_555), .Y(n_560) );
AND2x2_ASAP7_75t_L g603 ( .A(n_555), .B(n_559), .Y(n_603) );
NOR2xp33_ASAP7_75t_L g609 ( .A(n_555), .B(n_610), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_555), .B(n_630), .Y(n_657) );
AOI21xp33_ASAP7_75t_SL g556 ( .A1(n_557), .A2(n_560), .B(n_561), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_558), .B(n_630), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_558), .B(n_585), .Y(n_726) );
OR2x2_ASAP7_75t_L g598 ( .A(n_559), .B(n_577), .Y(n_598) );
AND2x2_ASAP7_75t_L g697 ( .A(n_559), .B(n_688), .Y(n_697) );
OAI22xp5_ASAP7_75t_SL g572 ( .A1(n_560), .A2(n_573), .B1(n_578), .B2(n_581), .Y(n_572) );
NOR2xp33_ASAP7_75t_L g605 ( .A(n_560), .B(n_606), .Y(n_605) );
OR2x2_ASAP7_75t_L g620 ( .A(n_562), .B(n_568), .Y(n_620) );
INVx1_ASAP7_75t_L g684 ( .A(n_562), .Y(n_684) );
AOI311xp33_ASAP7_75t_L g563 ( .A1(n_564), .A2(n_569), .A3(n_571), .B(n_572), .C(n_583), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_566), .B(n_567), .Y(n_565) );
AOI221xp5_ASAP7_75t_L g710 ( .A1(n_567), .A2(n_699), .B1(n_711), .B2(n_714), .C(n_716), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_567), .B(n_722), .Y(n_724) );
INVx2_ASAP7_75t_SL g567 ( .A(n_568), .Y(n_567) );
INVx1_ASAP7_75t_L g621 ( .A(n_569), .Y(n_621) );
AOI211xp5_ASAP7_75t_L g611 ( .A1(n_570), .A2(n_612), .B(n_613), .C(n_615), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_574), .B(n_576), .Y(n_573) );
O2A1O1Ixp33_ASAP7_75t_SL g680 ( .A1(n_574), .A2(n_576), .B(n_681), .C(n_682), .Y(n_680) );
INVx3_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_575), .B(n_649), .Y(n_715) );
INVx1_ASAP7_75t_SL g576 ( .A(n_577), .Y(n_576) );
OAI221xp5_ASAP7_75t_L g597 ( .A1(n_578), .A2(n_598), .B1(n_599), .B2(n_602), .C(n_604), .Y(n_597) );
INVx1_ASAP7_75t_SL g579 ( .A(n_580), .Y(n_579) );
AND2x2_ASAP7_75t_L g600 ( .A(n_580), .B(n_601), .Y(n_600) );
AND2x2_ASAP7_75t_L g683 ( .A(n_580), .B(n_684), .Y(n_683) );
INVx1_ASAP7_75t_SL g581 ( .A(n_582), .Y(n_581) );
NOR2xp33_ASAP7_75t_L g583 ( .A(n_584), .B(n_587), .Y(n_583) );
A2O1A1Ixp33_ASAP7_75t_L g641 ( .A1(n_584), .A2(n_642), .B(n_643), .C(n_647), .Y(n_641) );
NAND2xp5_ASAP7_75t_SL g584 ( .A(n_585), .B(n_586), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_585), .B(n_675), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_585), .B(n_688), .Y(n_687) );
OR2x2_ASAP7_75t_L g587 ( .A(n_588), .B(n_590), .Y(n_587) );
INVxp67_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
AND2x2_ASAP7_75t_L g607 ( .A(n_591), .B(n_608), .Y(n_607) );
INVx1_ASAP7_75t_SL g593 ( .A(n_594), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_595), .B(n_596), .Y(n_594) );
NOR2xp33_ASAP7_75t_L g666 ( .A(n_595), .B(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g709 ( .A(n_598), .Y(n_709) );
INVx1_ASAP7_75t_SL g599 ( .A(n_600), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_601), .B(n_630), .Y(n_629) );
AND2x2_ASAP7_75t_L g636 ( .A(n_601), .B(n_637), .Y(n_636) );
INVx1_ASAP7_75t_SL g713 ( .A(n_601), .Y(n_713) );
INVx1_ASAP7_75t_SL g602 ( .A(n_603), .Y(n_602) );
AND2x2_ASAP7_75t_L g654 ( .A(n_603), .B(n_630), .Y(n_654) );
INVx1_ASAP7_75t_SL g648 ( .A(n_610), .Y(n_648) );
INVx1_ASAP7_75t_L g625 ( .A(n_616), .Y(n_625) );
NAND3xp33_ASAP7_75t_SL g617 ( .A(n_618), .B(n_635), .C(n_651), .Y(n_617) );
AOI322xp5_ASAP7_75t_L g618 ( .A1(n_619), .A2(n_621), .A3(n_622), .B1(n_624), .B2(n_628), .C1(n_632), .C2(n_634), .Y(n_618) );
AOI211xp5_ASAP7_75t_L g671 ( .A1(n_619), .A2(n_672), .B(n_673), .C(n_680), .Y(n_671) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
OAI22xp5_ASAP7_75t_L g673 ( .A1(n_622), .A2(n_643), .B1(n_674), .B2(n_676), .Y(n_673) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
AND2x2_ASAP7_75t_L g632 ( .A(n_630), .B(n_633), .Y(n_632) );
AND2x2_ASAP7_75t_L g669 ( .A(n_630), .B(n_670), .Y(n_669) );
AOI32xp33_ASAP7_75t_L g720 ( .A1(n_630), .A2(n_721), .A3(n_722), .B1(n_723), .B2(n_725), .Y(n_720) );
INVx2_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
INVx1_ASAP7_75t_L g642 ( .A(n_633), .Y(n_642) );
AOI221xp5_ASAP7_75t_L g685 ( .A1(n_633), .A2(n_686), .B1(n_690), .B2(n_692), .C(n_695), .Y(n_685) );
AND2x2_ASAP7_75t_L g699 ( .A(n_633), .B(n_700), .Y(n_699) );
AND2x2_ASAP7_75t_L g702 ( .A(n_637), .B(n_703), .Y(n_702) );
OR2x2_ASAP7_75t_L g712 ( .A(n_637), .B(n_713), .Y(n_712) );
INVxp67_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
INVx2_ASAP7_75t_SL g643 ( .A(n_644), .Y(n_643) );
INVxp67_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
AND2x2_ASAP7_75t_L g703 ( .A(n_646), .B(n_667), .Y(n_703) );
AOI211xp5_ASAP7_75t_L g651 ( .A1(n_652), .A2(n_654), .B(n_655), .C(n_658), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
AOI21xp33_ASAP7_75t_L g658 ( .A1(n_659), .A2(n_660), .B(n_662), .Y(n_658) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
OAI211xp5_ASAP7_75t_SL g664 ( .A1(n_665), .A2(n_668), .B(n_671), .C(n_685), .Y(n_664) );
INVxp67_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
AND2x2_ASAP7_75t_L g677 ( .A(n_678), .B(n_679), .Y(n_677) );
NAND2xp5_ASAP7_75t_SL g693 ( .A(n_679), .B(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g694 ( .A(n_691), .Y(n_694) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
AOI21xp33_ASAP7_75t_L g695 ( .A1(n_696), .A2(n_698), .B(n_701), .Y(n_695) );
INVx1_ASAP7_75t_SL g696 ( .A(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
OAI211xp5_ASAP7_75t_SL g704 ( .A1(n_705), .A2(n_707), .B(n_710), .C(n_720), .Y(n_704) );
CKINVDCx20_ASAP7_75t_R g705 ( .A(n_706), .Y(n_705) );
NOR2xp33_ASAP7_75t_L g707 ( .A(n_708), .B(n_709), .Y(n_707) );
INVx1_ASAP7_75t_SL g711 ( .A(n_712), .Y(n_711) );
INVx1_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
AOI21xp33_ASAP7_75t_L g716 ( .A1(n_717), .A2(n_718), .B(n_719), .Y(n_716) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
INVx1_ASAP7_75t_SL g731 ( .A(n_732), .Y(n_731) );
INVx2_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
HB1xp67_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
AND2x2_ASAP7_75t_L g738 ( .A(n_739), .B(n_741), .Y(n_738) );
INVx1_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
OAI21xp5_ASAP7_75t_SL g742 ( .A1(n_743), .A2(n_748), .B(n_750), .Y(n_742) );
INVx1_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
INVx1_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
INVx1_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
CKINVDCx20_ASAP7_75t_R g753 ( .A(n_754), .Y(n_753) );
endmodule