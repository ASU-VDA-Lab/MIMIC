module fake_aes_943_n_1349 (n_303, n_117, n_219, n_44, n_133, n_149, n_289, n_220, n_81, n_69, n_214, n_267, n_204, n_221, n_249, n_185, n_22, n_203, n_57, n_88, n_52, n_244, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_284, n_107, n_158, n_278, n_60, n_300, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_240, n_254, n_9, n_161, n_262, n_10, n_177, n_130, n_189, n_103, n_239, n_19, n_87, n_137, n_180, n_292, n_104, n_277, n_160, n_98, n_74, n_206, n_276, n_154, n_272, n_7, n_29, n_285, n_195, n_165, n_146, n_45, n_85, n_250, n_237, n_181, n_101, n_62, n_255, n_36, n_47, n_215, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_217, n_139, n_229, n_230, n_274, n_16, n_13, n_198, n_169, n_193, n_273, n_282, n_252, n_152, n_113, n_241, n_95, n_124, n_156, n_238, n_297, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_247, n_197, n_201, n_242, n_260, n_6, n_4, n_304, n_127, n_291, n_170, n_294, n_40, n_111, n_157, n_296, n_79, n_202, n_210, n_38, n_64, n_142, n_184, n_245, n_265, n_191, n_264, n_281, n_232, n_200, n_46, n_31, n_208, n_211, n_58, n_122, n_187, n_138, n_126, n_275, n_178, n_118, n_258, n_253, n_32, n_0, n_179, n_84, n_131, n_112, n_266, n_55, n_205, n_12, n_86, n_143, n_213, n_235, n_243, n_295, n_182, n_263, n_166, n_162, n_186, n_75, n_163, n_226, n_105, n_159, n_174, n_227, n_248, n_268, n_231, n_72, n_136, n_298, n_283, n_299, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_256, n_67, n_77, n_216, n_20, n_2, n_147, n_199, n_54, n_148, n_293, n_123, n_83, n_172, n_28, n_48, n_100, n_212, n_305, n_228, n_92, n_11, n_223, n_251, n_25, n_30, n_59, n_236, n_150, n_218, n_168, n_194, n_3, n_287, n_18, n_110, n_261, n_301, n_66, n_134, n_222, n_234, n_1, n_164, n_233, n_271, n_82, n_106, n_175, n_15, n_173, n_190, n_286, n_302, n_145, n_270, n_246, n_153, n_61, n_259, n_290, n_280, n_21, n_99, n_109, n_93, n_132, n_288, n_151, n_51, n_140, n_207, n_257, n_224, n_96, n_269, n_225, n_39, n_279, n_1349);
input n_303;
input n_117;
input n_219;
input n_44;
input n_133;
input n_149;
input n_289;
input n_220;
input n_81;
input n_69;
input n_214;
input n_267;
input n_204;
input n_221;
input n_249;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_244;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_284;
input n_107;
input n_158;
input n_278;
input n_60;
input n_300;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_240;
input n_254;
input n_9;
input n_161;
input n_262;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_239;
input n_19;
input n_87;
input n_137;
input n_180;
input n_292;
input n_104;
input n_277;
input n_160;
input n_98;
input n_74;
input n_206;
input n_276;
input n_154;
input n_272;
input n_7;
input n_29;
input n_285;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_250;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_47;
input n_215;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_217;
input n_139;
input n_229;
input n_230;
input n_274;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_273;
input n_282;
input n_252;
input n_152;
input n_113;
input n_241;
input n_95;
input n_124;
input n_156;
input n_238;
input n_297;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_247;
input n_197;
input n_201;
input n_242;
input n_260;
input n_6;
input n_4;
input n_304;
input n_127;
input n_291;
input n_170;
input n_294;
input n_40;
input n_111;
input n_157;
input n_296;
input n_79;
input n_202;
input n_210;
input n_38;
input n_64;
input n_142;
input n_184;
input n_245;
input n_265;
input n_191;
input n_264;
input n_281;
input n_232;
input n_200;
input n_46;
input n_31;
input n_208;
input n_211;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_275;
input n_178;
input n_118;
input n_258;
input n_253;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_266;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_213;
input n_235;
input n_243;
input n_295;
input n_182;
input n_263;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_226;
input n_105;
input n_159;
input n_174;
input n_227;
input n_248;
input n_268;
input n_231;
input n_72;
input n_136;
input n_298;
input n_283;
input n_299;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_256;
input n_67;
input n_77;
input n_216;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_293;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_212;
input n_305;
input n_228;
input n_92;
input n_11;
input n_223;
input n_251;
input n_25;
input n_30;
input n_59;
input n_236;
input n_150;
input n_218;
input n_168;
input n_194;
input n_3;
input n_287;
input n_18;
input n_110;
input n_261;
input n_301;
input n_66;
input n_134;
input n_222;
input n_234;
input n_1;
input n_164;
input n_233;
input n_271;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_286;
input n_302;
input n_145;
input n_270;
input n_246;
input n_153;
input n_61;
input n_259;
input n_290;
input n_280;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_288;
input n_151;
input n_51;
input n_140;
input n_207;
input n_257;
input n_224;
input n_96;
input n_269;
input n_225;
input n_39;
input n_279;
output n_1349;
wire n_1309;
wire n_963;
wire n_1034;
wire n_949;
wire n_1277;
wire n_1312;
wire n_858;
wire n_646;
wire n_1334;
wire n_829;
wire n_1198;
wire n_667;
wire n_988;
wire n_311;
wire n_655;
wire n_1298;
wire n_903;
wire n_965;
wire n_918;
wire n_770;
wire n_1211;
wire n_878;
wire n_637;
wire n_564;
wire n_779;
wire n_528;
wire n_1128;
wire n_850;
wire n_672;
wire n_627;
wire n_1118;
wire n_1161;
wire n_1030;
wire n_807;
wire n_877;
wire n_545;
wire n_896;
wire n_334;
wire n_588;
wire n_1019;
wire n_940;
wire n_789;
wire n_1197;
wire n_1163;
wire n_387;
wire n_452;
wire n_518;
wire n_1336;
wire n_411;
wire n_1341;
wire n_860;
wire n_1208;
wire n_1201;
wire n_1342;
wire n_340;
wire n_373;
wire n_1194;
wire n_922;
wire n_465;
wire n_636;
wire n_914;
wire n_1005;
wire n_1097;
wire n_1125;
wire n_1017;
wire n_324;
wire n_773;
wire n_847;
wire n_668;
wire n_437;
wire n_680;
wire n_642;
wire n_1267;
wire n_830;
wire n_1112;
wire n_517;
wire n_1295;
wire n_1297;
wire n_502;
wire n_543;
wire n_312;
wire n_1159;
wire n_1250;
wire n_1002;
wire n_915;
wire n_367;
wire n_314;
wire n_999;
wire n_769;
wire n_624;
wire n_725;
wire n_1018;
wire n_979;
wire n_319;
wire n_499;
wire n_1033;
wire n_1063;
wire n_1010;
wire n_533;
wire n_490;
wire n_648;
wire n_613;
wire n_892;
wire n_571;
wire n_610;
wire n_771;
wire n_1337;
wire n_474;
wire n_402;
wire n_413;
wire n_676;
wire n_950;
wire n_995;
wire n_938;
wire n_331;
wire n_746;
wire n_1307;
wire n_619;
wire n_501;
wire n_699;
wire n_338;
wire n_551;
wire n_404;
wire n_1061;
wire n_509;
wire n_849;
wire n_864;
wire n_961;
wire n_1140;
wire n_611;
wire n_990;
wire n_800;
wire n_626;
wire n_1209;
wire n_926;
wire n_1274;
wire n_537;
wire n_660;
wire n_839;
wire n_1210;
wire n_1001;
wire n_1129;
wire n_450;
wire n_1099;
wire n_1328;
wire n_556;
wire n_1214;
wire n_379;
wire n_641;
wire n_966;
wire n_527;
wire n_797;
wire n_666;
wire n_1313;
wire n_954;
wire n_574;
wire n_822;
wire n_706;
wire n_823;
wire n_1181;
wire n_390;
wire n_514;
wire n_486;
wire n_568;
wire n_716;
wire n_899;
wire n_1066;
wire n_1251;
wire n_1199;
wire n_883;
wire n_573;
wire n_1308;
wire n_673;
wire n_1071;
wire n_1323;
wire n_1079;
wire n_315;
wire n_409;
wire n_1321;
wire n_677;
wire n_1242;
wire n_756;
wire n_1240;
wire n_1139;
wire n_577;
wire n_870;
wire n_1324;
wire n_790;
wire n_761;
wire n_1287;
wire n_472;
wire n_1100;
wire n_419;
wire n_1193;
wire n_1119;
wire n_825;
wire n_477;
wire n_815;
wire n_908;
wire n_429;
wire n_488;
wire n_821;
wire n_745;
wire n_684;
wire n_1281;
wire n_327;
wire n_1102;
wire n_723;
wire n_972;
wire n_997;
wire n_1244;
wire n_1184;
wire n_947;
wire n_620;
wire n_1141;
wire n_1213;
wire n_359;
wire n_1189;
wire n_1316;
wire n_923;
wire n_1205;
wire n_1172;
wire n_741;
wire n_1142;
wire n_1228;
wire n_831;
wire n_859;
wire n_1165;
wire n_1300;
wire n_930;
wire n_994;
wire n_410;
wire n_774;
wire n_1207;
wire n_377;
wire n_510;
wire n_1075;
wire n_1282;
wire n_493;
wire n_855;
wire n_722;
wire n_1083;
wire n_690;
wire n_1164;
wire n_451;
wire n_487;
wire n_748;
wire n_824;
wire n_793;
wire n_753;
wire n_355;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_1226;
wire n_1233;
wire n_1067;
wire n_866;
wire n_1108;
wire n_350;
wire n_433;
wire n_1311;
wire n_483;
wire n_395;
wire n_992;
wire n_361;
wire n_1077;
wire n_838;
wire n_705;
wire n_964;
wire n_590;
wire n_407;
wire n_1229;
wire n_792;
wire n_925;
wire n_1289;
wire n_957;
wire n_808;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_1306;
wire n_958;
wire n_468;
wire n_917;
wire n_523;
wire n_920;
wire n_1202;
wire n_1333;
wire n_911;
wire n_980;
wire n_817;
wire n_1056;
wire n_856;
wire n_1345;
wire n_661;
wire n_890;
wire n_787;
wire n_1015;
wire n_548;
wire n_1048;
wire n_973;
wire n_587;
wire n_476;
wire n_434;
wire n_489;
wire n_752;
wire n_1098;
wire n_1012;
wire n_461;
wire n_857;
wire n_1090;
wire n_786;
wire n_1121;
wire n_576;
wire n_1179;
wire n_796;
wire n_1216;
wire n_927;
wire n_840;
wire n_846;
wire n_968;
wire n_512;
wire n_1330;
wire n_586;
wire n_1246;
wire n_1276;
wire n_560;
wire n_697;
wire n_780;
wire n_447;
wire n_897;
wire n_1188;
wire n_580;
wire n_1009;
wire n_921;
wire n_854;
wire n_1011;
wire n_1155;
wire n_511;
wire n_467;
wire n_692;
wire n_644;
wire n_1116;
wire n_818;
wire n_738;
wire n_1225;
wire n_575;
wire n_711;
wire n_977;
wire n_884;
wire n_767;
wire n_393;
wire n_550;
wire n_826;
wire n_399;
wire n_1235;
wire n_1171;
wire n_459;
wire n_907;
wire n_310;
wire n_1062;
wire n_708;
wire n_1271;
wire n_307;
wire n_634;
wire n_696;
wire n_1203;
wire n_1013;
wire n_1000;
wire n_939;
wire n_953;
wire n_391;
wire n_478;
wire n_482;
wire n_394;
wire n_442;
wire n_485;
wire n_1248;
wire n_519;
wire n_329;
wire n_1020;
wire n_1106;
wire n_635;
wire n_731;
wire n_986;
wire n_507;
wire n_605;
wire n_704;
wire n_633;
wire n_873;
wire n_1322;
wire n_751;
wire n_1147;
wire n_466;
wire n_900;
wire n_952;
wire n_685;
wire n_308;
wire n_565;
wire n_1035;
wire n_475;
wire n_578;
wire n_542;
wire n_430;
wire n_943;
wire n_1326;
wire n_557;
wire n_842;
wire n_1269;
wire n_439;
wire n_614;
wire n_1346;
wire n_1107;
wire n_446;
wire n_423;
wire n_342;
wire n_799;
wire n_1050;
wire n_643;
wire n_874;
wire n_1049;
wire n_454;
wire n_687;
wire n_970;
wire n_984;
wire n_720;
wire n_806;
wire n_1157;
wire n_539;
wire n_1153;
wire n_317;
wire n_816;
wire n_522;
wire n_898;
wire n_1135;
wire n_669;
wire n_541;
wire n_363;
wire n_733;
wire n_894;
wire n_376;
wire n_744;
wire n_520;
wire n_681;
wire n_942;
wire n_1029;
wire n_508;
wire n_721;
wire n_1060;
wire n_438;
wire n_640;
wire n_1037;
wire n_686;
wire n_944;
wire n_1110;
wire n_498;
wire n_1069;
wire n_1123;
wire n_811;
wire n_530;
wire n_737;
wire n_1266;
wire n_795;
wire n_1232;
wire n_449;
wire n_734;
wire n_919;
wire n_763;
wire n_1174;
wire n_657;
wire n_583;
wire n_841;
wire n_582;
wire n_836;
wire n_561;
wire n_1096;
wire n_594;
wire n_531;
wire n_1136;
wire n_306;
wire n_1117;
wire n_1007;
wire n_424;
wire n_714;
wire n_932;
wire n_837;
wire n_1339;
wire n_1315;
wire n_867;
wire n_1070;
wire n_1270;
wire n_675;
wire n_504;
wire n_581;
wire n_698;
wire n_555;
wire n_834;
wire n_901;
wire n_727;
wire n_1038;
wire n_1162;
wire n_1103;
wire n_785;
wire n_375;
wire n_688;
wire n_323;
wire n_347;
wire n_515;
wire n_1290;
wire n_1234;
wire n_592;
wire n_1045;
wire n_1115;
wire n_521;
wire n_625;
wire n_585;
wire n_1190;
wire n_1237;
wire n_713;
wire n_457;
wire n_736;
wire n_606;
wire n_332;
wire n_1292;
wire n_421;
wire n_1148;
wire n_739;
wire n_1166;
wire n_987;
wire n_1086;
wire n_406;
wire n_1236;
wire n_791;
wire n_707;
wire n_603;
wire n_1261;
wire n_885;
wire n_500;
wire n_607;
wire n_496;
wire n_801;
wire n_1059;
wire n_309;
wire n_701;
wire n_612;
wire n_1032;
wire n_1284;
wire n_336;
wire n_464;
wire n_1243;
wire n_1196;
wire n_1338;
wire n_814;
wire n_985;
wire n_1191;
wire n_971;
wire n_904;
wire n_1301;
wire n_532;
wire n_400;
wire n_386;
wire n_432;
wire n_659;
wire n_1329;
wire n_316;
wire n_1185;
wire n_389;
wire n_436;
wire n_1217;
wire n_715;
wire n_330;
wire n_1087;
wire n_662;
wire n_617;
wire n_598;
wire n_732;
wire n_724;
wire n_599;
wire n_609;
wire n_909;
wire n_1273;
wire n_366;
wire n_1319;
wire n_596;
wire n_1215;
wire n_951;
wire n_321;
wire n_1024;
wire n_1016;
wire n_652;
wire n_333;
wire n_638;
wire n_563;
wire n_479;
wire n_623;
wire n_1222;
wire n_593;
wire n_872;
wire n_809;
wire n_1101;
wire n_1072;
wire n_865;
wire n_1064;
wire n_1254;
wire n_764;
wire n_426;
wire n_969;
wire n_417;
wire n_1253;
wire n_632;
wire n_1182;
wire n_828;
wire n_1138;
wire n_506;
wire n_381;
wire n_1255;
wire n_313;
wire n_322;
wire n_1299;
wire n_1332;
wire n_427;
wire n_703;
wire n_415;
wire n_1272;
wire n_928;
wire n_352;
wire n_882;
wire n_871;
wire n_803;
wire n_729;
wire n_805;
wire n_693;
wire n_1036;
wire n_1145;
wire n_651;
wire n_1303;
wire n_1320;
wire n_747;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_959;
wire n_719;
wire n_1206;
wire n_1257;
wire n_710;
wire n_1178;
wire n_546;
wire n_412;
wire n_664;
wire n_1249;
wire n_788;
wire n_403;
wire n_516;
wire n_549;
wire n_832;
wire n_996;
wire n_420;
wire n_1089;
wire n_1058;
wire n_388;
wire n_1082;
wire n_1052;
wire n_1055;
wire n_974;
wire n_591;
wire n_933;
wire n_1252;
wire n_416;
wire n_536;
wire n_1256;
wire n_1259;
wire n_1318;
wire n_956;
wire n_989;
wire n_754;
wire n_775;
wire n_616;
wire n_1227;
wire n_365;
wire n_495;
wire n_364;
wire n_566;
wire n_1144;
wire n_344;
wire n_503;
wire n_1279;
wire n_1152;
wire n_1068;
wire n_1149;
wire n_615;
wire n_1170;
wire n_804;
wire n_570;
wire n_1133;
wire n_1317;
wire n_440;
wire n_422;
wire n_679;
wire n_1131;
wire n_597;
wire n_1039;
wire n_835;
wire n_778;
wire n_1156;
wire n_1288;
wire n_1340;
wire n_1042;
wire n_1130;
wire n_584;
wire n_912;
wire n_1325;
wire n_1043;
wire n_1283;
wire n_346;
wire n_397;
wire n_1008;
wire n_1109;
wire n_1026;
wire n_1027;
wire n_1040;
wire n_569;
wire n_946;
wire n_960;
wire n_1168;
wire n_343;
wire n_458;
wire n_1084;
wire n_618;
wire n_341;
wire n_470;
wire n_1085;
wire n_1073;
wire n_868;
wire n_473;
wire n_991;
wire n_843;
wire n_1263;
wire n_538;
wire n_492;
wire n_1150;
wire n_1327;
wire n_368;
wire n_650;
wire n_469;
wire n_1187;
wire n_742;
wire n_913;
wire n_845;
wire n_891;
wire n_1134;
wire n_494;
wire n_372;
wire n_631;
wire n_934;
wire n_425;
wire n_562;
wire n_1192;
wire n_983;
wire n_781;
wire n_709;
wire n_1105;
wire n_408;
wire n_385;
wire n_1127;
wire n_1348;
wire n_1173;
wire n_663;
wire n_513;
wire n_1092;
wire n_1124;
wire n_1278;
wire n_998;
wire n_604;
wire n_1260;
wire n_755;
wire n_848;
wire n_1031;
wire n_1293;
wire n_1280;
wire n_1158;
wire n_328;
wire n_743;
wire n_757;
wire n_750;
wire n_448;
wire n_645;
wire n_348;
wire n_1022;
wire n_802;
wire n_353;
wire n_993;
wire n_1122;
wire n_1224;
wire n_383;
wire n_762;
wire n_981;
wire n_1095;
wire n_758;
wire n_544;
wire n_1175;
wire n_853;
wire n_765;
wire n_1177;
wire n_1310;
wire n_462;
wire n_1347;
wire n_783;
wire n_1074;
wire n_463;
wire n_1003;
wire n_678;
wire n_1200;
wire n_384;
wire n_978;
wire n_547;
wire n_1247;
wire n_628;
wire n_812;
wire n_777;
wire n_351;
wire n_401;
wire n_360;
wire n_345;
wire n_481;
wire n_443;
wire n_694;
wire n_1262;
wire n_1078;
wire n_702;
wire n_572;
wire n_1094;
wire n_1204;
wire n_392;
wire n_1169;
wire n_975;
wire n_326;
wire n_1081;
wire n_671;
wire n_540;
wire n_937;
wire n_1093;
wire n_955;
wire n_1275;
wire n_945;
wire n_554;
wire n_726;
wire n_712;
wire n_608;
wire n_567;
wire n_888;
wire n_529;
wire n_455;
wire n_1025;
wire n_1132;
wire n_630;
wire n_1180;
wire n_647;
wire n_844;
wire n_1160;
wire n_1245;
wire n_1195;
wire n_1241;
wire n_1302;
wire n_895;
wire n_798;
wire n_318;
wire n_887;
wire n_471;
wire n_1014;
wire n_665;
wire n_1154;
wire n_863;
wire n_1265;
wire n_730;
wire n_1212;
wire n_735;
wire n_1091;
wire n_784;
wire n_354;
wire n_1220;
wire n_893;
wire n_1028;
wire n_935;
wire n_910;
wire n_1046;
wire n_1183;
wire n_460;
wire n_813;
wire n_1076;
wire n_369;
wire n_1186;
wire n_1167;
wire n_674;
wire n_810;
wire n_982;
wire n_889;
wire n_689;
wire n_902;
wire n_1113;
wire n_1264;
wire n_760;
wire n_941;
wire n_362;
wire n_931;
wire n_827;
wire n_1218;
wire n_1343;
wire n_1041;
wire n_1080;
wire n_1126;
wire n_1151;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_1065;
wire n_622;
wire n_601;
wire n_1331;
wire n_1176;
wire n_649;
wire n_526;
wire n_1047;
wire n_320;
wire n_768;
wire n_869;
wire n_880;
wire n_621;
wire n_370;
wire n_589;
wire n_505;
wire n_682;
wire n_906;
wire n_357;
wire n_653;
wire n_881;
wire n_374;
wire n_718;
wire n_1238;
wire n_1114;
wire n_1286;
wire n_948;
wire n_1304;
wire n_1314;
wire n_717;
wire n_861;
wire n_654;
wire n_1221;
wire n_428;
wire n_794;
wire n_1268;
wire n_639;
wire n_1305;
wire n_552;
wire n_1023;
wire n_1057;
wire n_435;
wire n_1294;
wire n_1051;
wire n_1088;
wire n_851;
wire n_396;
wire n_445;
wire n_398;
wire n_656;
wire n_1230;
wire n_553;
wire n_325;
wire n_349;
wire n_1021;
wire n_749;
wire n_535;
wire n_1006;
wire n_1054;
wire n_1231;
wire n_358;
wire n_456;
wire n_962;
wire n_782;
wire n_524;
wire n_1044;
wire n_875;
wire n_497;
wire n_728;
wire n_339;
wire n_1239;
wire n_1335;
wire n_924;
wire n_378;
wire n_441;
wire n_1285;
wire n_1344;
wire n_335;
wire n_700;
wire n_534;
wire n_1296;
wire n_766;
wire n_602;
wire n_1143;
wire n_629;
wire n_1053;
wire n_1223;
wire n_967;
wire n_1258;
wire n_418;
wire n_380;
wire n_356;
wire n_600;
wire n_371;
wire n_820;
wire n_558;
wire n_670;
wire n_1004;
wire n_683;
wire n_929;
wire n_1111;
wire n_976;
wire n_695;
wire n_1104;
wire n_1120;
wire n_1219;
wire n_595;
wire n_759;
wire n_559;
wire n_480;
wire n_453;
wire n_833;
wire n_1146;
wire n_414;
wire n_1137;
wire n_916;
wire n_740;
wire n_772;
wire n_819;
wire n_405;
wire n_491;
wire n_1291;
BUFx3_ASAP7_75t_L g306 ( .A(n_175), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_141), .Y(n_307) );
INVx1_ASAP7_75t_SL g308 ( .A(n_174), .Y(n_308) );
INVx2_ASAP7_75t_L g309 ( .A(n_136), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_198), .Y(n_310) );
INVx2_ASAP7_75t_L g311 ( .A(n_294), .Y(n_311) );
CKINVDCx5p33_ASAP7_75t_R g312 ( .A(n_300), .Y(n_312) );
CKINVDCx20_ASAP7_75t_R g313 ( .A(n_285), .Y(n_313) );
BUFx3_ASAP7_75t_L g314 ( .A(n_295), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_103), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_227), .Y(n_316) );
CKINVDCx5p33_ASAP7_75t_R g317 ( .A(n_177), .Y(n_317) );
INVxp67_ASAP7_75t_SL g318 ( .A(n_49), .Y(n_318) );
HB1xp67_ASAP7_75t_L g319 ( .A(n_218), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_212), .Y(n_320) );
INVxp33_ASAP7_75t_L g321 ( .A(n_91), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_180), .Y(n_322) );
INVx2_ASAP7_75t_L g323 ( .A(n_296), .Y(n_323) );
BUFx10_ASAP7_75t_L g324 ( .A(n_43), .Y(n_324) );
INVx2_ASAP7_75t_L g325 ( .A(n_216), .Y(n_325) );
INVx2_ASAP7_75t_L g326 ( .A(n_40), .Y(n_326) );
BUFx6f_ASAP7_75t_L g327 ( .A(n_284), .Y(n_327) );
INVx1_ASAP7_75t_SL g328 ( .A(n_206), .Y(n_328) );
BUFx5_ASAP7_75t_L g329 ( .A(n_238), .Y(n_329) );
INVx2_ASAP7_75t_L g330 ( .A(n_43), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_228), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_213), .Y(n_332) );
OR2x2_ASAP7_75t_L g333 ( .A(n_149), .B(n_100), .Y(n_333) );
CKINVDCx5p33_ASAP7_75t_R g334 ( .A(n_193), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_118), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_15), .Y(n_336) );
CKINVDCx16_ASAP7_75t_R g337 ( .A(n_54), .Y(n_337) );
INVx2_ASAP7_75t_L g338 ( .A(n_225), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_36), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_18), .Y(n_340) );
INVxp67_ASAP7_75t_SL g341 ( .A(n_252), .Y(n_341) );
CKINVDCx14_ASAP7_75t_R g342 ( .A(n_205), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_131), .Y(n_343) );
CKINVDCx5p33_ASAP7_75t_R g344 ( .A(n_32), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_159), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_17), .Y(n_346) );
CKINVDCx20_ASAP7_75t_R g347 ( .A(n_219), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_163), .Y(n_348) );
CKINVDCx5p33_ASAP7_75t_R g349 ( .A(n_234), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_199), .Y(n_350) );
BUFx5_ASAP7_75t_L g351 ( .A(n_297), .Y(n_351) );
CKINVDCx5p33_ASAP7_75t_R g352 ( .A(n_214), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_268), .Y(n_353) );
BUFx10_ASAP7_75t_L g354 ( .A(n_200), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_292), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_178), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_190), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_223), .Y(n_358) );
CKINVDCx5p33_ASAP7_75t_R g359 ( .A(n_19), .Y(n_359) );
CKINVDCx5p33_ASAP7_75t_R g360 ( .A(n_293), .Y(n_360) );
CKINVDCx16_ASAP7_75t_R g361 ( .A(n_211), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_65), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_197), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_80), .Y(n_364) );
HB1xp67_ASAP7_75t_L g365 ( .A(n_170), .Y(n_365) );
CKINVDCx20_ASAP7_75t_R g366 ( .A(n_162), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_264), .Y(n_367) );
CKINVDCx5p33_ASAP7_75t_R g368 ( .A(n_210), .Y(n_368) );
INVx1_ASAP7_75t_SL g369 ( .A(n_109), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_286), .Y(n_370) );
INVxp67_ASAP7_75t_SL g371 ( .A(n_304), .Y(n_371) );
BUFx2_ASAP7_75t_SL g372 ( .A(n_103), .Y(n_372) );
INVx2_ASAP7_75t_L g373 ( .A(n_265), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_185), .Y(n_374) );
INVxp67_ASAP7_75t_SL g375 ( .A(n_251), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_165), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_22), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_146), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_261), .Y(n_379) );
INVxp67_ASAP7_75t_SL g380 ( .A(n_189), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_183), .Y(n_381) );
CKINVDCx20_ASAP7_75t_R g382 ( .A(n_275), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_241), .Y(n_383) );
CKINVDCx5p33_ASAP7_75t_R g384 ( .A(n_144), .Y(n_384) );
CKINVDCx5p33_ASAP7_75t_R g385 ( .A(n_2), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_117), .Y(n_386) );
CKINVDCx5p33_ASAP7_75t_R g387 ( .A(n_186), .Y(n_387) );
INVx2_ASAP7_75t_L g388 ( .A(n_271), .Y(n_388) );
INVxp67_ASAP7_75t_L g389 ( .A(n_68), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_224), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_105), .Y(n_391) );
INVx2_ASAP7_75t_L g392 ( .A(n_237), .Y(n_392) );
INVxp67_ASAP7_75t_SL g393 ( .A(n_158), .Y(n_393) );
CKINVDCx20_ASAP7_75t_R g394 ( .A(n_157), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_187), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_164), .Y(n_396) );
CKINVDCx20_ASAP7_75t_R g397 ( .A(n_208), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_263), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_41), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_118), .Y(n_400) );
CKINVDCx14_ASAP7_75t_R g401 ( .A(n_171), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_72), .Y(n_402) );
CKINVDCx20_ASAP7_75t_R g403 ( .A(n_76), .Y(n_403) );
INVx2_ASAP7_75t_L g404 ( .A(n_34), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_204), .Y(n_405) );
INVxp67_ASAP7_75t_SL g406 ( .A(n_96), .Y(n_406) );
BUFx6f_ASAP7_75t_L g407 ( .A(n_274), .Y(n_407) );
BUFx6f_ASAP7_75t_L g408 ( .A(n_99), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_131), .Y(n_409) );
XOR2xp5_ASAP7_75t_L g410 ( .A(n_188), .B(n_37), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_169), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_72), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_27), .Y(n_413) );
CKINVDCx5p33_ASAP7_75t_R g414 ( .A(n_47), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_24), .Y(n_415) );
CKINVDCx16_ASAP7_75t_R g416 ( .A(n_63), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_64), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_168), .Y(n_418) );
BUFx2_ASAP7_75t_L g419 ( .A(n_258), .Y(n_419) );
BUFx3_ASAP7_75t_L g420 ( .A(n_184), .Y(n_420) );
INVxp67_ASAP7_75t_L g421 ( .A(n_256), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_128), .Y(n_422) );
BUFx6f_ASAP7_75t_L g423 ( .A(n_182), .Y(n_423) );
CKINVDCx14_ASAP7_75t_R g424 ( .A(n_134), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_273), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_95), .Y(n_426) );
CKINVDCx20_ASAP7_75t_R g427 ( .A(n_92), .Y(n_427) );
BUFx2_ASAP7_75t_L g428 ( .A(n_181), .Y(n_428) );
CKINVDCx16_ASAP7_75t_R g429 ( .A(n_98), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_143), .Y(n_430) );
BUFx6f_ASAP7_75t_L g431 ( .A(n_260), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_46), .Y(n_432) );
CKINVDCx20_ASAP7_75t_R g433 ( .A(n_30), .Y(n_433) );
INVxp33_ASAP7_75t_SL g434 ( .A(n_58), .Y(n_434) );
BUFx2_ASAP7_75t_L g435 ( .A(n_83), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_25), .Y(n_436) );
INVx3_ASAP7_75t_L g437 ( .A(n_108), .Y(n_437) );
CKINVDCx5p33_ASAP7_75t_R g438 ( .A(n_255), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_122), .Y(n_439) );
INVx2_ASAP7_75t_L g440 ( .A(n_217), .Y(n_440) );
INVx2_ASAP7_75t_L g441 ( .A(n_4), .Y(n_441) );
CKINVDCx20_ASAP7_75t_R g442 ( .A(n_270), .Y(n_442) );
BUFx6f_ASAP7_75t_L g443 ( .A(n_25), .Y(n_443) );
CKINVDCx5p33_ASAP7_75t_R g444 ( .A(n_116), .Y(n_444) );
CKINVDCx5p33_ASAP7_75t_R g445 ( .A(n_226), .Y(n_445) );
CKINVDCx5p33_ASAP7_75t_R g446 ( .A(n_196), .Y(n_446) );
BUFx2_ASAP7_75t_L g447 ( .A(n_26), .Y(n_447) );
INVxp33_ASAP7_75t_SL g448 ( .A(n_35), .Y(n_448) );
CKINVDCx20_ASAP7_75t_R g449 ( .A(n_45), .Y(n_449) );
BUFx2_ASAP7_75t_SL g450 ( .A(n_176), .Y(n_450) );
BUFx2_ASAP7_75t_L g451 ( .A(n_114), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_230), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_109), .Y(n_453) );
INVx3_ASAP7_75t_L g454 ( .A(n_106), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_48), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_71), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_1), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_52), .Y(n_458) );
CKINVDCx5p33_ASAP7_75t_R g459 ( .A(n_107), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_66), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_2), .Y(n_461) );
CKINVDCx5p33_ASAP7_75t_R g462 ( .A(n_115), .Y(n_462) );
CKINVDCx5p33_ASAP7_75t_R g463 ( .A(n_281), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_51), .Y(n_464) );
CKINVDCx5p33_ASAP7_75t_R g465 ( .A(n_28), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_41), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_73), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_62), .Y(n_468) );
CKINVDCx5p33_ASAP7_75t_R g469 ( .A(n_128), .Y(n_469) );
CKINVDCx5p33_ASAP7_75t_R g470 ( .A(n_266), .Y(n_470) );
CKINVDCx20_ASAP7_75t_R g471 ( .A(n_5), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_50), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_97), .Y(n_473) );
CKINVDCx20_ASAP7_75t_R g474 ( .A(n_179), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_437), .Y(n_475) );
AND2x4_ASAP7_75t_L g476 ( .A(n_437), .B(n_0), .Y(n_476) );
OAI22xp5_ASAP7_75t_SL g477 ( .A1(n_403), .A2(n_3), .B1(n_0), .B2(n_1), .Y(n_477) );
BUFx6f_ASAP7_75t_L g478 ( .A(n_327), .Y(n_478) );
AOI22x1_ASAP7_75t_SL g479 ( .A1(n_403), .A2(n_5), .B1(n_3), .B2(n_4), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_454), .Y(n_480) );
CKINVDCx5p33_ASAP7_75t_R g481 ( .A(n_361), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_419), .B(n_6), .Y(n_482) );
AND2x2_ASAP7_75t_L g483 ( .A(n_321), .B(n_7), .Y(n_483) );
NOR2x1_ASAP7_75t_L g484 ( .A(n_454), .B(n_7), .Y(n_484) );
AND2x6_ASAP7_75t_L g485 ( .A(n_306), .B(n_133), .Y(n_485) );
INVx2_ASAP7_75t_L g486 ( .A(n_329), .Y(n_486) );
BUFx3_ASAP7_75t_L g487 ( .A(n_306), .Y(n_487) );
OA21x2_ASAP7_75t_L g488 ( .A1(n_309), .A2(n_137), .B(n_135), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_326), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_326), .Y(n_490) );
INVx4_ASAP7_75t_L g491 ( .A(n_428), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_321), .B(n_8), .Y(n_492) );
OAI22xp5_ASAP7_75t_SL g493 ( .A1(n_427), .A2(n_10), .B1(n_8), .B2(n_9), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_330), .Y(n_494) );
BUFx6f_ASAP7_75t_L g495 ( .A(n_327), .Y(n_495) );
BUFx6f_ASAP7_75t_L g496 ( .A(n_327), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_319), .B(n_9), .Y(n_497) );
CKINVDCx6p67_ASAP7_75t_R g498 ( .A(n_354), .Y(n_498) );
BUFx6f_ASAP7_75t_L g499 ( .A(n_327), .Y(n_499) );
INVx3_ASAP7_75t_L g500 ( .A(n_354), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_365), .B(n_10), .Y(n_501) );
AND2x2_ASAP7_75t_L g502 ( .A(n_435), .B(n_11), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_447), .B(n_11), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_451), .B(n_315), .Y(n_504) );
BUFx2_ASAP7_75t_L g505 ( .A(n_344), .Y(n_505) );
AND2x4_ASAP7_75t_SL g506 ( .A(n_354), .B(n_138), .Y(n_506) );
INVx4_ASAP7_75t_L g507 ( .A(n_314), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_330), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_404), .Y(n_509) );
BUFx6f_ASAP7_75t_L g510 ( .A(n_407), .Y(n_510) );
INVx2_ASAP7_75t_L g511 ( .A(n_329), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_404), .Y(n_512) );
AND2x2_ASAP7_75t_L g513 ( .A(n_337), .B(n_12), .Y(n_513) );
AND2x4_ASAP7_75t_L g514 ( .A(n_441), .B(n_12), .Y(n_514) );
INVx2_ASAP7_75t_L g515 ( .A(n_329), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_441), .Y(n_516) );
INVx2_ASAP7_75t_SL g517 ( .A(n_500), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_491), .B(n_344), .Y(n_518) );
OR2x2_ASAP7_75t_L g519 ( .A(n_505), .B(n_416), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_491), .B(n_444), .Y(n_520) );
NOR2xp33_ASAP7_75t_L g521 ( .A(n_491), .B(n_421), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_486), .Y(n_522) );
HB1xp67_ASAP7_75t_L g523 ( .A(n_505), .Y(n_523) );
BUFx10_ASAP7_75t_L g524 ( .A(n_506), .Y(n_524) );
INVx1_ASAP7_75t_SL g525 ( .A(n_498), .Y(n_525) );
AOI22xp33_ASAP7_75t_L g526 ( .A1(n_483), .A2(n_336), .B1(n_339), .B2(n_335), .Y(n_526) );
NOR2xp33_ASAP7_75t_L g527 ( .A(n_500), .B(n_307), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_486), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_500), .B(n_444), .Y(n_529) );
INVx5_ASAP7_75t_L g530 ( .A(n_485), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_486), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_498), .B(n_384), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_511), .Y(n_533) );
AND2x2_ASAP7_75t_SL g534 ( .A(n_506), .B(n_333), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_511), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_498), .B(n_384), .Y(n_536) );
CKINVDCx5p33_ASAP7_75t_R g537 ( .A(n_481), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_475), .B(n_438), .Y(n_538) );
BUFx6f_ASAP7_75t_L g539 ( .A(n_478), .Y(n_539) );
NOR2xp33_ASAP7_75t_L g540 ( .A(n_475), .B(n_480), .Y(n_540) );
NAND2xp5_ASAP7_75t_SL g541 ( .A(n_504), .B(n_438), .Y(n_541) );
AND2x2_ASAP7_75t_L g542 ( .A(n_483), .B(n_342), .Y(n_542) );
AOI22xp5_ASAP7_75t_L g543 ( .A1(n_502), .A2(n_434), .B1(n_448), .B2(n_429), .Y(n_543) );
AOI22xp5_ASAP7_75t_L g544 ( .A1(n_502), .A2(n_448), .B1(n_434), .B2(n_313), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_480), .B(n_445), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_511), .Y(n_546) );
INVx4_ASAP7_75t_L g547 ( .A(n_485), .Y(n_547) );
NOR2xp33_ASAP7_75t_L g548 ( .A(n_504), .B(n_310), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_515), .Y(n_549) );
NOR2xp33_ASAP7_75t_L g550 ( .A(n_507), .B(n_316), .Y(n_550) );
INVx3_ASAP7_75t_L g551 ( .A(n_476), .Y(n_551) );
AOI22xp33_ASAP7_75t_L g552 ( .A1(n_514), .A2(n_340), .B1(n_346), .B2(n_343), .Y(n_552) );
NAND2xp5_ASAP7_75t_SL g553 ( .A(n_476), .B(n_445), .Y(n_553) );
BUFx3_ASAP7_75t_L g554 ( .A(n_487), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_515), .Y(n_555) );
INVx3_ASAP7_75t_L g556 ( .A(n_476), .Y(n_556) );
NAND2xp5_ASAP7_75t_SL g557 ( .A(n_476), .B(n_446), .Y(n_557) );
NOR2xp33_ASAP7_75t_SL g558 ( .A(n_485), .B(n_313), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_542), .B(n_502), .Y(n_559) );
INVx2_ASAP7_75t_L g560 ( .A(n_554), .Y(n_560) );
NOR2xp33_ASAP7_75t_L g561 ( .A(n_529), .B(n_482), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_551), .Y(n_562) );
AOI22xp5_ASAP7_75t_L g563 ( .A1(n_534), .A2(n_513), .B1(n_492), .B2(n_482), .Y(n_563) );
AOI22xp5_ASAP7_75t_L g564 ( .A1(n_534), .A2(n_513), .B1(n_492), .B2(n_503), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_551), .Y(n_565) );
AND2x4_ASAP7_75t_L g566 ( .A(n_525), .B(n_506), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_548), .B(n_497), .Y(n_567) );
CKINVDCx5p33_ASAP7_75t_R g568 ( .A(n_537), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_518), .B(n_501), .Y(n_569) );
NOR2x2_ASAP7_75t_L g570 ( .A(n_544), .B(n_479), .Y(n_570) );
AOI22xp33_ASAP7_75t_L g571 ( .A1(n_556), .A2(n_514), .B1(n_485), .B2(n_515), .Y(n_571) );
INVx3_ASAP7_75t_L g572 ( .A(n_556), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_520), .B(n_501), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_521), .B(n_487), .Y(n_574) );
AOI22xp33_ASAP7_75t_L g575 ( .A1(n_556), .A2(n_514), .B1(n_485), .B2(n_484), .Y(n_575) );
BUFx6f_ASAP7_75t_L g576 ( .A(n_547), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_538), .B(n_487), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_545), .B(n_507), .Y(n_578) );
INVx2_ASAP7_75t_L g579 ( .A(n_517), .Y(n_579) );
NAND2x1p5_ASAP7_75t_L g580 ( .A(n_534), .B(n_514), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_532), .B(n_507), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_536), .B(n_507), .Y(n_582) );
OR2x6_ASAP7_75t_L g583 ( .A(n_519), .B(n_477), .Y(n_583) );
AOI22xp33_ASAP7_75t_SL g584 ( .A1(n_558), .A2(n_479), .B1(n_493), .B2(n_477), .Y(n_584) );
AOI22xp5_ASAP7_75t_L g585 ( .A1(n_543), .A2(n_503), .B1(n_347), .B2(n_382), .Y(n_585) );
AOI21xp5_ASAP7_75t_L g586 ( .A1(n_553), .A2(n_488), .B(n_484), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_541), .B(n_446), .Y(n_587) );
AOI22xp5_ASAP7_75t_L g588 ( .A1(n_543), .A2(n_347), .B1(n_382), .B2(n_366), .Y(n_588) );
O2A1O1Ixp33_ASAP7_75t_L g589 ( .A1(n_557), .A2(n_490), .B(n_494), .C(n_489), .Y(n_589) );
HB1xp67_ASAP7_75t_L g590 ( .A(n_523), .Y(n_590) );
BUFx3_ASAP7_75t_L g591 ( .A(n_537), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_517), .Y(n_592) );
NOR2xp33_ASAP7_75t_L g593 ( .A(n_527), .B(n_489), .Y(n_593) );
BUFx3_ASAP7_75t_L g594 ( .A(n_524), .Y(n_594) );
INVx2_ASAP7_75t_SL g595 ( .A(n_524), .Y(n_595) );
AOI21xp5_ASAP7_75t_L g596 ( .A1(n_550), .A2(n_488), .B(n_311), .Y(n_596) );
NOR2xp33_ASAP7_75t_L g597 ( .A(n_519), .B(n_342), .Y(n_597) );
AND2x2_ASAP7_75t_L g598 ( .A(n_544), .B(n_324), .Y(n_598) );
NOR2xp33_ASAP7_75t_L g599 ( .A(n_540), .B(n_490), .Y(n_599) );
NAND2xp5_ASAP7_75t_SL g600 ( .A(n_524), .B(n_312), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_552), .B(n_401), .Y(n_601) );
BUFx3_ASAP7_75t_L g602 ( .A(n_522), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_522), .Y(n_603) );
NOR2xp33_ASAP7_75t_L g604 ( .A(n_526), .B(n_401), .Y(n_604) );
BUFx3_ASAP7_75t_L g605 ( .A(n_528), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_528), .B(n_424), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_531), .B(n_424), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_531), .Y(n_608) );
NAND2xp5_ASAP7_75t_SL g609 ( .A(n_547), .B(n_317), .Y(n_609) );
AND2x2_ASAP7_75t_L g610 ( .A(n_533), .B(n_324), .Y(n_610) );
NOR2xp33_ASAP7_75t_L g611 ( .A(n_555), .B(n_508), .Y(n_611) );
INVxp67_ASAP7_75t_L g612 ( .A(n_555), .Y(n_612) );
AND2x2_ASAP7_75t_L g613 ( .A(n_533), .B(n_324), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_535), .B(n_516), .Y(n_614) );
OR2x2_ASAP7_75t_L g615 ( .A(n_546), .B(n_493), .Y(n_615) );
INVx8_ASAP7_75t_L g616 ( .A(n_530), .Y(n_616) );
BUFx5_ASAP7_75t_L g617 ( .A(n_549), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_549), .B(n_512), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_530), .B(n_508), .Y(n_619) );
BUFx6f_ASAP7_75t_SL g620 ( .A(n_539), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_530), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_530), .B(n_509), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_530), .B(n_509), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_530), .B(n_334), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_539), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_539), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_539), .B(n_349), .Y(n_627) );
NAND2xp5_ASAP7_75t_SL g628 ( .A(n_539), .B(n_352), .Y(n_628) );
INVx2_ASAP7_75t_L g629 ( .A(n_554), .Y(n_629) );
NAND2x1_ASAP7_75t_L g630 ( .A(n_551), .B(n_485), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_542), .B(n_360), .Y(n_631) );
AND2x4_ASAP7_75t_L g632 ( .A(n_525), .B(n_394), .Y(n_632) );
NOR2xp33_ASAP7_75t_L g633 ( .A(n_529), .B(n_320), .Y(n_633) );
INVx3_ASAP7_75t_L g634 ( .A(n_551), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_542), .B(n_368), .Y(n_635) );
INVx2_ASAP7_75t_L g636 ( .A(n_554), .Y(n_636) );
OR2x6_ASAP7_75t_L g637 ( .A(n_519), .B(n_372), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_542), .Y(n_638) );
AOI21xp5_ASAP7_75t_L g639 ( .A1(n_586), .A2(n_488), .B(n_371), .Y(n_639) );
NOR2xp33_ASAP7_75t_L g640 ( .A(n_564), .B(n_397), .Y(n_640) );
AOI21xp5_ASAP7_75t_L g641 ( .A1(n_586), .A2(n_488), .B(n_375), .Y(n_641) );
BUFx6f_ASAP7_75t_L g642 ( .A(n_616), .Y(n_642) );
OA22x2_ASAP7_75t_L g643 ( .A1(n_588), .A2(n_410), .B1(n_433), .B2(n_427), .Y(n_643) );
NOR2xp33_ASAP7_75t_R g644 ( .A(n_568), .B(n_442), .Y(n_644) );
NAND2xp5_ASAP7_75t_SL g645 ( .A(n_617), .B(n_442), .Y(n_645) );
AOI21xp5_ASAP7_75t_L g646 ( .A1(n_596), .A2(n_488), .B(n_380), .Y(n_646) );
NAND2xp5_ASAP7_75t_SL g647 ( .A(n_617), .B(n_474), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_572), .Y(n_648) );
AOI22xp33_ASAP7_75t_L g649 ( .A1(n_580), .A2(n_449), .B1(n_471), .B2(n_433), .Y(n_649) );
AOI33xp33_ASAP7_75t_L g650 ( .A1(n_584), .A2(n_377), .A3(n_364), .B1(n_391), .B2(n_386), .B3(n_362), .Y(n_650) );
AND2x4_ASAP7_75t_L g651 ( .A(n_594), .B(n_318), .Y(n_651) );
INVx2_ASAP7_75t_L g652 ( .A(n_602), .Y(n_652) );
AOI21xp5_ASAP7_75t_L g653 ( .A1(n_596), .A2(n_393), .B(n_341), .Y(n_653) );
AOI21xp5_ASAP7_75t_L g654 ( .A1(n_569), .A2(n_331), .B(n_322), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_567), .B(n_389), .Y(n_655) );
AOI21xp5_ASAP7_75t_L g656 ( .A1(n_573), .A2(n_345), .B(n_332), .Y(n_656) );
AOI21xp5_ASAP7_75t_L g657 ( .A1(n_581), .A2(n_350), .B(n_348), .Y(n_657) );
AOI22xp5_ASAP7_75t_L g658 ( .A1(n_563), .A2(n_474), .B1(n_385), .B2(n_414), .Y(n_658) );
INVxp67_ASAP7_75t_L g659 ( .A(n_590), .Y(n_659) );
AOI21xp5_ASAP7_75t_L g660 ( .A1(n_582), .A2(n_355), .B(n_353), .Y(n_660) );
INVx1_ASAP7_75t_L g661 ( .A(n_634), .Y(n_661) );
A2O1A1Ixp33_ASAP7_75t_L g662 ( .A1(n_561), .A2(n_400), .B(n_402), .C(n_399), .Y(n_662) );
NOR2xp33_ASAP7_75t_L g663 ( .A(n_637), .B(n_449), .Y(n_663) );
INVx2_ASAP7_75t_SL g664 ( .A(n_590), .Y(n_664) );
AND2x2_ASAP7_75t_L g665 ( .A(n_598), .B(n_471), .Y(n_665) );
AOI21xp5_ASAP7_75t_L g666 ( .A1(n_578), .A2(n_357), .B(n_356), .Y(n_666) );
NOR2xp33_ASAP7_75t_L g667 ( .A(n_637), .B(n_359), .Y(n_667) );
AOI22xp5_ASAP7_75t_L g668 ( .A1(n_561), .A2(n_485), .B1(n_406), .B2(n_412), .Y(n_668) );
OR2x6_ASAP7_75t_L g669 ( .A(n_632), .B(n_450), .Y(n_669) );
O2A1O1Ixp5_ASAP7_75t_L g670 ( .A1(n_630), .A2(n_309), .B(n_323), .C(n_311), .Y(n_670) );
NOR2xp33_ASAP7_75t_R g671 ( .A(n_591), .B(n_595), .Y(n_671) );
OAI22xp5_ASAP7_75t_L g672 ( .A1(n_580), .A2(n_409), .B1(n_415), .B2(n_413), .Y(n_672) );
INVx2_ASAP7_75t_L g673 ( .A(n_605), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_559), .B(n_459), .Y(n_674) );
BUFx6f_ASAP7_75t_L g675 ( .A(n_616), .Y(n_675) );
A2O1A1Ixp33_ASAP7_75t_SL g676 ( .A1(n_633), .A2(n_325), .B(n_338), .C(n_323), .Y(n_676) );
NOR2xp67_ASAP7_75t_L g677 ( .A(n_612), .B(n_139), .Y(n_677) );
NOR2xp33_ASAP7_75t_R g678 ( .A(n_632), .B(n_462), .Y(n_678) );
OR2x6_ASAP7_75t_L g679 ( .A(n_583), .B(n_417), .Y(n_679) );
OAI21xp5_ASAP7_75t_L g680 ( .A1(n_571), .A2(n_485), .B(n_363), .Y(n_680) );
AO21x2_ASAP7_75t_L g681 ( .A1(n_606), .A2(n_367), .B(n_358), .Y(n_681) );
BUFx2_ASAP7_75t_L g682 ( .A(n_637), .Y(n_682) );
AOI21xp5_ASAP7_75t_L g683 ( .A1(n_574), .A2(n_374), .B(n_370), .Y(n_683) );
AND2x2_ASAP7_75t_L g684 ( .A(n_585), .B(n_369), .Y(n_684) );
OAI22xp5_ASAP7_75t_SL g685 ( .A1(n_584), .A2(n_469), .B1(n_465), .B2(n_426), .Y(n_685) );
BUFx3_ASAP7_75t_L g686 ( .A(n_617), .Y(n_686) );
AOI21xp33_ASAP7_75t_L g687 ( .A1(n_604), .A2(n_328), .B(n_308), .Y(n_687) );
INVx2_ASAP7_75t_L g688 ( .A(n_562), .Y(n_688) );
AND2x6_ASAP7_75t_L g689 ( .A(n_566), .B(n_314), .Y(n_689) );
NOR2xp33_ASAP7_75t_L g690 ( .A(n_597), .B(n_422), .Y(n_690) );
OR2x6_ASAP7_75t_L g691 ( .A(n_583), .B(n_615), .Y(n_691) );
A2O1A1Ixp33_ASAP7_75t_L g692 ( .A1(n_633), .A2(n_436), .B(n_439), .C(n_432), .Y(n_692) );
BUFx12f_ASAP7_75t_L g693 ( .A(n_583), .Y(n_693) );
BUFx6f_ASAP7_75t_L g694 ( .A(n_616), .Y(n_694) );
INVx2_ASAP7_75t_L g695 ( .A(n_565), .Y(n_695) );
AOI22xp5_ASAP7_75t_L g696 ( .A1(n_610), .A2(n_613), .B1(n_566), .B2(n_638), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_599), .B(n_453), .Y(n_697) );
BUFx2_ASAP7_75t_L g698 ( .A(n_570), .Y(n_698) );
INVx4_ASAP7_75t_L g699 ( .A(n_620), .Y(n_699) );
NOR2xp33_ASAP7_75t_L g700 ( .A(n_587), .B(n_455), .Y(n_700) );
AOI22xp33_ASAP7_75t_L g701 ( .A1(n_603), .A2(n_485), .B1(n_457), .B2(n_458), .Y(n_701) );
INVx1_ASAP7_75t_L g702 ( .A(n_611), .Y(n_702) );
HB1xp67_ASAP7_75t_L g703 ( .A(n_614), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_599), .B(n_456), .Y(n_704) );
INVx1_ASAP7_75t_L g705 ( .A(n_611), .Y(n_705) );
AOI21xp5_ASAP7_75t_L g706 ( .A1(n_577), .A2(n_378), .B(n_376), .Y(n_706) );
CKINVDCx20_ASAP7_75t_R g707 ( .A(n_600), .Y(n_707) );
NAND2x1p5_ASAP7_75t_L g708 ( .A(n_608), .B(n_460), .Y(n_708) );
BUFx2_ASAP7_75t_L g709 ( .A(n_631), .Y(n_709) );
INVx4_ASAP7_75t_L g710 ( .A(n_620), .Y(n_710) );
BUFx6f_ASAP7_75t_L g711 ( .A(n_576), .Y(n_711) );
NOR2xp33_ASAP7_75t_L g712 ( .A(n_635), .B(n_461), .Y(n_712) );
INVx2_ASAP7_75t_L g713 ( .A(n_560), .Y(n_713) );
AOI21xp5_ASAP7_75t_L g714 ( .A1(n_607), .A2(n_381), .B(n_379), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_593), .B(n_464), .Y(n_715) );
OAI22xp5_ASAP7_75t_SL g716 ( .A1(n_601), .A2(n_467), .B1(n_468), .B2(n_466), .Y(n_716) );
NOR2xp33_ASAP7_75t_L g717 ( .A(n_592), .B(n_472), .Y(n_717) );
NAND2xp5_ASAP7_75t_SL g718 ( .A(n_576), .B(n_387), .Y(n_718) );
OAI22xp5_ASAP7_75t_L g719 ( .A1(n_571), .A2(n_473), .B1(n_443), .B2(n_408), .Y(n_719) );
BUFx5_ASAP7_75t_L g720 ( .A(n_621), .Y(n_720) );
OAI21xp5_ASAP7_75t_L g721 ( .A1(n_575), .A2(n_390), .B(n_383), .Y(n_721) );
INVx4_ASAP7_75t_L g722 ( .A(n_579), .Y(n_722) );
NOR2xp33_ASAP7_75t_SL g723 ( .A(n_589), .B(n_463), .Y(n_723) );
INVx1_ASAP7_75t_L g724 ( .A(n_618), .Y(n_724) );
BUFx8_ASAP7_75t_L g725 ( .A(n_629), .Y(n_725) );
INVx2_ASAP7_75t_L g726 ( .A(n_636), .Y(n_726) );
OR2x6_ASAP7_75t_L g727 ( .A(n_628), .B(n_408), .Y(n_727) );
OAI22xp5_ASAP7_75t_L g728 ( .A1(n_609), .A2(n_622), .B1(n_623), .B2(n_619), .Y(n_728) );
INVxp67_ASAP7_75t_L g729 ( .A(n_627), .Y(n_729) );
NOR2xp33_ASAP7_75t_L g730 ( .A(n_624), .B(n_470), .Y(n_730) );
AND2x4_ASAP7_75t_L g731 ( .A(n_625), .B(n_395), .Y(n_731) );
AOI21xp5_ASAP7_75t_L g732 ( .A1(n_626), .A2(n_398), .B(n_396), .Y(n_732) );
OR2x6_ASAP7_75t_L g733 ( .A(n_632), .B(n_408), .Y(n_733) );
BUFx2_ASAP7_75t_L g734 ( .A(n_590), .Y(n_734) );
OAI21x1_ASAP7_75t_L g735 ( .A1(n_596), .A2(n_338), .B(n_325), .Y(n_735) );
A2O1A1Ixp33_ASAP7_75t_L g736 ( .A1(n_561), .A2(n_411), .B(n_418), .C(n_405), .Y(n_736) );
O2A1O1Ixp33_ASAP7_75t_L g737 ( .A1(n_567), .A2(n_430), .B(n_452), .C(n_425), .Y(n_737) );
CKINVDCx5p33_ASAP7_75t_R g738 ( .A(n_568), .Y(n_738) );
O2A1O1Ixp5_ASAP7_75t_L g739 ( .A1(n_586), .A2(n_388), .B(n_392), .C(n_373), .Y(n_739) );
AOI21xp5_ASAP7_75t_L g740 ( .A1(n_586), .A2(n_388), .B(n_373), .Y(n_740) );
NOR2xp33_ASAP7_75t_R g741 ( .A(n_568), .B(n_13), .Y(n_741) );
BUFx3_ASAP7_75t_L g742 ( .A(n_591), .Y(n_742) );
A2O1A1Ixp33_ASAP7_75t_L g743 ( .A1(n_561), .A2(n_440), .B(n_392), .C(n_420), .Y(n_743) );
NAND2xp5_ASAP7_75t_SL g744 ( .A(n_617), .B(n_440), .Y(n_744) );
NAND2xp5_ASAP7_75t_L g745 ( .A(n_567), .B(n_443), .Y(n_745) );
NOR2xp33_ASAP7_75t_R g746 ( .A(n_568), .B(n_14), .Y(n_746) );
BUFx3_ASAP7_75t_L g747 ( .A(n_591), .Y(n_747) );
AND2x2_ASAP7_75t_L g748 ( .A(n_590), .B(n_443), .Y(n_748) );
AND2x6_ASAP7_75t_L g749 ( .A(n_594), .B(n_420), .Y(n_749) );
BUFx3_ASAP7_75t_L g750 ( .A(n_591), .Y(n_750) );
A2O1A1Ixp33_ASAP7_75t_L g751 ( .A1(n_561), .A2(n_423), .B(n_431), .C(n_407), .Y(n_751) );
AOI21xp5_ASAP7_75t_L g752 ( .A1(n_586), .A2(n_423), .B(n_407), .Y(n_752) );
NOR2xp33_ASAP7_75t_L g753 ( .A(n_640), .B(n_14), .Y(n_753) );
OAI211xp5_ASAP7_75t_L g754 ( .A1(n_687), .A2(n_423), .B(n_431), .C(n_407), .Y(n_754) );
A2O1A1Ixp33_ASAP7_75t_L g755 ( .A1(n_737), .A2(n_431), .B(n_423), .C(n_478), .Y(n_755) );
INVx1_ASAP7_75t_L g756 ( .A(n_748), .Y(n_756) );
AO31x2_ASAP7_75t_L g757 ( .A1(n_752), .A2(n_495), .A3(n_496), .B(n_478), .Y(n_757) );
AOI22xp33_ASAP7_75t_SL g758 ( .A1(n_644), .A2(n_351), .B1(n_329), .B2(n_20), .Y(n_758) );
AND2x4_ASAP7_75t_L g759 ( .A(n_664), .B(n_16), .Y(n_759) );
O2A1O1Ixp33_ASAP7_75t_SL g760 ( .A1(n_676), .A2(n_351), .B(n_329), .C(n_142), .Y(n_760) );
INVx1_ASAP7_75t_L g761 ( .A(n_708), .Y(n_761) );
A2O1A1Ixp33_ASAP7_75t_L g762 ( .A1(n_714), .A2(n_495), .B(n_496), .C(n_478), .Y(n_762) );
AOI21xp5_ASAP7_75t_SL g763 ( .A1(n_686), .A2(n_495), .B(n_478), .Y(n_763) );
AOI21xp5_ASAP7_75t_L g764 ( .A1(n_639), .A2(n_510), .B(n_496), .Y(n_764) );
AOI21xp5_ASAP7_75t_L g765 ( .A1(n_641), .A2(n_496), .B(n_495), .Y(n_765) );
OAI21xp5_ASAP7_75t_L g766 ( .A1(n_739), .A2(n_351), .B(n_329), .Y(n_766) );
A2O1A1Ixp33_ASAP7_75t_L g767 ( .A1(n_653), .A2(n_495), .B(n_499), .C(n_496), .Y(n_767) );
AND2x4_ASAP7_75t_L g768 ( .A(n_696), .B(n_21), .Y(n_768) );
AO31x2_ASAP7_75t_L g769 ( .A1(n_646), .A2(n_496), .A3(n_510), .B(n_499), .Y(n_769) );
NAND3xp33_ASAP7_75t_L g770 ( .A(n_690), .B(n_510), .C(n_499), .Y(n_770) );
NOR2xp33_ASAP7_75t_L g771 ( .A(n_663), .B(n_21), .Y(n_771) );
INVx3_ASAP7_75t_SL g772 ( .A(n_738), .Y(n_772) );
NOR2xp33_ASAP7_75t_L g773 ( .A(n_665), .B(n_23), .Y(n_773) );
AOI21xp5_ASAP7_75t_L g774 ( .A1(n_744), .A2(n_510), .B(n_499), .Y(n_774) );
AOI22xp5_ASAP7_75t_L g775 ( .A1(n_659), .A2(n_351), .B1(n_26), .B2(n_23), .Y(n_775) );
NAND3xp33_ASAP7_75t_L g776 ( .A(n_751), .B(n_351), .C(n_24), .Y(n_776) );
INVx2_ASAP7_75t_L g777 ( .A(n_688), .Y(n_777) );
INVx1_ASAP7_75t_L g778 ( .A(n_724), .Y(n_778) );
INVx2_ASAP7_75t_L g779 ( .A(n_695), .Y(n_779) );
OA21x2_ASAP7_75t_L g780 ( .A1(n_735), .A2(n_145), .B(n_140), .Y(n_780) );
OAI21x1_ASAP7_75t_L g781 ( .A1(n_740), .A2(n_148), .B(n_147), .Y(n_781) );
HB1xp67_ASAP7_75t_L g782 ( .A(n_733), .Y(n_782) );
OAI22x1_ASAP7_75t_L g783 ( .A1(n_698), .A2(n_29), .B1(n_27), .B2(n_28), .Y(n_783) );
O2A1O1Ixp33_ASAP7_75t_L g784 ( .A1(n_692), .A2(n_31), .B(n_29), .C(n_30), .Y(n_784) );
AND2x6_ASAP7_75t_SL g785 ( .A(n_691), .B(n_32), .Y(n_785) );
INVx1_ASAP7_75t_SL g786 ( .A(n_678), .Y(n_786) );
OAI21xp5_ASAP7_75t_L g787 ( .A1(n_670), .A2(n_151), .B(n_150), .Y(n_787) );
AOI221x1_ASAP7_75t_L g788 ( .A1(n_743), .A2(n_33), .B1(n_38), .B2(n_39), .C(n_40), .Y(n_788) );
AO31x2_ASAP7_75t_L g789 ( .A1(n_719), .A2(n_42), .A3(n_38), .B(n_39), .Y(n_789) );
BUFx2_ASAP7_75t_R g790 ( .A(n_742), .Y(n_790) );
BUFx3_ASAP7_75t_L g791 ( .A(n_725), .Y(n_791) );
O2A1O1Ixp33_ASAP7_75t_SL g792 ( .A1(n_736), .A2(n_153), .B(n_154), .C(n_152), .Y(n_792) );
AOI22xp33_ASAP7_75t_L g793 ( .A1(n_643), .A2(n_45), .B1(n_42), .B2(n_44), .Y(n_793) );
NOR2xp33_ASAP7_75t_L g794 ( .A(n_658), .B(n_44), .Y(n_794) );
A2O1A1Ixp33_ASAP7_75t_L g795 ( .A1(n_654), .A2(n_656), .B(n_712), .C(n_700), .Y(n_795) );
OAI21xp5_ASAP7_75t_L g796 ( .A1(n_680), .A2(n_156), .B(n_155), .Y(n_796) );
BUFx2_ASAP7_75t_L g797 ( .A(n_725), .Y(n_797) );
INVx1_ASAP7_75t_L g798 ( .A(n_745), .Y(n_798) );
CKINVDCx5p33_ASAP7_75t_R g799 ( .A(n_671), .Y(n_799) );
NAND2xp5_ASAP7_75t_L g800 ( .A(n_705), .B(n_47), .Y(n_800) );
INVx5_ASAP7_75t_L g801 ( .A(n_642), .Y(n_801) );
A2O1A1Ixp33_ASAP7_75t_L g802 ( .A1(n_666), .A2(n_52), .B(n_50), .C(n_51), .Y(n_802) );
AO31x2_ASAP7_75t_L g803 ( .A1(n_717), .A2(n_55), .A3(n_53), .B(n_54), .Y(n_803) );
NOR2x1_ASAP7_75t_R g804 ( .A(n_693), .B(n_53), .Y(n_804) );
OAI21xp5_ASAP7_75t_L g805 ( .A1(n_668), .A2(n_161), .B(n_160), .Y(n_805) );
A2O1A1Ixp33_ASAP7_75t_L g806 ( .A1(n_657), .A2(n_660), .B(n_721), .C(n_683), .Y(n_806) );
AND2x2_ASAP7_75t_L g807 ( .A(n_684), .B(n_55), .Y(n_807) );
HB1xp67_ASAP7_75t_L g808 ( .A(n_747), .Y(n_808) );
BUFx2_ASAP7_75t_L g809 ( .A(n_750), .Y(n_809) );
AOI22xp33_ASAP7_75t_L g810 ( .A1(n_679), .A2(n_58), .B1(n_56), .B2(n_57), .Y(n_810) );
AOI22xp33_ASAP7_75t_L g811 ( .A1(n_679), .A2(n_59), .B1(n_56), .B2(n_57), .Y(n_811) );
NOR2xp33_ASAP7_75t_L g812 ( .A(n_669), .B(n_59), .Y(n_812) );
NAND2xp5_ASAP7_75t_L g813 ( .A(n_650), .B(n_60), .Y(n_813) );
AO31x2_ASAP7_75t_L g814 ( .A1(n_728), .A2(n_62), .A3(n_60), .B(n_61), .Y(n_814) );
OAI22xp5_ASAP7_75t_L g815 ( .A1(n_645), .A2(n_61), .B1(n_63), .B2(n_64), .Y(n_815) );
BUFx2_ASAP7_75t_L g816 ( .A(n_689), .Y(n_816) );
NOR2xp33_ASAP7_75t_L g817 ( .A(n_669), .B(n_682), .Y(n_817) );
OAI21xp5_ASAP7_75t_L g818 ( .A1(n_668), .A2(n_167), .B(n_166), .Y(n_818) );
AO21x2_ASAP7_75t_L g819 ( .A1(n_677), .A2(n_173), .B(n_172), .Y(n_819) );
AND2x4_ASAP7_75t_L g820 ( .A(n_642), .B(n_67), .Y(n_820) );
O2A1O1Ixp33_ASAP7_75t_L g821 ( .A1(n_672), .A2(n_704), .B(n_697), .C(n_715), .Y(n_821) );
AOI221xp5_ASAP7_75t_L g822 ( .A1(n_655), .A2(n_69), .B1(n_70), .B2(n_71), .C(n_73), .Y(n_822) );
A2O1A1Ixp33_ASAP7_75t_L g823 ( .A1(n_706), .A2(n_69), .B(n_70), .C(n_74), .Y(n_823) );
AOI221xp5_ASAP7_75t_SL g824 ( .A1(n_716), .A2(n_685), .B1(n_729), .B2(n_674), .C(n_647), .Y(n_824) );
CKINVDCx20_ASAP7_75t_R g825 ( .A(n_741), .Y(n_825) );
AND2x4_ASAP7_75t_L g826 ( .A(n_675), .B(n_74), .Y(n_826) );
AOI22xp33_ASAP7_75t_L g827 ( .A1(n_691), .A2(n_75), .B1(n_76), .B2(n_77), .Y(n_827) );
INVxp67_ASAP7_75t_L g828 ( .A(n_709), .Y(n_828) );
AO31x2_ASAP7_75t_L g829 ( .A1(n_732), .A2(n_78), .A3(n_79), .B(n_80), .Y(n_829) );
AOI22xp5_ASAP7_75t_L g830 ( .A1(n_649), .A2(n_667), .B1(n_707), .B2(n_689), .Y(n_830) );
HB1xp67_ASAP7_75t_L g831 ( .A(n_699), .Y(n_831) );
INVx2_ASAP7_75t_SL g832 ( .A(n_710), .Y(n_832) );
CKINVDCx5p33_ASAP7_75t_R g833 ( .A(n_746), .Y(n_833) );
NAND2xp5_ASAP7_75t_L g834 ( .A(n_689), .B(n_79), .Y(n_834) );
INVx2_ASAP7_75t_L g835 ( .A(n_713), .Y(n_835) );
INVx2_ASAP7_75t_L g836 ( .A(n_726), .Y(n_836) );
INVx2_ASAP7_75t_L g837 ( .A(n_711), .Y(n_837) );
INVx1_ASAP7_75t_L g838 ( .A(n_652), .Y(n_838) );
NAND2xp5_ASAP7_75t_L g839 ( .A(n_689), .B(n_81), .Y(n_839) );
AOI21xp5_ASAP7_75t_L g840 ( .A1(n_648), .A2(n_192), .B(n_191), .Y(n_840) );
AND2x2_ASAP7_75t_L g841 ( .A(n_651), .B(n_82), .Y(n_841) );
INVx1_ASAP7_75t_L g842 ( .A(n_673), .Y(n_842) );
NOR2xp33_ASAP7_75t_L g843 ( .A(n_651), .B(n_82), .Y(n_843) );
INVx2_ASAP7_75t_SL g844 ( .A(n_710), .Y(n_844) );
AOI22xp33_ASAP7_75t_L g845 ( .A1(n_681), .A2(n_84), .B1(n_85), .B2(n_86), .Y(n_845) );
NAND2xp5_ASAP7_75t_SL g846 ( .A(n_675), .B(n_86), .Y(n_846) );
O2A1O1Ixp33_ASAP7_75t_SL g847 ( .A1(n_661), .A2(n_233), .B(n_303), .C(n_302), .Y(n_847) );
O2A1O1Ixp33_ASAP7_75t_L g848 ( .A1(n_718), .A2(n_87), .B(n_88), .C(n_89), .Y(n_848) );
INVx4_ASAP7_75t_L g849 ( .A(n_694), .Y(n_849) );
AOI21xp5_ASAP7_75t_L g850 ( .A1(n_681), .A2(n_195), .B(n_194), .Y(n_850) );
OAI22xp5_ASAP7_75t_L g851 ( .A1(n_731), .A2(n_90), .B1(n_91), .B2(n_92), .Y(n_851) );
INVx1_ASAP7_75t_L g852 ( .A(n_722), .Y(n_852) );
BUFx12f_ASAP7_75t_L g853 ( .A(n_749), .Y(n_853) );
BUFx8_ASAP7_75t_L g854 ( .A(n_749), .Y(n_854) );
BUFx8_ASAP7_75t_L g855 ( .A(n_749), .Y(n_855) );
OAI21x1_ASAP7_75t_SL g856 ( .A1(n_722), .A2(n_93), .B(n_94), .Y(n_856) );
O2A1O1Ixp33_ASAP7_75t_SL g857 ( .A1(n_730), .A2(n_236), .B(n_301), .C(n_299), .Y(n_857) );
A2O1A1Ixp33_ASAP7_75t_L g858 ( .A1(n_723), .A2(n_93), .B(n_94), .C(n_95), .Y(n_858) );
A2O1A1Ixp33_ASAP7_75t_L g859 ( .A1(n_701), .A2(n_711), .B(n_694), .C(n_749), .Y(n_859) );
CKINVDCx5p33_ASAP7_75t_R g860 ( .A(n_727), .Y(n_860) );
OAI21x1_ASAP7_75t_L g861 ( .A1(n_720), .A2(n_243), .B(n_298), .Y(n_861) );
O2A1O1Ixp33_ASAP7_75t_L g862 ( .A1(n_720), .A2(n_101), .B(n_102), .C(n_104), .Y(n_862) );
AOI22xp5_ASAP7_75t_SL g863 ( .A1(n_698), .A2(n_101), .B1(n_102), .B2(n_104), .Y(n_863) );
A2O1A1Ixp33_ASAP7_75t_L g864 ( .A1(n_737), .A2(n_107), .B(n_108), .C(n_110), .Y(n_864) );
A2O1A1Ixp33_ASAP7_75t_L g865 ( .A1(n_737), .A2(n_110), .B(n_111), .C(n_112), .Y(n_865) );
INVx2_ASAP7_75t_SL g866 ( .A(n_725), .Y(n_866) );
NAND3xp33_ASAP7_75t_L g867 ( .A(n_690), .B(n_111), .C(n_112), .Y(n_867) );
BUFx6f_ASAP7_75t_L g868 ( .A(n_642), .Y(n_868) );
AO31x2_ASAP7_75t_L g869 ( .A1(n_752), .A2(n_113), .A3(n_114), .B(n_116), .Y(n_869) );
AO31x2_ASAP7_75t_L g870 ( .A1(n_752), .A2(n_113), .A3(n_117), .B(n_119), .Y(n_870) );
O2A1O1Ixp33_ASAP7_75t_L g871 ( .A1(n_662), .A2(n_119), .B(n_120), .C(n_121), .Y(n_871) );
INVx1_ASAP7_75t_L g872 ( .A(n_703), .Y(n_872) );
NOR2xp33_ASAP7_75t_L g873 ( .A(n_830), .B(n_122), .Y(n_873) );
BUFx6f_ASAP7_75t_L g874 ( .A(n_868), .Y(n_874) );
OAI21xp5_ASAP7_75t_L g875 ( .A1(n_806), .A2(n_795), .B(n_821), .Y(n_875) );
NAND2xp5_ASAP7_75t_L g876 ( .A(n_778), .B(n_123), .Y(n_876) );
INVx2_ASAP7_75t_L g877 ( .A(n_777), .Y(n_877) );
AO31x2_ASAP7_75t_L g878 ( .A1(n_788), .A2(n_124), .A3(n_125), .B(n_126), .Y(n_878) );
AND2x4_ASAP7_75t_L g879 ( .A(n_761), .B(n_126), .Y(n_879) );
OAI21xp5_ASAP7_75t_L g880 ( .A1(n_766), .A2(n_127), .B(n_129), .Y(n_880) );
INVx2_ASAP7_75t_L g881 ( .A(n_779), .Y(n_881) );
CKINVDCx5p33_ASAP7_75t_R g882 ( .A(n_791), .Y(n_882) );
HB1xp67_ASAP7_75t_L g883 ( .A(n_797), .Y(n_883) );
BUFx8_ASAP7_75t_L g884 ( .A(n_866), .Y(n_884) );
INVx1_ASAP7_75t_L g885 ( .A(n_872), .Y(n_885) );
AOI221xp5_ASAP7_75t_L g886 ( .A1(n_773), .A2(n_130), .B1(n_132), .B2(n_201), .C(n_202), .Y(n_886) );
AOI22xp33_ASAP7_75t_L g887 ( .A1(n_768), .A2(n_203), .B1(n_207), .B2(n_209), .Y(n_887) );
INVx4_ASAP7_75t_L g888 ( .A(n_801), .Y(n_888) );
NAND2xp5_ASAP7_75t_L g889 ( .A(n_807), .B(n_305), .Y(n_889) );
INVx1_ASAP7_75t_L g890 ( .A(n_759), .Y(n_890) );
NAND2xp5_ASAP7_75t_L g891 ( .A(n_768), .B(n_215), .Y(n_891) );
INVx1_ASAP7_75t_L g892 ( .A(n_759), .Y(n_892) );
AOI21xp5_ASAP7_75t_SL g893 ( .A1(n_859), .A2(n_220), .B(n_221), .Y(n_893) );
NAND2x1p5_ASAP7_75t_L g894 ( .A(n_801), .B(n_222), .Y(n_894) );
HB1xp67_ASAP7_75t_L g895 ( .A(n_828), .Y(n_895) );
INVx1_ASAP7_75t_L g896 ( .A(n_813), .Y(n_896) );
AOI211xp5_ASAP7_75t_L g897 ( .A1(n_804), .A2(n_812), .B(n_794), .C(n_771), .Y(n_897) );
INVx5_ASAP7_75t_L g898 ( .A(n_868), .Y(n_898) );
HB1xp67_ASAP7_75t_L g899 ( .A(n_801), .Y(n_899) );
INVx3_ASAP7_75t_L g900 ( .A(n_868), .Y(n_900) );
AND2x2_ASAP7_75t_L g901 ( .A(n_841), .B(n_229), .Y(n_901) );
AO21x2_ASAP7_75t_L g902 ( .A1(n_787), .A2(n_231), .B(n_232), .Y(n_902) );
BUFx6f_ASAP7_75t_SL g903 ( .A(n_832), .Y(n_903) );
OAI22xp33_ASAP7_75t_L g904 ( .A1(n_860), .A2(n_235), .B1(n_239), .B2(n_240), .Y(n_904) );
OAI21xp5_ASAP7_75t_L g905 ( .A1(n_800), .A2(n_242), .B(n_244), .Y(n_905) );
OR2x2_ASAP7_75t_L g906 ( .A(n_786), .B(n_245), .Y(n_906) );
AND2x2_ASAP7_75t_L g907 ( .A(n_793), .B(n_246), .Y(n_907) );
BUFx8_ASAP7_75t_L g908 ( .A(n_809), .Y(n_908) );
O2A1O1Ixp33_ASAP7_75t_L g909 ( .A1(n_864), .A2(n_247), .B(n_248), .C(n_249), .Y(n_909) );
AND2x4_ASAP7_75t_L g910 ( .A(n_849), .B(n_250), .Y(n_910) );
OAI211xp5_ASAP7_75t_L g911 ( .A1(n_758), .A2(n_253), .B(n_254), .C(n_257), .Y(n_911) );
NOR2xp67_ASAP7_75t_L g912 ( .A(n_853), .B(n_849), .Y(n_912) );
AND2x2_ASAP7_75t_L g913 ( .A(n_843), .B(n_259), .Y(n_913) );
AND2x4_ASAP7_75t_L g914 ( .A(n_852), .B(n_262), .Y(n_914) );
INVx2_ASAP7_75t_L g915 ( .A(n_835), .Y(n_915) );
INVx2_ASAP7_75t_L g916 ( .A(n_836), .Y(n_916) );
O2A1O1Ixp33_ASAP7_75t_L g917 ( .A1(n_865), .A2(n_267), .B(n_269), .C(n_272), .Y(n_917) );
INVx4_ASAP7_75t_SL g918 ( .A(n_772), .Y(n_918) );
AOI22xp33_ASAP7_75t_L g919 ( .A1(n_782), .A2(n_276), .B1(n_277), .B2(n_278), .Y(n_919) );
INVx1_ASAP7_75t_L g920 ( .A(n_838), .Y(n_920) );
AND2x2_ASAP7_75t_L g921 ( .A(n_808), .B(n_279), .Y(n_921) );
INVx2_ASAP7_75t_L g922 ( .A(n_756), .Y(n_922) );
INVx1_ASAP7_75t_L g923 ( .A(n_842), .Y(n_923) );
CKINVDCx20_ASAP7_75t_R g924 ( .A(n_799), .Y(n_924) );
NAND2xp5_ASAP7_75t_L g925 ( .A(n_817), .B(n_280), .Y(n_925) );
AOI21xp5_ASAP7_75t_L g926 ( .A1(n_798), .A2(n_282), .B(n_283), .Y(n_926) );
AO21x2_ASAP7_75t_L g927 ( .A1(n_760), .A2(n_287), .B(n_288), .Y(n_927) );
AO22x1_ASAP7_75t_L g928 ( .A1(n_854), .A2(n_289), .B1(n_290), .B2(n_291), .Y(n_928) );
OA21x2_ASAP7_75t_L g929 ( .A1(n_796), .A2(n_767), .B(n_781), .Y(n_929) );
NAND2xp5_ASAP7_75t_L g930 ( .A(n_820), .B(n_826), .Y(n_930) );
OAI21xp5_ASAP7_75t_L g931 ( .A1(n_805), .A2(n_818), .B(n_850), .Y(n_931) );
NAND2xp5_ASAP7_75t_L g932 ( .A(n_820), .B(n_826), .Y(n_932) );
AND2x2_ASAP7_75t_L g933 ( .A(n_831), .B(n_863), .Y(n_933) );
INVx1_ASAP7_75t_L g934 ( .A(n_803), .Y(n_934) );
OA21x2_ASAP7_75t_L g935 ( .A1(n_861), .A2(n_762), .B(n_776), .Y(n_935) );
INVx1_ASAP7_75t_L g936 ( .A(n_803), .Y(n_936) );
NAND2xp5_ASAP7_75t_L g937 ( .A(n_855), .B(n_844), .Y(n_937) );
INVx1_ASAP7_75t_L g938 ( .A(n_803), .Y(n_938) );
AND2x2_ASAP7_75t_SL g939 ( .A(n_816), .B(n_855), .Y(n_939) );
BUFx6f_ASAP7_75t_L g940 ( .A(n_837), .Y(n_940) );
AOI22xp5_ASAP7_75t_L g941 ( .A1(n_815), .A2(n_851), .B1(n_822), .B2(n_775), .Y(n_941) );
OAI22xp5_ASAP7_75t_L g942 ( .A1(n_845), .A2(n_834), .B1(n_839), .B2(n_867), .Y(n_942) );
A2O1A1Ixp33_ASAP7_75t_L g943 ( .A1(n_871), .A2(n_784), .B(n_848), .C(n_862), .Y(n_943) );
INVx1_ASAP7_75t_L g944 ( .A(n_856), .Y(n_944) );
AOI222xp33_ASAP7_75t_L g945 ( .A1(n_783), .A2(n_827), .B1(n_811), .B2(n_810), .C1(n_825), .C2(n_833), .Y(n_945) );
A2O1A1Ixp33_ASAP7_75t_L g946 ( .A1(n_755), .A2(n_858), .B(n_823), .C(n_802), .Y(n_946) );
AOI21xp5_ASAP7_75t_L g947 ( .A1(n_774), .A2(n_857), .B(n_792), .Y(n_947) );
NAND2x1p5_ASAP7_75t_L g948 ( .A(n_790), .B(n_846), .Y(n_948) );
OA21x2_ASAP7_75t_L g949 ( .A1(n_770), .A2(n_754), .B(n_840), .Y(n_949) );
BUFx8_ASAP7_75t_L g950 ( .A(n_785), .Y(n_950) );
INVx1_ASAP7_75t_L g951 ( .A(n_814), .Y(n_951) );
AOI21xp5_ASAP7_75t_L g952 ( .A1(n_780), .A2(n_847), .B(n_819), .Y(n_952) );
INVx1_ASAP7_75t_L g953 ( .A(n_814), .Y(n_953) );
INVx2_ASAP7_75t_L g954 ( .A(n_870), .Y(n_954) );
AOI21xp33_ASAP7_75t_SL g955 ( .A1(n_789), .A2(n_829), .B(n_869), .Y(n_955) );
AOI21xp5_ASAP7_75t_L g956 ( .A1(n_763), .A2(n_769), .B(n_757), .Y(n_956) );
INVx1_ASAP7_75t_L g957 ( .A(n_869), .Y(n_957) );
OAI21x1_ASAP7_75t_L g958 ( .A1(n_769), .A2(n_757), .B(n_869), .Y(n_958) );
INVx2_ASAP7_75t_L g959 ( .A(n_870), .Y(n_959) );
INVx1_ASAP7_75t_SL g960 ( .A(n_870), .Y(n_960) );
NAND2xp5_ASAP7_75t_L g961 ( .A(n_789), .B(n_829), .Y(n_961) );
INVx1_ASAP7_75t_L g962 ( .A(n_829), .Y(n_962) );
OAI211xp5_ASAP7_75t_L g963 ( .A1(n_793), .A2(n_584), .B(n_758), .C(n_678), .Y(n_963) );
BUFx3_ASAP7_75t_L g964 ( .A(n_791), .Y(n_964) );
OA21x2_ASAP7_75t_L g965 ( .A1(n_766), .A2(n_735), .B(n_752), .Y(n_965) );
OA21x2_ASAP7_75t_L g966 ( .A1(n_766), .A2(n_735), .B(n_752), .Y(n_966) );
INVx1_ASAP7_75t_L g967 ( .A(n_778), .Y(n_967) );
OR2x2_ASAP7_75t_L g968 ( .A(n_828), .B(n_734), .Y(n_968) );
HB1xp67_ASAP7_75t_L g969 ( .A(n_791), .Y(n_969) );
OAI21x1_ASAP7_75t_L g970 ( .A1(n_764), .A2(n_735), .B(n_765), .Y(n_970) );
AOI22xp33_ASAP7_75t_SL g971 ( .A1(n_768), .A2(n_644), .B1(n_678), .B2(n_632), .Y(n_971) );
AO31x2_ASAP7_75t_L g972 ( .A1(n_788), .A2(n_752), .A3(n_646), .B(n_639), .Y(n_972) );
AOI22xp33_ASAP7_75t_L g973 ( .A1(n_768), .A2(n_583), .B1(n_679), .B2(n_643), .Y(n_973) );
INVx1_ASAP7_75t_L g974 ( .A(n_778), .Y(n_974) );
OA21x2_ASAP7_75t_L g975 ( .A1(n_766), .A2(n_735), .B(n_752), .Y(n_975) );
NAND2xp5_ASAP7_75t_L g976 ( .A(n_778), .B(n_703), .Y(n_976) );
INVx1_ASAP7_75t_L g977 ( .A(n_778), .Y(n_977) );
INVx2_ASAP7_75t_L g978 ( .A(n_778), .Y(n_978) );
A2O1A1Ixp33_ASAP7_75t_L g979 ( .A1(n_821), .A2(n_795), .B(n_806), .C(n_753), .Y(n_979) );
AOI21xp5_ASAP7_75t_L g980 ( .A1(n_764), .A2(n_752), .B(n_646), .Y(n_980) );
INVx2_ASAP7_75t_L g981 ( .A(n_778), .Y(n_981) );
OAI221xp5_ASAP7_75t_L g982 ( .A1(n_824), .A2(n_584), .B1(n_583), .B2(n_585), .C(n_637), .Y(n_982) );
INVx2_ASAP7_75t_L g983 ( .A(n_778), .Y(n_983) );
INVx3_ASAP7_75t_L g984 ( .A(n_801), .Y(n_984) );
NAND2xp5_ASAP7_75t_L g985 ( .A(n_778), .B(n_702), .Y(n_985) );
NAND2xp5_ASAP7_75t_L g986 ( .A(n_778), .B(n_703), .Y(n_986) );
NAND2xp5_ASAP7_75t_L g987 ( .A(n_778), .B(n_703), .Y(n_987) );
INVx3_ASAP7_75t_L g988 ( .A(n_801), .Y(n_988) );
AO21x2_ASAP7_75t_L g989 ( .A1(n_766), .A2(n_752), .B(n_764), .Y(n_989) );
CKINVDCx5p33_ASAP7_75t_R g990 ( .A(n_791), .Y(n_990) );
INVx3_ASAP7_75t_L g991 ( .A(n_801), .Y(n_991) );
NAND2xp5_ASAP7_75t_L g992 ( .A(n_778), .B(n_703), .Y(n_992) );
NAND2x1p5_ASAP7_75t_L g993 ( .A(n_791), .B(n_801), .Y(n_993) );
AOI22xp33_ASAP7_75t_SL g994 ( .A1(n_768), .A2(n_644), .B1(n_678), .B2(n_632), .Y(n_994) );
AOI21xp5_ASAP7_75t_L g995 ( .A1(n_764), .A2(n_752), .B(n_646), .Y(n_995) );
INVx1_ASAP7_75t_L g996 ( .A(n_778), .Y(n_996) );
AOI21xp5_ASAP7_75t_L g997 ( .A1(n_764), .A2(n_752), .B(n_646), .Y(n_997) );
OA21x2_ASAP7_75t_L g998 ( .A1(n_875), .A2(n_952), .B(n_961), .Y(n_998) );
OA21x2_ASAP7_75t_L g999 ( .A1(n_875), .A2(n_956), .B(n_979), .Y(n_999) );
AND2x2_ASAP7_75t_L g1000 ( .A(n_877), .B(n_881), .Y(n_1000) );
OA21x2_ASAP7_75t_L g1001 ( .A1(n_951), .A2(n_953), .B(n_957), .Y(n_1001) );
AND2x4_ASAP7_75t_L g1002 ( .A(n_898), .B(n_914), .Y(n_1002) );
INVx2_ASAP7_75t_L g1003 ( .A(n_970), .Y(n_1003) );
INVx1_ASAP7_75t_L g1004 ( .A(n_885), .Y(n_1004) );
HB1xp67_ASAP7_75t_L g1005 ( .A(n_895), .Y(n_1005) );
INVx4_ASAP7_75t_L g1006 ( .A(n_888), .Y(n_1006) );
BUFx3_ASAP7_75t_L g1007 ( .A(n_993), .Y(n_1007) );
AND2x2_ASAP7_75t_L g1008 ( .A(n_915), .B(n_916), .Y(n_1008) );
AND2x2_ASAP7_75t_L g1009 ( .A(n_896), .B(n_978), .Y(n_1009) );
INVx1_ASAP7_75t_L g1010 ( .A(n_962), .Y(n_1010) );
INVx1_ASAP7_75t_L g1011 ( .A(n_934), .Y(n_1011) );
OR2x2_ASAP7_75t_L g1012 ( .A(n_976), .B(n_986), .Y(n_1012) );
AND2x2_ASAP7_75t_L g1013 ( .A(n_981), .B(n_983), .Y(n_1013) );
HB1xp67_ASAP7_75t_L g1014 ( .A(n_987), .Y(n_1014) );
NAND2xp5_ASAP7_75t_L g1015 ( .A(n_985), .B(n_992), .Y(n_1015) );
INVx1_ASAP7_75t_L g1016 ( .A(n_936), .Y(n_1016) );
INVx5_ASAP7_75t_L g1017 ( .A(n_874), .Y(n_1017) );
OAI21xp5_ASAP7_75t_L g1018 ( .A1(n_943), .A2(n_946), .B(n_941), .Y(n_1018) );
OR2x2_ASAP7_75t_L g1019 ( .A(n_938), .B(n_930), .Y(n_1019) );
AO21x2_ASAP7_75t_L g1020 ( .A1(n_955), .A2(n_931), .B(n_954), .Y(n_1020) );
BUFx2_ASAP7_75t_SL g1021 ( .A(n_912), .Y(n_1021) );
INVx1_ASAP7_75t_L g1022 ( .A(n_959), .Y(n_1022) );
OR2x6_ASAP7_75t_L g1023 ( .A(n_914), .B(n_932), .Y(n_1023) );
AOI22xp33_ASAP7_75t_L g1024 ( .A1(n_982), .A2(n_945), .B1(n_994), .B2(n_971), .Y(n_1024) );
INVx1_ASAP7_75t_L g1025 ( .A(n_967), .Y(n_1025) );
INVx1_ASAP7_75t_L g1026 ( .A(n_974), .Y(n_1026) );
INVx1_ASAP7_75t_L g1027 ( .A(n_977), .Y(n_1027) );
OA21x2_ASAP7_75t_L g1028 ( .A1(n_931), .A2(n_960), .B(n_997), .Y(n_1028) );
INVx1_ASAP7_75t_L g1029 ( .A(n_996), .Y(n_1029) );
INVx4_ASAP7_75t_L g1030 ( .A(n_888), .Y(n_1030) );
AO21x2_ASAP7_75t_L g1031 ( .A1(n_955), .A2(n_995), .B(n_980), .Y(n_1031) );
INVxp67_ASAP7_75t_L g1032 ( .A(n_968), .Y(n_1032) );
NAND2xp5_ASAP7_75t_L g1033 ( .A(n_985), .B(n_973), .Y(n_1033) );
AOI21x1_ASAP7_75t_L g1034 ( .A1(n_947), .A2(n_929), .B(n_935), .Y(n_1034) );
INVx2_ASAP7_75t_L g1035 ( .A(n_922), .Y(n_1035) );
INVx2_ASAP7_75t_SL g1036 ( .A(n_908), .Y(n_1036) );
INVx1_ASAP7_75t_L g1037 ( .A(n_944), .Y(n_1037) );
BUFx3_ASAP7_75t_L g1038 ( .A(n_884), .Y(n_1038) );
AND2x2_ASAP7_75t_L g1039 ( .A(n_920), .B(n_923), .Y(n_1039) );
INVx2_ASAP7_75t_SL g1040 ( .A(n_908), .Y(n_1040) );
OR2x6_ASAP7_75t_L g1041 ( .A(n_894), .B(n_910), .Y(n_1041) );
NOR2xp33_ASAP7_75t_L g1042 ( .A(n_883), .B(n_933), .Y(n_1042) );
OAI22xp5_ASAP7_75t_L g1043 ( .A1(n_941), .A2(n_963), .B1(n_897), .B2(n_891), .Y(n_1043) );
AO21x2_ASAP7_75t_L g1044 ( .A1(n_880), .A2(n_927), .B(n_989), .Y(n_1044) );
INVx1_ASAP7_75t_L g1045 ( .A(n_876), .Y(n_1045) );
AND2x2_ASAP7_75t_L g1046 ( .A(n_873), .B(n_890), .Y(n_1046) );
HB1xp67_ASAP7_75t_L g1047 ( .A(n_899), .Y(n_1047) );
NAND2xp5_ASAP7_75t_L g1048 ( .A(n_897), .B(n_945), .Y(n_1048) );
HB1xp67_ASAP7_75t_L g1049 ( .A(n_984), .Y(n_1049) );
INVx1_ASAP7_75t_L g1050 ( .A(n_878), .Y(n_1050) );
BUFx3_ASAP7_75t_L g1051 ( .A(n_884), .Y(n_1051) );
INVx1_ASAP7_75t_SL g1052 ( .A(n_964), .Y(n_1052) );
AND2x2_ASAP7_75t_L g1053 ( .A(n_892), .B(n_879), .Y(n_1053) );
OR2x6_ASAP7_75t_L g1054 ( .A(n_910), .B(n_948), .Y(n_1054) );
AO21x2_ASAP7_75t_L g1055 ( .A1(n_942), .A2(n_902), .B(n_905), .Y(n_1055) );
OAI33xp33_ASAP7_75t_L g1056 ( .A1(n_942), .A2(n_906), .A3(n_904), .B1(n_937), .B2(n_889), .B3(n_925), .Y(n_1056) );
OAI21x1_ASAP7_75t_L g1057 ( .A1(n_965), .A2(n_975), .B(n_966), .Y(n_1057) );
OR2x2_ASAP7_75t_L g1058 ( .A(n_984), .B(n_988), .Y(n_1058) );
OAI22xp5_ASAP7_75t_L g1059 ( .A1(n_887), .A2(n_879), .B1(n_939), .B2(n_901), .Y(n_1059) );
BUFx3_ASAP7_75t_L g1060 ( .A(n_898), .Y(n_1060) );
INVx2_ASAP7_75t_L g1061 ( .A(n_972), .Y(n_1061) );
HB1xp67_ASAP7_75t_L g1062 ( .A(n_988), .Y(n_1062) );
HB1xp67_ASAP7_75t_L g1063 ( .A(n_991), .Y(n_1063) );
HB1xp67_ASAP7_75t_L g1064 ( .A(n_991), .Y(n_1064) );
INVx2_ASAP7_75t_L g1065 ( .A(n_972), .Y(n_1065) );
NOR2xp33_ASAP7_75t_L g1066 ( .A(n_969), .B(n_882), .Y(n_1066) );
INVx2_ASAP7_75t_L g1067 ( .A(n_972), .Y(n_1067) );
AND2x2_ASAP7_75t_L g1068 ( .A(n_900), .B(n_898), .Y(n_1068) );
BUFx2_ASAP7_75t_L g1069 ( .A(n_900), .Y(n_1069) );
AND2x2_ASAP7_75t_L g1070 ( .A(n_921), .B(n_913), .Y(n_1070) );
INVx1_ASAP7_75t_L g1071 ( .A(n_940), .Y(n_1071) );
HB1xp67_ASAP7_75t_L g1072 ( .A(n_903), .Y(n_1072) );
INVx1_ASAP7_75t_L g1073 ( .A(n_903), .Y(n_1073) );
BUFx2_ASAP7_75t_L g1074 ( .A(n_940), .Y(n_1074) );
OAI33xp33_ASAP7_75t_L g1075 ( .A1(n_990), .A2(n_917), .A3(n_909), .B1(n_950), .B2(n_918), .B3(n_886), .Y(n_1075) );
OAI21xp5_ASAP7_75t_L g1076 ( .A1(n_907), .A2(n_911), .B(n_926), .Y(n_1076) );
OR2x2_ASAP7_75t_L g1077 ( .A(n_949), .B(n_928), .Y(n_1077) );
INVxp33_ASAP7_75t_L g1078 ( .A(n_918), .Y(n_1078) );
INVx1_ASAP7_75t_L g1079 ( .A(n_893), .Y(n_1079) );
INVx3_ASAP7_75t_L g1080 ( .A(n_950), .Y(n_1080) );
OA21x2_ASAP7_75t_L g1081 ( .A1(n_919), .A2(n_875), .B(n_958), .Y(n_1081) );
INVx2_ASAP7_75t_L g1082 ( .A(n_924), .Y(n_1082) );
AOI211xp5_ASAP7_75t_L g1083 ( .A1(n_982), .A2(n_963), .B(n_685), .C(n_804), .Y(n_1083) );
BUFx4f_ASAP7_75t_SL g1084 ( .A(n_884), .Y(n_1084) );
AND2x2_ASAP7_75t_L g1085 ( .A(n_877), .B(n_768), .Y(n_1085) );
NAND2xp5_ASAP7_75t_L g1086 ( .A(n_985), .B(n_778), .Y(n_1086) );
HB1xp67_ASAP7_75t_L g1087 ( .A(n_895), .Y(n_1087) );
AND2x4_ASAP7_75t_L g1088 ( .A(n_898), .B(n_914), .Y(n_1088) );
OA21x2_ASAP7_75t_L g1089 ( .A1(n_875), .A2(n_958), .B(n_952), .Y(n_1089) );
INVx1_ASAP7_75t_L g1090 ( .A(n_885), .Y(n_1090) );
OR2x6_ASAP7_75t_L g1091 ( .A(n_914), .B(n_930), .Y(n_1091) );
AND2x2_ASAP7_75t_L g1092 ( .A(n_877), .B(n_768), .Y(n_1092) );
AND2x2_ASAP7_75t_L g1093 ( .A(n_877), .B(n_768), .Y(n_1093) );
AND2x2_ASAP7_75t_L g1094 ( .A(n_877), .B(n_768), .Y(n_1094) );
AO21x2_ASAP7_75t_L g1095 ( .A1(n_955), .A2(n_875), .B(n_952), .Y(n_1095) );
AND2x2_ASAP7_75t_L g1096 ( .A(n_877), .B(n_768), .Y(n_1096) );
AND2x2_ASAP7_75t_L g1097 ( .A(n_877), .B(n_768), .Y(n_1097) );
AND2x2_ASAP7_75t_L g1098 ( .A(n_877), .B(n_768), .Y(n_1098) );
INVx1_ASAP7_75t_L g1099 ( .A(n_962), .Y(n_1099) );
OA21x2_ASAP7_75t_L g1100 ( .A1(n_875), .A2(n_958), .B(n_952), .Y(n_1100) );
INVx1_ASAP7_75t_L g1101 ( .A(n_962), .Y(n_1101) );
OR2x2_ASAP7_75t_L g1102 ( .A(n_1019), .B(n_1033), .Y(n_1102) );
AND2x4_ASAP7_75t_SL g1103 ( .A(n_1041), .B(n_1002), .Y(n_1103) );
AND2x2_ASAP7_75t_L g1104 ( .A(n_1013), .B(n_1010), .Y(n_1104) );
AND2x2_ASAP7_75t_L g1105 ( .A(n_1013), .B(n_1010), .Y(n_1105) );
INVx1_ASAP7_75t_L g1106 ( .A(n_1099), .Y(n_1106) );
BUFx6f_ASAP7_75t_L g1107 ( .A(n_1017), .Y(n_1107) );
HB1xp67_ASAP7_75t_L g1108 ( .A(n_1014), .Y(n_1108) );
HB1xp67_ASAP7_75t_L g1109 ( .A(n_1005), .Y(n_1109) );
INVxp67_ASAP7_75t_SL g1110 ( .A(n_1002), .Y(n_1110) );
AND2x2_ASAP7_75t_L g1111 ( .A(n_1101), .B(n_1011), .Y(n_1111) );
AND2x4_ASAP7_75t_SL g1112 ( .A(n_1041), .B(n_1002), .Y(n_1112) );
AND2x2_ASAP7_75t_L g1113 ( .A(n_1011), .B(n_1016), .Y(n_1113) );
OR2x2_ASAP7_75t_L g1114 ( .A(n_1019), .B(n_1012), .Y(n_1114) );
NAND2x1p5_ASAP7_75t_L g1115 ( .A(n_1088), .B(n_1017), .Y(n_1115) );
INVx1_ASAP7_75t_L g1116 ( .A(n_1016), .Y(n_1116) );
INVx3_ASAP7_75t_SL g1117 ( .A(n_1038), .Y(n_1117) );
AOI22xp33_ASAP7_75t_L g1118 ( .A1(n_1048), .A2(n_1024), .B1(n_1043), .B2(n_1018), .Y(n_1118) );
AOI222xp33_ASAP7_75t_L g1119 ( .A1(n_1084), .A2(n_1046), .B1(n_1042), .B2(n_1051), .C1(n_1038), .C2(n_1045), .Y(n_1119) );
AND2x2_ASAP7_75t_L g1120 ( .A(n_1039), .B(n_1025), .Y(n_1120) );
AND2x2_ASAP7_75t_L g1121 ( .A(n_1039), .B(n_1025), .Y(n_1121) );
AND2x2_ASAP7_75t_L g1122 ( .A(n_1027), .B(n_1029), .Y(n_1122) );
OAI21xp33_ASAP7_75t_L g1123 ( .A1(n_1083), .A2(n_1015), .B(n_1054), .Y(n_1123) );
INVx1_ASAP7_75t_L g1124 ( .A(n_1001), .Y(n_1124) );
INVxp67_ASAP7_75t_SL g1125 ( .A(n_1088), .Y(n_1125) );
AND2x2_ASAP7_75t_L g1126 ( .A(n_1027), .B(n_1029), .Y(n_1126) );
NOR2xp33_ASAP7_75t_L g1127 ( .A(n_1082), .B(n_1052), .Y(n_1127) );
AND2x2_ASAP7_75t_L g1128 ( .A(n_1037), .B(n_1035), .Y(n_1128) );
AOI22xp33_ASAP7_75t_L g1129 ( .A1(n_1054), .A2(n_1059), .B1(n_1056), .B2(n_1023), .Y(n_1129) );
INVx1_ASAP7_75t_SL g1130 ( .A(n_1058), .Y(n_1130) );
INVx1_ASAP7_75t_L g1131 ( .A(n_1001), .Y(n_1131) );
NAND2xp5_ASAP7_75t_L g1132 ( .A(n_1009), .B(n_1086), .Y(n_1132) );
INVx2_ASAP7_75t_L g1133 ( .A(n_1022), .Y(n_1133) );
BUFx3_ASAP7_75t_L g1134 ( .A(n_1088), .Y(n_1134) );
NAND2xp5_ASAP7_75t_L g1135 ( .A(n_1004), .B(n_1090), .Y(n_1135) );
INVx1_ASAP7_75t_L g1136 ( .A(n_1001), .Y(n_1136) );
AND2x2_ASAP7_75t_L g1137 ( .A(n_999), .B(n_1000), .Y(n_1137) );
INVxp67_ASAP7_75t_SL g1138 ( .A(n_1087), .Y(n_1138) );
AND2x2_ASAP7_75t_L g1139 ( .A(n_999), .B(n_1000), .Y(n_1139) );
AND2x2_ASAP7_75t_L g1140 ( .A(n_999), .B(n_1008), .Y(n_1140) );
NAND2xp5_ASAP7_75t_L g1141 ( .A(n_1032), .B(n_1026), .Y(n_1141) );
INVxp67_ASAP7_75t_SL g1142 ( .A(n_1047), .Y(n_1142) );
AND2x2_ASAP7_75t_L g1143 ( .A(n_1050), .B(n_1061), .Y(n_1143) );
NAND2xp5_ASAP7_75t_L g1144 ( .A(n_1085), .B(n_1092), .Y(n_1144) );
AND2x2_ASAP7_75t_L g1145 ( .A(n_1050), .B(n_1065), .Y(n_1145) );
INVx2_ASAP7_75t_SL g1146 ( .A(n_1017), .Y(n_1146) );
NAND2xp5_ASAP7_75t_L g1147 ( .A(n_1085), .B(n_1092), .Y(n_1147) );
AND2x2_ASAP7_75t_L g1148 ( .A(n_1067), .B(n_1093), .Y(n_1148) );
INVx1_ASAP7_75t_L g1149 ( .A(n_1031), .Y(n_1149) );
AOI22xp33_ASAP7_75t_L g1150 ( .A1(n_1054), .A2(n_1023), .B1(n_1091), .B2(n_1097), .Y(n_1150) );
OR2x2_ASAP7_75t_L g1151 ( .A(n_1049), .B(n_1062), .Y(n_1151) );
HB1xp67_ASAP7_75t_L g1152 ( .A(n_1063), .Y(n_1152) );
AND2x2_ASAP7_75t_L g1153 ( .A(n_1093), .B(n_1094), .Y(n_1153) );
NAND2xp5_ASAP7_75t_L g1154 ( .A(n_1094), .B(n_1096), .Y(n_1154) );
AND2x2_ASAP7_75t_L g1155 ( .A(n_1096), .B(n_1097), .Y(n_1155) );
AND2x2_ASAP7_75t_L g1156 ( .A(n_1098), .B(n_998), .Y(n_1156) );
OR2x2_ASAP7_75t_L g1157 ( .A(n_1064), .B(n_1058), .Y(n_1157) );
NAND2xp5_ASAP7_75t_L g1158 ( .A(n_1098), .B(n_1053), .Y(n_1158) );
INVx4_ASAP7_75t_L g1159 ( .A(n_1041), .Y(n_1159) );
BUFx3_ASAP7_75t_L g1160 ( .A(n_1017), .Y(n_1160) );
INVxp67_ASAP7_75t_SL g1161 ( .A(n_1069), .Y(n_1161) );
AND2x2_ASAP7_75t_L g1162 ( .A(n_998), .B(n_1020), .Y(n_1162) );
NOR2xp33_ASAP7_75t_L g1163 ( .A(n_1082), .B(n_1066), .Y(n_1163) );
AND2x2_ASAP7_75t_L g1164 ( .A(n_998), .B(n_1020), .Y(n_1164) );
OAI22xp5_ASAP7_75t_L g1165 ( .A1(n_1041), .A2(n_1091), .B1(n_1023), .B2(n_1070), .Y(n_1165) );
AND2x2_ASAP7_75t_L g1166 ( .A(n_1095), .B(n_1028), .Y(n_1166) );
AND2x2_ASAP7_75t_L g1167 ( .A(n_1095), .B(n_1071), .Y(n_1167) );
NAND2xp5_ASAP7_75t_L g1168 ( .A(n_1053), .B(n_1070), .Y(n_1168) );
OR2x6_ASAP7_75t_L g1169 ( .A(n_1077), .B(n_1091), .Y(n_1169) );
OR2x2_ASAP7_75t_L g1170 ( .A(n_1114), .B(n_1100), .Y(n_1170) );
INVx1_ASAP7_75t_L g1171 ( .A(n_1122), .Y(n_1171) );
OR2x2_ASAP7_75t_L g1172 ( .A(n_1114), .B(n_1100), .Y(n_1172) );
INVx1_ASAP7_75t_L g1173 ( .A(n_1122), .Y(n_1173) );
AND2x2_ASAP7_75t_L g1174 ( .A(n_1137), .B(n_1100), .Y(n_1174) );
AND2x2_ASAP7_75t_L g1175 ( .A(n_1137), .B(n_1089), .Y(n_1175) );
INVx1_ASAP7_75t_L g1176 ( .A(n_1126), .Y(n_1176) );
OR2x2_ASAP7_75t_L g1177 ( .A(n_1102), .B(n_1089), .Y(n_1177) );
NAND2x1p5_ASAP7_75t_L g1178 ( .A(n_1159), .B(n_1030), .Y(n_1178) );
INVx1_ASAP7_75t_SL g1179 ( .A(n_1117), .Y(n_1179) );
AOI22xp33_ASAP7_75t_L g1180 ( .A1(n_1123), .A2(n_1075), .B1(n_1091), .B2(n_1023), .Y(n_1180) );
OR2x2_ASAP7_75t_L g1181 ( .A(n_1102), .B(n_1089), .Y(n_1181) );
NAND2xp5_ASAP7_75t_L g1182 ( .A(n_1120), .B(n_1073), .Y(n_1182) );
NAND2xp5_ASAP7_75t_L g1183 ( .A(n_1120), .B(n_1030), .Y(n_1183) );
INVx1_ASAP7_75t_SL g1184 ( .A(n_1117), .Y(n_1184) );
AND2x2_ASAP7_75t_L g1185 ( .A(n_1139), .B(n_1140), .Y(n_1185) );
NAND2xp5_ASAP7_75t_L g1186 ( .A(n_1121), .B(n_1030), .Y(n_1186) );
AND2x4_ASAP7_75t_L g1187 ( .A(n_1156), .B(n_1003), .Y(n_1187) );
NAND2x1p5_ASAP7_75t_L g1188 ( .A(n_1159), .B(n_1006), .Y(n_1188) );
AND2x2_ASAP7_75t_L g1189 ( .A(n_1139), .B(n_1081), .Y(n_1189) );
NAND2xp5_ASAP7_75t_L g1190 ( .A(n_1121), .B(n_1104), .Y(n_1190) );
INVx1_ASAP7_75t_L g1191 ( .A(n_1106), .Y(n_1191) );
NAND2xp5_ASAP7_75t_L g1192 ( .A(n_1104), .B(n_1069), .Y(n_1192) );
INVx1_ASAP7_75t_L g1193 ( .A(n_1106), .Y(n_1193) );
HB1xp67_ASAP7_75t_L g1194 ( .A(n_1108), .Y(n_1194) );
AND2x2_ASAP7_75t_L g1195 ( .A(n_1156), .B(n_1057), .Y(n_1195) );
AND2x2_ASAP7_75t_L g1196 ( .A(n_1148), .B(n_1057), .Y(n_1196) );
BUFx2_ASAP7_75t_L g1197 ( .A(n_1161), .Y(n_1197) );
INVx1_ASAP7_75t_L g1198 ( .A(n_1126), .Y(n_1198) );
NAND2xp5_ASAP7_75t_L g1199 ( .A(n_1105), .B(n_1072), .Y(n_1199) );
CKINVDCx16_ASAP7_75t_R g1200 ( .A(n_1160), .Y(n_1200) );
INVx1_ASAP7_75t_L g1201 ( .A(n_1116), .Y(n_1201) );
NAND2xp33_ASAP7_75t_SL g1202 ( .A(n_1159), .B(n_1078), .Y(n_1202) );
AND2x2_ASAP7_75t_L g1203 ( .A(n_1111), .B(n_1055), .Y(n_1203) );
NAND2x1p5_ASAP7_75t_L g1204 ( .A(n_1159), .B(n_1017), .Y(n_1204) );
AND2x2_ASAP7_75t_L g1205 ( .A(n_1113), .B(n_1055), .Y(n_1205) );
AND2x2_ASAP7_75t_L g1206 ( .A(n_1113), .B(n_1055), .Y(n_1206) );
AND2x2_ASAP7_75t_SL g1207 ( .A(n_1103), .B(n_1077), .Y(n_1207) );
NOR2xp33_ASAP7_75t_L g1208 ( .A(n_1163), .B(n_1036), .Y(n_1208) );
NAND2xp5_ASAP7_75t_L g1209 ( .A(n_1105), .B(n_1021), .Y(n_1209) );
NAND2xp5_ASAP7_75t_L g1210 ( .A(n_1132), .B(n_1074), .Y(n_1210) );
AND2x4_ASAP7_75t_SL g1211 ( .A(n_1107), .B(n_1040), .Y(n_1211) );
NAND2xp5_ASAP7_75t_L g1212 ( .A(n_1153), .B(n_1155), .Y(n_1212) );
AND2x2_ASAP7_75t_L g1213 ( .A(n_1153), .B(n_1034), .Y(n_1213) );
AND2x2_ASAP7_75t_L g1214 ( .A(n_1155), .B(n_1034), .Y(n_1214) );
AND2x2_ASAP7_75t_L g1215 ( .A(n_1167), .B(n_1044), .Y(n_1215) );
AND2x2_ASAP7_75t_L g1216 ( .A(n_1167), .B(n_1044), .Y(n_1216) );
OR2x2_ASAP7_75t_L g1217 ( .A(n_1185), .B(n_1109), .Y(n_1217) );
AND2x2_ASAP7_75t_L g1218 ( .A(n_1185), .B(n_1162), .Y(n_1218) );
INVx1_ASAP7_75t_L g1219 ( .A(n_1191), .Y(n_1219) );
OR2x2_ASAP7_75t_L g1220 ( .A(n_1170), .B(n_1138), .Y(n_1220) );
INVx1_ASAP7_75t_SL g1221 ( .A(n_1179), .Y(n_1221) );
AND2x2_ASAP7_75t_L g1222 ( .A(n_1195), .B(n_1162), .Y(n_1222) );
AND2x2_ASAP7_75t_L g1223 ( .A(n_1195), .B(n_1164), .Y(n_1223) );
NAND2xp5_ASAP7_75t_L g1224 ( .A(n_1171), .B(n_1142), .Y(n_1224) );
OR2x2_ASAP7_75t_L g1225 ( .A(n_1170), .B(n_1130), .Y(n_1225) );
INVx1_ASAP7_75t_L g1226 ( .A(n_1191), .Y(n_1226) );
AND2x2_ASAP7_75t_L g1227 ( .A(n_1213), .B(n_1164), .Y(n_1227) );
INVx1_ASAP7_75t_L g1228 ( .A(n_1194), .Y(n_1228) );
NAND2xp5_ASAP7_75t_L g1229 ( .A(n_1173), .B(n_1152), .Y(n_1229) );
INVx1_ASAP7_75t_L g1230 ( .A(n_1193), .Y(n_1230) );
NOR2xp33_ASAP7_75t_L g1231 ( .A(n_1208), .B(n_1036), .Y(n_1231) );
AND2x2_ASAP7_75t_L g1232 ( .A(n_1213), .B(n_1166), .Y(n_1232) );
AND2x2_ASAP7_75t_L g1233 ( .A(n_1214), .B(n_1166), .Y(n_1233) );
INVx1_ASAP7_75t_L g1234 ( .A(n_1201), .Y(n_1234) );
AND2x2_ASAP7_75t_L g1235 ( .A(n_1214), .B(n_1143), .Y(n_1235) );
AND2x2_ASAP7_75t_L g1236 ( .A(n_1196), .B(n_1145), .Y(n_1236) );
NAND2xp5_ASAP7_75t_L g1237 ( .A(n_1176), .B(n_1141), .Y(n_1237) );
NAND4xp25_ASAP7_75t_L g1238 ( .A(n_1180), .B(n_1118), .C(n_1123), .D(n_1129), .Y(n_1238) );
INVx1_ASAP7_75t_L g1239 ( .A(n_1201), .Y(n_1239) );
OR2x2_ASAP7_75t_L g1240 ( .A(n_1172), .B(n_1190), .Y(n_1240) );
NAND2x1p5_ASAP7_75t_L g1241 ( .A(n_1207), .B(n_1160), .Y(n_1241) );
AOI22xp33_ASAP7_75t_L g1242 ( .A1(n_1183), .A2(n_1165), .B1(n_1119), .B2(n_1169), .Y(n_1242) );
INVx2_ASAP7_75t_SL g1243 ( .A(n_1200), .Y(n_1243) );
NAND2xp5_ASAP7_75t_L g1244 ( .A(n_1198), .B(n_1130), .Y(n_1244) );
OR2x2_ASAP7_75t_L g1245 ( .A(n_1172), .B(n_1133), .Y(n_1245) );
AND2x2_ASAP7_75t_L g1246 ( .A(n_1174), .B(n_1124), .Y(n_1246) );
AND2x2_ASAP7_75t_L g1247 ( .A(n_1174), .B(n_1124), .Y(n_1247) );
NAND2xp5_ASAP7_75t_L g1248 ( .A(n_1212), .B(n_1168), .Y(n_1248) );
AND2x2_ASAP7_75t_L g1249 ( .A(n_1175), .B(n_1131), .Y(n_1249) );
NAND2xp5_ASAP7_75t_L g1250 ( .A(n_1182), .B(n_1135), .Y(n_1250) );
AND2x2_ASAP7_75t_L g1251 ( .A(n_1175), .B(n_1131), .Y(n_1251) );
HB1xp67_ASAP7_75t_L g1252 ( .A(n_1197), .Y(n_1252) );
NAND2xp5_ASAP7_75t_L g1253 ( .A(n_1210), .B(n_1128), .Y(n_1253) );
AND2x2_ASAP7_75t_L g1254 ( .A(n_1189), .B(n_1136), .Y(n_1254) );
NOR2x1_ASAP7_75t_L g1255 ( .A(n_1184), .B(n_1080), .Y(n_1255) );
OR2x2_ASAP7_75t_L g1256 ( .A(n_1177), .B(n_1157), .Y(n_1256) );
NAND2xp5_ASAP7_75t_L g1257 ( .A(n_1246), .B(n_1203), .Y(n_1257) );
OR2x2_ASAP7_75t_L g1258 ( .A(n_1240), .B(n_1181), .Y(n_1258) );
INVxp67_ASAP7_75t_L g1259 ( .A(n_1255), .Y(n_1259) );
INVx1_ASAP7_75t_L g1260 ( .A(n_1219), .Y(n_1260) );
AND2x2_ASAP7_75t_L g1261 ( .A(n_1232), .B(n_1189), .Y(n_1261) );
INVx1_ASAP7_75t_L g1262 ( .A(n_1226), .Y(n_1262) );
INVx1_ASAP7_75t_L g1263 ( .A(n_1226), .Y(n_1263) );
AND2x4_ASAP7_75t_L g1264 ( .A(n_1247), .B(n_1187), .Y(n_1264) );
AOI22xp5_ASAP7_75t_L g1265 ( .A1(n_1238), .A2(n_1127), .B1(n_1186), .B2(n_1209), .Y(n_1265) );
AND2x2_ASAP7_75t_L g1266 ( .A(n_1232), .B(n_1215), .Y(n_1266) );
NAND2xp5_ASAP7_75t_L g1267 ( .A(n_1249), .B(n_1205), .Y(n_1267) );
HB1xp67_ASAP7_75t_L g1268 ( .A(n_1252), .Y(n_1268) );
OAI22xp5_ASAP7_75t_L g1269 ( .A1(n_1242), .A2(n_1207), .B1(n_1178), .B2(n_1188), .Y(n_1269) );
AOI21xp33_ASAP7_75t_L g1270 ( .A1(n_1228), .A2(n_1151), .B(n_1199), .Y(n_1270) );
AND2x2_ASAP7_75t_L g1271 ( .A(n_1233), .B(n_1215), .Y(n_1271) );
INVx1_ASAP7_75t_L g1272 ( .A(n_1230), .Y(n_1272) );
INVx1_ASAP7_75t_L g1273 ( .A(n_1230), .Y(n_1273) );
AND2x2_ASAP7_75t_L g1274 ( .A(n_1233), .B(n_1216), .Y(n_1274) );
INVx1_ASAP7_75t_L g1275 ( .A(n_1234), .Y(n_1275) );
INVx1_ASAP7_75t_SL g1276 ( .A(n_1221), .Y(n_1276) );
INVx1_ASAP7_75t_L g1277 ( .A(n_1234), .Y(n_1277) );
AOI221x1_ASAP7_75t_L g1278 ( .A1(n_1231), .A2(n_1202), .B1(n_1079), .B2(n_1080), .C(n_1149), .Y(n_1278) );
NAND2xp5_ASAP7_75t_L g1279 ( .A(n_1249), .B(n_1206), .Y(n_1279) );
INVx1_ASAP7_75t_L g1280 ( .A(n_1239), .Y(n_1280) );
AND2x2_ASAP7_75t_L g1281 ( .A(n_1227), .B(n_1216), .Y(n_1281) );
AND2x2_ASAP7_75t_L g1282 ( .A(n_1227), .B(n_1206), .Y(n_1282) );
NOR2xp33_ASAP7_75t_L g1283 ( .A(n_1276), .B(n_1217), .Y(n_1283) );
INVx1_ASAP7_75t_L g1284 ( .A(n_1258), .Y(n_1284) );
A2O1A1Ixp33_ASAP7_75t_L g1285 ( .A1(n_1269), .A2(n_1243), .B(n_1211), .C(n_1103), .Y(n_1285) );
OAI31xp33_ASAP7_75t_L g1286 ( .A1(n_1259), .A2(n_1243), .A3(n_1241), .B(n_1211), .Y(n_1286) );
AND2x2_ASAP7_75t_L g1287 ( .A(n_1261), .B(n_1218), .Y(n_1287) );
AOI221xp5_ASAP7_75t_L g1288 ( .A1(n_1270), .A2(n_1229), .B1(n_1248), .B2(n_1237), .C(n_1250), .Y(n_1288) );
XNOR2x1_ASAP7_75t_L g1289 ( .A(n_1265), .B(n_1241), .Y(n_1289) );
INVx1_ASAP7_75t_L g1290 ( .A(n_1258), .Y(n_1290) );
AOI21xp5_ASAP7_75t_L g1291 ( .A1(n_1278), .A2(n_1188), .B(n_1178), .Y(n_1291) );
HB1xp67_ASAP7_75t_L g1292 ( .A(n_1268), .Y(n_1292) );
INVx1_ASAP7_75t_L g1293 ( .A(n_1260), .Y(n_1293) );
AND2x2_ASAP7_75t_L g1294 ( .A(n_1261), .B(n_1218), .Y(n_1294) );
OAI22xp5_ASAP7_75t_L g1295 ( .A1(n_1264), .A2(n_1188), .B1(n_1178), .B2(n_1220), .Y(n_1295) );
NAND2xp5_ASAP7_75t_L g1296 ( .A(n_1282), .B(n_1251), .Y(n_1296) );
NAND2xp5_ASAP7_75t_L g1297 ( .A(n_1282), .B(n_1251), .Y(n_1297) );
NAND2xp5_ASAP7_75t_L g1298 ( .A(n_1266), .B(n_1222), .Y(n_1298) );
INVx1_ASAP7_75t_L g1299 ( .A(n_1262), .Y(n_1299) );
INVx1_ASAP7_75t_L g1300 ( .A(n_1262), .Y(n_1300) );
INVxp67_ASAP7_75t_L g1301 ( .A(n_1292), .Y(n_1301) );
INVx1_ASAP7_75t_L g1302 ( .A(n_1284), .Y(n_1302) );
INVx1_ASAP7_75t_L g1303 ( .A(n_1290), .Y(n_1303) );
NOR2xp33_ASAP7_75t_L g1304 ( .A(n_1283), .B(n_1257), .Y(n_1304) );
AOI21xp5_ASAP7_75t_L g1305 ( .A1(n_1285), .A2(n_1264), .B(n_1224), .Y(n_1305) );
OAI21xp33_ASAP7_75t_L g1306 ( .A1(n_1289), .A2(n_1264), .B(n_1271), .Y(n_1306) );
AND2x2_ASAP7_75t_L g1307 ( .A(n_1287), .B(n_1271), .Y(n_1307) );
AOI22xp5_ASAP7_75t_L g1308 ( .A1(n_1289), .A2(n_1254), .B1(n_1274), .B2(n_1281), .Y(n_1308) );
OAI211xp5_ASAP7_75t_L g1309 ( .A1(n_1286), .A2(n_1150), .B(n_1110), .C(n_1125), .Y(n_1309) );
OAI31xp33_ASAP7_75t_L g1310 ( .A1(n_1295), .A2(n_1281), .A3(n_1274), .B(n_1103), .Y(n_1310) );
NOR2x1_ASAP7_75t_L g1311 ( .A(n_1291), .B(n_1160), .Y(n_1311) );
AOI22xp5_ASAP7_75t_L g1312 ( .A1(n_1288), .A2(n_1254), .B1(n_1223), .B2(n_1235), .Y(n_1312) );
INVx2_ASAP7_75t_L g1313 ( .A(n_1293), .Y(n_1313) );
INVx3_ASAP7_75t_L g1314 ( .A(n_1293), .Y(n_1314) );
AOI22xp5_ASAP7_75t_L g1315 ( .A1(n_1306), .A2(n_1294), .B1(n_1300), .B2(n_1299), .Y(n_1315) );
INVx1_ASAP7_75t_L g1316 ( .A(n_1301), .Y(n_1316) );
XNOR2xp5_ASAP7_75t_L g1317 ( .A(n_1308), .B(n_1112), .Y(n_1317) );
AOI211xp5_ASAP7_75t_L g1318 ( .A1(n_1309), .A2(n_1256), .B(n_1294), .C(n_1225), .Y(n_1318) );
NOR2xp33_ASAP7_75t_R g1319 ( .A(n_1304), .B(n_1007), .Y(n_1319) );
NAND4xp25_ASAP7_75t_L g1320 ( .A(n_1310), .B(n_1134), .C(n_1158), .D(n_1144), .Y(n_1320) );
AND2x2_ASAP7_75t_L g1321 ( .A(n_1307), .B(n_1298), .Y(n_1321) );
AOI221xp5_ASAP7_75t_L g1322 ( .A1(n_1312), .A2(n_1297), .B1(n_1296), .B2(n_1267), .C(n_1279), .Y(n_1322) );
AOI221xp5_ASAP7_75t_L g1323 ( .A1(n_1304), .A2(n_1263), .B1(n_1280), .B2(n_1277), .C(n_1275), .Y(n_1323) );
NOR4xp25_ASAP7_75t_L g1324 ( .A(n_1302), .B(n_1263), .C(n_1280), .D(n_1277), .Y(n_1324) );
NAND5xp2_ASAP7_75t_L g1325 ( .A(n_1318), .B(n_1305), .C(n_1204), .D(n_1115), .E(n_1079), .Y(n_1325) );
NAND2xp5_ASAP7_75t_L g1326 ( .A(n_1322), .B(n_1303), .Y(n_1326) );
AND2x4_ASAP7_75t_L g1327 ( .A(n_1316), .B(n_1311), .Y(n_1327) );
NOR3xp33_ASAP7_75t_SL g1328 ( .A(n_1320), .B(n_1076), .C(n_1244), .Y(n_1328) );
NAND2xp5_ASAP7_75t_L g1329 ( .A(n_1323), .B(n_1314), .Y(n_1329) );
OAI211xp5_ASAP7_75t_SL g1330 ( .A1(n_1315), .A2(n_1314), .B(n_1313), .C(n_1256), .Y(n_1330) );
AOI211x1_ASAP7_75t_L g1331 ( .A1(n_1319), .A2(n_1275), .B(n_1273), .C(n_1272), .Y(n_1331) );
NOR2x1_ASAP7_75t_L g1332 ( .A(n_1317), .B(n_1060), .Y(n_1332) );
INVx1_ASAP7_75t_L g1333 ( .A(n_1326), .Y(n_1333) );
NOR2x1_ASAP7_75t_L g1334 ( .A(n_1332), .B(n_1060), .Y(n_1334) );
OAI211xp5_ASAP7_75t_SL g1335 ( .A1(n_1329), .A2(n_1324), .B(n_1146), .C(n_1225), .Y(n_1335) );
NOR3xp33_ASAP7_75t_L g1336 ( .A(n_1325), .B(n_1321), .C(n_1068), .Y(n_1336) );
INVx1_ASAP7_75t_L g1337 ( .A(n_1327), .Y(n_1337) );
AND2x4_ASAP7_75t_L g1338 ( .A(n_1337), .B(n_1328), .Y(n_1338) );
OR2x2_ASAP7_75t_L g1339 ( .A(n_1333), .B(n_1245), .Y(n_1339) );
OR3x1_ASAP7_75t_L g1340 ( .A(n_1335), .B(n_1330), .C(n_1331), .Y(n_1340) );
INVx2_ASAP7_75t_L g1341 ( .A(n_1334), .Y(n_1341) );
INVx2_ASAP7_75t_L g1342 ( .A(n_1339), .Y(n_1342) );
NAND3xp33_ASAP7_75t_L g1343 ( .A(n_1338), .B(n_1336), .C(n_1273), .Y(n_1343) );
CKINVDCx20_ASAP7_75t_R g1344 ( .A(n_1342), .Y(n_1344) );
OAI21xp5_ASAP7_75t_L g1345 ( .A1(n_1343), .A2(n_1341), .B(n_1340), .Y(n_1345) );
INVxp33_ASAP7_75t_SL g1346 ( .A(n_1345), .Y(n_1346) );
AOI21xp33_ASAP7_75t_L g1347 ( .A1(n_1346), .A2(n_1344), .B(n_1272), .Y(n_1347) );
AO221x2_ASAP7_75t_L g1348 ( .A1(n_1347), .A2(n_1147), .B1(n_1154), .B2(n_1253), .C(n_1192), .Y(n_1348) );
AOI22xp5_ASAP7_75t_L g1349 ( .A1(n_1348), .A2(n_1107), .B1(n_1134), .B2(n_1236), .Y(n_1349) );
endmodule