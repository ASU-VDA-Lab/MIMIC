module fake_netlist_1_9035_n_714 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_714);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_714;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_383;
wire n_288;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_462;
wire n_232;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_307;
wire n_191;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_699;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_522;
wire n_264;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_363;
wire n_409;
wire n_315;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_428;
wire n_364;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_109;
wire n_99;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVxp33_ASAP7_75t_SL g81 ( .A(n_21), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_67), .Y(n_82) );
CKINVDCx5p33_ASAP7_75t_R g83 ( .A(n_48), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_46), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_76), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_66), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_19), .Y(n_87) );
INVxp67_ASAP7_75t_SL g88 ( .A(n_13), .Y(n_88) );
INVx2_ASAP7_75t_L g89 ( .A(n_22), .Y(n_89) );
HB1xp67_ASAP7_75t_L g90 ( .A(n_53), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_70), .Y(n_91) );
CKINVDCx5p33_ASAP7_75t_R g92 ( .A(n_79), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_71), .Y(n_93) );
CKINVDCx5p33_ASAP7_75t_R g94 ( .A(n_18), .Y(n_94) );
INVxp67_ASAP7_75t_SL g95 ( .A(n_35), .Y(n_95) );
CKINVDCx20_ASAP7_75t_R g96 ( .A(n_44), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_30), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_34), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_33), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_75), .Y(n_100) );
INVx2_ASAP7_75t_L g101 ( .A(n_28), .Y(n_101) );
CKINVDCx5p33_ASAP7_75t_R g102 ( .A(n_58), .Y(n_102) );
CKINVDCx20_ASAP7_75t_R g103 ( .A(n_18), .Y(n_103) );
INVxp67_ASAP7_75t_L g104 ( .A(n_57), .Y(n_104) );
INVxp33_ASAP7_75t_L g105 ( .A(n_29), .Y(n_105) );
CKINVDCx20_ASAP7_75t_R g106 ( .A(n_15), .Y(n_106) );
INVxp67_ASAP7_75t_L g107 ( .A(n_36), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_1), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_20), .Y(n_109) );
INVx3_ASAP7_75t_L g110 ( .A(n_2), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_39), .Y(n_111) );
BUFx3_ASAP7_75t_L g112 ( .A(n_23), .Y(n_112) );
CKINVDCx16_ASAP7_75t_R g113 ( .A(n_42), .Y(n_113) );
INVxp33_ASAP7_75t_L g114 ( .A(n_14), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_20), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_69), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_11), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_80), .Y(n_118) );
CKINVDCx5p33_ASAP7_75t_R g119 ( .A(n_5), .Y(n_119) );
OR2x2_ASAP7_75t_L g120 ( .A(n_13), .B(n_47), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_10), .Y(n_121) );
CKINVDCx20_ASAP7_75t_R g122 ( .A(n_12), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_74), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_62), .Y(n_124) );
BUFx6f_ASAP7_75t_L g125 ( .A(n_19), .Y(n_125) );
NOR2xp33_ASAP7_75t_L g126 ( .A(n_12), .B(n_24), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_32), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_16), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_5), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_77), .Y(n_130) );
BUFx6f_ASAP7_75t_L g131 ( .A(n_112), .Y(n_131) );
BUFx6f_ASAP7_75t_L g132 ( .A(n_112), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_110), .Y(n_133) );
BUFx6f_ASAP7_75t_L g134 ( .A(n_125), .Y(n_134) );
BUFx6f_ASAP7_75t_L g135 ( .A(n_125), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_110), .Y(n_136) );
NOR2x1_ASAP7_75t_L g137 ( .A(n_110), .B(n_40), .Y(n_137) );
CKINVDCx5p33_ASAP7_75t_R g138 ( .A(n_113), .Y(n_138) );
INVx2_ASAP7_75t_L g139 ( .A(n_89), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_90), .Y(n_140) );
HB1xp67_ASAP7_75t_L g141 ( .A(n_94), .Y(n_141) );
NAND2xp33_ASAP7_75t_SL g142 ( .A(n_114), .B(n_0), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_86), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_86), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_91), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_91), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_93), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_93), .Y(n_148) );
BUFx8_ASAP7_75t_L g149 ( .A(n_120), .Y(n_149) );
NAND2x1_ASAP7_75t_L g150 ( .A(n_87), .B(n_0), .Y(n_150) );
OA21x2_ASAP7_75t_L g151 ( .A1(n_97), .A2(n_130), .B(n_98), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_94), .B(n_1), .Y(n_152) );
INVx2_ASAP7_75t_L g153 ( .A(n_89), .Y(n_153) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_125), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_87), .Y(n_155) );
BUFx6f_ASAP7_75t_L g156 ( .A(n_125), .Y(n_156) );
OAI22xp5_ASAP7_75t_SL g157 ( .A1(n_103), .A2(n_2), .B1(n_3), .B2(n_4), .Y(n_157) );
INVx3_ASAP7_75t_L g158 ( .A(n_125), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_128), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_128), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_119), .B(n_3), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_129), .Y(n_162) );
INVx6_ASAP7_75t_L g163 ( .A(n_120), .Y(n_163) );
BUFx2_ASAP7_75t_L g164 ( .A(n_119), .Y(n_164) );
NOR2xp33_ASAP7_75t_L g165 ( .A(n_82), .B(n_4), .Y(n_165) );
AND2x2_ASAP7_75t_L g166 ( .A(n_105), .B(n_6), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_129), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_108), .B(n_109), .Y(n_168) );
INVx2_ASAP7_75t_L g169 ( .A(n_101), .Y(n_169) );
INVxp67_ASAP7_75t_L g170 ( .A(n_115), .Y(n_170) );
BUFx6f_ASAP7_75t_L g171 ( .A(n_101), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_117), .B(n_6), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_121), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_130), .Y(n_174) );
INVx5_ASAP7_75t_L g175 ( .A(n_81), .Y(n_175) );
AND3x4_ASAP7_75t_L g176 ( .A(n_137), .B(n_122), .C(n_106), .Y(n_176) );
AND2x6_ASAP7_75t_L g177 ( .A(n_166), .B(n_97), .Y(n_177) );
AND2x2_ASAP7_75t_SL g178 ( .A(n_166), .B(n_127), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_171), .Y(n_179) );
BUFx6f_ASAP7_75t_L g180 ( .A(n_171), .Y(n_180) );
AND2x4_ASAP7_75t_L g181 ( .A(n_140), .B(n_127), .Y(n_181) );
INVx2_ASAP7_75t_L g182 ( .A(n_171), .Y(n_182) );
AND2x4_ASAP7_75t_L g183 ( .A(n_133), .B(n_98), .Y(n_183) );
OR2x6_ASAP7_75t_SL g184 ( .A(n_138), .B(n_83), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_164), .B(n_83), .Y(n_185) );
AND2x4_ASAP7_75t_L g186 ( .A(n_136), .B(n_124), .Y(n_186) );
BUFx3_ASAP7_75t_L g187 ( .A(n_131), .Y(n_187) );
AND2x4_ASAP7_75t_L g188 ( .A(n_175), .B(n_124), .Y(n_188) );
AND2x2_ASAP7_75t_L g189 ( .A(n_164), .B(n_92), .Y(n_189) );
INVx4_ASAP7_75t_L g190 ( .A(n_163), .Y(n_190) );
INVx2_ASAP7_75t_L g191 ( .A(n_171), .Y(n_191) );
NOR2xp33_ASAP7_75t_L g192 ( .A(n_175), .B(n_104), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_171), .Y(n_193) );
AND2x4_ASAP7_75t_L g194 ( .A(n_175), .B(n_88), .Y(n_194) );
INVxp67_ASAP7_75t_L g195 ( .A(n_141), .Y(n_195) );
INVx1_ASAP7_75t_L g196 ( .A(n_151), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_151), .Y(n_197) );
BUFx3_ASAP7_75t_L g198 ( .A(n_131), .Y(n_198) );
NOR2xp33_ASAP7_75t_L g199 ( .A(n_175), .B(n_107), .Y(n_199) );
AND2x2_ASAP7_75t_L g200 ( .A(n_170), .B(n_92), .Y(n_200) );
NOR2xp33_ASAP7_75t_L g201 ( .A(n_175), .B(n_81), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_155), .Y(n_202) );
NOR2xp33_ASAP7_75t_L g203 ( .A(n_163), .B(n_100), .Y(n_203) );
AND2x2_ASAP7_75t_L g204 ( .A(n_163), .B(n_102), .Y(n_204) );
INVxp33_ASAP7_75t_L g205 ( .A(n_152), .Y(n_205) );
INVx1_ASAP7_75t_L g206 ( .A(n_151), .Y(n_206) );
INVx2_ASAP7_75t_L g207 ( .A(n_131), .Y(n_207) );
INVx4_ASAP7_75t_L g208 ( .A(n_163), .Y(n_208) );
INVx2_ASAP7_75t_L g209 ( .A(n_131), .Y(n_209) );
AND2x6_ASAP7_75t_L g210 ( .A(n_143), .B(n_84), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_151), .Y(n_211) );
OR2x2_ASAP7_75t_L g212 ( .A(n_138), .B(n_102), .Y(n_212) );
XNOR2xp5_ASAP7_75t_L g213 ( .A(n_157), .B(n_96), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_174), .B(n_111), .Y(n_214) );
INVxp67_ASAP7_75t_L g215 ( .A(n_149), .Y(n_215) );
AND2x2_ASAP7_75t_SL g216 ( .A(n_161), .B(n_126), .Y(n_216) );
OR2x6_ASAP7_75t_L g217 ( .A(n_150), .B(n_123), .Y(n_217) );
INVx2_ASAP7_75t_L g218 ( .A(n_131), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_139), .Y(n_219) );
INVx2_ASAP7_75t_L g220 ( .A(n_132), .Y(n_220) );
INVx2_ASAP7_75t_L g221 ( .A(n_132), .Y(n_221) );
INVx1_ASAP7_75t_L g222 ( .A(n_139), .Y(n_222) );
CKINVDCx16_ASAP7_75t_R g223 ( .A(n_142), .Y(n_223) );
BUFx10_ASAP7_75t_L g224 ( .A(n_143), .Y(n_224) );
INVx2_ASAP7_75t_L g225 ( .A(n_132), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_153), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_159), .Y(n_227) );
AND2x4_ASAP7_75t_L g228 ( .A(n_144), .B(n_147), .Y(n_228) );
AND2x2_ASAP7_75t_L g229 ( .A(n_160), .B(n_95), .Y(n_229) );
HB1xp67_ASAP7_75t_L g230 ( .A(n_149), .Y(n_230) );
NAND2xp5_ASAP7_75t_SL g231 ( .A(n_144), .B(n_118), .Y(n_231) );
INVx4_ASAP7_75t_SL g232 ( .A(n_132), .Y(n_232) );
INVx2_ASAP7_75t_L g233 ( .A(n_132), .Y(n_233) );
INVx4_ASAP7_75t_L g234 ( .A(n_158), .Y(n_234) );
AND2x2_ASAP7_75t_L g235 ( .A(n_162), .B(n_116), .Y(n_235) );
CKINVDCx5p33_ASAP7_75t_R g236 ( .A(n_149), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_153), .Y(n_237) );
AND2x2_ASAP7_75t_L g238 ( .A(n_167), .B(n_99), .Y(n_238) );
AND2x2_ASAP7_75t_L g239 ( .A(n_173), .B(n_85), .Y(n_239) );
AND2x2_ASAP7_75t_L g240 ( .A(n_145), .B(n_7), .Y(n_240) );
INVx2_ASAP7_75t_L g241 ( .A(n_134), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_169), .Y(n_242) );
AND2x4_ASAP7_75t_L g243 ( .A(n_145), .B(n_7), .Y(n_243) );
OAI22xp5_ASAP7_75t_L g244 ( .A1(n_146), .A2(n_8), .B1(n_9), .B2(n_10), .Y(n_244) );
BUFx8_ASAP7_75t_L g245 ( .A(n_189), .Y(n_245) );
AND2x4_ASAP7_75t_L g246 ( .A(n_194), .B(n_150), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_228), .Y(n_247) );
BUFx3_ASAP7_75t_L g248 ( .A(n_224), .Y(n_248) );
AOI22xp33_ASAP7_75t_L g249 ( .A1(n_178), .A2(n_142), .B1(n_148), .B2(n_146), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_228), .B(n_147), .Y(n_250) );
BUFx3_ASAP7_75t_L g251 ( .A(n_224), .Y(n_251) );
BUFx6f_ASAP7_75t_L g252 ( .A(n_224), .Y(n_252) );
INVx5_ASAP7_75t_L g253 ( .A(n_210), .Y(n_253) );
AND2x4_ASAP7_75t_L g254 ( .A(n_194), .B(n_148), .Y(n_254) );
HB1xp67_ASAP7_75t_L g255 ( .A(n_189), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_228), .B(n_165), .Y(n_256) );
AOI22xp33_ASAP7_75t_L g257 ( .A1(n_178), .A2(n_172), .B1(n_169), .B2(n_168), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_243), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_243), .Y(n_259) );
INVx2_ASAP7_75t_L g260 ( .A(n_207), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_200), .B(n_158), .Y(n_261) );
AND2x6_ASAP7_75t_SL g262 ( .A(n_217), .B(n_8), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_243), .Y(n_263) );
INVx5_ASAP7_75t_L g264 ( .A(n_210), .Y(n_264) );
AND2x4_ASAP7_75t_L g265 ( .A(n_194), .B(n_9), .Y(n_265) );
AOI22xp33_ASAP7_75t_L g266 ( .A1(n_177), .A2(n_158), .B1(n_156), .B2(n_154), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_219), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_219), .Y(n_268) );
OAI21xp33_ASAP7_75t_SL g269 ( .A1(n_196), .A2(n_11), .B(n_14), .Y(n_269) );
NAND3xp33_ASAP7_75t_SL g270 ( .A(n_176), .B(n_15), .C(n_16), .Y(n_270) );
INVx2_ASAP7_75t_L g271 ( .A(n_207), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_200), .B(n_156), .Y(n_272) );
INVx2_ASAP7_75t_L g273 ( .A(n_209), .Y(n_273) );
NOR2xp33_ASAP7_75t_L g274 ( .A(n_205), .B(n_55), .Y(n_274) );
INVx2_ASAP7_75t_L g275 ( .A(n_209), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_204), .B(n_156), .Y(n_276) );
BUFx3_ASAP7_75t_L g277 ( .A(n_210), .Y(n_277) );
INVx2_ASAP7_75t_L g278 ( .A(n_218), .Y(n_278) );
NAND2xp5_ASAP7_75t_SL g279 ( .A(n_181), .B(n_156), .Y(n_279) );
AND2x4_ASAP7_75t_L g280 ( .A(n_217), .B(n_181), .Y(n_280) );
AOI22xp33_ASAP7_75t_L g281 ( .A1(n_177), .A2(n_156), .B1(n_154), .B2(n_135), .Y(n_281) );
BUFx6f_ASAP7_75t_L g282 ( .A(n_187), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_204), .B(n_154), .Y(n_283) );
AOI22xp5_ASAP7_75t_L g284 ( .A1(n_177), .A2(n_135), .B1(n_134), .B2(n_154), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_222), .Y(n_285) );
AOI22xp33_ASAP7_75t_L g286 ( .A1(n_177), .A2(n_135), .B1(n_134), .B2(n_154), .Y(n_286) );
INVx2_ASAP7_75t_L g287 ( .A(n_218), .Y(n_287) );
INVx2_ASAP7_75t_L g288 ( .A(n_220), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_222), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_226), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_181), .B(n_135), .Y(n_291) );
CKINVDCx5p33_ASAP7_75t_R g292 ( .A(n_236), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_226), .Y(n_293) );
AND2x2_ASAP7_75t_L g294 ( .A(n_229), .B(n_17), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_237), .Y(n_295) );
INVx2_ASAP7_75t_L g296 ( .A(n_220), .Y(n_296) );
BUFx2_ASAP7_75t_L g297 ( .A(n_177), .Y(n_297) );
INVx2_ASAP7_75t_L g298 ( .A(n_221), .Y(n_298) );
BUFx3_ASAP7_75t_L g299 ( .A(n_210), .Y(n_299) );
INVx1_ASAP7_75t_SL g300 ( .A(n_212), .Y(n_300) );
NAND2x1p5_ASAP7_75t_L g301 ( .A(n_240), .B(n_135), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_237), .Y(n_302) );
AOI22xp33_ASAP7_75t_L g303 ( .A1(n_177), .A2(n_134), .B1(n_17), .B2(n_26), .Y(n_303) );
NOR2xp67_ASAP7_75t_L g304 ( .A(n_242), .B(n_25), .Y(n_304) );
BUFx3_ASAP7_75t_L g305 ( .A(n_210), .Y(n_305) );
INVx2_ASAP7_75t_L g306 ( .A(n_221), .Y(n_306) );
HB1xp67_ASAP7_75t_L g307 ( .A(n_195), .Y(n_307) );
INVx3_ASAP7_75t_L g308 ( .A(n_242), .Y(n_308) );
INVx2_ASAP7_75t_L g309 ( .A(n_225), .Y(n_309) );
AND2x6_ASAP7_75t_L g310 ( .A(n_196), .B(n_134), .Y(n_310) );
AOI22xp33_ASAP7_75t_L g311 ( .A1(n_240), .A2(n_27), .B1(n_31), .B2(n_37), .Y(n_311) );
INVx3_ASAP7_75t_L g312 ( .A(n_188), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_229), .B(n_38), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_197), .Y(n_314) );
INVx2_ASAP7_75t_L g315 ( .A(n_225), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_197), .Y(n_316) );
CKINVDCx5p33_ASAP7_75t_R g317 ( .A(n_236), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_190), .B(n_41), .Y(n_318) );
CKINVDCx11_ASAP7_75t_R g319 ( .A(n_262), .Y(n_319) );
AND2x2_ASAP7_75t_L g320 ( .A(n_280), .B(n_230), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_308), .Y(n_321) );
BUFx3_ASAP7_75t_L g322 ( .A(n_248), .Y(n_322) );
INVx2_ASAP7_75t_L g323 ( .A(n_314), .Y(n_323) );
AOI22xp33_ASAP7_75t_L g324 ( .A1(n_265), .A2(n_210), .B1(n_216), .B2(n_217), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_254), .B(n_202), .Y(n_325) );
AND2x4_ASAP7_75t_L g326 ( .A(n_280), .B(n_215), .Y(n_326) );
BUFx6f_ASAP7_75t_L g327 ( .A(n_252), .Y(n_327) );
AND2x4_ASAP7_75t_L g328 ( .A(n_280), .B(n_183), .Y(n_328) );
AOI22xp33_ASAP7_75t_L g329 ( .A1(n_265), .A2(n_216), .B1(n_217), .B2(n_190), .Y(n_329) );
BUFx6f_ASAP7_75t_L g330 ( .A(n_252), .Y(n_330) );
INVx2_ASAP7_75t_L g331 ( .A(n_314), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_254), .B(n_227), .Y(n_332) );
INVx2_ASAP7_75t_L g333 ( .A(n_316), .Y(n_333) );
BUFx12f_ASAP7_75t_L g334 ( .A(n_245), .Y(n_334) );
BUFx12f_ASAP7_75t_L g335 ( .A(n_245), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_308), .Y(n_336) );
INVx3_ASAP7_75t_L g337 ( .A(n_248), .Y(n_337) );
INVx2_ASAP7_75t_L g338 ( .A(n_316), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_308), .Y(n_339) );
AOI21xp5_ASAP7_75t_L g340 ( .A1(n_250), .A2(n_206), .B(n_211), .Y(n_340) );
INVx3_ASAP7_75t_L g341 ( .A(n_251), .Y(n_341) );
NAND2xp5_ASAP7_75t_SL g342 ( .A(n_251), .B(n_212), .Y(n_342) );
BUFx3_ASAP7_75t_L g343 ( .A(n_252), .Y(n_343) );
BUFx2_ASAP7_75t_L g344 ( .A(n_280), .Y(n_344) );
INVxp67_ASAP7_75t_SL g345 ( .A(n_252), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_267), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_267), .Y(n_347) );
O2A1O1Ixp33_ASAP7_75t_L g348 ( .A1(n_255), .A2(n_244), .B(n_185), .C(n_214), .Y(n_348) );
INVx5_ASAP7_75t_L g349 ( .A(n_252), .Y(n_349) );
HB1xp67_ASAP7_75t_L g350 ( .A(n_307), .Y(n_350) );
INVx2_ASAP7_75t_L g351 ( .A(n_268), .Y(n_351) );
INVx4_ASAP7_75t_L g352 ( .A(n_277), .Y(n_352) );
INVx2_ASAP7_75t_L g353 ( .A(n_268), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_285), .Y(n_354) );
INVxp67_ASAP7_75t_L g355 ( .A(n_245), .Y(n_355) );
AOI22xp5_ASAP7_75t_L g356 ( .A1(n_258), .A2(n_223), .B1(n_183), .B2(n_186), .Y(n_356) );
INVx2_ASAP7_75t_SL g357 ( .A(n_265), .Y(n_357) );
INVx3_ASAP7_75t_L g358 ( .A(n_277), .Y(n_358) );
BUFx2_ASAP7_75t_L g359 ( .A(n_297), .Y(n_359) );
AOI22xp33_ASAP7_75t_L g360 ( .A1(n_265), .A2(n_190), .B1(n_208), .B2(n_186), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_285), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_254), .B(n_208), .Y(n_362) );
INVx2_ASAP7_75t_L g363 ( .A(n_289), .Y(n_363) );
INVx4_ASAP7_75t_L g364 ( .A(n_299), .Y(n_364) );
OR2x6_ASAP7_75t_L g365 ( .A(n_297), .B(n_208), .Y(n_365) );
INVx2_ASAP7_75t_L g366 ( .A(n_289), .Y(n_366) );
NAND2x1p5_ASAP7_75t_L g367 ( .A(n_299), .B(n_188), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_290), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_254), .B(n_183), .Y(n_369) );
INVx2_ASAP7_75t_SL g370 ( .A(n_305), .Y(n_370) );
INVx2_ASAP7_75t_L g371 ( .A(n_290), .Y(n_371) );
OAI21xp33_ASAP7_75t_L g372 ( .A1(n_258), .A2(n_206), .B(n_211), .Y(n_372) );
AND2x2_ASAP7_75t_L g373 ( .A(n_300), .B(n_238), .Y(n_373) );
INVx3_ASAP7_75t_L g374 ( .A(n_305), .Y(n_374) );
NOR2xp33_ASAP7_75t_L g375 ( .A(n_246), .B(n_184), .Y(n_375) );
OAI22xp5_ASAP7_75t_L g376 ( .A1(n_324), .A2(n_263), .B1(n_259), .B2(n_302), .Y(n_376) );
INVxp33_ASAP7_75t_L g377 ( .A(n_350), .Y(n_377) );
NAND2xp5_ASAP7_75t_SL g378 ( .A(n_322), .B(n_253), .Y(n_378) );
BUFx2_ASAP7_75t_L g379 ( .A(n_328), .Y(n_379) );
INVx3_ASAP7_75t_L g380 ( .A(n_349), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_351), .B(n_294), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_351), .Y(n_382) );
BUFx3_ASAP7_75t_L g383 ( .A(n_349), .Y(n_383) );
OAI21xp5_ASAP7_75t_L g384 ( .A1(n_340), .A2(n_269), .B(n_263), .Y(n_384) );
AO31x2_ASAP7_75t_L g385 ( .A1(n_351), .A2(n_302), .A3(n_295), .B(n_293), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_353), .Y(n_386) );
O2A1O1Ixp33_ASAP7_75t_SL g387 ( .A1(n_323), .A2(n_318), .B(n_313), .C(n_295), .Y(n_387) );
AND2x2_ASAP7_75t_L g388 ( .A(n_373), .B(n_294), .Y(n_388) );
AND2x4_ASAP7_75t_SL g389 ( .A(n_328), .B(n_247), .Y(n_389) );
INVx2_ASAP7_75t_SL g390 ( .A(n_349), .Y(n_390) );
AOI22xp33_ASAP7_75t_L g391 ( .A1(n_373), .A2(n_176), .B1(n_246), .B2(n_249), .Y(n_391) );
AO221x2_ASAP7_75t_L g392 ( .A1(n_353), .A2(n_269), .B1(n_259), .B2(n_293), .C(n_247), .Y(n_392) );
INVx2_ASAP7_75t_SL g393 ( .A(n_349), .Y(n_393) );
OR2x2_ASAP7_75t_L g394 ( .A(n_320), .B(n_292), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_353), .B(n_246), .Y(n_395) );
INVx2_ASAP7_75t_L g396 ( .A(n_323), .Y(n_396) );
AOI22xp33_ASAP7_75t_L g397 ( .A1(n_328), .A2(n_246), .B1(n_270), .B2(n_312), .Y(n_397) );
AOI22xp5_ASAP7_75t_L g398 ( .A1(n_357), .A2(n_257), .B1(n_256), .B2(n_203), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_363), .Y(n_399) );
AND2x2_ASAP7_75t_L g400 ( .A(n_328), .B(n_363), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_363), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_366), .Y(n_402) );
INVx1_ASAP7_75t_SL g403 ( .A(n_349), .Y(n_403) );
HB1xp67_ASAP7_75t_L g404 ( .A(n_349), .Y(n_404) );
AOI22xp33_ASAP7_75t_L g405 ( .A1(n_375), .A2(n_312), .B1(n_188), .B2(n_292), .Y(n_405) );
AND2x2_ASAP7_75t_L g406 ( .A(n_366), .B(n_235), .Y(n_406) );
AND2x2_ASAP7_75t_L g407 ( .A(n_366), .B(n_235), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_371), .Y(n_408) );
AOI22xp33_ASAP7_75t_L g409 ( .A1(n_344), .A2(n_326), .B1(n_320), .B2(n_357), .Y(n_409) );
AOI22xp33_ASAP7_75t_L g410 ( .A1(n_371), .A2(n_186), .B1(n_312), .B2(n_239), .Y(n_410) );
INVx2_ASAP7_75t_L g411 ( .A(n_396), .Y(n_411) );
INVx2_ASAP7_75t_L g412 ( .A(n_396), .Y(n_412) );
BUFx12f_ASAP7_75t_L g413 ( .A(n_390), .Y(n_413) );
NAND2xp5_ASAP7_75t_SL g414 ( .A(n_403), .B(n_322), .Y(n_414) );
AOI221xp5_ASAP7_75t_L g415 ( .A1(n_391), .A2(n_348), .B1(n_239), .B2(n_355), .C(n_317), .Y(n_415) );
AOI211xp5_ASAP7_75t_SL g416 ( .A1(n_404), .A2(n_274), .B(n_337), .C(n_341), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_388), .B(n_406), .Y(n_417) );
OAI21xp33_ASAP7_75t_L g418 ( .A1(n_398), .A2(n_329), .B(n_356), .Y(n_418) );
NAND2x1p5_ASAP7_75t_L g419 ( .A(n_383), .B(n_327), .Y(n_419) );
OAI22xp5_ASAP7_75t_L g420 ( .A1(n_381), .A2(n_360), .B1(n_356), .B2(n_371), .Y(n_420) );
BUFx4f_ASAP7_75t_SL g421 ( .A(n_383), .Y(n_421) );
INVx2_ASAP7_75t_L g422 ( .A(n_396), .Y(n_422) );
OAI21xp5_ASAP7_75t_SL g423 ( .A1(n_397), .A2(n_213), .B(n_342), .Y(n_423) );
AND2x2_ASAP7_75t_L g424 ( .A(n_406), .B(n_323), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_382), .Y(n_425) );
INVx3_ASAP7_75t_L g426 ( .A(n_383), .Y(n_426) );
AOI222xp33_ASAP7_75t_L g427 ( .A1(n_388), .A2(n_319), .B1(n_334), .B2(n_335), .C1(n_213), .C2(n_238), .Y(n_427) );
AOI221xp5_ASAP7_75t_L g428 ( .A1(n_377), .A2(n_317), .B1(n_326), .B2(n_325), .C(n_332), .Y(n_428) );
OAI22xp5_ASAP7_75t_L g429 ( .A1(n_381), .A2(n_338), .B1(n_333), .B2(n_331), .Y(n_429) );
INVx3_ASAP7_75t_L g430 ( .A(n_380), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_382), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_386), .Y(n_432) );
AOI21xp5_ASAP7_75t_L g433 ( .A1(n_387), .A2(n_372), .B(n_333), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_386), .Y(n_434) );
AOI221xp5_ASAP7_75t_L g435 ( .A1(n_376), .A2(n_326), .B1(n_325), .B2(n_332), .C(n_369), .Y(n_435) );
AOI22xp33_ASAP7_75t_L g436 ( .A1(n_392), .A2(n_335), .B1(n_334), .B2(n_344), .Y(n_436) );
AOI22xp33_ASAP7_75t_SL g437 ( .A1(n_392), .A2(n_334), .B1(n_335), .B2(n_326), .Y(n_437) );
NAND3xp33_ASAP7_75t_L g438 ( .A(n_392), .B(n_311), .C(n_303), .Y(n_438) );
INVx1_ASAP7_75t_SL g439 ( .A(n_403), .Y(n_439) );
AO21x2_ASAP7_75t_L g440 ( .A1(n_384), .A2(n_304), .B(n_372), .Y(n_440) );
AO21x2_ASAP7_75t_L g441 ( .A1(n_433), .A2(n_384), .B(n_376), .Y(n_441) );
INVx2_ASAP7_75t_L g442 ( .A(n_411), .Y(n_442) );
INVx2_ASAP7_75t_L g443 ( .A(n_411), .Y(n_443) );
OAI22xp33_ASAP7_75t_L g444 ( .A1(n_435), .A2(n_399), .B1(n_408), .B2(n_401), .Y(n_444) );
HB1xp67_ASAP7_75t_L g445 ( .A(n_412), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_425), .Y(n_446) );
OAI221xp5_ASAP7_75t_L g447 ( .A1(n_423), .A2(n_405), .B1(n_394), .B2(n_409), .C(n_410), .Y(n_447) );
OAI22xp5_ASAP7_75t_L g448 ( .A1(n_437), .A2(n_394), .B1(n_408), .B2(n_399), .Y(n_448) );
OAI222xp33_ASAP7_75t_L g449 ( .A1(n_436), .A2(n_402), .B1(n_401), .B2(n_390), .C1(n_393), .C2(n_404), .Y(n_449) );
AOI31xp33_ASAP7_75t_L g450 ( .A1(n_427), .A2(n_390), .A3(n_393), .B(n_184), .Y(n_450) );
AOI21xp5_ASAP7_75t_L g451 ( .A1(n_429), .A2(n_392), .B(n_402), .Y(n_451) );
AND2x2_ASAP7_75t_L g452 ( .A(n_424), .B(n_407), .Y(n_452) );
OAI21xp5_ASAP7_75t_L g453 ( .A1(n_438), .A2(n_398), .B(n_410), .Y(n_453) );
INVx1_ASAP7_75t_SL g454 ( .A(n_421), .Y(n_454) );
AOI21xp5_ASAP7_75t_L g455 ( .A1(n_440), .A2(n_392), .B(n_338), .Y(n_455) );
OR2x6_ASAP7_75t_L g456 ( .A(n_413), .B(n_393), .Y(n_456) );
AOI221xp5_ASAP7_75t_L g457 ( .A1(n_415), .A2(n_407), .B1(n_261), .B2(n_400), .C(n_231), .Y(n_457) );
OAI31xp33_ASAP7_75t_L g458 ( .A1(n_423), .A2(n_389), .A3(n_379), .B(n_400), .Y(n_458) );
AND2x4_ASAP7_75t_L g459 ( .A(n_424), .B(n_385), .Y(n_459) );
OAI31xp33_ASAP7_75t_L g460 ( .A1(n_418), .A2(n_389), .A3(n_379), .B(n_201), .Y(n_460) );
BUFx2_ASAP7_75t_L g461 ( .A(n_413), .Y(n_461) );
AND2x4_ASAP7_75t_L g462 ( .A(n_425), .B(n_385), .Y(n_462) );
AND2x2_ASAP7_75t_L g463 ( .A(n_417), .B(n_389), .Y(n_463) );
AND2x2_ASAP7_75t_L g464 ( .A(n_427), .B(n_395), .Y(n_464) );
OAI33xp33_ASAP7_75t_L g465 ( .A1(n_420), .A2(n_272), .A3(n_283), .B1(n_276), .B2(n_291), .B3(n_395), .Y(n_465) );
AOI22xp33_ASAP7_75t_L g466 ( .A1(n_418), .A2(n_346), .B1(n_354), .B2(n_347), .Y(n_466) );
NAND3xp33_ASAP7_75t_L g467 ( .A(n_416), .B(n_192), .C(n_199), .Y(n_467) );
OAI21xp33_ASAP7_75t_SL g468 ( .A1(n_431), .A2(n_380), .B(n_346), .Y(n_468) );
AOI221xp5_ASAP7_75t_L g469 ( .A1(n_428), .A2(n_369), .B1(n_354), .B2(n_361), .C(n_368), .Y(n_469) );
AOI22xp33_ASAP7_75t_SL g470 ( .A1(n_431), .A2(n_380), .B1(n_361), .B2(n_347), .Y(n_470) );
OAI22xp5_ASAP7_75t_L g471 ( .A1(n_432), .A2(n_368), .B1(n_338), .B2(n_333), .Y(n_471) );
AOI221xp5_ASAP7_75t_L g472 ( .A1(n_432), .A2(n_279), .B1(n_362), .B2(n_339), .C(n_336), .Y(n_472) );
OAI21xp33_ASAP7_75t_L g473 ( .A1(n_438), .A2(n_301), .B(n_198), .Y(n_473) );
NAND3xp33_ASAP7_75t_L g474 ( .A(n_434), .B(n_304), .C(n_180), .Y(n_474) );
NAND4xp25_ASAP7_75t_L g475 ( .A(n_434), .B(n_266), .C(n_187), .D(n_198), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_412), .Y(n_476) );
OAI33xp33_ASAP7_75t_L g477 ( .A1(n_414), .A2(n_179), .A3(n_193), .B1(n_233), .B2(n_182), .B3(n_191), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_422), .Y(n_478) );
NAND2xp5_ASAP7_75t_SL g479 ( .A(n_450), .B(n_439), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_462), .Y(n_480) );
NOR3xp33_ASAP7_75t_L g481 ( .A(n_447), .B(n_430), .C(n_426), .Y(n_481) );
OR2x2_ASAP7_75t_L g482 ( .A(n_459), .B(n_422), .Y(n_482) );
AND2x2_ASAP7_75t_SL g483 ( .A(n_462), .B(n_426), .Y(n_483) );
OAI31xp33_ASAP7_75t_L g484 ( .A1(n_448), .A2(n_439), .A3(n_426), .B(n_380), .Y(n_484) );
AOI22xp33_ASAP7_75t_L g485 ( .A1(n_458), .A2(n_430), .B1(n_359), .B2(n_365), .Y(n_485) );
AOI33xp33_ASAP7_75t_L g486 ( .A1(n_464), .A2(n_193), .A3(n_179), .B1(n_233), .B2(n_182), .B3(n_191), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_462), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_446), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_445), .Y(n_489) );
AND2x2_ASAP7_75t_L g490 ( .A(n_459), .B(n_385), .Y(n_490) );
AND2x2_ASAP7_75t_L g491 ( .A(n_459), .B(n_385), .Y(n_491) );
NAND3xp33_ASAP7_75t_L g492 ( .A(n_470), .B(n_180), .C(n_430), .Y(n_492) );
OR2x2_ASAP7_75t_L g493 ( .A(n_445), .B(n_385), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_476), .Y(n_494) );
BUFx3_ASAP7_75t_L g495 ( .A(n_456), .Y(n_495) );
AND2x2_ASAP7_75t_L g496 ( .A(n_452), .B(n_385), .Y(n_496) );
INVx2_ASAP7_75t_L g497 ( .A(n_442), .Y(n_497) );
AND2x2_ASAP7_75t_SL g498 ( .A(n_461), .B(n_359), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_463), .B(n_331), .Y(n_499) );
NOR2x1_ASAP7_75t_L g500 ( .A(n_456), .B(n_322), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_478), .Y(n_501) );
AND2x2_ASAP7_75t_L g502 ( .A(n_442), .B(n_440), .Y(n_502) );
AND3x1_ASAP7_75t_L g503 ( .A(n_469), .B(n_337), .C(n_341), .Y(n_503) );
AOI211xp5_ASAP7_75t_L g504 ( .A1(n_444), .A2(n_180), .B(n_378), .C(n_337), .Y(n_504) );
HB1xp67_ASAP7_75t_L g505 ( .A(n_443), .Y(n_505) );
AND2x4_ASAP7_75t_SL g506 ( .A(n_443), .B(n_331), .Y(n_506) );
INVx2_ASAP7_75t_L g507 ( .A(n_441), .Y(n_507) );
INVx2_ASAP7_75t_L g508 ( .A(n_441), .Y(n_508) );
OR2x2_ASAP7_75t_L g509 ( .A(n_453), .B(n_419), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_468), .Y(n_510) );
NAND3xp33_ASAP7_75t_SL g511 ( .A(n_454), .B(n_419), .C(n_367), .Y(n_511) );
AND2x2_ASAP7_75t_L g512 ( .A(n_466), .B(n_440), .Y(n_512) );
AOI221xp5_ASAP7_75t_L g513 ( .A1(n_444), .A2(n_301), .B1(n_336), .B2(n_339), .C(n_321), .Y(n_513) );
AND2x2_ASAP7_75t_L g514 ( .A(n_466), .B(n_419), .Y(n_514) );
OR2x2_ASAP7_75t_L g515 ( .A(n_455), .B(n_301), .Y(n_515) );
INVx4_ASAP7_75t_L g516 ( .A(n_470), .Y(n_516) );
OAI221xp5_ASAP7_75t_L g517 ( .A1(n_457), .A2(n_281), .B1(n_286), .B2(n_284), .C(n_367), .Y(n_517) );
OAI31xp33_ASAP7_75t_L g518 ( .A1(n_449), .A2(n_367), .A3(n_337), .B(n_341), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_451), .Y(n_519) );
AOI222xp33_ASAP7_75t_L g520 ( .A1(n_465), .A2(n_321), .B1(n_232), .B2(n_341), .C1(n_310), .C2(n_343), .Y(n_520) );
OR2x2_ASAP7_75t_L g521 ( .A(n_471), .B(n_343), .Y(n_521) );
AND2x2_ASAP7_75t_L g522 ( .A(n_473), .B(n_327), .Y(n_522) );
AOI22xp33_ASAP7_75t_L g523 ( .A1(n_460), .A2(n_365), .B1(n_343), .B2(n_327), .Y(n_523) );
AOI211x1_ASAP7_75t_L g524 ( .A1(n_475), .A2(n_43), .B(n_45), .C(n_49), .Y(n_524) );
HB1xp67_ASAP7_75t_L g525 ( .A(n_472), .Y(n_525) );
OAI21xp33_ASAP7_75t_L g526 ( .A1(n_467), .A2(n_180), .B(n_241), .Y(n_526) );
OR2x2_ASAP7_75t_L g527 ( .A(n_474), .B(n_365), .Y(n_527) );
AND2x4_ASAP7_75t_SL g528 ( .A(n_477), .B(n_327), .Y(n_528) );
INVx2_ASAP7_75t_L g529 ( .A(n_445), .Y(n_529) );
OAI33xp33_ASAP7_75t_L g530 ( .A1(n_448), .A2(n_241), .A3(n_315), .B1(n_309), .B2(n_306), .B3(n_298), .Y(n_530) );
INVx2_ASAP7_75t_L g531 ( .A(n_445), .Y(n_531) );
AND2x2_ASAP7_75t_L g532 ( .A(n_490), .B(n_180), .Y(n_532) );
INVx1_ASAP7_75t_SL g533 ( .A(n_506), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_488), .Y(n_534) );
AND2x2_ASAP7_75t_L g535 ( .A(n_490), .B(n_50), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_496), .B(n_327), .Y(n_536) );
AND2x2_ASAP7_75t_L g537 ( .A(n_491), .B(n_51), .Y(n_537) );
OR2x2_ASAP7_75t_L g538 ( .A(n_482), .B(n_365), .Y(n_538) );
AND2x2_ASAP7_75t_L g539 ( .A(n_491), .B(n_52), .Y(n_539) );
AND2x2_ASAP7_75t_L g540 ( .A(n_480), .B(n_54), .Y(n_540) );
NAND3xp33_ASAP7_75t_L g541 ( .A(n_524), .B(n_330), .C(n_365), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_488), .Y(n_542) );
AND2x2_ASAP7_75t_L g543 ( .A(n_480), .B(n_56), .Y(n_543) );
AND2x2_ASAP7_75t_L g544 ( .A(n_487), .B(n_59), .Y(n_544) );
AND2x2_ASAP7_75t_L g545 ( .A(n_487), .B(n_60), .Y(n_545) );
OR2x2_ASAP7_75t_L g546 ( .A(n_493), .B(n_330), .Y(n_546) );
INVx2_ASAP7_75t_L g547 ( .A(n_497), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_494), .Y(n_548) );
OR2x2_ASAP7_75t_L g549 ( .A(n_493), .B(n_330), .Y(n_549) );
AND2x2_ASAP7_75t_L g550 ( .A(n_519), .B(n_61), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_501), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_489), .Y(n_552) );
HB1xp67_ASAP7_75t_L g553 ( .A(n_505), .Y(n_553) );
OAI322xp33_ASAP7_75t_L g554 ( .A1(n_516), .A2(n_271), .A3(n_309), .B1(n_306), .B2(n_298), .C1(n_296), .C2(n_288), .Y(n_554) );
OR2x2_ASAP7_75t_L g555 ( .A(n_531), .B(n_330), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_489), .Y(n_556) );
AND2x2_ASAP7_75t_L g557 ( .A(n_519), .B(n_63), .Y(n_557) );
XNOR2xp5_ASAP7_75t_L g558 ( .A(n_498), .B(n_370), .Y(n_558) );
NOR2xp33_ASAP7_75t_L g559 ( .A(n_516), .B(n_64), .Y(n_559) );
AOI21xp5_ASAP7_75t_L g560 ( .A1(n_504), .A2(n_330), .B(n_345), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_525), .B(n_65), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_529), .Y(n_562) );
OAI31xp33_ASAP7_75t_L g563 ( .A1(n_479), .A2(n_370), .A3(n_374), .B(n_358), .Y(n_563) );
AND2x2_ASAP7_75t_L g564 ( .A(n_529), .B(n_68), .Y(n_564) );
AND2x2_ASAP7_75t_L g565 ( .A(n_531), .B(n_72), .Y(n_565) );
AND2x4_ASAP7_75t_L g566 ( .A(n_510), .B(n_73), .Y(n_566) );
OR2x2_ASAP7_75t_L g567 ( .A(n_499), .B(n_78), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_516), .B(n_232), .Y(n_568) );
AOI31xp33_ASAP7_75t_L g569 ( .A1(n_503), .A2(n_352), .A3(n_364), .B(n_273), .Y(n_569) );
AND2x2_ASAP7_75t_L g570 ( .A(n_483), .B(n_232), .Y(n_570) );
AND2x2_ASAP7_75t_L g571 ( .A(n_483), .B(n_232), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_510), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_509), .Y(n_573) );
INVx1_ASAP7_75t_SL g574 ( .A(n_498), .Y(n_574) );
OAI21xp33_ASAP7_75t_SL g575 ( .A1(n_484), .A2(n_364), .B(n_352), .Y(n_575) );
AND2x4_ASAP7_75t_L g576 ( .A(n_514), .B(n_364), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_481), .B(n_310), .Y(n_577) );
INVx2_ASAP7_75t_L g578 ( .A(n_502), .Y(n_578) );
AND2x2_ASAP7_75t_L g579 ( .A(n_514), .B(n_287), .Y(n_579) );
AND2x4_ASAP7_75t_L g580 ( .A(n_502), .B(n_364), .Y(n_580) );
OAI22xp33_ASAP7_75t_SL g581 ( .A1(n_495), .A2(n_352), .B1(n_358), .B2(n_374), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_511), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_486), .B(n_310), .Y(n_583) );
OR2x2_ASAP7_75t_L g584 ( .A(n_521), .B(n_352), .Y(n_584) );
AND2x2_ASAP7_75t_L g585 ( .A(n_512), .B(n_278), .Y(n_585) );
OAI22xp5_ASAP7_75t_L g586 ( .A1(n_485), .A2(n_358), .B1(n_374), .B2(n_253), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_551), .Y(n_587) );
INVx2_ASAP7_75t_SL g588 ( .A(n_533), .Y(n_588) );
NAND3xp33_ASAP7_75t_L g589 ( .A(n_582), .B(n_520), .C(n_507), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_534), .Y(n_590) );
AND2x4_ASAP7_75t_L g591 ( .A(n_572), .B(n_507), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_552), .B(n_508), .Y(n_592) );
NAND2xp5_ASAP7_75t_SL g593 ( .A(n_574), .B(n_492), .Y(n_593) );
OAI31xp33_ASAP7_75t_SL g594 ( .A1(n_559), .A2(n_500), .A3(n_513), .B(n_526), .Y(n_594) );
OR2x2_ASAP7_75t_L g595 ( .A(n_553), .B(n_515), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_542), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_556), .B(n_508), .Y(n_597) );
INVx1_ASAP7_75t_SL g598 ( .A(n_546), .Y(n_598) );
NOR3xp33_ASAP7_75t_L g599 ( .A(n_561), .B(n_530), .C(n_527), .Y(n_599) );
OAI21xp33_ASAP7_75t_L g600 ( .A1(n_559), .A2(n_523), .B(n_528), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_548), .B(n_521), .Y(n_601) );
OAI211xp5_ASAP7_75t_L g602 ( .A1(n_575), .A2(n_518), .B(n_527), .C(n_517), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_562), .B(n_522), .Y(n_603) );
AND2x4_ASAP7_75t_L g604 ( .A(n_573), .B(n_522), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_578), .B(n_310), .Y(n_605) );
HB1xp67_ASAP7_75t_L g606 ( .A(n_549), .Y(n_606) );
AND2x2_ASAP7_75t_L g607 ( .A(n_532), .B(n_282), .Y(n_607) );
NOR2xp67_ASAP7_75t_L g608 ( .A(n_566), .B(n_253), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_585), .B(n_310), .Y(n_609) );
OAI21xp5_ASAP7_75t_L g610 ( .A1(n_569), .A2(n_310), .B(n_315), .Y(n_610) );
INVxp67_ASAP7_75t_SL g611 ( .A(n_555), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_585), .B(n_275), .Y(n_612) );
AOI21xp5_ASAP7_75t_L g613 ( .A1(n_554), .A2(n_374), .B(n_358), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_547), .B(n_273), .Y(n_614) );
OR2x2_ASAP7_75t_L g615 ( .A(n_536), .B(n_296), .Y(n_615) );
AOI22xp33_ASAP7_75t_L g616 ( .A1(n_576), .A2(n_282), .B1(n_260), .B2(n_275), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_535), .B(n_260), .Y(n_617) );
NAND2xp5_ASAP7_75t_SL g618 ( .A(n_566), .B(n_253), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_550), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_535), .B(n_288), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_550), .Y(n_621) );
NOR2xp33_ASAP7_75t_SL g622 ( .A(n_566), .B(n_253), .Y(n_622) );
INVxp67_ASAP7_75t_L g623 ( .A(n_537), .Y(n_623) );
OR2x2_ASAP7_75t_L g624 ( .A(n_579), .B(n_234), .Y(n_624) );
XNOR2x2_ASAP7_75t_L g625 ( .A(n_558), .B(n_253), .Y(n_625) );
AO211x2_ASAP7_75t_L g626 ( .A1(n_541), .A2(n_264), .B(n_234), .C(n_282), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_557), .Y(n_627) );
NAND3xp33_ASAP7_75t_L g628 ( .A(n_563), .B(n_282), .C(n_234), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_587), .Y(n_629) );
OAI221xp5_ASAP7_75t_L g630 ( .A1(n_594), .A2(n_568), .B1(n_577), .B2(n_567), .C(n_539), .Y(n_630) );
AND2x4_ASAP7_75t_L g631 ( .A(n_604), .B(n_576), .Y(n_631) );
O2A1O1Ixp33_ASAP7_75t_L g632 ( .A1(n_599), .A2(n_581), .B(n_539), .C(n_586), .Y(n_632) );
AOI21xp5_ASAP7_75t_L g633 ( .A1(n_610), .A2(n_560), .B(n_557), .Y(n_633) );
INVxp67_ASAP7_75t_SL g634 ( .A(n_606), .Y(n_634) );
INVx2_ASAP7_75t_SL g635 ( .A(n_588), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_590), .Y(n_636) );
XOR2x1_ASAP7_75t_L g637 ( .A(n_626), .B(n_545), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_596), .Y(n_638) );
A2O1A1Ixp33_ASAP7_75t_L g639 ( .A1(n_600), .A2(n_570), .B(n_571), .C(n_543), .Y(n_639) );
OR2x2_ASAP7_75t_L g640 ( .A(n_611), .B(n_580), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_595), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_592), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_597), .Y(n_643) );
AOI211x1_ASAP7_75t_L g644 ( .A1(n_602), .A2(n_540), .B(n_543), .C(n_545), .Y(n_644) );
HB1xp67_ASAP7_75t_L g645 ( .A(n_598), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_597), .Y(n_646) );
BUFx2_ASAP7_75t_L g647 ( .A(n_604), .Y(n_647) );
NAND2x1p5_ASAP7_75t_L g648 ( .A(n_608), .B(n_565), .Y(n_648) );
A2O1A1Ixp33_ASAP7_75t_L g649 ( .A1(n_622), .A2(n_571), .B(n_570), .C(n_544), .Y(n_649) );
OAI31xp33_ASAP7_75t_L g650 ( .A1(n_618), .A2(n_544), .A3(n_538), .B(n_584), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_603), .Y(n_651) );
OAI21xp33_ASAP7_75t_L g652 ( .A1(n_589), .A2(n_564), .B(n_565), .Y(n_652) );
INVx1_ASAP7_75t_L g653 ( .A(n_603), .Y(n_653) );
A2O1A1Ixp33_ASAP7_75t_SL g654 ( .A1(n_610), .A2(n_583), .B(n_282), .C(n_264), .Y(n_654) );
INVx1_ASAP7_75t_SL g655 ( .A(n_624), .Y(n_655) );
INVx1_ASAP7_75t_SL g656 ( .A(n_615), .Y(n_656) );
AOI21xp33_ASAP7_75t_SL g657 ( .A1(n_623), .A2(n_264), .B(n_593), .Y(n_657) );
INVx2_ASAP7_75t_L g658 ( .A(n_591), .Y(n_658) );
NOR2x1_ASAP7_75t_L g659 ( .A(n_628), .B(n_625), .Y(n_659) );
NOR2xp33_ASAP7_75t_L g660 ( .A(n_601), .B(n_627), .Y(n_660) );
OAI22xp33_ASAP7_75t_L g661 ( .A1(n_621), .A2(n_619), .B1(n_620), .B2(n_617), .Y(n_661) );
INVx1_ASAP7_75t_L g662 ( .A(n_612), .Y(n_662) );
A2O1A1Ixp33_ASAP7_75t_L g663 ( .A1(n_613), .A2(n_616), .B(n_607), .C(n_609), .Y(n_663) );
XOR2x2_ASAP7_75t_L g664 ( .A(n_614), .B(n_605), .Y(n_664) );
XOR2xp5_ASAP7_75t_L g665 ( .A(n_605), .B(n_213), .Y(n_665) );
XOR2x2_ASAP7_75t_L g666 ( .A(n_625), .B(n_176), .Y(n_666) );
XNOR2xp5_ASAP7_75t_L g667 ( .A(n_588), .B(n_176), .Y(n_667) );
INVx1_ASAP7_75t_L g668 ( .A(n_587), .Y(n_668) );
HB1xp67_ASAP7_75t_L g669 ( .A(n_611), .Y(n_669) );
XOR2xp5_ASAP7_75t_L g670 ( .A(n_606), .B(n_213), .Y(n_670) );
INVx1_ASAP7_75t_L g671 ( .A(n_587), .Y(n_671) );
AOI22x1_ASAP7_75t_SL g672 ( .A1(n_625), .A2(n_574), .B1(n_427), .B2(n_454), .Y(n_672) );
AOI21xp33_ASAP7_75t_L g673 ( .A1(n_589), .A2(n_450), .B(n_561), .Y(n_673) );
INVxp67_ASAP7_75t_L g674 ( .A(n_589), .Y(n_674) );
XOR2xp5_ASAP7_75t_L g675 ( .A(n_606), .B(n_213), .Y(n_675) );
OAI221xp5_ASAP7_75t_SL g676 ( .A1(n_674), .A2(n_630), .B1(n_650), .B2(n_639), .C(n_632), .Y(n_676) );
AOI211xp5_ASAP7_75t_L g677 ( .A1(n_673), .A2(n_674), .B(n_661), .C(n_667), .Y(n_677) );
OAI32xp33_ASAP7_75t_L g678 ( .A1(n_669), .A2(n_645), .A3(n_673), .B1(n_640), .B2(n_648), .Y(n_678) );
INVx2_ASAP7_75t_SL g679 ( .A(n_645), .Y(n_679) );
INVx1_ASAP7_75t_SL g680 ( .A(n_635), .Y(n_680) );
INVxp33_ASAP7_75t_SL g681 ( .A(n_672), .Y(n_681) );
CKINVDCx20_ASAP7_75t_L g682 ( .A(n_666), .Y(n_682) );
O2A1O1Ixp33_ASAP7_75t_SL g683 ( .A1(n_639), .A2(n_649), .B(n_634), .C(n_657), .Y(n_683) );
INVx1_ASAP7_75t_L g684 ( .A(n_642), .Y(n_684) );
AOI21xp5_ASAP7_75t_L g685 ( .A1(n_659), .A2(n_634), .B(n_649), .Y(n_685) );
INVx2_ASAP7_75t_SL g686 ( .A(n_647), .Y(n_686) );
AOI22x1_ASAP7_75t_L g687 ( .A1(n_675), .A2(n_670), .B1(n_633), .B2(n_648), .Y(n_687) );
INVx1_ASAP7_75t_L g688 ( .A(n_646), .Y(n_688) );
INVx2_ASAP7_75t_L g689 ( .A(n_658), .Y(n_689) );
AND2x2_ASAP7_75t_L g690 ( .A(n_653), .B(n_651), .Y(n_690) );
AND2x2_ASAP7_75t_L g691 ( .A(n_686), .B(n_631), .Y(n_691) );
NAND2xp5_ASAP7_75t_SL g692 ( .A(n_685), .B(n_644), .Y(n_692) );
XNOR2xp5_ASAP7_75t_L g693 ( .A(n_687), .B(n_664), .Y(n_693) );
OA22x2_ASAP7_75t_L g694 ( .A1(n_680), .A2(n_641), .B1(n_631), .B2(n_652), .Y(n_694) );
INVx1_ASAP7_75t_SL g695 ( .A(n_679), .Y(n_695) );
O2A1O1Ixp33_ASAP7_75t_L g696 ( .A1(n_681), .A2(n_654), .B(n_663), .C(n_671), .Y(n_696) );
AOI22xp5_ASAP7_75t_L g697 ( .A1(n_681), .A2(n_660), .B1(n_655), .B2(n_656), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_679), .B(n_643), .Y(n_698) );
OAI211xp5_ASAP7_75t_SL g699 ( .A1(n_677), .A2(n_662), .B(n_668), .C(n_629), .Y(n_699) );
OAI211xp5_ASAP7_75t_SL g700 ( .A1(n_692), .A2(n_683), .B(n_682), .C(n_686), .Y(n_700) );
OAI21xp5_ASAP7_75t_L g701 ( .A1(n_693), .A2(n_676), .B(n_687), .Y(n_701) );
NOR3xp33_ASAP7_75t_L g702 ( .A(n_699), .B(n_678), .C(n_682), .Y(n_702) );
OAI21xp5_ASAP7_75t_L g703 ( .A1(n_696), .A2(n_688), .B(n_684), .Y(n_703) );
AOI221xp5_ASAP7_75t_L g704 ( .A1(n_695), .A2(n_690), .B1(n_689), .B2(n_636), .C(n_638), .Y(n_704) );
NOR2x1p5_ASAP7_75t_L g705 ( .A(n_700), .B(n_637), .Y(n_705) );
INVxp67_ASAP7_75t_L g706 ( .A(n_701), .Y(n_706) );
AOI22xp5_ASAP7_75t_SL g707 ( .A1(n_703), .A2(n_694), .B1(n_695), .B2(n_691), .Y(n_707) );
OAI22xp5_ASAP7_75t_L g708 ( .A1(n_705), .A2(n_702), .B1(n_697), .B2(n_704), .Y(n_708) );
AO22x2_ASAP7_75t_L g709 ( .A1(n_706), .A2(n_698), .B1(n_665), .B2(n_689), .Y(n_709) );
INVx1_ASAP7_75t_L g710 ( .A(n_709), .Y(n_710) );
INVx1_ASAP7_75t_L g711 ( .A(n_708), .Y(n_711) );
INVxp67_ASAP7_75t_L g712 ( .A(n_710), .Y(n_712) );
INVx1_ASAP7_75t_L g713 ( .A(n_712), .Y(n_713) );
AOI21xp5_ASAP7_75t_L g714 ( .A1(n_713), .A2(n_711), .B(n_707), .Y(n_714) );
endmodule