module real_jpeg_11430_n_9 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_9);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;

output n_9;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_10;
wire n_114;
wire n_68;
wire n_78;
wire n_83;
wire n_104;
wire n_64;
wire n_11;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_13;
wire n_113;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_94;
wire n_26;
wire n_19;
wire n_17;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_103;
wire n_57;
wire n_43;
wire n_84;
wire n_82;
wire n_111;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_0),
.Y(n_53)
);

BUFx4f_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

AOI22xp33_ASAP7_75t_SL g21 ( 
.A1(n_3),
.A2(n_22),
.B1(n_23),
.B2(n_25),
.Y(n_21)
);

CKINVDCx14_ASAP7_75t_R g25 ( 
.A(n_3),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_3),
.A2(n_17),
.B1(n_18),
.B2(n_25),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_3),
.A2(n_25),
.B1(n_35),
.B2(n_36),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx12_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx2_ASAP7_75t_L g65 ( 
.A(n_6),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g27 ( 
.A1(n_7),
.A2(n_22),
.B1(n_23),
.B2(n_28),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_7),
.A2(n_17),
.B1(n_18),
.B2(n_28),
.Y(n_43)
);

O2A1O1Ixp33_ASAP7_75t_L g48 ( 
.A1(n_7),
.A2(n_19),
.B(n_22),
.C(n_49),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_7),
.A2(n_28),
.B1(n_35),
.B2(n_36),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_7),
.B(n_63),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_7),
.B(n_34),
.C(n_36),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_7),
.B(n_74),
.Y(n_90)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

XNOR2xp5_ASAP7_75t_L g9 ( 
.A(n_10),
.B(n_82),
.Y(n_9)
);

NAND2xp5_ASAP7_75t_SL g10 ( 
.A(n_11),
.B(n_81),
.Y(n_10)
);

INVxp67_ASAP7_75t_L g11 ( 
.A(n_12),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_57),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_13),
.B(n_57),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_31),
.C(n_46),
.Y(n_13)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_14),
.A2(n_15),
.B1(n_31),
.B2(n_99),
.Y(n_113)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

OAI21xp5_ASAP7_75t_L g15 ( 
.A1(n_16),
.A2(n_21),
.B(n_26),
.Y(n_15)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_16),
.B(n_30),
.Y(n_29)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_16),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_SL g16 ( 
.A1(n_17),
.A2(n_18),
.B1(n_19),
.B2(n_20),
.Y(n_16)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_17),
.A2(n_18),
.B1(n_34),
.B2(n_39),
.Y(n_45)
);

OAI21xp33_ASAP7_75t_L g49 ( 
.A1(n_17),
.A2(n_20),
.B(n_28),
.Y(n_49)
);

INVx4_ASAP7_75t_SL g17 ( 
.A(n_18),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_18),
.B(n_87),
.Y(n_86)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_19),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_19),
.A2(n_20),
.B1(n_22),
.B2(n_23),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_21),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_22),
.A2(n_23),
.B1(n_65),
.B2(n_66),
.Y(n_64)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_29),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_27),
.A2(n_29),
.B1(n_73),
.B2(n_74),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_28),
.B(n_56),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_28),
.B(n_32),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_31),
.B(n_86),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_31),
.A2(n_86),
.B1(n_98),
.B2(n_99),
.Y(n_97)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_31),
.Y(n_99)
);

OA21x2_ASAP7_75t_L g31 ( 
.A1(n_32),
.A2(n_40),
.B(n_42),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

NOR2x1_ASAP7_75t_L g44 ( 
.A(n_33),
.B(n_45),
.Y(n_44)
);

AO22x1_ASAP7_75t_SL g78 ( 
.A1(n_33),
.A2(n_41),
.B1(n_43),
.B2(n_44),
.Y(n_78)
);

AO22x1_ASAP7_75t_L g33 ( 
.A1(n_34),
.A2(n_35),
.B1(n_36),
.B2(n_39),
.Y(n_33)
);

INVx13_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_35),
.B(n_103),
.Y(n_102)
);

INVx3_ASAP7_75t_SL g35 ( 
.A(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_36),
.B(n_56),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_44),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_46),
.A2(n_47),
.B1(n_112),
.B2(n_113),
.Y(n_111)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

XOR2xp5_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_50),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_48),
.B(n_50),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_52),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_51),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_51),
.A2(n_55),
.B1(n_56),
.B2(n_69),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_54),
.Y(n_52)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_53),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_54),
.B(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_L g68 ( 
.A1(n_56),
.A2(n_69),
.B(n_70),
.Y(n_68)
);

XOR2xp5_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_76),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_59),
.A2(n_60),
.B1(n_72),
.B2(n_75),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_62),
.B1(n_67),
.B2(n_68),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_65),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_67),
.B(n_97),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_67),
.B(n_97),
.Y(n_107)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_68),
.B(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_72),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_77),
.A2(n_78),
.B1(n_79),
.B2(n_80),
.Y(n_76)
);

CKINVDCx14_ASAP7_75t_R g79 ( 
.A(n_77),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_78),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_78),
.A2(n_80),
.B1(n_90),
.B2(n_91),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_78),
.B(n_91),
.C(n_93),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_109),
.B(n_114),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_95),
.B(n_108),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_88),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_85),
.B(n_88),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_86),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_89),
.A2(n_92),
.B1(n_93),
.B2(n_94),
.Y(n_88)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_89),
.Y(n_94)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_90),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_93),
.B(n_105),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_93),
.B(n_105),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_100),
.B(n_107),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_101),
.A2(n_104),
.B(n_106),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_111),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_110),
.B(n_111),
.Y(n_114)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);


endmodule