module fake_ariane_2293_n_2045 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_195, n_38, n_47, n_110, n_153, n_18, n_197, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_198, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_194, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_2045);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_195;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_198;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_194;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_2045;

wire n_913;
wire n_1681;
wire n_1507;
wire n_1486;
wire n_1938;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_2002;
wire n_1463;
wire n_1238;
wire n_2011;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_2013;
wire n_1566;
wire n_717;
wire n_2006;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_214;
wire n_2042;
wire n_1853;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_1985;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1909;
wire n_1184;
wire n_1961;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1979;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_1944;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_1988;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_1977;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_1850;
wire n_238;
wire n_365;
wire n_2004;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_1917;
wire n_1924;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_2043;
wire n_780;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_225;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_2038;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_851;
wire n_212;
wire n_355;
wire n_444;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_2015;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_1880;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1970;
wire n_1920;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1911;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_1914;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_2019;
wire n_698;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_1992;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_1913;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_2041;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_552;
wire n_348;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1951;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_1943;
wire n_1802;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_1868;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_1901;
wire n_647;
wire n_2027;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_1939;
wire n_1906;
wire n_529;
wire n_1899;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_677;
wire n_604;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_2023;
wire n_1278;
wire n_707;
wire n_983;
wire n_699;
wire n_590;
wire n_727;
wire n_301;
wire n_1726;
wire n_1945;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_2031;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_1963;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_2033;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_1883;
wire n_1969;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_888;
wire n_845;
wire n_1649;
wire n_1677;
wire n_1927;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_1957;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_534;
wire n_1791;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_2008;
wire n_454;
wire n_298;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1966;
wire n_1243;
wire n_1400;
wire n_342;
wire n_2035;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1993;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1897;
wire n_1161;
wire n_811;
wire n_624;
wire n_876;
wire n_791;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_2026;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_1929;
wire n_1950;
wire n_805;
wire n_2032;
wire n_295;
wire n_1658;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1997;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_463;
wire n_1524;
wire n_1476;
wire n_1733;
wire n_1856;
wire n_2016;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_1971;
wire n_586;
wire n_1324;
wire n_1429;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_2022;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_2001;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_2044;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_2020;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_1881;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_1958;
wire n_467;
wire n_1511;
wire n_1422;
wire n_1965;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_2036;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_2003;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1955;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_1960;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_1978;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_526;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_1986;
wire n_540;
wire n_216;
wire n_692;
wire n_1857;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_2018;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_493;
wire n_1311;
wire n_1956;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_2014;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_508;
wire n_1679;
wire n_1952;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_1980;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_1998;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_2028;
wire n_919;
wire n_1663;
wire n_1625;
wire n_1926;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1904;
wire n_2000;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_898;
wire n_857;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1937;
wire n_2012;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_761;
wire n_733;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_1865;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_1792;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1727;
wire n_1991;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_2034;
wire n_1845;
wire n_1934;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_2005;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_1866;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_1964;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_1982;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_1946;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_1732;
wire n_415;
wire n_1967;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_1126;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_1102;
wire n_719;
wire n_263;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1905;
wire n_1569;
wire n_548;
wire n_289;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_1925;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_1228;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_411;
wire n_484;
wire n_849;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_1989;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2037;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_184),
.Y(n_199)
);

BUFx3_ASAP7_75t_L g200 ( 
.A(n_143),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_182),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_80),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_30),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_74),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_102),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_57),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_31),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_123),
.Y(n_208)
);

BUFx8_ASAP7_75t_SL g209 ( 
.A(n_167),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_89),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_18),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_31),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_139),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_154),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_36),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_186),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_73),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_49),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_101),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_161),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_87),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_47),
.Y(n_222)
);

BUFx3_ASAP7_75t_L g223 ( 
.A(n_162),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_16),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_77),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_64),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_97),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_153),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_152),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_50),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_73),
.Y(n_231)
);

BUFx3_ASAP7_75t_L g232 ( 
.A(n_2),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_15),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_18),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_9),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_35),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_138),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_49),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_44),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_128),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_45),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_107),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_27),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_190),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_100),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_36),
.Y(n_246)
);

BUFx3_ASAP7_75t_L g247 ( 
.A(n_98),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_157),
.Y(n_248)
);

BUFx8_ASAP7_75t_SL g249 ( 
.A(n_195),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_115),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_20),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_60),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_172),
.Y(n_253)
);

BUFx8_ASAP7_75t_SL g254 ( 
.A(n_151),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_196),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_176),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_30),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_173),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_112),
.Y(n_259)
);

BUFx5_ASAP7_75t_L g260 ( 
.A(n_12),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_75),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_26),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_91),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_159),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_133),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_44),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_53),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_12),
.Y(n_268)
);

BUFx10_ASAP7_75t_L g269 ( 
.A(n_13),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_171),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_179),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_7),
.Y(n_272)
);

INVx1_ASAP7_75t_SL g273 ( 
.A(n_28),
.Y(n_273)
);

CKINVDCx16_ASAP7_75t_R g274 ( 
.A(n_116),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_170),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_38),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_189),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_22),
.Y(n_278)
);

HB1xp67_ASAP7_75t_L g279 ( 
.A(n_109),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_95),
.Y(n_280)
);

BUFx6f_ASAP7_75t_L g281 ( 
.A(n_32),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_66),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_110),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_15),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_50),
.Y(n_285)
);

CKINVDCx14_ASAP7_75t_R g286 ( 
.A(n_32),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_177),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_96),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_137),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_57),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_38),
.Y(n_291)
);

BUFx10_ASAP7_75t_L g292 ( 
.A(n_59),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_84),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_194),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_13),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_4),
.Y(n_296)
);

INVxp33_ASAP7_75t_L g297 ( 
.A(n_85),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_60),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_6),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_175),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_99),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_20),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_16),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_136),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_27),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_26),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_8),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_46),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_191),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_24),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_78),
.Y(n_311)
);

BUFx6f_ASAP7_75t_L g312 ( 
.A(n_19),
.Y(n_312)
);

HB1xp67_ASAP7_75t_L g313 ( 
.A(n_193),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_163),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_3),
.Y(n_315)
);

INVx1_ASAP7_75t_SL g316 ( 
.A(n_120),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_144),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_3),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_74),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_34),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_125),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_39),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_37),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_147),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_59),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_168),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_83),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_141),
.Y(n_328)
);

INVx1_ASAP7_75t_SL g329 ( 
.A(n_127),
.Y(n_329)
);

BUFx6f_ASAP7_75t_L g330 ( 
.A(n_180),
.Y(n_330)
);

HB1xp67_ASAP7_75t_SL g331 ( 
.A(n_134),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_197),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_68),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_183),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_29),
.Y(n_335)
);

BUFx3_ASAP7_75t_L g336 ( 
.A(n_140),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_42),
.Y(n_337)
);

CKINVDCx16_ASAP7_75t_R g338 ( 
.A(n_124),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_119),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_43),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_158),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_63),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_126),
.Y(n_343)
);

INVx1_ASAP7_75t_SL g344 ( 
.A(n_43),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_29),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_72),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_24),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_90),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_25),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_113),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_63),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_129),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_40),
.Y(n_353)
);

BUFx2_ASAP7_75t_L g354 ( 
.A(n_35),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_121),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_28),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_130),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_132),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_69),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_88),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_41),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_33),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_174),
.Y(n_363)
);

INVx1_ASAP7_75t_SL g364 ( 
.A(n_25),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_55),
.Y(n_365)
);

BUFx5_ASAP7_75t_L g366 ( 
.A(n_169),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_51),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_146),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_148),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_46),
.Y(n_370)
);

BUFx6f_ASAP7_75t_L g371 ( 
.A(n_156),
.Y(n_371)
);

BUFx10_ASAP7_75t_L g372 ( 
.A(n_53),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_69),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_75),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_86),
.Y(n_375)
);

BUFx3_ASAP7_75t_L g376 ( 
.A(n_187),
.Y(n_376)
);

HB1xp67_ASAP7_75t_L g377 ( 
.A(n_58),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_68),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_1),
.Y(n_379)
);

INVxp67_ASAP7_75t_L g380 ( 
.A(n_72),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_70),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_5),
.Y(n_382)
);

INVx2_ASAP7_75t_SL g383 ( 
.A(n_142),
.Y(n_383)
);

INVx2_ASAP7_75t_SL g384 ( 
.A(n_2),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_39),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_108),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_62),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_103),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_79),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_64),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_58),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_81),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_1),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_56),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_33),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_0),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_260),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_260),
.Y(n_398)
);

HB1xp67_ASAP7_75t_L g399 ( 
.A(n_354),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_260),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_209),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_286),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_260),
.Y(n_403)
);

INVxp67_ASAP7_75t_L g404 ( 
.A(n_354),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_260),
.Y(n_405)
);

INVxp67_ASAP7_75t_L g406 ( 
.A(n_377),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_260),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_208),
.Y(n_408)
);

CKINVDCx16_ASAP7_75t_R g409 ( 
.A(n_216),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_260),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_260),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_277),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_201),
.Y(n_413)
);

HB1xp67_ASAP7_75t_L g414 ( 
.A(n_232),
.Y(n_414)
);

INVxp67_ASAP7_75t_L g415 ( 
.A(n_204),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_300),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_201),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_363),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_214),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_249),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_214),
.Y(n_421)
);

INVxp67_ASAP7_75t_SL g422 ( 
.A(n_232),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_254),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_375),
.Y(n_424)
);

INVxp33_ASAP7_75t_SL g425 ( 
.A(n_206),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_219),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_279),
.B(n_0),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_207),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_219),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_217),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_220),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_222),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_204),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_396),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_226),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_224),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_230),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_220),
.B(n_4),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_225),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_225),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_228),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_228),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_240),
.Y(n_443)
);

INVxp33_ASAP7_75t_L g444 ( 
.A(n_211),
.Y(n_444)
);

CKINVDCx16_ASAP7_75t_R g445 ( 
.A(n_274),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_231),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_240),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_242),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_234),
.Y(n_449)
);

HB1xp67_ASAP7_75t_L g450 ( 
.A(n_236),
.Y(n_450)
);

CKINVDCx20_ASAP7_75t_R g451 ( 
.A(n_239),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_238),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_242),
.Y(n_453)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_267),
.Y(n_454)
);

CKINVDCx14_ASAP7_75t_R g455 ( 
.A(n_269),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_284),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_244),
.Y(n_457)
);

HB1xp67_ASAP7_75t_L g458 ( 
.A(n_243),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_246),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_262),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_244),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_281),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_250),
.Y(n_463)
);

HB1xp67_ASAP7_75t_L g464 ( 
.A(n_276),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_278),
.Y(n_465)
);

NOR2xp67_ASAP7_75t_L g466 ( 
.A(n_384),
.B(n_5),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_250),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_296),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_264),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_282),
.Y(n_470)
);

BUFx6f_ASAP7_75t_SL g471 ( 
.A(n_200),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_285),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g473 ( 
.A(n_308),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_264),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_290),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_275),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_275),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_291),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_287),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_333),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_295),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_302),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_287),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_303),
.Y(n_484)
);

CKINVDCx20_ASAP7_75t_R g485 ( 
.A(n_385),
.Y(n_485)
);

CKINVDCx20_ASAP7_75t_R g486 ( 
.A(n_387),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_293),
.B(n_6),
.Y(n_487)
);

CKINVDCx20_ASAP7_75t_R g488 ( 
.A(n_338),
.Y(n_488)
);

CKINVDCx20_ASAP7_75t_R g489 ( 
.A(n_200),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_293),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_334),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_305),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_306),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_307),
.Y(n_494)
);

OR2x2_ASAP7_75t_L g495 ( 
.A(n_203),
.B(n_266),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_315),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_334),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_341),
.Y(n_498)
);

INVxp67_ASAP7_75t_L g499 ( 
.A(n_211),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_397),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_397),
.Y(n_501)
);

BUFx2_ASAP7_75t_L g502 ( 
.A(n_488),
.Y(n_502)
);

INVx3_ASAP7_75t_L g503 ( 
.A(n_407),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_398),
.Y(n_504)
);

BUFx6f_ASAP7_75t_L g505 ( 
.A(n_407),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_413),
.B(n_313),
.Y(n_506)
);

AND2x4_ASAP7_75t_L g507 ( 
.A(n_413),
.B(n_384),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_462),
.Y(n_508)
);

BUFx6f_ASAP7_75t_L g509 ( 
.A(n_398),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_422),
.B(n_425),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_462),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_400),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_400),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_403),
.Y(n_514)
);

OR2x6_ASAP7_75t_L g515 ( 
.A(n_427),
.B(n_203),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_403),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_405),
.Y(n_517)
);

AND2x4_ASAP7_75t_L g518 ( 
.A(n_417),
.B(n_266),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_405),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_410),
.Y(n_520)
);

BUFx6f_ASAP7_75t_L g521 ( 
.A(n_410),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_411),
.Y(n_522)
);

AND2x2_ASAP7_75t_L g523 ( 
.A(n_417),
.B(n_298),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_411),
.Y(n_524)
);

INVx6_ASAP7_75t_L g525 ( 
.A(n_495),
.Y(n_525)
);

BUFx8_ASAP7_75t_L g526 ( 
.A(n_471),
.Y(n_526)
);

AOI22xp5_ASAP7_75t_L g527 ( 
.A1(n_404),
.A2(n_406),
.B1(n_399),
.B2(n_402),
.Y(n_527)
);

AND2x2_ASAP7_75t_L g528 ( 
.A(n_419),
.B(n_298),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_450),
.B(n_297),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_419),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_421),
.Y(n_531)
);

INVxp67_ASAP7_75t_L g532 ( 
.A(n_458),
.Y(n_532)
);

INVx3_ASAP7_75t_L g533 ( 
.A(n_421),
.Y(n_533)
);

OA21x2_ASAP7_75t_L g534 ( 
.A1(n_426),
.A2(n_350),
.B(n_341),
.Y(n_534)
);

BUFx6f_ASAP7_75t_L g535 ( 
.A(n_426),
.Y(n_535)
);

XOR2xp5_ASAP7_75t_L g536 ( 
.A(n_436),
.B(n_320),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_429),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_429),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_SL g539 ( 
.A(n_409),
.B(n_269),
.Y(n_539)
);

BUFx2_ASAP7_75t_L g540 ( 
.A(n_428),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_431),
.Y(n_541)
);

INVx3_ASAP7_75t_L g542 ( 
.A(n_431),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_439),
.B(n_440),
.Y(n_543)
);

HB1xp67_ASAP7_75t_L g544 ( 
.A(n_414),
.Y(n_544)
);

HB1xp67_ASAP7_75t_L g545 ( 
.A(n_430),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_439),
.Y(n_546)
);

INVx2_ASAP7_75t_SL g547 ( 
.A(n_440),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_441),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_424),
.Y(n_549)
);

AND2x2_ASAP7_75t_L g550 ( 
.A(n_441),
.B(n_335),
.Y(n_550)
);

BUFx2_ASAP7_75t_L g551 ( 
.A(n_432),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_442),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_442),
.Y(n_553)
);

AND2x4_ASAP7_75t_L g554 ( 
.A(n_443),
.B(n_335),
.Y(n_554)
);

BUFx2_ASAP7_75t_L g555 ( 
.A(n_435),
.Y(n_555)
);

AND2x4_ASAP7_75t_L g556 ( 
.A(n_443),
.B(n_281),
.Y(n_556)
);

INVx3_ASAP7_75t_L g557 ( 
.A(n_447),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_447),
.B(n_448),
.Y(n_558)
);

BUFx6f_ASAP7_75t_L g559 ( 
.A(n_448),
.Y(n_559)
);

NAND2x1p5_ASAP7_75t_L g560 ( 
.A(n_453),
.B(n_223),
.Y(n_560)
);

NAND3xp33_ASAP7_75t_L g561 ( 
.A(n_438),
.B(n_215),
.C(n_212),
.Y(n_561)
);

BUFx2_ASAP7_75t_L g562 ( 
.A(n_446),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_453),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_457),
.Y(n_564)
);

BUFx6f_ASAP7_75t_L g565 ( 
.A(n_457),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_SL g566 ( 
.A(n_445),
.B(n_383),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_461),
.B(n_350),
.Y(n_567)
);

INVxp67_ASAP7_75t_L g568 ( 
.A(n_464),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_SL g569 ( 
.A(n_449),
.B(n_383),
.Y(n_569)
);

BUFx6f_ASAP7_75t_L g570 ( 
.A(n_461),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_463),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_463),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_467),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_467),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_L g575 ( 
.A(n_452),
.B(n_352),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_469),
.B(n_474),
.Y(n_576)
);

INVx6_ASAP7_75t_L g577 ( 
.A(n_495),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_469),
.B(n_352),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_474),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_SL g580 ( 
.A(n_510),
.B(n_459),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_SL g581 ( 
.A(n_510),
.B(n_460),
.Y(n_581)
);

OR2x6_ASAP7_75t_L g582 ( 
.A(n_515),
.B(n_466),
.Y(n_582)
);

BUFx6f_ASAP7_75t_SL g583 ( 
.A(n_515),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_514),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_SL g585 ( 
.A(n_575),
.B(n_465),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_535),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_535),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_514),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_514),
.Y(n_589)
);

NOR2xp33_ASAP7_75t_L g590 ( 
.A(n_525),
.B(n_455),
.Y(n_590)
);

BUFx3_ASAP7_75t_L g591 ( 
.A(n_526),
.Y(n_591)
);

BUFx3_ASAP7_75t_L g592 ( 
.A(n_526),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_535),
.Y(n_593)
);

NOR2xp33_ASAP7_75t_L g594 ( 
.A(n_525),
.B(n_470),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_SL g595 ( 
.A(n_529),
.B(n_472),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_547),
.B(n_476),
.Y(n_596)
);

AND2x2_ASAP7_75t_SL g597 ( 
.A(n_534),
.B(n_202),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_535),
.Y(n_598)
);

OR2x2_ASAP7_75t_L g599 ( 
.A(n_544),
.B(n_475),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_535),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_519),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_535),
.Y(n_602)
);

INVxp67_ASAP7_75t_SL g603 ( 
.A(n_543),
.Y(n_603)
);

BUFx4f_ASAP7_75t_L g604 ( 
.A(n_535),
.Y(n_604)
);

OR2x6_ASAP7_75t_L g605 ( 
.A(n_515),
.B(n_476),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_559),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_L g607 ( 
.A(n_525),
.B(n_478),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_559),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_SL g609 ( 
.A(n_529),
.B(n_481),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_547),
.B(n_477),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_519),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_559),
.Y(n_612)
);

BUFx3_ASAP7_75t_L g613 ( 
.A(n_526),
.Y(n_613)
);

BUFx6f_ASAP7_75t_L g614 ( 
.A(n_505),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_SL g615 ( 
.A(n_540),
.B(n_482),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_SL g616 ( 
.A(n_540),
.B(n_484),
.Y(n_616)
);

NAND3xp33_ASAP7_75t_L g617 ( 
.A(n_561),
.B(n_493),
.C(n_492),
.Y(n_617)
);

INVx3_ASAP7_75t_L g618 ( 
.A(n_559),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_559),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_559),
.Y(n_620)
);

OA22x2_ASAP7_75t_L g621 ( 
.A1(n_515),
.A2(n_499),
.B1(n_415),
.B2(n_479),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_SL g622 ( 
.A(n_551),
.B(n_494),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_547),
.B(n_477),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_519),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_559),
.Y(n_625)
);

AOI22xp33_ASAP7_75t_L g626 ( 
.A1(n_561),
.A2(n_487),
.B1(n_444),
.B2(n_483),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_533),
.B(n_479),
.Y(n_627)
);

AND2x2_ASAP7_75t_L g628 ( 
.A(n_523),
.B(n_528),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_524),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_524),
.Y(n_630)
);

CKINVDCx16_ASAP7_75t_R g631 ( 
.A(n_539),
.Y(n_631)
);

NAND3xp33_ASAP7_75t_L g632 ( 
.A(n_532),
.B(n_496),
.C(n_490),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_533),
.B(n_483),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_524),
.Y(n_634)
);

BUFx8_ASAP7_75t_SL g635 ( 
.A(n_549),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_565),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_565),
.Y(n_637)
);

AND2x2_ASAP7_75t_L g638 ( 
.A(n_523),
.B(n_528),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_503),
.Y(n_639)
);

CKINVDCx20_ASAP7_75t_R g640 ( 
.A(n_551),
.Y(n_640)
);

BUFx6f_ASAP7_75t_L g641 ( 
.A(n_505),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_503),
.Y(n_642)
);

INVx4_ASAP7_75t_L g643 ( 
.A(n_533),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_503),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_565),
.Y(n_645)
);

INVxp67_ASAP7_75t_SL g646 ( 
.A(n_543),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_503),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_565),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_509),
.Y(n_649)
);

NAND2xp33_ASAP7_75t_L g650 ( 
.A(n_545),
.B(n_565),
.Y(n_650)
);

AOI22xp5_ASAP7_75t_L g651 ( 
.A1(n_515),
.A2(n_273),
.B1(n_364),
.B2(n_344),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_509),
.Y(n_652)
);

INVx4_ASAP7_75t_L g653 ( 
.A(n_533),
.Y(n_653)
);

BUFx3_ASAP7_75t_L g654 ( 
.A(n_526),
.Y(n_654)
);

NOR2xp33_ASAP7_75t_L g655 ( 
.A(n_525),
.B(n_489),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_542),
.B(n_490),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_565),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_509),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_565),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_SL g660 ( 
.A(n_555),
.B(n_401),
.Y(n_660)
);

INVx4_ASAP7_75t_L g661 ( 
.A(n_542),
.Y(n_661)
);

INVx4_ASAP7_75t_L g662 ( 
.A(n_542),
.Y(n_662)
);

AOI22xp5_ASAP7_75t_L g663 ( 
.A1(n_515),
.A2(n_380),
.B1(n_337),
.B2(n_340),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_570),
.Y(n_664)
);

AND2x4_ASAP7_75t_L g665 ( 
.A(n_507),
.B(n_491),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_570),
.Y(n_666)
);

NAND2xp33_ASAP7_75t_L g667 ( 
.A(n_545),
.B(n_281),
.Y(n_667)
);

INVx3_ASAP7_75t_L g668 ( 
.A(n_570),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_542),
.B(n_491),
.Y(n_669)
);

AOI22xp33_ASAP7_75t_L g670 ( 
.A1(n_525),
.A2(n_498),
.B1(n_497),
.B2(n_471),
.Y(n_670)
);

OR2x6_ASAP7_75t_L g671 ( 
.A(n_560),
.B(n_497),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_557),
.B(n_498),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_526),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_SL g674 ( 
.A(n_555),
.B(n_420),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_557),
.B(n_433),
.Y(n_675)
);

INVx3_ASAP7_75t_L g676 ( 
.A(n_570),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_557),
.B(n_434),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_557),
.B(n_316),
.Y(n_678)
);

AND2x2_ASAP7_75t_L g679 ( 
.A(n_523),
.B(n_269),
.Y(n_679)
);

NOR2xp33_ASAP7_75t_L g680 ( 
.A(n_577),
.B(n_471),
.Y(n_680)
);

OR2x2_ASAP7_75t_L g681 ( 
.A(n_544),
.B(n_423),
.Y(n_681)
);

BUFx6f_ASAP7_75t_L g682 ( 
.A(n_505),
.Y(n_682)
);

INVx4_ASAP7_75t_L g683 ( 
.A(n_570),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_509),
.Y(n_684)
);

BUFx6f_ASAP7_75t_L g685 ( 
.A(n_505),
.Y(n_685)
);

INVx3_ASAP7_75t_L g686 ( 
.A(n_570),
.Y(n_686)
);

AND2x2_ASAP7_75t_L g687 ( 
.A(n_528),
.B(n_292),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_570),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_577),
.B(n_329),
.Y(n_689)
);

INVx5_ASAP7_75t_L g690 ( 
.A(n_509),
.Y(n_690)
);

BUFx2_ASAP7_75t_L g691 ( 
.A(n_562),
.Y(n_691)
);

BUFx8_ASAP7_75t_SL g692 ( 
.A(n_502),
.Y(n_692)
);

AND2x2_ASAP7_75t_L g693 ( 
.A(n_550),
.B(n_292),
.Y(n_693)
);

AOI22xp33_ASAP7_75t_L g694 ( 
.A1(n_577),
.A2(n_268),
.B1(n_212),
.B2(n_310),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_537),
.Y(n_695)
);

BUFx6f_ASAP7_75t_L g696 ( 
.A(n_505),
.Y(n_696)
);

CKINVDCx20_ASAP7_75t_R g697 ( 
.A(n_562),
.Y(n_697)
);

INVx2_ASAP7_75t_SL g698 ( 
.A(n_577),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_537),
.Y(n_699)
);

INVx3_ASAP7_75t_L g700 ( 
.A(n_509),
.Y(n_700)
);

NAND2xp33_ASAP7_75t_L g701 ( 
.A(n_558),
.B(n_281),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_577),
.B(n_357),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_537),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_509),
.Y(n_704)
);

OAI22xp5_ASAP7_75t_L g705 ( 
.A1(n_532),
.A2(n_345),
.B1(n_346),
.B2(n_351),
.Y(n_705)
);

BUFx6f_ASAP7_75t_L g706 ( 
.A(n_505),
.Y(n_706)
);

BUFx6f_ASAP7_75t_L g707 ( 
.A(n_505),
.Y(n_707)
);

INVx3_ASAP7_75t_L g708 ( 
.A(n_521),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_530),
.B(n_357),
.Y(n_709)
);

INVx2_ASAP7_75t_SL g710 ( 
.A(n_560),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_548),
.Y(n_711)
);

OR2x2_ASAP7_75t_L g712 ( 
.A(n_527),
.B(n_215),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_548),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_SL g714 ( 
.A(n_568),
.B(n_322),
.Y(n_714)
);

AND2x2_ASAP7_75t_SL g715 ( 
.A(n_534),
.B(n_202),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_521),
.Y(n_716)
);

AND2x2_ASAP7_75t_SL g717 ( 
.A(n_534),
.B(n_263),
.Y(n_717)
);

INVx4_ASAP7_75t_L g718 ( 
.A(n_521),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_530),
.B(n_360),
.Y(n_719)
);

BUFx2_ASAP7_75t_L g720 ( 
.A(n_568),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_548),
.Y(n_721)
);

INVx2_ASAP7_75t_SL g722 ( 
.A(n_560),
.Y(n_722)
);

AND2x2_ASAP7_75t_L g723 ( 
.A(n_550),
.B(n_292),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_502),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_536),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_521),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_552),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_552),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_552),
.Y(n_729)
);

BUFx4f_ASAP7_75t_L g730 ( 
.A(n_534),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_563),
.Y(n_731)
);

AOI22xp33_ASAP7_75t_L g732 ( 
.A1(n_507),
.A2(n_560),
.B1(n_534),
.B2(n_506),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_603),
.B(n_531),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_646),
.B(n_531),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_594),
.B(n_538),
.Y(n_735)
);

NOR3xp33_ASAP7_75t_L g736 ( 
.A(n_632),
.B(n_569),
.C(n_558),
.Y(n_736)
);

NOR2xp33_ASAP7_75t_L g737 ( 
.A(n_607),
.B(n_566),
.Y(n_737)
);

BUFx6f_ASAP7_75t_SL g738 ( 
.A(n_591),
.Y(n_738)
);

NOR2xp33_ASAP7_75t_L g739 ( 
.A(n_595),
.B(n_539),
.Y(n_739)
);

OR2x6_ASAP7_75t_L g740 ( 
.A(n_691),
.B(n_507),
.Y(n_740)
);

NOR3xp33_ASAP7_75t_L g741 ( 
.A(n_617),
.B(n_576),
.C(n_506),
.Y(n_741)
);

AOI22xp33_ASAP7_75t_L g742 ( 
.A1(n_597),
.A2(n_507),
.B1(n_554),
.B2(n_518),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_695),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_665),
.B(n_538),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_665),
.B(n_541),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_SL g746 ( 
.A(n_698),
.B(n_507),
.Y(n_746)
);

NOR2xp33_ASAP7_75t_L g747 ( 
.A(n_609),
.B(n_500),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_665),
.B(n_541),
.Y(n_748)
);

AO22x2_ASAP7_75t_L g749 ( 
.A1(n_712),
.A2(n_536),
.B1(n_233),
.B2(n_235),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_SL g750 ( 
.A(n_698),
.B(n_576),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_695),
.Y(n_751)
);

INVxp67_ASAP7_75t_SL g752 ( 
.A(n_730),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_584),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_SL g754 ( 
.A(n_720),
.B(n_546),
.Y(n_754)
);

AND2x2_ASAP7_75t_L g755 ( 
.A(n_720),
.B(n_691),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_665),
.B(n_546),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_699),
.Y(n_757)
);

O2A1O1Ixp33_ASAP7_75t_L g758 ( 
.A1(n_627),
.A2(n_501),
.B(n_504),
.C(n_500),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_SL g759 ( 
.A(n_643),
.B(n_653),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_590),
.B(n_553),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_584),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_689),
.B(n_553),
.Y(n_762)
);

INVx4_ASAP7_75t_L g763 ( 
.A(n_591),
.Y(n_763)
);

AND2x6_ASAP7_75t_L g764 ( 
.A(n_592),
.B(n_613),
.Y(n_764)
);

NOR2xp33_ASAP7_75t_L g765 ( 
.A(n_580),
.B(n_501),
.Y(n_765)
);

INVxp67_ASAP7_75t_L g766 ( 
.A(n_655),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_679),
.B(n_687),
.Y(n_767)
);

BUFx6f_ASAP7_75t_L g768 ( 
.A(n_614),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_703),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_679),
.B(n_572),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_588),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_SL g772 ( 
.A(n_663),
.B(n_572),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_687),
.B(n_573),
.Y(n_773)
);

AOI22xp5_ASAP7_75t_L g774 ( 
.A1(n_605),
.A2(n_574),
.B1(n_573),
.B2(n_564),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_SL g775 ( 
.A(n_663),
.B(n_574),
.Y(n_775)
);

OR2x2_ASAP7_75t_L g776 ( 
.A(n_599),
.B(n_527),
.Y(n_776)
);

BUFx6f_ASAP7_75t_L g777 ( 
.A(n_614),
.Y(n_777)
);

NAND2x1_ASAP7_75t_L g778 ( 
.A(n_643),
.B(n_563),
.Y(n_778)
);

NOR2xp33_ASAP7_75t_R g779 ( 
.A(n_673),
.B(n_408),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_SL g780 ( 
.A(n_599),
.B(n_567),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_SL g781 ( 
.A(n_693),
.B(n_567),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_693),
.B(n_563),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_703),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_711),
.Y(n_784)
);

NOR2xp33_ASAP7_75t_L g785 ( 
.A(n_581),
.B(n_504),
.Y(n_785)
);

NOR2xp33_ASAP7_75t_L g786 ( 
.A(n_585),
.B(n_512),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_SL g787 ( 
.A(n_643),
.B(n_512),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_723),
.B(n_564),
.Y(n_788)
);

BUFx6f_ASAP7_75t_L g789 ( 
.A(n_614),
.Y(n_789)
);

NOR2xp33_ASAP7_75t_L g790 ( 
.A(n_653),
.B(n_513),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_723),
.B(n_680),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_SL g792 ( 
.A(n_670),
.B(n_578),
.Y(n_792)
);

NAND2xp33_ASAP7_75t_L g793 ( 
.A(n_596),
.B(n_513),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_588),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_589),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_589),
.Y(n_796)
);

NAND2xp33_ASAP7_75t_L g797 ( 
.A(n_610),
.B(n_516),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_628),
.B(n_564),
.Y(n_798)
);

BUFx6f_ASAP7_75t_L g799 ( 
.A(n_614),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_713),
.Y(n_800)
);

BUFx12f_ASAP7_75t_L g801 ( 
.A(n_724),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_601),
.Y(n_802)
);

AOI22xp33_ASAP7_75t_L g803 ( 
.A1(n_597),
.A2(n_717),
.B1(n_715),
.B2(n_621),
.Y(n_803)
);

INVxp67_ASAP7_75t_L g804 ( 
.A(n_635),
.Y(n_804)
);

BUFx3_ASAP7_75t_L g805 ( 
.A(n_640),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_601),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_628),
.B(n_571),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_SL g808 ( 
.A(n_621),
.B(n_578),
.Y(n_808)
);

AND2x6_ASAP7_75t_L g809 ( 
.A(n_592),
.B(n_613),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_SL g810 ( 
.A(n_621),
.B(n_579),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_SL g811 ( 
.A(n_651),
.B(n_653),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_638),
.B(n_571),
.Y(n_812)
);

OR2x2_ASAP7_75t_L g813 ( 
.A(n_681),
.B(n_550),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_638),
.B(n_571),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_661),
.B(n_579),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_SL g816 ( 
.A(n_651),
.B(n_579),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_611),
.Y(n_817)
);

OR2x6_ASAP7_75t_L g818 ( 
.A(n_605),
.B(n_518),
.Y(n_818)
);

AO22x2_ASAP7_75t_L g819 ( 
.A1(n_712),
.A2(n_272),
.B1(n_218),
.B2(n_233),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_SL g820 ( 
.A(n_661),
.B(n_518),
.Y(n_820)
);

AND2x4_ASAP7_75t_SL g821 ( 
.A(n_697),
.B(n_412),
.Y(n_821)
);

NOR2xp33_ASAP7_75t_L g822 ( 
.A(n_661),
.B(n_516),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_SL g823 ( 
.A(n_662),
.B(n_517),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_662),
.B(n_517),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_713),
.Y(n_825)
);

INVx2_ASAP7_75t_L g826 ( 
.A(n_611),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_SL g827 ( 
.A(n_662),
.B(n_520),
.Y(n_827)
);

INVxp33_ASAP7_75t_L g828 ( 
.A(n_692),
.Y(n_828)
);

INVx2_ASAP7_75t_SL g829 ( 
.A(n_681),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_721),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_732),
.B(n_520),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_678),
.B(n_522),
.Y(n_832)
);

BUFx3_ASAP7_75t_L g833 ( 
.A(n_724),
.Y(n_833)
);

INVx2_ASAP7_75t_SL g834 ( 
.A(n_631),
.Y(n_834)
);

O2A1O1Ixp33_ASAP7_75t_L g835 ( 
.A1(n_633),
.A2(n_522),
.B(n_235),
.C(n_218),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_SL g836 ( 
.A(n_710),
.B(n_518),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_623),
.B(n_518),
.Y(n_837)
);

AND2x2_ASAP7_75t_L g838 ( 
.A(n_631),
.B(n_416),
.Y(n_838)
);

OAI22xp5_ASAP7_75t_L g839 ( 
.A1(n_605),
.A2(n_370),
.B1(n_353),
.B2(n_356),
.Y(n_839)
);

INVxp67_ASAP7_75t_SL g840 ( 
.A(n_730),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_702),
.B(n_554),
.Y(n_841)
);

NOR2xp33_ASAP7_75t_L g842 ( 
.A(n_714),
.B(n_521),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_721),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_727),
.Y(n_844)
);

AND2x2_ASAP7_75t_L g845 ( 
.A(n_626),
.B(n_418),
.Y(n_845)
);

INVx2_ASAP7_75t_SL g846 ( 
.A(n_582),
.Y(n_846)
);

AOI22xp33_ASAP7_75t_L g847 ( 
.A1(n_597),
.A2(n_554),
.B1(n_556),
.B2(n_241),
.Y(n_847)
);

INVx2_ASAP7_75t_SL g848 ( 
.A(n_582),
.Y(n_848)
);

NOR2xp33_ASAP7_75t_L g849 ( 
.A(n_605),
.B(n_521),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_675),
.B(n_554),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_677),
.B(n_554),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_SL g852 ( 
.A(n_710),
.B(n_556),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_727),
.Y(n_853)
);

NAND2xp33_ASAP7_75t_L g854 ( 
.A(n_722),
.B(n_521),
.Y(n_854)
);

OR2x2_ASAP7_75t_L g855 ( 
.A(n_615),
.B(n_437),
.Y(n_855)
);

OR2x6_ASAP7_75t_L g856 ( 
.A(n_605),
.B(n_556),
.Y(n_856)
);

BUFx6f_ASAP7_75t_L g857 ( 
.A(n_614),
.Y(n_857)
);

NOR2xp33_ASAP7_75t_L g858 ( 
.A(n_582),
.B(n_556),
.Y(n_858)
);

INVxp67_ASAP7_75t_SL g859 ( 
.A(n_730),
.Y(n_859)
);

AND2x2_ASAP7_75t_L g860 ( 
.A(n_616),
.B(n_451),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_SL g861 ( 
.A(n_722),
.B(n_556),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_SL g862 ( 
.A(n_715),
.B(n_360),
.Y(n_862)
);

INVx2_ASAP7_75t_L g863 ( 
.A(n_624),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_728),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_SL g865 ( 
.A(n_622),
.B(n_359),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_656),
.B(n_369),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_728),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_SL g868 ( 
.A(n_673),
.B(n_654),
.Y(n_868)
);

OR2x2_ASAP7_75t_L g869 ( 
.A(n_705),
.B(n_454),
.Y(n_869)
);

NOR2xp33_ASAP7_75t_L g870 ( 
.A(n_582),
.B(n_361),
.Y(n_870)
);

NOR2xp33_ASAP7_75t_L g871 ( 
.A(n_582),
.B(n_365),
.Y(n_871)
);

AND2x2_ASAP7_75t_L g872 ( 
.A(n_660),
.B(n_456),
.Y(n_872)
);

INVxp67_ASAP7_75t_L g873 ( 
.A(n_674),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_624),
.Y(n_874)
);

NOR2x1p5_ASAP7_75t_L g875 ( 
.A(n_654),
.B(n_367),
.Y(n_875)
);

NOR2xp33_ASAP7_75t_SL g876 ( 
.A(n_583),
.B(n_671),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_669),
.B(n_369),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_672),
.B(n_386),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_629),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_729),
.Y(n_880)
);

AOI22xp5_ASAP7_75t_L g881 ( 
.A1(n_650),
.A2(n_386),
.B1(n_388),
.B2(n_389),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_SL g882 ( 
.A(n_694),
.B(n_373),
.Y(n_882)
);

BUFx5_ASAP7_75t_L g883 ( 
.A(n_715),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_639),
.B(n_388),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_SL g885 ( 
.A(n_604),
.B(n_381),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_729),
.Y(n_886)
);

NOR2xp33_ASAP7_75t_L g887 ( 
.A(n_671),
.B(n_382),
.Y(n_887)
);

AOI22xp33_ASAP7_75t_L g888 ( 
.A1(n_717),
.A2(n_252),
.B1(n_396),
.B2(n_395),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_731),
.Y(n_889)
);

INVx8_ASAP7_75t_L g890 ( 
.A(n_583),
.Y(n_890)
);

NOR2xp33_ASAP7_75t_L g891 ( 
.A(n_671),
.B(n_390),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_639),
.B(n_389),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_642),
.B(n_241),
.Y(n_893)
);

INVxp67_ASAP7_75t_L g894 ( 
.A(n_725),
.Y(n_894)
);

BUFx6f_ASAP7_75t_L g895 ( 
.A(n_641),
.Y(n_895)
);

HB1xp67_ASAP7_75t_L g896 ( 
.A(n_671),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_642),
.B(n_251),
.Y(n_897)
);

AND2x2_ASAP7_75t_L g898 ( 
.A(n_671),
.B(n_468),
.Y(n_898)
);

BUFx6f_ASAP7_75t_SL g899 ( 
.A(n_717),
.Y(n_899)
);

AO221x1_ASAP7_75t_L g900 ( 
.A1(n_583),
.A2(n_281),
.B1(n_312),
.B2(n_268),
.C(n_342),
.Y(n_900)
);

AND2x2_ASAP7_75t_L g901 ( 
.A(n_725),
.B(n_473),
.Y(n_901)
);

NOR2xp33_ASAP7_75t_L g902 ( 
.A(n_718),
.B(n_391),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_644),
.B(n_251),
.Y(n_903)
);

INVx2_ASAP7_75t_L g904 ( 
.A(n_753),
.Y(n_904)
);

AND2x2_ASAP7_75t_L g905 ( 
.A(n_755),
.B(n_480),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_761),
.Y(n_906)
);

AOI21xp5_ASAP7_75t_L g907 ( 
.A1(n_759),
.A2(n_604),
.B(n_649),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_766),
.B(n_731),
.Y(n_908)
);

AND2x2_ASAP7_75t_SL g909 ( 
.A(n_876),
.B(n_667),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_SL g910 ( 
.A(n_883),
.B(n_641),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_737),
.B(n_644),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_737),
.B(n_647),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_771),
.Y(n_913)
);

AOI21xp5_ASAP7_75t_L g914 ( 
.A1(n_759),
.A2(n_604),
.B(n_649),
.Y(n_914)
);

INVx4_ASAP7_75t_L g915 ( 
.A(n_818),
.Y(n_915)
);

INVx1_ASAP7_75t_SL g916 ( 
.A(n_821),
.Y(n_916)
);

AOI21xp5_ASAP7_75t_L g917 ( 
.A1(n_790),
.A2(n_658),
.B(n_652),
.Y(n_917)
);

AOI21xp5_ASAP7_75t_L g918 ( 
.A1(n_790),
.A2(n_658),
.B(n_652),
.Y(n_918)
);

AOI21xp5_ASAP7_75t_L g919 ( 
.A1(n_822),
.A2(n_704),
.B(n_684),
.Y(n_919)
);

AOI21xp5_ASAP7_75t_L g920 ( 
.A1(n_822),
.A2(n_704),
.B(n_684),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_791),
.B(n_647),
.Y(n_921)
);

OAI21xp33_ASAP7_75t_L g922 ( 
.A1(n_735),
.A2(n_394),
.B(n_393),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_743),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_770),
.B(n_629),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_773),
.B(n_630),
.Y(n_925)
);

O2A1O1Ixp5_ASAP7_75t_L g926 ( 
.A1(n_885),
.A2(n_683),
.B(n_719),
.C(n_709),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_767),
.B(n_630),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_781),
.B(n_634),
.Y(n_928)
);

HB1xp67_ASAP7_75t_L g929 ( 
.A(n_818),
.Y(n_929)
);

OAI22xp5_ASAP7_75t_L g930 ( 
.A1(n_803),
.A2(n_718),
.B1(n_683),
.B2(n_700),
.Y(n_930)
);

INVx3_ASAP7_75t_L g931 ( 
.A(n_763),
.Y(n_931)
);

INVx4_ASAP7_75t_L g932 ( 
.A(n_818),
.Y(n_932)
);

NOR3xp33_ASAP7_75t_L g933 ( 
.A(n_829),
.B(n_257),
.C(n_252),
.Y(n_933)
);

AOI21xp5_ASAP7_75t_L g934 ( 
.A1(n_824),
.A2(n_726),
.B(n_716),
.Y(n_934)
);

HB1xp67_ASAP7_75t_L g935 ( 
.A(n_856),
.Y(n_935)
);

HB1xp67_ASAP7_75t_L g936 ( 
.A(n_856),
.Y(n_936)
);

AOI21xp5_ASAP7_75t_L g937 ( 
.A1(n_815),
.A2(n_726),
.B(n_716),
.Y(n_937)
);

AOI21xp5_ASAP7_75t_L g938 ( 
.A1(n_787),
.A2(n_708),
.B(n_700),
.Y(n_938)
);

AOI21xp5_ASAP7_75t_L g939 ( 
.A1(n_787),
.A2(n_708),
.B(n_700),
.Y(n_939)
);

AND2x4_ASAP7_75t_L g940 ( 
.A(n_856),
.B(n_683),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_751),
.Y(n_941)
);

AOI21x1_ASAP7_75t_L g942 ( 
.A1(n_823),
.A2(n_827),
.B(n_862),
.Y(n_942)
);

INVx2_ASAP7_75t_L g943 ( 
.A(n_794),
.Y(n_943)
);

CKINVDCx14_ASAP7_75t_R g944 ( 
.A(n_779),
.Y(n_944)
);

AO21x1_ASAP7_75t_L g945 ( 
.A1(n_862),
.A2(n_831),
.B(n_752),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_782),
.B(n_788),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_741),
.B(n_634),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_741),
.B(n_708),
.Y(n_948)
);

INVx2_ASAP7_75t_L g949 ( 
.A(n_795),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_SL g950 ( 
.A(n_883),
.B(n_641),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_780),
.B(n_718),
.Y(n_951)
);

INVx2_ASAP7_75t_L g952 ( 
.A(n_796),
.Y(n_952)
);

OR2x6_ASAP7_75t_L g953 ( 
.A(n_890),
.B(n_586),
.Y(n_953)
);

OAI21xp5_ASAP7_75t_L g954 ( 
.A1(n_823),
.A2(n_587),
.B(n_586),
.Y(n_954)
);

OAI22x1_ASAP7_75t_L g955 ( 
.A1(n_776),
.A2(n_485),
.B1(n_486),
.B2(n_299),
.Y(n_955)
);

BUFx2_ASAP7_75t_L g956 ( 
.A(n_805),
.Y(n_956)
);

AOI22xp5_ASAP7_75t_L g957 ( 
.A1(n_739),
.A2(n_618),
.B1(n_668),
.B2(n_676),
.Y(n_957)
);

AOI21xp5_ASAP7_75t_L g958 ( 
.A1(n_827),
.A2(n_593),
.B(n_587),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_757),
.Y(n_959)
);

A2O1A1Ixp33_ASAP7_75t_L g960 ( 
.A1(n_888),
.A2(n_325),
.B(n_257),
.C(n_323),
.Y(n_960)
);

OAI22xp5_ASAP7_75t_L g961 ( 
.A1(n_803),
.A2(n_888),
.B1(n_847),
.B2(n_745),
.Y(n_961)
);

AOI21xp5_ASAP7_75t_L g962 ( 
.A1(n_832),
.A2(n_598),
.B(n_593),
.Y(n_962)
);

NOR3xp33_ASAP7_75t_L g963 ( 
.A(n_739),
.B(n_272),
.C(n_261),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_760),
.B(n_618),
.Y(n_964)
);

AOI33xp33_ASAP7_75t_L g965 ( 
.A1(n_845),
.A2(n_299),
.A3(n_310),
.B1(n_261),
.B2(n_318),
.B3(n_319),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_SL g966 ( 
.A(n_883),
.B(n_641),
.Y(n_966)
);

NOR2xp67_ASAP7_75t_L g967 ( 
.A(n_804),
.B(n_618),
.Y(n_967)
);

INVx2_ASAP7_75t_L g968 ( 
.A(n_802),
.Y(n_968)
);

AOI21xp5_ASAP7_75t_L g969 ( 
.A1(n_752),
.A2(n_600),
.B(n_598),
.Y(n_969)
);

AOI21xp5_ASAP7_75t_L g970 ( 
.A1(n_840),
.A2(n_602),
.B(n_600),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_SL g971 ( 
.A(n_883),
.B(n_641),
.Y(n_971)
);

AOI21xp5_ASAP7_75t_L g972 ( 
.A1(n_840),
.A2(n_606),
.B(n_602),
.Y(n_972)
);

AOI21xp5_ASAP7_75t_L g973 ( 
.A1(n_859),
.A2(n_608),
.B(n_606),
.Y(n_973)
);

AOI21xp5_ASAP7_75t_L g974 ( 
.A1(n_859),
.A2(n_612),
.B(n_608),
.Y(n_974)
);

AOI22xp5_ASAP7_75t_L g975 ( 
.A1(n_887),
.A2(n_668),
.B1(n_676),
.B2(n_686),
.Y(n_975)
);

NOR2xp33_ASAP7_75t_L g976 ( 
.A(n_754),
.B(n_668),
.Y(n_976)
);

NAND2x1_ASAP7_75t_L g977 ( 
.A(n_768),
.B(n_676),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_747),
.B(n_686),
.Y(n_978)
);

AOI21xp5_ASAP7_75t_L g979 ( 
.A1(n_733),
.A2(n_619),
.B(n_612),
.Y(n_979)
);

AOI21xp5_ASAP7_75t_L g980 ( 
.A1(n_734),
.A2(n_620),
.B(n_619),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_747),
.B(n_686),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_769),
.Y(n_982)
);

OAI21xp5_ASAP7_75t_L g983 ( 
.A1(n_758),
.A2(n_625),
.B(n_620),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_765),
.B(n_625),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_765),
.B(n_636),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_785),
.B(n_636),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_SL g987 ( 
.A(n_883),
.B(n_682),
.Y(n_987)
);

AOI21xp5_ASAP7_75t_L g988 ( 
.A1(n_793),
.A2(n_645),
.B(n_637),
.Y(n_988)
);

AOI22xp5_ASAP7_75t_L g989 ( 
.A1(n_887),
.A2(n_666),
.B1(n_637),
.B2(n_664),
.Y(n_989)
);

NOR2xp33_ASAP7_75t_L g990 ( 
.A(n_786),
.B(n_645),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_785),
.B(n_648),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_786),
.B(n_648),
.Y(n_992)
);

AOI21xp5_ASAP7_75t_L g993 ( 
.A1(n_797),
.A2(n_659),
.B(n_657),
.Y(n_993)
);

OAI22xp5_ASAP7_75t_L g994 ( 
.A1(n_847),
.A2(n_744),
.B1(n_756),
.B2(n_748),
.Y(n_994)
);

AOI21xp5_ASAP7_75t_L g995 ( 
.A1(n_778),
.A2(n_659),
.B(n_657),
.Y(n_995)
);

OAI21xp5_ASAP7_75t_L g996 ( 
.A1(n_820),
.A2(n_666),
.B(n_664),
.Y(n_996)
);

O2A1O1Ixp33_ASAP7_75t_L g997 ( 
.A1(n_811),
.A2(n_349),
.B(n_362),
.C(n_395),
.Y(n_997)
);

BUFx4f_ASAP7_75t_L g998 ( 
.A(n_801),
.Y(n_998)
);

OAI21xp5_ASAP7_75t_L g999 ( 
.A1(n_798),
.A2(n_688),
.B(n_690),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_783),
.Y(n_1000)
);

AOI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_762),
.A2(n_854),
.B(n_812),
.Y(n_1001)
);

AND2x4_ASAP7_75t_L g1002 ( 
.A(n_875),
.B(n_688),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_772),
.B(n_682),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_784),
.Y(n_1004)
);

INVx2_ASAP7_75t_L g1005 ( 
.A(n_806),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_775),
.B(n_807),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_SL g1007 ( 
.A(n_883),
.B(n_682),
.Y(n_1007)
);

AOI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_814),
.A2(n_707),
.B(n_685),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_800),
.Y(n_1009)
);

AND2x2_ASAP7_75t_L g1010 ( 
.A(n_813),
.B(n_372),
.Y(n_1010)
);

O2A1O1Ixp33_ASAP7_75t_L g1011 ( 
.A1(n_750),
.A2(n_347),
.B(n_379),
.C(n_378),
.Y(n_1011)
);

BUFx12f_ASAP7_75t_L g1012 ( 
.A(n_833),
.Y(n_1012)
);

AND2x2_ASAP7_75t_L g1013 ( 
.A(n_740),
.B(n_372),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_816),
.B(n_682),
.Y(n_1014)
);

AOI21xp5_ASAP7_75t_L g1015 ( 
.A1(n_850),
.A2(n_707),
.B(n_685),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_736),
.B(n_742),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_736),
.B(n_682),
.Y(n_1017)
);

INVx2_ASAP7_75t_L g1018 ( 
.A(n_817),
.Y(n_1018)
);

OAI21xp33_ASAP7_75t_L g1019 ( 
.A1(n_902),
.A2(n_319),
.B(n_318),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_SL g1020 ( 
.A(n_849),
.B(n_685),
.Y(n_1020)
);

AOI21x1_ASAP7_75t_L g1021 ( 
.A1(n_884),
.A2(n_511),
.B(n_508),
.Y(n_1021)
);

AOI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_851),
.A2(n_837),
.B(n_830),
.Y(n_1022)
);

NOR2xp33_ASAP7_75t_L g1023 ( 
.A(n_740),
.B(n_685),
.Y(n_1023)
);

OAI22xp5_ASAP7_75t_L g1024 ( 
.A1(n_774),
.A2(n_707),
.B1(n_706),
.B2(n_696),
.Y(n_1024)
);

AOI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_825),
.A2(n_696),
.B(n_685),
.Y(n_1025)
);

AOI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_843),
.A2(n_707),
.B(n_706),
.Y(n_1026)
);

AOI21xp5_ASAP7_75t_L g1027 ( 
.A1(n_844),
.A2(n_864),
.B(n_853),
.Y(n_1027)
);

AOI22xp5_ASAP7_75t_L g1028 ( 
.A1(n_891),
.A2(n_899),
.B1(n_871),
.B2(n_870),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_742),
.B(n_696),
.Y(n_1029)
);

NOR2xp33_ASAP7_75t_SL g1030 ( 
.A(n_894),
.B(n_372),
.Y(n_1030)
);

AOI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_867),
.A2(n_706),
.B(n_696),
.Y(n_1031)
);

O2A1O1Ixp33_ASAP7_75t_SL g1032 ( 
.A1(n_880),
.A2(n_349),
.B(n_379),
.C(n_378),
.Y(n_1032)
);

BUFx6f_ASAP7_75t_L g1033 ( 
.A(n_768),
.Y(n_1033)
);

AND2x2_ASAP7_75t_L g1034 ( 
.A(n_740),
.B(n_323),
.Y(n_1034)
);

INVx2_ASAP7_75t_SL g1035 ( 
.A(n_901),
.Y(n_1035)
);

AOI21xp5_ASAP7_75t_L g1036 ( 
.A1(n_886),
.A2(n_889),
.B(n_842),
.Y(n_1036)
);

AOI21xp5_ASAP7_75t_L g1037 ( 
.A1(n_842),
.A2(n_707),
.B(n_706),
.Y(n_1037)
);

AOI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_746),
.A2(n_706),
.B(n_696),
.Y(n_1038)
);

INVx2_ASAP7_75t_L g1039 ( 
.A(n_826),
.Y(n_1039)
);

AOI21xp5_ASAP7_75t_L g1040 ( 
.A1(n_841),
.A2(n_690),
.B(n_701),
.Y(n_1040)
);

AND2x2_ASAP7_75t_L g1041 ( 
.A(n_898),
.B(n_325),
.Y(n_1041)
);

NOR2xp33_ASAP7_75t_L g1042 ( 
.A(n_873),
.B(n_690),
.Y(n_1042)
);

A2O1A1Ixp33_ASAP7_75t_L g1043 ( 
.A1(n_891),
.A2(n_871),
.B(n_870),
.C(n_849),
.Y(n_1043)
);

INVxp67_ASAP7_75t_L g1044 ( 
.A(n_838),
.Y(n_1044)
);

NOR2xp33_ASAP7_75t_L g1045 ( 
.A(n_834),
.B(n_690),
.Y(n_1045)
);

AOI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_902),
.A2(n_690),
.B(n_311),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_SL g1047 ( 
.A(n_768),
.B(n_777),
.Y(n_1047)
);

AND2x2_ASAP7_75t_L g1048 ( 
.A(n_819),
.B(n_342),
.Y(n_1048)
);

NOR2xp67_ASAP7_75t_L g1049 ( 
.A(n_855),
.B(n_690),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_SL g1050 ( 
.A(n_768),
.B(n_366),
.Y(n_1050)
);

OAI22xp5_ASAP7_75t_L g1051 ( 
.A1(n_899),
.A2(n_347),
.B1(n_362),
.B2(n_374),
.Y(n_1051)
);

OAI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_808),
.A2(n_301),
.B(n_263),
.Y(n_1052)
);

AOI21xp5_ASAP7_75t_L g1053 ( 
.A1(n_777),
.A2(n_304),
.B(n_205),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_SL g1054 ( 
.A(n_777),
.B(n_366),
.Y(n_1054)
);

INVx2_ASAP7_75t_L g1055 ( 
.A(n_863),
.Y(n_1055)
);

AOI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_777),
.A2(n_309),
.B(n_210),
.Y(n_1056)
);

NAND2x1p5_ASAP7_75t_L g1057 ( 
.A(n_846),
.B(n_848),
.Y(n_1057)
);

O2A1O1Ixp33_ASAP7_75t_L g1058 ( 
.A1(n_839),
.A2(n_374),
.B(n_271),
.C(n_301),
.Y(n_1058)
);

INVx2_ASAP7_75t_L g1059 ( 
.A(n_874),
.Y(n_1059)
);

AO21x1_ASAP7_75t_L g1060 ( 
.A1(n_792),
.A2(n_271),
.B(n_508),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_858),
.B(n_508),
.Y(n_1061)
);

AOI21xp5_ASAP7_75t_L g1062 ( 
.A1(n_789),
.A2(n_857),
.B(n_799),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_858),
.B(n_511),
.Y(n_1063)
);

INVxp67_ASAP7_75t_L g1064 ( 
.A(n_860),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_836),
.B(n_511),
.Y(n_1065)
);

AOI21xp5_ASAP7_75t_L g1066 ( 
.A1(n_789),
.A2(n_392),
.B(n_199),
.Y(n_1066)
);

AOI22xp5_ASAP7_75t_L g1067 ( 
.A1(n_896),
.A2(n_331),
.B1(n_213),
.B2(n_368),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_896),
.B(n_312),
.Y(n_1068)
);

OAI21xp5_ASAP7_75t_L g1069 ( 
.A1(n_810),
.A2(n_294),
.B(n_229),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_764),
.B(n_312),
.Y(n_1070)
);

AOI21x1_ASAP7_75t_L g1071 ( 
.A1(n_892),
.A2(n_366),
.B(n_371),
.Y(n_1071)
);

BUFx2_ASAP7_75t_L g1072 ( 
.A(n_779),
.Y(n_1072)
);

BUFx2_ASAP7_75t_L g1073 ( 
.A(n_869),
.Y(n_1073)
);

A2O1A1Ixp33_ASAP7_75t_L g1074 ( 
.A1(n_835),
.A2(n_312),
.B(n_247),
.C(n_223),
.Y(n_1074)
);

AOI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_789),
.A2(n_221),
.B(n_248),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_893),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_SL g1077 ( 
.A(n_789),
.B(n_366),
.Y(n_1077)
);

AOI21xp5_ASAP7_75t_L g1078 ( 
.A1(n_799),
.A2(n_314),
.B(n_237),
.Y(n_1078)
);

INVx5_ASAP7_75t_L g1079 ( 
.A(n_764),
.Y(n_1079)
);

AOI21xp5_ASAP7_75t_L g1080 ( 
.A1(n_799),
.A2(n_317),
.B(n_245),
.Y(n_1080)
);

AND2x4_ASAP7_75t_L g1081 ( 
.A(n_763),
.B(n_247),
.Y(n_1081)
);

OAI321xp33_ASAP7_75t_L g1082 ( 
.A1(n_881),
.A2(n_312),
.A3(n_227),
.B1(n_330),
.B2(n_371),
.C(n_11),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_764),
.B(n_253),
.Y(n_1083)
);

AND2x2_ASAP7_75t_SL g1084 ( 
.A(n_799),
.B(n_227),
.Y(n_1084)
);

AOI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_857),
.A2(n_326),
.B(n_255),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_SL g1086 ( 
.A(n_857),
.B(n_366),
.Y(n_1086)
);

NAND2x1p5_ASAP7_75t_L g1087 ( 
.A(n_852),
.B(n_376),
.Y(n_1087)
);

NOR2xp33_ASAP7_75t_L g1088 ( 
.A(n_865),
.B(n_7),
.Y(n_1088)
);

OAI21x1_ASAP7_75t_SL g1089 ( 
.A1(n_897),
.A2(n_8),
.B(n_9),
.Y(n_1089)
);

AOI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_857),
.A2(n_327),
.B(n_256),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_764),
.B(n_258),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_764),
.B(n_809),
.Y(n_1092)
);

AOI21xp5_ASAP7_75t_L g1093 ( 
.A1(n_895),
.A2(n_328),
.B(n_259),
.Y(n_1093)
);

NOR2xp33_ASAP7_75t_L g1094 ( 
.A(n_868),
.B(n_10),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_903),
.Y(n_1095)
);

AOI21xp5_ASAP7_75t_SL g1096 ( 
.A1(n_1043),
.A2(n_895),
.B(n_861),
.Y(n_1096)
);

CKINVDCx6p67_ASAP7_75t_R g1097 ( 
.A(n_1012),
.Y(n_1097)
);

OAI22xp5_ASAP7_75t_L g1098 ( 
.A1(n_1043),
.A2(n_866),
.B1(n_878),
.B2(n_877),
.Y(n_1098)
);

INVx2_ASAP7_75t_L g1099 ( 
.A(n_904),
.Y(n_1099)
);

AO22x1_ASAP7_75t_L g1100 ( 
.A1(n_1072),
.A2(n_963),
.B1(n_828),
.B2(n_905),
.Y(n_1100)
);

AOI21xp5_ASAP7_75t_L g1101 ( 
.A1(n_1022),
.A2(n_895),
.B(n_879),
.Y(n_1101)
);

OAI21xp5_ASAP7_75t_L g1102 ( 
.A1(n_1036),
.A2(n_882),
.B(n_809),
.Y(n_1102)
);

NOR2xp33_ASAP7_75t_SL g1103 ( 
.A(n_1084),
.B(n_890),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_923),
.Y(n_1104)
);

OAI21xp5_ASAP7_75t_L g1105 ( 
.A1(n_1017),
.A2(n_809),
.B(n_900),
.Y(n_1105)
);

INVx2_ASAP7_75t_SL g1106 ( 
.A(n_998),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_941),
.Y(n_1107)
);

INVx2_ASAP7_75t_L g1108 ( 
.A(n_904),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_946),
.B(n_890),
.Y(n_1109)
);

NOR3xp33_ASAP7_75t_L g1110 ( 
.A(n_1088),
.B(n_872),
.C(n_376),
.Y(n_1110)
);

OR2x2_ASAP7_75t_L g1111 ( 
.A(n_1073),
.B(n_749),
.Y(n_1111)
);

AND2x2_ASAP7_75t_L g1112 ( 
.A(n_1041),
.B(n_1010),
.Y(n_1112)
);

AO21x1_ASAP7_75t_L g1113 ( 
.A1(n_947),
.A2(n_819),
.B(n_895),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_1016),
.B(n_819),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_SL g1115 ( 
.A(n_1030),
.B(n_1035),
.Y(n_1115)
);

INVx2_ASAP7_75t_L g1116 ( 
.A(n_1059),
.Y(n_1116)
);

INVx2_ASAP7_75t_L g1117 ( 
.A(n_1059),
.Y(n_1117)
);

OR2x2_ASAP7_75t_L g1118 ( 
.A(n_1064),
.B(n_749),
.Y(n_1118)
);

OR2x6_ASAP7_75t_L g1119 ( 
.A(n_956),
.B(n_749),
.Y(n_1119)
);

BUFx6f_ASAP7_75t_L g1120 ( 
.A(n_1033),
.Y(n_1120)
);

AOI21x1_ASAP7_75t_L g1121 ( 
.A1(n_1071),
.A2(n_366),
.B(n_336),
.Y(n_1121)
);

BUFx3_ASAP7_75t_L g1122 ( 
.A(n_998),
.Y(n_1122)
);

A2O1A1Ixp33_ASAP7_75t_SL g1123 ( 
.A1(n_976),
.A2(n_10),
.B(n_11),
.C(n_14),
.Y(n_1123)
);

A2O1A1Ixp33_ASAP7_75t_L g1124 ( 
.A1(n_990),
.A2(n_336),
.B(n_265),
.C(n_270),
.Y(n_1124)
);

INVx2_ASAP7_75t_L g1125 ( 
.A(n_906),
.Y(n_1125)
);

NOR2xp33_ASAP7_75t_L g1126 ( 
.A(n_1044),
.B(n_738),
.Y(n_1126)
);

O2A1O1Ixp33_ASAP7_75t_L g1127 ( 
.A1(n_1088),
.A2(n_14),
.B(n_17),
.C(n_19),
.Y(n_1127)
);

AND2x4_ASAP7_75t_L g1128 ( 
.A(n_915),
.B(n_809),
.Y(n_1128)
);

OR2x6_ASAP7_75t_L g1129 ( 
.A(n_915),
.B(n_738),
.Y(n_1129)
);

INVx2_ASAP7_75t_L g1130 ( 
.A(n_913),
.Y(n_1130)
);

INVx2_ASAP7_75t_L g1131 ( 
.A(n_943),
.Y(n_1131)
);

BUFx6f_ASAP7_75t_L g1132 ( 
.A(n_1033),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_959),
.Y(n_1133)
);

O2A1O1Ixp33_ASAP7_75t_L g1134 ( 
.A1(n_963),
.A2(n_17),
.B(n_21),
.C(n_22),
.Y(n_1134)
);

A2O1A1Ixp33_ASAP7_75t_L g1135 ( 
.A1(n_990),
.A2(n_332),
.B(n_280),
.C(n_283),
.Y(n_1135)
);

NOR2xp33_ASAP7_75t_L g1136 ( 
.A(n_1028),
.B(n_288),
.Y(n_1136)
);

AOI22xp5_ASAP7_75t_L g1137 ( 
.A1(n_961),
.A2(n_809),
.B1(n_343),
.B2(n_339),
.Y(n_1137)
);

AOI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_1001),
.A2(n_289),
.B(n_358),
.Y(n_1138)
);

AOI221xp5_ASAP7_75t_L g1139 ( 
.A1(n_933),
.A2(n_355),
.B1(n_348),
.B2(n_324),
.C(n_321),
.Y(n_1139)
);

CKINVDCx20_ASAP7_75t_R g1140 ( 
.A(n_944),
.Y(n_1140)
);

NOR2x1_ASAP7_75t_L g1141 ( 
.A(n_1049),
.B(n_371),
.Y(n_1141)
);

INVx1_ASAP7_75t_SL g1142 ( 
.A(n_916),
.Y(n_1142)
);

AOI21xp5_ASAP7_75t_L g1143 ( 
.A1(n_999),
.A2(n_371),
.B(n_330),
.Y(n_1143)
);

CKINVDCx16_ASAP7_75t_R g1144 ( 
.A(n_944),
.Y(n_1144)
);

O2A1O1Ixp33_ASAP7_75t_L g1145 ( 
.A1(n_922),
.A2(n_21),
.B(n_23),
.C(n_34),
.Y(n_1145)
);

BUFx6f_ASAP7_75t_L g1146 ( 
.A(n_1033),
.Y(n_1146)
);

NOR2xp33_ASAP7_75t_L g1147 ( 
.A(n_932),
.B(n_23),
.Y(n_1147)
);

AOI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_964),
.A2(n_371),
.B(n_330),
.Y(n_1148)
);

A2O1A1Ixp33_ASAP7_75t_L g1149 ( 
.A1(n_1058),
.A2(n_330),
.B(n_227),
.C(n_366),
.Y(n_1149)
);

BUFx12f_ASAP7_75t_L g1150 ( 
.A(n_1034),
.Y(n_1150)
);

A2O1A1Ixp33_ASAP7_75t_L g1151 ( 
.A1(n_1094),
.A2(n_330),
.B(n_227),
.C(n_366),
.Y(n_1151)
);

BUFx6f_ASAP7_75t_L g1152 ( 
.A(n_1033),
.Y(n_1152)
);

BUFx12f_ASAP7_75t_L g1153 ( 
.A(n_1013),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_1006),
.B(n_37),
.Y(n_1154)
);

INVx4_ASAP7_75t_L g1155 ( 
.A(n_953),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_SL g1156 ( 
.A(n_940),
.B(n_227),
.Y(n_1156)
);

OAI21xp33_ASAP7_75t_L g1157 ( 
.A1(n_1019),
.A2(n_40),
.B(n_41),
.Y(n_1157)
);

AOI21xp5_ASAP7_75t_L g1158 ( 
.A1(n_1008),
.A2(n_105),
.B(n_192),
.Y(n_1158)
);

BUFx6f_ASAP7_75t_L g1159 ( 
.A(n_953),
.Y(n_1159)
);

NOR2xp33_ASAP7_75t_L g1160 ( 
.A(n_932),
.B(n_42),
.Y(n_1160)
);

INVxp67_ASAP7_75t_L g1161 ( 
.A(n_1094),
.Y(n_1161)
);

BUFx2_ASAP7_75t_L g1162 ( 
.A(n_929),
.Y(n_1162)
);

INVx2_ASAP7_75t_L g1163 ( 
.A(n_949),
.Y(n_1163)
);

INVx2_ASAP7_75t_L g1164 ( 
.A(n_952),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_911),
.B(n_45),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_L g1166 ( 
.A(n_912),
.B(n_47),
.Y(n_1166)
);

BUFx6f_ASAP7_75t_L g1167 ( 
.A(n_953),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_SL g1168 ( 
.A(n_940),
.B(n_48),
.Y(n_1168)
);

AO21x1_ASAP7_75t_L g1169 ( 
.A1(n_1020),
.A2(n_111),
.B(n_188),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_982),
.Y(n_1170)
);

AND2x2_ASAP7_75t_L g1171 ( 
.A(n_1048),
.B(n_933),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_L g1172 ( 
.A(n_1076),
.B(n_48),
.Y(n_1172)
);

CKINVDCx5p33_ASAP7_75t_R g1173 ( 
.A(n_955),
.Y(n_1173)
);

AOI21xp5_ASAP7_75t_L g1174 ( 
.A1(n_1015),
.A2(n_106),
.B(n_185),
.Y(n_1174)
);

BUFx2_ASAP7_75t_L g1175 ( 
.A(n_929),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_1000),
.Y(n_1176)
);

AOI21xp5_ASAP7_75t_L g1177 ( 
.A1(n_992),
.A2(n_104),
.B(n_181),
.Y(n_1177)
);

AOI21x1_ASAP7_75t_L g1178 ( 
.A1(n_1021),
.A2(n_94),
.B(n_178),
.Y(n_1178)
);

AOI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_984),
.A2(n_93),
.B(n_166),
.Y(n_1179)
);

INVxp67_ASAP7_75t_L g1180 ( 
.A(n_1051),
.Y(n_1180)
);

AND2x2_ASAP7_75t_L g1181 ( 
.A(n_935),
.B(n_51),
.Y(n_1181)
);

AND2x4_ASAP7_75t_SL g1182 ( 
.A(n_935),
.B(n_52),
.Y(n_1182)
);

AND2x2_ASAP7_75t_L g1183 ( 
.A(n_936),
.B(n_52),
.Y(n_1183)
);

BUFx6f_ASAP7_75t_L g1184 ( 
.A(n_1079),
.Y(n_1184)
);

AOI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_985),
.A2(n_114),
.B(n_165),
.Y(n_1185)
);

AO32x2_ASAP7_75t_L g1186 ( 
.A1(n_1024),
.A2(n_54),
.A3(n_55),
.B1(n_56),
.B2(n_61),
.Y(n_1186)
);

INVx2_ASAP7_75t_L g1187 ( 
.A(n_968),
.Y(n_1187)
);

AOI21xp5_ASAP7_75t_L g1188 ( 
.A1(n_986),
.A2(n_117),
.B(n_164),
.Y(n_1188)
);

AO21x1_ASAP7_75t_L g1189 ( 
.A1(n_1020),
.A2(n_92),
.B(n_160),
.Y(n_1189)
);

NAND2x1p5_ASAP7_75t_L g1190 ( 
.A(n_1079),
.B(n_82),
.Y(n_1190)
);

NOR2xp33_ASAP7_75t_L g1191 ( 
.A(n_936),
.B(n_54),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_1095),
.B(n_994),
.Y(n_1192)
);

INVx2_ASAP7_75t_L g1193 ( 
.A(n_1005),
.Y(n_1193)
);

A2O1A1Ixp33_ASAP7_75t_SL g1194 ( 
.A1(n_976),
.A2(n_61),
.B(n_62),
.C(n_65),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_SL g1195 ( 
.A(n_1084),
.B(n_65),
.Y(n_1195)
);

AOI21xp5_ASAP7_75t_L g1196 ( 
.A1(n_991),
.A2(n_131),
.B(n_155),
.Y(n_1196)
);

INVx2_ASAP7_75t_L g1197 ( 
.A(n_1018),
.Y(n_1197)
);

CKINVDCx8_ASAP7_75t_R g1198 ( 
.A(n_1002),
.Y(n_1198)
);

AOI21xp5_ASAP7_75t_L g1199 ( 
.A1(n_937),
.A2(n_981),
.B(n_978),
.Y(n_1199)
);

A2O1A1Ixp33_ASAP7_75t_L g1200 ( 
.A1(n_960),
.A2(n_66),
.B(n_67),
.C(n_70),
.Y(n_1200)
);

A2O1A1Ixp33_ASAP7_75t_L g1201 ( 
.A1(n_960),
.A2(n_67),
.B(n_71),
.C(n_76),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_SL g1202 ( 
.A(n_1023),
.B(n_71),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_1004),
.Y(n_1203)
);

NOR2xp33_ASAP7_75t_L g1204 ( 
.A(n_908),
.B(n_76),
.Y(n_1204)
);

INVx2_ASAP7_75t_L g1205 ( 
.A(n_1039),
.Y(n_1205)
);

AND2x2_ASAP7_75t_L g1206 ( 
.A(n_965),
.B(n_198),
.Y(n_1206)
);

INVx2_ASAP7_75t_L g1207 ( 
.A(n_1055),
.Y(n_1207)
);

AOI21xp5_ASAP7_75t_L g1208 ( 
.A1(n_917),
.A2(n_118),
.B(n_122),
.Y(n_1208)
);

INVx3_ASAP7_75t_SL g1209 ( 
.A(n_1002),
.Y(n_1209)
);

O2A1O1Ixp33_ASAP7_75t_L g1210 ( 
.A1(n_1032),
.A2(n_135),
.B(n_145),
.C(n_149),
.Y(n_1210)
);

NOR2xp33_ASAP7_75t_L g1211 ( 
.A(n_1067),
.B(n_150),
.Y(n_1211)
);

AOI21xp5_ASAP7_75t_L g1212 ( 
.A1(n_918),
.A2(n_919),
.B(n_920),
.Y(n_1212)
);

NOR2x1_ASAP7_75t_L g1213 ( 
.A(n_967),
.B(n_931),
.Y(n_1213)
);

AOI22x1_ASAP7_75t_L g1214 ( 
.A1(n_938),
.A2(n_939),
.B1(n_995),
.B2(n_914),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_SL g1215 ( 
.A(n_1023),
.B(n_931),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_927),
.B(n_924),
.Y(n_1216)
);

NOR2xp33_ASAP7_75t_L g1217 ( 
.A(n_1009),
.B(n_951),
.Y(n_1217)
);

INVx2_ASAP7_75t_SL g1218 ( 
.A(n_1081),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_925),
.B(n_921),
.Y(n_1219)
);

BUFx6f_ASAP7_75t_L g1220 ( 
.A(n_1079),
.Y(n_1220)
);

INVx3_ASAP7_75t_L g1221 ( 
.A(n_1079),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_928),
.Y(n_1222)
);

INVx8_ASAP7_75t_L g1223 ( 
.A(n_1081),
.Y(n_1223)
);

AOI221xp5_ASAP7_75t_L g1224 ( 
.A1(n_1082),
.A2(n_1032),
.B1(n_997),
.B2(n_1011),
.C(n_1027),
.Y(n_1224)
);

INVx1_ASAP7_75t_SL g1225 ( 
.A(n_1029),
.Y(n_1225)
);

BUFx3_ASAP7_75t_L g1226 ( 
.A(n_1057),
.Y(n_1226)
);

BUFx6f_ASAP7_75t_L g1227 ( 
.A(n_1057),
.Y(n_1227)
);

CKINVDCx8_ASAP7_75t_R g1228 ( 
.A(n_1042),
.Y(n_1228)
);

NOR2xp33_ASAP7_75t_SL g1229 ( 
.A(n_909),
.B(n_1092),
.Y(n_1229)
);

BUFx6f_ASAP7_75t_L g1230 ( 
.A(n_977),
.Y(n_1230)
);

NAND2xp33_ASAP7_75t_SL g1231 ( 
.A(n_948),
.B(n_965),
.Y(n_1231)
);

O2A1O1Ixp33_ASAP7_75t_L g1232 ( 
.A1(n_1089),
.A2(n_1074),
.B(n_996),
.C(n_983),
.Y(n_1232)
);

INVx2_ASAP7_75t_L g1233 ( 
.A(n_1065),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_SL g1234 ( 
.A(n_1042),
.B(n_909),
.Y(n_1234)
);

BUFx2_ASAP7_75t_L g1235 ( 
.A(n_1087),
.Y(n_1235)
);

NOR2xp33_ASAP7_75t_R g1236 ( 
.A(n_942),
.B(n_1083),
.Y(n_1236)
);

NAND2xp33_ASAP7_75t_L g1237 ( 
.A(n_975),
.B(n_957),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_1061),
.B(n_1063),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_945),
.B(n_1052),
.Y(n_1239)
);

AOI21xp5_ASAP7_75t_L g1240 ( 
.A1(n_934),
.A2(n_1031),
.B(n_1026),
.Y(n_1240)
);

CKINVDCx5p33_ASAP7_75t_R g1241 ( 
.A(n_1045),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_L g1242 ( 
.A(n_1003),
.B(n_989),
.Y(n_1242)
);

A2O1A1Ixp33_ASAP7_75t_L g1243 ( 
.A1(n_1045),
.A2(n_1069),
.B(n_926),
.C(n_962),
.Y(n_1243)
);

NOR3xp33_ASAP7_75t_SL g1244 ( 
.A(n_1074),
.B(n_1093),
.C(n_1090),
.Y(n_1244)
);

AOI21xp5_ASAP7_75t_L g1245 ( 
.A1(n_1025),
.A2(n_907),
.B(n_1037),
.Y(n_1245)
);

INVx2_ASAP7_75t_L g1246 ( 
.A(n_1014),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1068),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1087),
.Y(n_1248)
);

A2O1A1Ixp33_ASAP7_75t_L g1249 ( 
.A1(n_969),
.A2(n_974),
.B(n_973),
.C(n_972),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_954),
.Y(n_1250)
);

NOR2xp33_ASAP7_75t_L g1251 ( 
.A(n_1047),
.B(n_1054),
.Y(n_1251)
);

INVx1_ASAP7_75t_SL g1252 ( 
.A(n_1070),
.Y(n_1252)
);

OAI22x1_ASAP7_75t_L g1253 ( 
.A1(n_1050),
.A2(n_1054),
.B1(n_1086),
.B2(n_1077),
.Y(n_1253)
);

AOI21xp5_ASAP7_75t_L g1254 ( 
.A1(n_1062),
.A2(n_910),
.B(n_1007),
.Y(n_1254)
);

AOI21xp5_ASAP7_75t_L g1255 ( 
.A1(n_910),
.A2(n_1007),
.B(n_950),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_L g1256 ( 
.A(n_979),
.B(n_980),
.Y(n_1256)
);

BUFx6f_ASAP7_75t_L g1257 ( 
.A(n_1047),
.Y(n_1257)
);

NOR2xp33_ASAP7_75t_L g1258 ( 
.A(n_1050),
.B(n_1086),
.Y(n_1258)
);

OAI22xp5_ASAP7_75t_L g1259 ( 
.A1(n_930),
.A2(n_970),
.B1(n_958),
.B2(n_988),
.Y(n_1259)
);

OAI21x1_ASAP7_75t_L g1260 ( 
.A1(n_1240),
.A2(n_950),
.B(n_966),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1104),
.Y(n_1261)
);

OA21x2_ASAP7_75t_L g1262 ( 
.A1(n_1245),
.A2(n_1060),
.B(n_1077),
.Y(n_1262)
);

INVx8_ASAP7_75t_L g1263 ( 
.A(n_1223),
.Y(n_1263)
);

OA21x2_ASAP7_75t_L g1264 ( 
.A1(n_1199),
.A2(n_1239),
.B(n_1256),
.Y(n_1264)
);

OAI21x1_ASAP7_75t_L g1265 ( 
.A1(n_1214),
.A2(n_966),
.B(n_971),
.Y(n_1265)
);

AO21x2_ASAP7_75t_L g1266 ( 
.A1(n_1239),
.A2(n_971),
.B(n_987),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1107),
.Y(n_1267)
);

AO31x2_ASAP7_75t_L g1268 ( 
.A1(n_1113),
.A2(n_1243),
.A3(n_1259),
.B(n_1256),
.Y(n_1268)
);

AOI21xp5_ASAP7_75t_L g1269 ( 
.A1(n_1098),
.A2(n_987),
.B(n_1038),
.Y(n_1269)
);

INVx4_ASAP7_75t_L g1270 ( 
.A(n_1122),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_L g1271 ( 
.A(n_1112),
.B(n_1066),
.Y(n_1271)
);

O2A1O1Ixp33_ASAP7_75t_L g1272 ( 
.A1(n_1161),
.A2(n_1040),
.B(n_993),
.C(n_1046),
.Y(n_1272)
);

AO31x2_ASAP7_75t_L g1273 ( 
.A1(n_1259),
.A2(n_1091),
.A3(n_1056),
.B(n_1075),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_SL g1274 ( 
.A(n_1241),
.B(n_1053),
.Y(n_1274)
);

NOR2x1_ASAP7_75t_SL g1275 ( 
.A(n_1184),
.B(n_1078),
.Y(n_1275)
);

AOI21xp5_ASAP7_75t_L g1276 ( 
.A1(n_1098),
.A2(n_1080),
.B(n_1085),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1133),
.Y(n_1277)
);

AO31x2_ASAP7_75t_L g1278 ( 
.A1(n_1253),
.A2(n_1143),
.A3(n_1249),
.B(n_1212),
.Y(n_1278)
);

AOI21xp5_ASAP7_75t_L g1279 ( 
.A1(n_1192),
.A2(n_1238),
.B(n_1237),
.Y(n_1279)
);

NOR2xp33_ASAP7_75t_L g1280 ( 
.A(n_1209),
.B(n_1180),
.Y(n_1280)
);

OAI21x1_ASAP7_75t_SL g1281 ( 
.A1(n_1192),
.A2(n_1232),
.B(n_1154),
.Y(n_1281)
);

BUFx3_ASAP7_75t_L g1282 ( 
.A(n_1140),
.Y(n_1282)
);

AOI21xp5_ASAP7_75t_L g1283 ( 
.A1(n_1238),
.A2(n_1216),
.B(n_1096),
.Y(n_1283)
);

INVx2_ASAP7_75t_SL g1284 ( 
.A(n_1144),
.Y(n_1284)
);

NAND3xp33_ASAP7_75t_L g1285 ( 
.A(n_1127),
.B(n_1204),
.C(n_1134),
.Y(n_1285)
);

NOR2xp33_ASAP7_75t_L g1286 ( 
.A(n_1109),
.B(n_1115),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_L g1287 ( 
.A(n_1171),
.B(n_1114),
.Y(n_1287)
);

AO31x2_ASAP7_75t_L g1288 ( 
.A1(n_1254),
.A2(n_1151),
.A3(n_1255),
.B(n_1148),
.Y(n_1288)
);

AOI22xp5_ASAP7_75t_L g1289 ( 
.A1(n_1231),
.A2(n_1157),
.B1(n_1136),
.B2(n_1211),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_L g1290 ( 
.A(n_1114),
.B(n_1109),
.Y(n_1290)
);

AOI21xp5_ASAP7_75t_L g1291 ( 
.A1(n_1216),
.A2(n_1219),
.B(n_1101),
.Y(n_1291)
);

A2O1A1Ixp33_ASAP7_75t_L g1292 ( 
.A1(n_1224),
.A2(n_1110),
.B(n_1217),
.C(n_1137),
.Y(n_1292)
);

OAI21xp5_ASAP7_75t_L g1293 ( 
.A1(n_1154),
.A2(n_1242),
.B(n_1165),
.Y(n_1293)
);

A2O1A1Ixp33_ASAP7_75t_L g1294 ( 
.A1(n_1145),
.A2(n_1139),
.B(n_1165),
.C(n_1166),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1170),
.Y(n_1295)
);

OR2x2_ASAP7_75t_L g1296 ( 
.A(n_1111),
.B(n_1118),
.Y(n_1296)
);

O2A1O1Ixp33_ASAP7_75t_SL g1297 ( 
.A1(n_1135),
.A2(n_1166),
.B(n_1234),
.C(n_1124),
.Y(n_1297)
);

A2O1A1Ixp33_ASAP7_75t_L g1298 ( 
.A1(n_1139),
.A2(n_1172),
.B(n_1258),
.C(n_1195),
.Y(n_1298)
);

AND2x2_ASAP7_75t_L g1299 ( 
.A(n_1181),
.B(n_1183),
.Y(n_1299)
);

AO22x2_ASAP7_75t_L g1300 ( 
.A1(n_1225),
.A2(n_1119),
.B1(n_1246),
.B2(n_1206),
.Y(n_1300)
);

AND2x2_ASAP7_75t_L g1301 ( 
.A(n_1162),
.B(n_1175),
.Y(n_1301)
);

NOR2xp33_ASAP7_75t_L g1302 ( 
.A(n_1198),
.B(n_1150),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1176),
.Y(n_1303)
);

O2A1O1Ixp33_ASAP7_75t_L g1304 ( 
.A1(n_1200),
.A2(n_1201),
.B(n_1194),
.C(n_1123),
.Y(n_1304)
);

BUFx3_ASAP7_75t_L g1305 ( 
.A(n_1097),
.Y(n_1305)
);

OAI21xp5_ASAP7_75t_L g1306 ( 
.A1(n_1242),
.A2(n_1250),
.B(n_1251),
.Y(n_1306)
);

BUFx6f_ASAP7_75t_L g1307 ( 
.A(n_1159),
.Y(n_1307)
);

O2A1O1Ixp33_ASAP7_75t_L g1308 ( 
.A1(n_1168),
.A2(n_1202),
.B(n_1172),
.C(n_1191),
.Y(n_1308)
);

AOI21xp5_ASAP7_75t_L g1309 ( 
.A1(n_1219),
.A2(n_1208),
.B(n_1188),
.Y(n_1309)
);

AOI21xp5_ASAP7_75t_L g1310 ( 
.A1(n_1177),
.A2(n_1196),
.B(n_1185),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_L g1311 ( 
.A(n_1222),
.B(n_1142),
.Y(n_1311)
);

AO31x2_ASAP7_75t_L g1312 ( 
.A1(n_1169),
.A2(n_1189),
.A3(n_1247),
.B(n_1149),
.Y(n_1312)
);

O2A1O1Ixp33_ASAP7_75t_L g1313 ( 
.A1(n_1210),
.A2(n_1160),
.B(n_1147),
.C(n_1203),
.Y(n_1313)
);

OAI22xp33_ASAP7_75t_L g1314 ( 
.A1(n_1119),
.A2(n_1103),
.B1(n_1153),
.B2(n_1228),
.Y(n_1314)
);

AOI21xp5_ASAP7_75t_L g1315 ( 
.A1(n_1179),
.A2(n_1103),
.B(n_1102),
.Y(n_1315)
);

A2O1A1Ixp33_ASAP7_75t_L g1316 ( 
.A1(n_1105),
.A2(n_1102),
.B(n_1248),
.C(n_1244),
.Y(n_1316)
);

AND2x4_ASAP7_75t_L g1317 ( 
.A(n_1129),
.B(n_1128),
.Y(n_1317)
);

INVx2_ASAP7_75t_SL g1318 ( 
.A(n_1223),
.Y(n_1318)
);

AO32x2_ASAP7_75t_L g1319 ( 
.A1(n_1155),
.A2(n_1186),
.A3(n_1218),
.B1(n_1225),
.B2(n_1119),
.Y(n_1319)
);

BUFx10_ASAP7_75t_L g1320 ( 
.A(n_1106),
.Y(n_1320)
);

OAI21x1_ASAP7_75t_L g1321 ( 
.A1(n_1121),
.A2(n_1178),
.B(n_1158),
.Y(n_1321)
);

AND2x4_ASAP7_75t_L g1322 ( 
.A(n_1129),
.B(n_1128),
.Y(n_1322)
);

OA21x2_ASAP7_75t_L g1323 ( 
.A1(n_1105),
.A2(n_1174),
.B(n_1252),
.Y(n_1323)
);

INVx2_ASAP7_75t_L g1324 ( 
.A(n_1108),
.Y(n_1324)
);

OAI21xp5_ASAP7_75t_L g1325 ( 
.A1(n_1138),
.A2(n_1215),
.B(n_1229),
.Y(n_1325)
);

NAND2xp5_ASAP7_75t_L g1326 ( 
.A(n_1142),
.B(n_1100),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_L g1327 ( 
.A(n_1126),
.B(n_1226),
.Y(n_1327)
);

AOI22xp5_ASAP7_75t_L g1328 ( 
.A1(n_1229),
.A2(n_1235),
.B1(n_1156),
.B2(n_1182),
.Y(n_1328)
);

AO32x2_ASAP7_75t_L g1329 ( 
.A1(n_1155),
.A2(n_1186),
.A3(n_1236),
.B1(n_1173),
.B2(n_1257),
.Y(n_1329)
);

AO31x2_ASAP7_75t_L g1330 ( 
.A1(n_1116),
.A2(n_1117),
.A3(n_1233),
.B(n_1125),
.Y(n_1330)
);

OAI21x1_ASAP7_75t_L g1331 ( 
.A1(n_1190),
.A2(n_1141),
.B(n_1221),
.Y(n_1331)
);

NOR2xp33_ASAP7_75t_L g1332 ( 
.A(n_1227),
.B(n_1129),
.Y(n_1332)
);

O2A1O1Ixp33_ASAP7_75t_L g1333 ( 
.A1(n_1213),
.A2(n_1190),
.B(n_1130),
.C(n_1131),
.Y(n_1333)
);

O2A1O1Ixp33_ASAP7_75t_L g1334 ( 
.A1(n_1163),
.A2(n_1193),
.B(n_1187),
.C(n_1197),
.Y(n_1334)
);

BUFx12f_ASAP7_75t_L g1335 ( 
.A(n_1159),
.Y(n_1335)
);

AND2x2_ASAP7_75t_L g1336 ( 
.A(n_1186),
.B(n_1227),
.Y(n_1336)
);

OAI21x1_ASAP7_75t_L g1337 ( 
.A1(n_1221),
.A2(n_1207),
.B(n_1205),
.Y(n_1337)
);

OAI21xp33_ASAP7_75t_SL g1338 ( 
.A1(n_1252),
.A2(n_1164),
.B(n_1132),
.Y(n_1338)
);

NOR2xp33_ASAP7_75t_L g1339 ( 
.A(n_1227),
.B(n_1167),
.Y(n_1339)
);

A2O1A1Ixp33_ASAP7_75t_L g1340 ( 
.A1(n_1257),
.A2(n_1220),
.B(n_1184),
.C(n_1230),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1257),
.Y(n_1341)
);

INVxp67_ASAP7_75t_L g1342 ( 
.A(n_1159),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_SL g1343 ( 
.A(n_1167),
.B(n_1120),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_L g1344 ( 
.A(n_1167),
.B(n_1120),
.Y(n_1344)
);

AOI21xp5_ASAP7_75t_L g1345 ( 
.A1(n_1132),
.A2(n_1146),
.B(n_1152),
.Y(n_1345)
);

INVx1_ASAP7_75t_SL g1346 ( 
.A(n_1132),
.Y(n_1346)
);

OAI22x1_ASAP7_75t_L g1347 ( 
.A1(n_1146),
.A2(n_1152),
.B1(n_1184),
.B2(n_1220),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1146),
.Y(n_1348)
);

INVx2_ASAP7_75t_L g1349 ( 
.A(n_1152),
.Y(n_1349)
);

BUFx3_ASAP7_75t_L g1350 ( 
.A(n_1230),
.Y(n_1350)
);

OA21x2_ASAP7_75t_L g1351 ( 
.A1(n_1220),
.A2(n_1245),
.B(n_1240),
.Y(n_1351)
);

INVxp67_ASAP7_75t_L g1352 ( 
.A(n_1230),
.Y(n_1352)
);

NAND3xp33_ASAP7_75t_SL g1353 ( 
.A(n_1139),
.B(n_549),
.C(n_640),
.Y(n_1353)
);

AO31x2_ASAP7_75t_L g1354 ( 
.A1(n_1113),
.A2(n_1060),
.A3(n_1239),
.B(n_945),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_L g1355 ( 
.A(n_1112),
.B(n_755),
.Y(n_1355)
);

AOI21xp5_ASAP7_75t_L g1356 ( 
.A1(n_1256),
.A2(n_1098),
.B(n_1199),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_L g1357 ( 
.A(n_1112),
.B(n_755),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1104),
.Y(n_1358)
);

AO31x2_ASAP7_75t_L g1359 ( 
.A1(n_1113),
.A2(n_1060),
.A3(n_1239),
.B(n_945),
.Y(n_1359)
);

NOR2xp33_ASAP7_75t_L g1360 ( 
.A(n_1161),
.B(n_549),
.Y(n_1360)
);

AND2x4_ASAP7_75t_L g1361 ( 
.A(n_1129),
.B(n_915),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1104),
.Y(n_1362)
);

BUFx3_ASAP7_75t_L g1363 ( 
.A(n_1122),
.Y(n_1363)
);

AOI22xp33_ASAP7_75t_L g1364 ( 
.A1(n_1119),
.A2(n_749),
.B1(n_845),
.B2(n_1073),
.Y(n_1364)
);

NAND2xp33_ASAP7_75t_SL g1365 ( 
.A(n_1241),
.B(n_1106),
.Y(n_1365)
);

BUFx3_ASAP7_75t_L g1366 ( 
.A(n_1122),
.Y(n_1366)
);

OAI21xp5_ASAP7_75t_L g1367 ( 
.A1(n_1192),
.A2(n_1098),
.B(n_1001),
.Y(n_1367)
);

INVx1_ASAP7_75t_SL g1368 ( 
.A(n_1142),
.Y(n_1368)
);

OAI21x1_ASAP7_75t_L g1369 ( 
.A1(n_1240),
.A2(n_1245),
.B(n_1214),
.Y(n_1369)
);

AOI22xp5_ASAP7_75t_L g1370 ( 
.A1(n_1180),
.A2(n_1161),
.B1(n_963),
.B2(n_737),
.Y(n_1370)
);

INVx3_ASAP7_75t_L g1371 ( 
.A(n_1128),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1104),
.Y(n_1372)
);

NOR2xp33_ASAP7_75t_L g1373 ( 
.A(n_1161),
.B(n_549),
.Y(n_1373)
);

CKINVDCx5p33_ASAP7_75t_R g1374 ( 
.A(n_1144),
.Y(n_1374)
);

INVx4_ASAP7_75t_L g1375 ( 
.A(n_1122),
.Y(n_1375)
);

CKINVDCx5p33_ASAP7_75t_R g1376 ( 
.A(n_1144),
.Y(n_1376)
);

A2O1A1Ixp33_ASAP7_75t_L g1377 ( 
.A1(n_1161),
.A2(n_737),
.B(n_1043),
.C(n_739),
.Y(n_1377)
);

NAND3xp33_ASAP7_75t_L g1378 ( 
.A(n_1127),
.B(n_737),
.C(n_1161),
.Y(n_1378)
);

INVxp67_ASAP7_75t_L g1379 ( 
.A(n_1112),
.Y(n_1379)
);

INVx3_ASAP7_75t_L g1380 ( 
.A(n_1128),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_L g1381 ( 
.A(n_1112),
.B(n_755),
.Y(n_1381)
);

INVx4_ASAP7_75t_L g1382 ( 
.A(n_1122),
.Y(n_1382)
);

AOI21xp5_ASAP7_75t_L g1383 ( 
.A1(n_1256),
.A2(n_1098),
.B(n_1199),
.Y(n_1383)
);

O2A1O1Ixp33_ASAP7_75t_SL g1384 ( 
.A1(n_1135),
.A2(n_1043),
.B(n_1166),
.C(n_1165),
.Y(n_1384)
);

AND2x2_ASAP7_75t_L g1385 ( 
.A(n_1112),
.B(n_755),
.Y(n_1385)
);

INVx2_ASAP7_75t_L g1386 ( 
.A(n_1099),
.Y(n_1386)
);

AOI21xp5_ASAP7_75t_L g1387 ( 
.A1(n_1256),
.A2(n_1098),
.B(n_1199),
.Y(n_1387)
);

AO21x1_ASAP7_75t_L g1388 ( 
.A1(n_1098),
.A2(n_1234),
.B(n_1192),
.Y(n_1388)
);

A2O1A1Ixp33_ASAP7_75t_L g1389 ( 
.A1(n_1161),
.A2(n_737),
.B(n_1043),
.C(n_739),
.Y(n_1389)
);

A2O1A1Ixp33_ASAP7_75t_L g1390 ( 
.A1(n_1161),
.A2(n_737),
.B(n_1043),
.C(n_739),
.Y(n_1390)
);

O2A1O1Ixp33_ASAP7_75t_SL g1391 ( 
.A1(n_1135),
.A2(n_1043),
.B(n_1166),
.C(n_1165),
.Y(n_1391)
);

OAI21x1_ASAP7_75t_L g1392 ( 
.A1(n_1240),
.A2(n_1245),
.B(n_1214),
.Y(n_1392)
);

NAND2xp5_ASAP7_75t_L g1393 ( 
.A(n_1112),
.B(n_755),
.Y(n_1393)
);

OAI21x1_ASAP7_75t_L g1394 ( 
.A1(n_1240),
.A2(n_1245),
.B(n_1214),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_SL g1395 ( 
.A(n_1241),
.B(n_1228),
.Y(n_1395)
);

AND2x2_ASAP7_75t_L g1396 ( 
.A(n_1112),
.B(n_755),
.Y(n_1396)
);

NAND2xp5_ASAP7_75t_L g1397 ( 
.A(n_1112),
.B(n_755),
.Y(n_1397)
);

AO22x2_ASAP7_75t_L g1398 ( 
.A1(n_1111),
.A2(n_1114),
.B1(n_1118),
.B2(n_1171),
.Y(n_1398)
);

HB1xp67_ASAP7_75t_L g1399 ( 
.A(n_1162),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1104),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_L g1401 ( 
.A(n_1216),
.B(n_1219),
.Y(n_1401)
);

BUFx6f_ASAP7_75t_L g1402 ( 
.A(n_1159),
.Y(n_1402)
);

OAI21xp5_ASAP7_75t_L g1403 ( 
.A1(n_1192),
.A2(n_1098),
.B(n_1001),
.Y(n_1403)
);

OR2x6_ASAP7_75t_SL g1404 ( 
.A(n_1241),
.B(n_725),
.Y(n_1404)
);

A2O1A1Ixp33_ASAP7_75t_L g1405 ( 
.A1(n_1161),
.A2(n_737),
.B(n_1043),
.C(n_739),
.Y(n_1405)
);

AND2x2_ASAP7_75t_SL g1406 ( 
.A(n_1103),
.B(n_631),
.Y(n_1406)
);

BUFx12f_ASAP7_75t_L g1407 ( 
.A(n_1106),
.Y(n_1407)
);

O2A1O1Ixp33_ASAP7_75t_L g1408 ( 
.A1(n_1161),
.A2(n_737),
.B(n_609),
.C(n_595),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1104),
.Y(n_1409)
);

OAI21x1_ASAP7_75t_L g1410 ( 
.A1(n_1240),
.A2(n_1245),
.B(n_1214),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_L g1411 ( 
.A(n_1112),
.B(n_755),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_SL g1412 ( 
.A(n_1241),
.B(n_1228),
.Y(n_1412)
);

OAI21x1_ASAP7_75t_L g1413 ( 
.A1(n_1240),
.A2(n_1245),
.B(n_1214),
.Y(n_1413)
);

AO31x2_ASAP7_75t_L g1414 ( 
.A1(n_1113),
.A2(n_1060),
.A3(n_1239),
.B(n_945),
.Y(n_1414)
);

NOR2xp67_ASAP7_75t_SL g1415 ( 
.A(n_1122),
.B(n_801),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_L g1416 ( 
.A(n_1112),
.B(n_755),
.Y(n_1416)
);

A2O1A1Ixp33_ASAP7_75t_L g1417 ( 
.A1(n_1161),
.A2(n_737),
.B(n_1043),
.C(n_739),
.Y(n_1417)
);

O2A1O1Ixp33_ASAP7_75t_L g1418 ( 
.A1(n_1161),
.A2(n_737),
.B(n_609),
.C(n_595),
.Y(n_1418)
);

AND2x4_ASAP7_75t_L g1419 ( 
.A(n_1129),
.B(n_915),
.Y(n_1419)
);

O2A1O1Ixp33_ASAP7_75t_L g1420 ( 
.A1(n_1161),
.A2(n_737),
.B(n_609),
.C(n_595),
.Y(n_1420)
);

OAI21xp33_ASAP7_75t_L g1421 ( 
.A1(n_1204),
.A2(n_575),
.B(n_1019),
.Y(n_1421)
);

OAI21x1_ASAP7_75t_L g1422 ( 
.A1(n_1240),
.A2(n_1245),
.B(n_1214),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1104),
.Y(n_1423)
);

BUFx8_ASAP7_75t_L g1424 ( 
.A(n_1122),
.Y(n_1424)
);

INVx1_ASAP7_75t_SL g1425 ( 
.A(n_1142),
.Y(n_1425)
);

AOI21xp5_ASAP7_75t_L g1426 ( 
.A1(n_1256),
.A2(n_1098),
.B(n_1199),
.Y(n_1426)
);

NAND2x1p5_ASAP7_75t_L g1427 ( 
.A(n_1122),
.B(n_998),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1261),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1267),
.Y(n_1429)
);

OAI22xp5_ASAP7_75t_L g1430 ( 
.A1(n_1370),
.A2(n_1289),
.B1(n_1378),
.B2(n_1285),
.Y(n_1430)
);

BUFx12f_ASAP7_75t_L g1431 ( 
.A(n_1424),
.Y(n_1431)
);

CKINVDCx11_ASAP7_75t_R g1432 ( 
.A(n_1404),
.Y(n_1432)
);

BUFx6f_ASAP7_75t_L g1433 ( 
.A(n_1263),
.Y(n_1433)
);

OAI22xp5_ASAP7_75t_L g1434 ( 
.A1(n_1370),
.A2(n_1289),
.B1(n_1378),
.B2(n_1285),
.Y(n_1434)
);

INVx4_ASAP7_75t_L g1435 ( 
.A(n_1263),
.Y(n_1435)
);

AOI22xp33_ASAP7_75t_L g1436 ( 
.A1(n_1364),
.A2(n_1421),
.B1(n_1300),
.B2(n_1398),
.Y(n_1436)
);

INVx1_ASAP7_75t_SL g1437 ( 
.A(n_1368),
.Y(n_1437)
);

INVx6_ASAP7_75t_L g1438 ( 
.A(n_1263),
.Y(n_1438)
);

OAI22xp33_ASAP7_75t_L g1439 ( 
.A1(n_1355),
.A2(n_1357),
.B1(n_1397),
.B2(n_1393),
.Y(n_1439)
);

AOI22xp33_ASAP7_75t_SL g1440 ( 
.A1(n_1300),
.A2(n_1406),
.B1(n_1326),
.B2(n_1398),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1277),
.Y(n_1441)
);

AOI22xp33_ASAP7_75t_SL g1442 ( 
.A1(n_1336),
.A2(n_1299),
.B1(n_1401),
.B2(n_1287),
.Y(n_1442)
);

BUFx12f_ASAP7_75t_L g1443 ( 
.A(n_1424),
.Y(n_1443)
);

AOI22xp33_ASAP7_75t_L g1444 ( 
.A1(n_1421),
.A2(n_1353),
.B1(n_1296),
.B2(n_1314),
.Y(n_1444)
);

AOI22xp33_ASAP7_75t_L g1445 ( 
.A1(n_1388),
.A2(n_1271),
.B1(n_1396),
.B2(n_1385),
.Y(n_1445)
);

BUFx6f_ASAP7_75t_L g1446 ( 
.A(n_1335),
.Y(n_1446)
);

CKINVDCx11_ASAP7_75t_R g1447 ( 
.A(n_1407),
.Y(n_1447)
);

AOI22xp33_ASAP7_75t_SL g1448 ( 
.A1(n_1401),
.A2(n_1293),
.B1(n_1329),
.B2(n_1319),
.Y(n_1448)
);

AOI22xp33_ASAP7_75t_L g1449 ( 
.A1(n_1379),
.A2(n_1293),
.B1(n_1290),
.B2(n_1373),
.Y(n_1449)
);

OAI22xp5_ASAP7_75t_L g1450 ( 
.A1(n_1377),
.A2(n_1405),
.B1(n_1417),
.B2(n_1390),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1295),
.Y(n_1451)
);

NOR2xp33_ASAP7_75t_L g1452 ( 
.A(n_1360),
.B(n_1395),
.Y(n_1452)
);

BUFx8_ASAP7_75t_L g1453 ( 
.A(n_1305),
.Y(n_1453)
);

BUFx6f_ASAP7_75t_L g1454 ( 
.A(n_1363),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1303),
.Y(n_1455)
);

NAND2xp33_ASAP7_75t_SL g1456 ( 
.A(n_1415),
.B(n_1412),
.Y(n_1456)
);

AOI22xp33_ASAP7_75t_L g1457 ( 
.A1(n_1381),
.A2(n_1411),
.B1(n_1416),
.B2(n_1286),
.Y(n_1457)
);

OAI21xp5_ASAP7_75t_L g1458 ( 
.A1(n_1389),
.A2(n_1292),
.B(n_1279),
.Y(n_1458)
);

INVx4_ASAP7_75t_L g1459 ( 
.A(n_1427),
.Y(n_1459)
);

BUFx6f_ASAP7_75t_L g1460 ( 
.A(n_1366),
.Y(n_1460)
);

AOI22xp33_ASAP7_75t_SL g1461 ( 
.A1(n_1329),
.A2(n_1319),
.B1(n_1281),
.B2(n_1323),
.Y(n_1461)
);

CKINVDCx11_ASAP7_75t_R g1462 ( 
.A(n_1320),
.Y(n_1462)
);

OAI22xp33_ASAP7_75t_L g1463 ( 
.A1(n_1328),
.A2(n_1280),
.B1(n_1284),
.B2(n_1327),
.Y(n_1463)
);

AOI22xp33_ASAP7_75t_L g1464 ( 
.A1(n_1324),
.A2(n_1386),
.B1(n_1283),
.B2(n_1425),
.Y(n_1464)
);

AOI22xp33_ASAP7_75t_L g1465 ( 
.A1(n_1368),
.A2(n_1425),
.B1(n_1328),
.B2(n_1274),
.Y(n_1465)
);

INVx11_ASAP7_75t_L g1466 ( 
.A(n_1365),
.Y(n_1466)
);

AND2x2_ASAP7_75t_L g1467 ( 
.A(n_1301),
.B(n_1399),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1358),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1362),
.Y(n_1469)
);

AOI22xp33_ASAP7_75t_L g1470 ( 
.A1(n_1311),
.A2(n_1423),
.B1(n_1400),
.B2(n_1372),
.Y(n_1470)
);

OAI22xp5_ASAP7_75t_L g1471 ( 
.A1(n_1298),
.A2(n_1294),
.B1(n_1367),
.B2(n_1403),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1409),
.Y(n_1472)
);

AOI22xp33_ASAP7_75t_L g1473 ( 
.A1(n_1302),
.A2(n_1341),
.B1(n_1306),
.B2(n_1282),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1330),
.Y(n_1474)
);

BUFx8_ASAP7_75t_SL g1475 ( 
.A(n_1374),
.Y(n_1475)
);

INVx6_ASAP7_75t_L g1476 ( 
.A(n_1270),
.Y(n_1476)
);

INVx1_ASAP7_75t_SL g1477 ( 
.A(n_1344),
.Y(n_1477)
);

NAND2x1p5_ASAP7_75t_L g1478 ( 
.A(n_1371),
.B(n_1380),
.Y(n_1478)
);

OR2x2_ASAP7_75t_L g1479 ( 
.A(n_1306),
.B(n_1342),
.Y(n_1479)
);

AOI22xp33_ASAP7_75t_L g1480 ( 
.A1(n_1317),
.A2(n_1322),
.B1(n_1325),
.B2(n_1419),
.Y(n_1480)
);

BUFx6f_ASAP7_75t_L g1481 ( 
.A(n_1307),
.Y(n_1481)
);

BUFx12f_ASAP7_75t_L g1482 ( 
.A(n_1376),
.Y(n_1482)
);

INVx6_ASAP7_75t_L g1483 ( 
.A(n_1270),
.Y(n_1483)
);

AOI22xp33_ASAP7_75t_SL g1484 ( 
.A1(n_1329),
.A2(n_1319),
.B1(n_1323),
.B2(n_1338),
.Y(n_1484)
);

AOI22xp33_ASAP7_75t_SL g1485 ( 
.A1(n_1367),
.A2(n_1403),
.B1(n_1322),
.B2(n_1317),
.Y(n_1485)
);

AOI22xp33_ASAP7_75t_L g1486 ( 
.A1(n_1325),
.A2(n_1361),
.B1(n_1419),
.B2(n_1338),
.Y(n_1486)
);

INVx4_ASAP7_75t_L g1487 ( 
.A(n_1375),
.Y(n_1487)
);

CKINVDCx6p67_ASAP7_75t_R g1488 ( 
.A(n_1375),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1334),
.Y(n_1489)
);

CKINVDCx11_ASAP7_75t_R g1490 ( 
.A(n_1320),
.Y(n_1490)
);

BUFx4f_ASAP7_75t_L g1491 ( 
.A(n_1361),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_L g1492 ( 
.A(n_1291),
.B(n_1268),
.Y(n_1492)
);

AOI22xp33_ASAP7_75t_L g1493 ( 
.A1(n_1350),
.A2(n_1371),
.B1(n_1380),
.B2(n_1266),
.Y(n_1493)
);

INVx8_ASAP7_75t_L g1494 ( 
.A(n_1402),
.Y(n_1494)
);

AOI22xp33_ASAP7_75t_L g1495 ( 
.A1(n_1266),
.A2(n_1332),
.B1(n_1402),
.B2(n_1339),
.Y(n_1495)
);

AOI22xp33_ASAP7_75t_SL g1496 ( 
.A1(n_1315),
.A2(n_1402),
.B1(n_1313),
.B2(n_1308),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_L g1497 ( 
.A(n_1268),
.B(n_1316),
.Y(n_1497)
);

INVx3_ASAP7_75t_SL g1498 ( 
.A(n_1382),
.Y(n_1498)
);

AOI22xp5_ASAP7_75t_SL g1499 ( 
.A1(n_1318),
.A2(n_1382),
.B1(n_1352),
.B2(n_1347),
.Y(n_1499)
);

NOR2x1_ASAP7_75t_SL g1500 ( 
.A(n_1343),
.B(n_1348),
.Y(n_1500)
);

AOI22xp33_ASAP7_75t_L g1501 ( 
.A1(n_1276),
.A2(n_1309),
.B1(n_1337),
.B2(n_1349),
.Y(n_1501)
);

AOI22xp33_ASAP7_75t_SL g1502 ( 
.A1(n_1275),
.A2(n_1297),
.B1(n_1387),
.B2(n_1356),
.Y(n_1502)
);

BUFx8_ASAP7_75t_L g1503 ( 
.A(n_1408),
.Y(n_1503)
);

BUFx6f_ASAP7_75t_L g1504 ( 
.A(n_1331),
.Y(n_1504)
);

AOI22xp33_ASAP7_75t_SL g1505 ( 
.A1(n_1383),
.A2(n_1426),
.B1(n_1391),
.B2(n_1384),
.Y(n_1505)
);

INVx2_ASAP7_75t_SL g1506 ( 
.A(n_1346),
.Y(n_1506)
);

NAND2xp5_ASAP7_75t_L g1507 ( 
.A(n_1268),
.B(n_1264),
.Y(n_1507)
);

BUFx3_ASAP7_75t_L g1508 ( 
.A(n_1346),
.Y(n_1508)
);

OAI22xp5_ASAP7_75t_L g1509 ( 
.A1(n_1418),
.A2(n_1420),
.B1(n_1304),
.B2(n_1269),
.Y(n_1509)
);

OAI22xp5_ASAP7_75t_L g1510 ( 
.A1(n_1310),
.A2(n_1264),
.B1(n_1272),
.B2(n_1340),
.Y(n_1510)
);

AOI22xp33_ASAP7_75t_L g1511 ( 
.A1(n_1262),
.A2(n_1260),
.B1(n_1345),
.B2(n_1351),
.Y(n_1511)
);

AOI22xp33_ASAP7_75t_L g1512 ( 
.A1(n_1262),
.A2(n_1351),
.B1(n_1265),
.B2(n_1321),
.Y(n_1512)
);

INVx6_ASAP7_75t_L g1513 ( 
.A(n_1333),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1354),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1354),
.Y(n_1515)
);

BUFx4f_ASAP7_75t_SL g1516 ( 
.A(n_1273),
.Y(n_1516)
);

INVx4_ASAP7_75t_L g1517 ( 
.A(n_1273),
.Y(n_1517)
);

NAND2xp5_ASAP7_75t_L g1518 ( 
.A(n_1354),
.B(n_1359),
.Y(n_1518)
);

AOI22xp33_ASAP7_75t_SL g1519 ( 
.A1(n_1312),
.A2(n_1414),
.B1(n_1359),
.B2(n_1422),
.Y(n_1519)
);

OAI22xp5_ASAP7_75t_L g1520 ( 
.A1(n_1278),
.A2(n_1273),
.B1(n_1312),
.B2(n_1288),
.Y(n_1520)
);

BUFx8_ASAP7_75t_SL g1521 ( 
.A(n_1278),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_L g1522 ( 
.A(n_1414),
.B(n_1278),
.Y(n_1522)
);

OAI22xp5_ASAP7_75t_L g1523 ( 
.A1(n_1312),
.A2(n_1288),
.B1(n_1369),
.B2(n_1392),
.Y(n_1523)
);

INVx6_ASAP7_75t_L g1524 ( 
.A(n_1288),
.Y(n_1524)
);

AOI22xp33_ASAP7_75t_L g1525 ( 
.A1(n_1394),
.A2(n_749),
.B1(n_1119),
.B2(n_1364),
.Y(n_1525)
);

BUFx2_ASAP7_75t_L g1526 ( 
.A(n_1410),
.Y(n_1526)
);

AOI22xp33_ASAP7_75t_L g1527 ( 
.A1(n_1413),
.A2(n_749),
.B1(n_1119),
.B2(n_1364),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1261),
.Y(n_1528)
);

OAI22xp33_ASAP7_75t_L g1529 ( 
.A1(n_1289),
.A2(n_1370),
.B1(n_1028),
.B2(n_1030),
.Y(n_1529)
);

INVxp67_ASAP7_75t_SL g1530 ( 
.A(n_1399),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1261),
.Y(n_1531)
);

AOI22xp33_ASAP7_75t_SL g1532 ( 
.A1(n_1300),
.A2(n_749),
.B1(n_1119),
.B2(n_408),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_L g1533 ( 
.A(n_1401),
.B(n_1306),
.Y(n_1533)
);

CKINVDCx5p33_ASAP7_75t_R g1534 ( 
.A(n_1424),
.Y(n_1534)
);

INVx3_ASAP7_75t_SL g1535 ( 
.A(n_1374),
.Y(n_1535)
);

INVx1_ASAP7_75t_SL g1536 ( 
.A(n_1368),
.Y(n_1536)
);

AOI22xp33_ASAP7_75t_L g1537 ( 
.A1(n_1364),
.A2(n_749),
.B1(n_1119),
.B2(n_955),
.Y(n_1537)
);

CKINVDCx11_ASAP7_75t_R g1538 ( 
.A(n_1404),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1261),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1261),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1261),
.Y(n_1541)
);

CKINVDCx20_ASAP7_75t_R g1542 ( 
.A(n_1424),
.Y(n_1542)
);

AOI22xp33_ASAP7_75t_L g1543 ( 
.A1(n_1364),
.A2(n_749),
.B1(n_1119),
.B2(n_955),
.Y(n_1543)
);

AOI22xp33_ASAP7_75t_SL g1544 ( 
.A1(n_1300),
.A2(n_749),
.B1(n_1119),
.B2(n_408),
.Y(n_1544)
);

CKINVDCx20_ASAP7_75t_R g1545 ( 
.A(n_1424),
.Y(n_1545)
);

NAND2xp5_ASAP7_75t_L g1546 ( 
.A(n_1401),
.B(n_1306),
.Y(n_1546)
);

INVx2_ASAP7_75t_SL g1547 ( 
.A(n_1424),
.Y(n_1547)
);

AOI22xp33_ASAP7_75t_L g1548 ( 
.A1(n_1364),
.A2(n_749),
.B1(n_1119),
.B2(n_955),
.Y(n_1548)
);

AOI22xp33_ASAP7_75t_L g1549 ( 
.A1(n_1364),
.A2(n_749),
.B1(n_1119),
.B2(n_955),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1261),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1261),
.Y(n_1551)
);

OAI22xp5_ASAP7_75t_L g1552 ( 
.A1(n_1370),
.A2(n_1289),
.B1(n_1378),
.B2(n_1285),
.Y(n_1552)
);

CKINVDCx11_ASAP7_75t_R g1553 ( 
.A(n_1404),
.Y(n_1553)
);

CKINVDCx5p33_ASAP7_75t_R g1554 ( 
.A(n_1424),
.Y(n_1554)
);

OAI22xp33_ASAP7_75t_L g1555 ( 
.A1(n_1289),
.A2(n_1370),
.B1(n_1028),
.B2(n_1030),
.Y(n_1555)
);

CKINVDCx20_ASAP7_75t_R g1556 ( 
.A(n_1424),
.Y(n_1556)
);

BUFx2_ASAP7_75t_SL g1557 ( 
.A(n_1270),
.Y(n_1557)
);

INVx4_ASAP7_75t_L g1558 ( 
.A(n_1263),
.Y(n_1558)
);

BUFx8_ASAP7_75t_L g1559 ( 
.A(n_1407),
.Y(n_1559)
);

HB1xp67_ASAP7_75t_L g1560 ( 
.A(n_1399),
.Y(n_1560)
);

OAI21xp5_ASAP7_75t_SL g1561 ( 
.A1(n_1289),
.A2(n_1285),
.B(n_1370),
.Y(n_1561)
);

INVx1_ASAP7_75t_SL g1562 ( 
.A(n_1368),
.Y(n_1562)
);

BUFx6f_ASAP7_75t_L g1563 ( 
.A(n_1263),
.Y(n_1563)
);

CKINVDCx11_ASAP7_75t_R g1564 ( 
.A(n_1404),
.Y(n_1564)
);

OAI22xp5_ASAP7_75t_L g1565 ( 
.A1(n_1370),
.A2(n_1289),
.B1(n_1378),
.B2(n_1285),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1261),
.Y(n_1566)
);

INVx3_ASAP7_75t_L g1567 ( 
.A(n_1263),
.Y(n_1567)
);

BUFx6f_ASAP7_75t_L g1568 ( 
.A(n_1263),
.Y(n_1568)
);

AOI22xp33_ASAP7_75t_L g1569 ( 
.A1(n_1364),
.A2(n_749),
.B1(n_1119),
.B2(n_955),
.Y(n_1569)
);

AOI22xp33_ASAP7_75t_SL g1570 ( 
.A1(n_1300),
.A2(n_749),
.B1(n_1119),
.B2(n_408),
.Y(n_1570)
);

AOI22xp5_ASAP7_75t_L g1571 ( 
.A1(n_1289),
.A2(n_1421),
.B1(n_697),
.B2(n_640),
.Y(n_1571)
);

INVx4_ASAP7_75t_L g1572 ( 
.A(n_1263),
.Y(n_1572)
);

BUFx2_ASAP7_75t_SL g1573 ( 
.A(n_1270),
.Y(n_1573)
);

BUFx2_ASAP7_75t_L g1574 ( 
.A(n_1365),
.Y(n_1574)
);

CKINVDCx11_ASAP7_75t_R g1575 ( 
.A(n_1404),
.Y(n_1575)
);

OAI22xp5_ASAP7_75t_L g1576 ( 
.A1(n_1370),
.A2(n_1289),
.B1(n_1378),
.B2(n_1285),
.Y(n_1576)
);

BUFx3_ASAP7_75t_L g1577 ( 
.A(n_1424),
.Y(n_1577)
);

AOI22xp33_ASAP7_75t_SL g1578 ( 
.A1(n_1300),
.A2(n_749),
.B1(n_1119),
.B2(n_408),
.Y(n_1578)
);

INVx8_ASAP7_75t_L g1579 ( 
.A(n_1263),
.Y(n_1579)
);

CKINVDCx5p33_ASAP7_75t_R g1580 ( 
.A(n_1424),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1474),
.Y(n_1581)
);

NAND2x1p5_ASAP7_75t_L g1582 ( 
.A(n_1491),
.B(n_1479),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_L g1583 ( 
.A(n_1437),
.B(n_1536),
.Y(n_1583)
);

AO21x2_ASAP7_75t_L g1584 ( 
.A1(n_1518),
.A2(n_1520),
.B(n_1522),
.Y(n_1584)
);

O2A1O1Ixp5_ASAP7_75t_L g1585 ( 
.A1(n_1430),
.A2(n_1552),
.B(n_1565),
.C(n_1434),
.Y(n_1585)
);

INVx2_ASAP7_75t_SL g1586 ( 
.A(n_1560),
.Y(n_1586)
);

OAI21x1_ASAP7_75t_L g1587 ( 
.A1(n_1523),
.A2(n_1510),
.B(n_1512),
.Y(n_1587)
);

AND2x4_ASAP7_75t_L g1588 ( 
.A(n_1504),
.B(n_1497),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1497),
.B(n_1461),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1514),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1515),
.Y(n_1591)
);

CKINVDCx16_ASAP7_75t_R g1592 ( 
.A(n_1431),
.Y(n_1592)
);

OAI21x1_ASAP7_75t_L g1593 ( 
.A1(n_1523),
.A2(n_1510),
.B(n_1520),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1428),
.Y(n_1594)
);

OR2x2_ASAP7_75t_L g1595 ( 
.A(n_1437),
.B(n_1536),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1429),
.Y(n_1596)
);

INVxp33_ASAP7_75t_SL g1597 ( 
.A(n_1534),
.Y(n_1597)
);

OR2x2_ASAP7_75t_L g1598 ( 
.A(n_1562),
.B(n_1507),
.Y(n_1598)
);

BUFx6f_ASAP7_75t_L g1599 ( 
.A(n_1491),
.Y(n_1599)
);

HB1xp67_ASAP7_75t_L g1600 ( 
.A(n_1530),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_L g1601 ( 
.A(n_1562),
.B(n_1533),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1441),
.Y(n_1602)
);

AOI22xp33_ASAP7_75t_L g1603 ( 
.A1(n_1532),
.A2(n_1544),
.B1(n_1578),
.B2(n_1570),
.Y(n_1603)
);

AO21x2_ASAP7_75t_L g1604 ( 
.A1(n_1518),
.A2(n_1522),
.B(n_1507),
.Y(n_1604)
);

INVx4_ASAP7_75t_L g1605 ( 
.A(n_1466),
.Y(n_1605)
);

AND2x2_ASAP7_75t_L g1606 ( 
.A(n_1448),
.B(n_1451),
.Y(n_1606)
);

OAI21x1_ASAP7_75t_L g1607 ( 
.A1(n_1501),
.A2(n_1511),
.B(n_1458),
.Y(n_1607)
);

CKINVDCx11_ASAP7_75t_R g1608 ( 
.A(n_1542),
.Y(n_1608)
);

AO21x2_ASAP7_75t_L g1609 ( 
.A1(n_1492),
.A2(n_1471),
.B(n_1458),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1455),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1468),
.Y(n_1611)
);

OAI21x1_ASAP7_75t_L g1612 ( 
.A1(n_1492),
.A2(n_1471),
.B(n_1450),
.Y(n_1612)
);

INVx2_ASAP7_75t_L g1613 ( 
.A(n_1469),
.Y(n_1613)
);

AOI22xp33_ASAP7_75t_L g1614 ( 
.A1(n_1537),
.A2(n_1569),
.B1(n_1543),
.B2(n_1549),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_1472),
.B(n_1528),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1531),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1539),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1540),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_L g1619 ( 
.A(n_1533),
.B(n_1546),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1541),
.Y(n_1620)
);

HB1xp67_ASAP7_75t_L g1621 ( 
.A(n_1467),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1550),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1551),
.Y(n_1623)
);

INVx2_ASAP7_75t_L g1624 ( 
.A(n_1566),
.Y(n_1624)
);

O2A1O1Ixp5_ASAP7_75t_L g1625 ( 
.A1(n_1430),
.A2(n_1552),
.B(n_1576),
.C(n_1434),
.Y(n_1625)
);

INVx3_ASAP7_75t_L g1626 ( 
.A(n_1524),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1546),
.Y(n_1627)
);

AO21x2_ASAP7_75t_L g1628 ( 
.A1(n_1565),
.A2(n_1576),
.B(n_1529),
.Y(n_1628)
);

BUFx3_ASAP7_75t_L g1629 ( 
.A(n_1476),
.Y(n_1629)
);

OA21x2_ASAP7_75t_L g1630 ( 
.A1(n_1526),
.A2(n_1464),
.B(n_1561),
.Y(n_1630)
);

OAI21x1_ASAP7_75t_L g1631 ( 
.A1(n_1450),
.A2(n_1509),
.B(n_1493),
.Y(n_1631)
);

AND2x2_ASAP7_75t_L g1632 ( 
.A(n_1485),
.B(n_1442),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1516),
.Y(n_1633)
);

NAND2xp5_ASAP7_75t_L g1634 ( 
.A(n_1449),
.B(n_1439),
.Y(n_1634)
);

INVx2_ASAP7_75t_SL g1635 ( 
.A(n_1504),
.Y(n_1635)
);

INVxp67_ASAP7_75t_SL g1636 ( 
.A(n_1519),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_L g1637 ( 
.A(n_1457),
.B(n_1470),
.Y(n_1637)
);

OAI21x1_ASAP7_75t_SL g1638 ( 
.A1(n_1509),
.A2(n_1500),
.B(n_1444),
.Y(n_1638)
);

CKINVDCx20_ASAP7_75t_R g1639 ( 
.A(n_1545),
.Y(n_1639)
);

INVx3_ASAP7_75t_L g1640 ( 
.A(n_1517),
.Y(n_1640)
);

AND2x2_ASAP7_75t_L g1641 ( 
.A(n_1485),
.B(n_1484),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1504),
.Y(n_1642)
);

HB1xp67_ASAP7_75t_L g1643 ( 
.A(n_1477),
.Y(n_1643)
);

AND2x2_ASAP7_75t_L g1644 ( 
.A(n_1445),
.B(n_1517),
.Y(n_1644)
);

OR2x2_ASAP7_75t_L g1645 ( 
.A(n_1477),
.B(n_1436),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1521),
.Y(n_1646)
);

AND2x2_ASAP7_75t_L g1647 ( 
.A(n_1473),
.B(n_1505),
.Y(n_1647)
);

OR2x2_ASAP7_75t_L g1648 ( 
.A(n_1465),
.B(n_1463),
.Y(n_1648)
);

INVx2_ASAP7_75t_L g1649 ( 
.A(n_1489),
.Y(n_1649)
);

OR2x2_ASAP7_75t_L g1650 ( 
.A(n_1486),
.B(n_1571),
.Y(n_1650)
);

INVxp33_ASAP7_75t_L g1651 ( 
.A(n_1454),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1502),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1513),
.Y(n_1653)
);

AND2x2_ASAP7_75t_L g1654 ( 
.A(n_1496),
.B(n_1480),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1513),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1440),
.B(n_1478),
.Y(n_1656)
);

INVx2_ASAP7_75t_L g1657 ( 
.A(n_1513),
.Y(n_1657)
);

HB1xp67_ASAP7_75t_L g1658 ( 
.A(n_1508),
.Y(n_1658)
);

BUFx2_ASAP7_75t_L g1659 ( 
.A(n_1574),
.Y(n_1659)
);

AO21x2_ASAP7_75t_L g1660 ( 
.A1(n_1555),
.A2(n_1495),
.B(n_1503),
.Y(n_1660)
);

INVx2_ASAP7_75t_L g1661 ( 
.A(n_1506),
.Y(n_1661)
);

BUFx8_ASAP7_75t_L g1662 ( 
.A(n_1443),
.Y(n_1662)
);

AOI221xp5_ASAP7_75t_L g1663 ( 
.A1(n_1525),
.A2(n_1527),
.B1(n_1548),
.B2(n_1456),
.C(n_1452),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1499),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1478),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1503),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1481),
.Y(n_1667)
);

NOR2x1_ASAP7_75t_L g1668 ( 
.A(n_1487),
.B(n_1459),
.Y(n_1668)
);

INVx4_ASAP7_75t_SL g1669 ( 
.A(n_1438),
.Y(n_1669)
);

OAI21xp33_ASAP7_75t_SL g1670 ( 
.A1(n_1487),
.A2(n_1572),
.B(n_1558),
.Y(n_1670)
);

AOI22xp5_ASAP7_75t_L g1671 ( 
.A1(n_1432),
.A2(n_1538),
.B1(n_1564),
.B2(n_1575),
.Y(n_1671)
);

OR2x6_ASAP7_75t_L g1672 ( 
.A(n_1494),
.B(n_1579),
.Y(n_1672)
);

AND2x2_ASAP7_75t_L g1673 ( 
.A(n_1557),
.B(n_1573),
.Y(n_1673)
);

AND2x2_ASAP7_75t_L g1674 ( 
.A(n_1483),
.B(n_1498),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1567),
.Y(n_1675)
);

HB1xp67_ASAP7_75t_L g1676 ( 
.A(n_1454),
.Y(n_1676)
);

BUFx2_ASAP7_75t_L g1677 ( 
.A(n_1567),
.Y(n_1677)
);

BUFx2_ASAP7_75t_L g1678 ( 
.A(n_1488),
.Y(n_1678)
);

HB1xp67_ASAP7_75t_L g1679 ( 
.A(n_1460),
.Y(n_1679)
);

INVx2_ASAP7_75t_L g1680 ( 
.A(n_1460),
.Y(n_1680)
);

BUFx6f_ASAP7_75t_L g1681 ( 
.A(n_1433),
.Y(n_1681)
);

INVx1_ASAP7_75t_SL g1682 ( 
.A(n_1462),
.Y(n_1682)
);

INVx2_ASAP7_75t_L g1683 ( 
.A(n_1459),
.Y(n_1683)
);

OR2x6_ASAP7_75t_L g1684 ( 
.A(n_1579),
.B(n_1446),
.Y(n_1684)
);

AND2x2_ASAP7_75t_L g1685 ( 
.A(n_1553),
.B(n_1547),
.Y(n_1685)
);

AOI22xp33_ASAP7_75t_SL g1686 ( 
.A1(n_1446),
.A2(n_1559),
.B1(n_1577),
.B2(n_1453),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1433),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1563),
.Y(n_1688)
);

AO21x1_ASAP7_75t_SL g1689 ( 
.A1(n_1579),
.A2(n_1435),
.B(n_1558),
.Y(n_1689)
);

BUFx2_ASAP7_75t_L g1690 ( 
.A(n_1659),
.Y(n_1690)
);

AND2x2_ASAP7_75t_L g1691 ( 
.A(n_1609),
.B(n_1535),
.Y(n_1691)
);

AOI21xp5_ASAP7_75t_L g1692 ( 
.A1(n_1585),
.A2(n_1435),
.B(n_1572),
.Y(n_1692)
);

A2O1A1Ixp33_ASAP7_75t_L g1693 ( 
.A1(n_1625),
.A2(n_1568),
.B(n_1580),
.C(n_1554),
.Y(n_1693)
);

AND2x2_ASAP7_75t_L g1694 ( 
.A(n_1621),
.B(n_1490),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1594),
.Y(n_1695)
);

AND2x2_ASAP7_75t_L g1696 ( 
.A(n_1659),
.B(n_1482),
.Y(n_1696)
);

AO32x2_ASAP7_75t_L g1697 ( 
.A1(n_1586),
.A2(n_1453),
.A3(n_1559),
.B1(n_1447),
.B2(n_1475),
.Y(n_1697)
);

NAND2xp5_ASAP7_75t_L g1698 ( 
.A(n_1601),
.B(n_1556),
.Y(n_1698)
);

OAI22xp5_ASAP7_75t_SL g1699 ( 
.A1(n_1671),
.A2(n_1592),
.B1(n_1686),
.B2(n_1639),
.Y(n_1699)
);

OR2x6_ASAP7_75t_L g1700 ( 
.A(n_1633),
.B(n_1588),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1594),
.Y(n_1701)
);

INVx4_ASAP7_75t_L g1702 ( 
.A(n_1628),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1596),
.Y(n_1703)
);

AOI22xp33_ASAP7_75t_L g1704 ( 
.A1(n_1641),
.A2(n_1603),
.B1(n_1632),
.B2(n_1589),
.Y(n_1704)
);

AND2x2_ASAP7_75t_L g1705 ( 
.A(n_1609),
.B(n_1589),
.Y(n_1705)
);

NAND2xp5_ASAP7_75t_L g1706 ( 
.A(n_1600),
.B(n_1627),
.Y(n_1706)
);

NAND2xp33_ASAP7_75t_L g1707 ( 
.A(n_1668),
.B(n_1647),
.Y(n_1707)
);

A2O1A1Ixp33_ASAP7_75t_L g1708 ( 
.A1(n_1634),
.A2(n_1647),
.B(n_1654),
.C(n_1650),
.Y(n_1708)
);

O2A1O1Ixp33_ASAP7_75t_L g1709 ( 
.A1(n_1628),
.A2(n_1652),
.B(n_1638),
.C(n_1648),
.Y(n_1709)
);

OA21x2_ASAP7_75t_L g1710 ( 
.A1(n_1593),
.A2(n_1587),
.B(n_1612),
.Y(n_1710)
);

NOR2xp33_ASAP7_75t_L g1711 ( 
.A(n_1628),
.B(n_1653),
.Y(n_1711)
);

O2A1O1Ixp33_ASAP7_75t_L g1712 ( 
.A1(n_1652),
.A2(n_1638),
.B(n_1648),
.C(n_1650),
.Y(n_1712)
);

AND2x2_ASAP7_75t_L g1713 ( 
.A(n_1627),
.B(n_1615),
.Y(n_1713)
);

AND2x2_ASAP7_75t_L g1714 ( 
.A(n_1615),
.B(n_1612),
.Y(n_1714)
);

OA21x2_ASAP7_75t_L g1715 ( 
.A1(n_1593),
.A2(n_1587),
.B(n_1607),
.Y(n_1715)
);

INVxp67_ASAP7_75t_L g1716 ( 
.A(n_1658),
.Y(n_1716)
);

AND2x2_ASAP7_75t_L g1717 ( 
.A(n_1596),
.B(n_1602),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_L g1718 ( 
.A(n_1619),
.B(n_1595),
.Y(n_1718)
);

OAI21xp5_ASAP7_75t_L g1719 ( 
.A1(n_1631),
.A2(n_1653),
.B(n_1655),
.Y(n_1719)
);

OAI21xp5_ASAP7_75t_L g1720 ( 
.A1(n_1631),
.A2(n_1655),
.B(n_1654),
.Y(n_1720)
);

BUFx6f_ASAP7_75t_L g1721 ( 
.A(n_1689),
.Y(n_1721)
);

BUFx4f_ASAP7_75t_SL g1722 ( 
.A(n_1662),
.Y(n_1722)
);

AO32x1_ASAP7_75t_L g1723 ( 
.A1(n_1586),
.A2(n_1641),
.A3(n_1649),
.B1(n_1632),
.B2(n_1606),
.Y(n_1723)
);

AND2x4_ASAP7_75t_L g1724 ( 
.A(n_1626),
.B(n_1598),
.Y(n_1724)
);

OR2x2_ASAP7_75t_L g1725 ( 
.A(n_1595),
.B(n_1583),
.Y(n_1725)
);

AND2x2_ASAP7_75t_L g1726 ( 
.A(n_1676),
.B(n_1679),
.Y(n_1726)
);

AOI22xp5_ASAP7_75t_L g1727 ( 
.A1(n_1663),
.A2(n_1657),
.B1(n_1664),
.B2(n_1660),
.Y(n_1727)
);

OAI22xp5_ASAP7_75t_L g1728 ( 
.A1(n_1657),
.A2(n_1671),
.B1(n_1664),
.B2(n_1637),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1610),
.Y(n_1729)
);

OAI21xp5_ASAP7_75t_L g1730 ( 
.A1(n_1607),
.A2(n_1630),
.B(n_1670),
.Y(n_1730)
);

CKINVDCx5p33_ASAP7_75t_R g1731 ( 
.A(n_1608),
.Y(n_1731)
);

AOI22xp5_ASAP7_75t_L g1732 ( 
.A1(n_1660),
.A2(n_1636),
.B1(n_1656),
.B2(n_1606),
.Y(n_1732)
);

AND2x2_ASAP7_75t_L g1733 ( 
.A(n_1611),
.B(n_1616),
.Y(n_1733)
);

OAI221xp5_ASAP7_75t_L g1734 ( 
.A1(n_1666),
.A2(n_1630),
.B1(n_1614),
.B2(n_1683),
.C(n_1642),
.Y(n_1734)
);

OA21x2_ASAP7_75t_L g1735 ( 
.A1(n_1649),
.A2(n_1591),
.B(n_1590),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1617),
.Y(n_1736)
);

A2O1A1Ixp33_ASAP7_75t_L g1737 ( 
.A1(n_1644),
.A2(n_1656),
.B(n_1666),
.C(n_1646),
.Y(n_1737)
);

OA21x2_ASAP7_75t_L g1738 ( 
.A1(n_1590),
.A2(n_1591),
.B(n_1581),
.Y(n_1738)
);

OAI21xp5_ASAP7_75t_L g1739 ( 
.A1(n_1630),
.A2(n_1670),
.B(n_1668),
.Y(n_1739)
);

AOI221xp5_ASAP7_75t_L g1740 ( 
.A1(n_1617),
.A2(n_1618),
.B1(n_1623),
.B2(n_1622),
.C(n_1620),
.Y(n_1740)
);

AND2x2_ASAP7_75t_L g1741 ( 
.A(n_1618),
.B(n_1620),
.Y(n_1741)
);

AND2x2_ASAP7_75t_L g1742 ( 
.A(n_1622),
.B(n_1623),
.Y(n_1742)
);

AND2x2_ASAP7_75t_L g1743 ( 
.A(n_1613),
.B(n_1624),
.Y(n_1743)
);

OR2x2_ASAP7_75t_L g1744 ( 
.A(n_1643),
.B(n_1661),
.Y(n_1744)
);

OAI22xp5_ASAP7_75t_L g1745 ( 
.A1(n_1684),
.A2(n_1582),
.B1(n_1672),
.B2(n_1605),
.Y(n_1745)
);

AOI21xp5_ASAP7_75t_L g1746 ( 
.A1(n_1630),
.A2(n_1660),
.B(n_1640),
.Y(n_1746)
);

AOI22xp5_ASAP7_75t_L g1747 ( 
.A1(n_1644),
.A2(n_1646),
.B1(n_1680),
.B2(n_1683),
.Y(n_1747)
);

A2O1A1Ixp33_ASAP7_75t_L g1748 ( 
.A1(n_1645),
.A2(n_1599),
.B(n_1673),
.C(n_1651),
.Y(n_1748)
);

AOI221xp5_ASAP7_75t_L g1749 ( 
.A1(n_1581),
.A2(n_1584),
.B1(n_1642),
.B2(n_1645),
.C(n_1680),
.Y(n_1749)
);

BUFx2_ASAP7_75t_L g1750 ( 
.A(n_1629),
.Y(n_1750)
);

AOI221xp5_ASAP7_75t_L g1751 ( 
.A1(n_1584),
.A2(n_1604),
.B1(n_1665),
.B2(n_1685),
.C(n_1635),
.Y(n_1751)
);

AND2x2_ASAP7_75t_L g1752 ( 
.A(n_1604),
.B(n_1640),
.Y(n_1752)
);

INVx1_ASAP7_75t_SL g1753 ( 
.A(n_1678),
.Y(n_1753)
);

AOI22xp33_ASAP7_75t_L g1754 ( 
.A1(n_1704),
.A2(n_1685),
.B1(n_1599),
.B2(n_1662),
.Y(n_1754)
);

AND2x2_ASAP7_75t_L g1755 ( 
.A(n_1714),
.B(n_1675),
.Y(n_1755)
);

OR2x2_ASAP7_75t_L g1756 ( 
.A(n_1705),
.B(n_1667),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1738),
.Y(n_1757)
);

INVx2_ASAP7_75t_L g1758 ( 
.A(n_1738),
.Y(n_1758)
);

INVx2_ASAP7_75t_L g1759 ( 
.A(n_1738),
.Y(n_1759)
);

INVxp67_ASAP7_75t_SL g1760 ( 
.A(n_1711),
.Y(n_1760)
);

HB1xp67_ASAP7_75t_L g1761 ( 
.A(n_1714),
.Y(n_1761)
);

INVx2_ASAP7_75t_L g1762 ( 
.A(n_1735),
.Y(n_1762)
);

BUFx6f_ASAP7_75t_L g1763 ( 
.A(n_1710),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1695),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1701),
.Y(n_1765)
);

HB1xp67_ASAP7_75t_L g1766 ( 
.A(n_1752),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1703),
.Y(n_1767)
);

HB1xp67_ASAP7_75t_L g1768 ( 
.A(n_1752),
.Y(n_1768)
);

AOI221xp5_ASAP7_75t_L g1769 ( 
.A1(n_1708),
.A2(n_1682),
.B1(n_1592),
.B2(n_1688),
.C(n_1687),
.Y(n_1769)
);

AOI22xp5_ASAP7_75t_L g1770 ( 
.A1(n_1708),
.A2(n_1599),
.B1(n_1582),
.B2(n_1665),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1729),
.Y(n_1771)
);

NAND2xp5_ASAP7_75t_L g1772 ( 
.A(n_1691),
.B(n_1713),
.Y(n_1772)
);

AND2x4_ASAP7_75t_L g1773 ( 
.A(n_1700),
.B(n_1669),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1736),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1717),
.Y(n_1775)
);

INVx1_ASAP7_75t_SL g1776 ( 
.A(n_1750),
.Y(n_1776)
);

NAND2xp5_ASAP7_75t_L g1777 ( 
.A(n_1718),
.B(n_1677),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1717),
.Y(n_1778)
);

HB1xp67_ASAP7_75t_L g1779 ( 
.A(n_1706),
.Y(n_1779)
);

INVx4_ASAP7_75t_L g1780 ( 
.A(n_1721),
.Y(n_1780)
);

AND2x2_ASAP7_75t_L g1781 ( 
.A(n_1715),
.B(n_1677),
.Y(n_1781)
);

INVx1_ASAP7_75t_SL g1782 ( 
.A(n_1690),
.Y(n_1782)
);

HB1xp67_ASAP7_75t_L g1783 ( 
.A(n_1733),
.Y(n_1783)
);

INVxp67_ASAP7_75t_L g1784 ( 
.A(n_1711),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1764),
.Y(n_1785)
);

NAND2xp5_ASAP7_75t_L g1786 ( 
.A(n_1779),
.B(n_1741),
.Y(n_1786)
);

CKINVDCx5p33_ASAP7_75t_R g1787 ( 
.A(n_1776),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1764),
.Y(n_1788)
);

NAND3xp33_ASAP7_75t_L g1789 ( 
.A(n_1784),
.B(n_1702),
.C(n_1709),
.Y(n_1789)
);

AND2x4_ASAP7_75t_L g1790 ( 
.A(n_1773),
.B(n_1739),
.Y(n_1790)
);

BUFx12f_ASAP7_75t_L g1791 ( 
.A(n_1773),
.Y(n_1791)
);

INVx2_ASAP7_75t_L g1792 ( 
.A(n_1762),
.Y(n_1792)
);

HB1xp67_ASAP7_75t_L g1793 ( 
.A(n_1766),
.Y(n_1793)
);

AND2x2_ASAP7_75t_L g1794 ( 
.A(n_1761),
.B(n_1730),
.Y(n_1794)
);

INVx2_ASAP7_75t_L g1795 ( 
.A(n_1762),
.Y(n_1795)
);

AND2x2_ASAP7_75t_L g1796 ( 
.A(n_1761),
.B(n_1702),
.Y(n_1796)
);

OAI22xp5_ASAP7_75t_L g1797 ( 
.A1(n_1769),
.A2(n_1727),
.B1(n_1732),
.B2(n_1693),
.Y(n_1797)
);

OR2x6_ASAP7_75t_L g1798 ( 
.A(n_1773),
.B(n_1746),
.Y(n_1798)
);

AOI31xp33_ASAP7_75t_L g1799 ( 
.A1(n_1769),
.A2(n_1728),
.A3(n_1751),
.B(n_1693),
.Y(n_1799)
);

AOI21xp5_ASAP7_75t_L g1800 ( 
.A1(n_1760),
.A2(n_1707),
.B(n_1723),
.Y(n_1800)
);

NAND2xp5_ASAP7_75t_L g1801 ( 
.A(n_1784),
.B(n_1742),
.Y(n_1801)
);

AOI22xp33_ASAP7_75t_L g1802 ( 
.A1(n_1770),
.A2(n_1734),
.B1(n_1720),
.B2(n_1749),
.Y(n_1802)
);

NOR2xp33_ASAP7_75t_L g1803 ( 
.A(n_1776),
.B(n_1731),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1764),
.Y(n_1804)
);

AO21x2_ASAP7_75t_L g1805 ( 
.A1(n_1757),
.A2(n_1719),
.B(n_1748),
.Y(n_1805)
);

AND2x2_ASAP7_75t_L g1806 ( 
.A(n_1783),
.B(n_1716),
.Y(n_1806)
);

OR2x2_ASAP7_75t_L g1807 ( 
.A(n_1783),
.B(n_1725),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1765),
.Y(n_1808)
);

AND2x2_ASAP7_75t_L g1809 ( 
.A(n_1772),
.B(n_1726),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1765),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1767),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1767),
.Y(n_1812)
);

AOI22xp33_ASAP7_75t_L g1813 ( 
.A1(n_1770),
.A2(n_1699),
.B1(n_1747),
.B2(n_1724),
.Y(n_1813)
);

AND2x2_ASAP7_75t_L g1814 ( 
.A(n_1772),
.B(n_1694),
.Y(n_1814)
);

AOI33xp33_ASAP7_75t_L g1815 ( 
.A1(n_1782),
.A2(n_1753),
.A3(n_1712),
.B1(n_1740),
.B2(n_1696),
.B3(n_1674),
.Y(n_1815)
);

AND2x2_ASAP7_75t_L g1816 ( 
.A(n_1782),
.B(n_1700),
.Y(n_1816)
);

OR2x2_ASAP7_75t_L g1817 ( 
.A(n_1756),
.B(n_1744),
.Y(n_1817)
);

NAND2xp5_ASAP7_75t_L g1818 ( 
.A(n_1760),
.B(n_1743),
.Y(n_1818)
);

AND2x4_ASAP7_75t_L g1819 ( 
.A(n_1773),
.B(n_1700),
.Y(n_1819)
);

BUFx6f_ASAP7_75t_L g1820 ( 
.A(n_1763),
.Y(n_1820)
);

AND2x2_ASAP7_75t_L g1821 ( 
.A(n_1766),
.B(n_1724),
.Y(n_1821)
);

INVx4_ASAP7_75t_L g1822 ( 
.A(n_1780),
.Y(n_1822)
);

AOI21xp5_ASAP7_75t_L g1823 ( 
.A1(n_1781),
.A2(n_1723),
.B(n_1737),
.Y(n_1823)
);

NAND2xp5_ASAP7_75t_L g1824 ( 
.A(n_1786),
.B(n_1768),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1785),
.Y(n_1825)
);

AND2x2_ASAP7_75t_L g1826 ( 
.A(n_1794),
.B(n_1755),
.Y(n_1826)
);

OR2x2_ASAP7_75t_L g1827 ( 
.A(n_1801),
.B(n_1777),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1785),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1788),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1788),
.Y(n_1830)
);

NAND5xp2_ASAP7_75t_L g1831 ( 
.A(n_1803),
.B(n_1692),
.C(n_1597),
.D(n_1722),
.E(n_1754),
.Y(n_1831)
);

OR2x2_ASAP7_75t_L g1832 ( 
.A(n_1801),
.B(n_1775),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1804),
.Y(n_1833)
);

AND2x4_ASAP7_75t_L g1834 ( 
.A(n_1819),
.B(n_1773),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1804),
.Y(n_1835)
);

INVx2_ASAP7_75t_L g1836 ( 
.A(n_1792),
.Y(n_1836)
);

AND2x2_ASAP7_75t_L g1837 ( 
.A(n_1794),
.B(n_1755),
.Y(n_1837)
);

AND2x2_ASAP7_75t_L g1838 ( 
.A(n_1794),
.B(n_1755),
.Y(n_1838)
);

INVx2_ASAP7_75t_L g1839 ( 
.A(n_1792),
.Y(n_1839)
);

AND2x2_ASAP7_75t_L g1840 ( 
.A(n_1796),
.B(n_1781),
.Y(n_1840)
);

AND2x2_ASAP7_75t_L g1841 ( 
.A(n_1796),
.B(n_1781),
.Y(n_1841)
);

NAND2xp5_ASAP7_75t_L g1842 ( 
.A(n_1808),
.B(n_1771),
.Y(n_1842)
);

NAND2xp5_ASAP7_75t_L g1843 ( 
.A(n_1808),
.B(n_1774),
.Y(n_1843)
);

AND2x4_ASAP7_75t_SL g1844 ( 
.A(n_1790),
.B(n_1721),
.Y(n_1844)
);

AND2x2_ASAP7_75t_L g1845 ( 
.A(n_1821),
.B(n_1775),
.Y(n_1845)
);

BUFx2_ASAP7_75t_L g1846 ( 
.A(n_1791),
.Y(n_1846)
);

INVx2_ASAP7_75t_L g1847 ( 
.A(n_1792),
.Y(n_1847)
);

OR2x2_ASAP7_75t_L g1848 ( 
.A(n_1807),
.B(n_1777),
.Y(n_1848)
);

NAND2xp5_ASAP7_75t_L g1849 ( 
.A(n_1810),
.B(n_1774),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1811),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1811),
.Y(n_1851)
);

INVx1_ASAP7_75t_SL g1852 ( 
.A(n_1787),
.Y(n_1852)
);

INVx2_ASAP7_75t_L g1853 ( 
.A(n_1795),
.Y(n_1853)
);

AND2x2_ASAP7_75t_L g1854 ( 
.A(n_1821),
.B(n_1778),
.Y(n_1854)
);

INVx4_ASAP7_75t_L g1855 ( 
.A(n_1822),
.Y(n_1855)
);

HB1xp67_ASAP7_75t_L g1856 ( 
.A(n_1812),
.Y(n_1856)
);

AND2x2_ASAP7_75t_L g1857 ( 
.A(n_1846),
.B(n_1816),
.Y(n_1857)
);

NAND2xp5_ASAP7_75t_L g1858 ( 
.A(n_1826),
.B(n_1815),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_1856),
.Y(n_1859)
);

AND2x2_ASAP7_75t_L g1860 ( 
.A(n_1846),
.B(n_1816),
.Y(n_1860)
);

OR2x6_ASAP7_75t_L g1861 ( 
.A(n_1855),
.B(n_1797),
.Y(n_1861)
);

INVx1_ASAP7_75t_L g1862 ( 
.A(n_1856),
.Y(n_1862)
);

NOR2x1p5_ASAP7_75t_L g1863 ( 
.A(n_1855),
.B(n_1731),
.Y(n_1863)
);

AND2x4_ASAP7_75t_SL g1864 ( 
.A(n_1834),
.B(n_1822),
.Y(n_1864)
);

AND2x2_ASAP7_75t_L g1865 ( 
.A(n_1826),
.B(n_1814),
.Y(n_1865)
);

BUFx2_ASAP7_75t_L g1866 ( 
.A(n_1855),
.Y(n_1866)
);

INVxp67_ASAP7_75t_SL g1867 ( 
.A(n_1842),
.Y(n_1867)
);

NAND2xp33_ASAP7_75t_L g1868 ( 
.A(n_1852),
.B(n_1806),
.Y(n_1868)
);

AND2x2_ASAP7_75t_L g1869 ( 
.A(n_1826),
.B(n_1814),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1825),
.Y(n_1870)
);

HB1xp67_ASAP7_75t_L g1871 ( 
.A(n_1842),
.Y(n_1871)
);

NOR2x1p5_ASAP7_75t_L g1872 ( 
.A(n_1855),
.B(n_1605),
.Y(n_1872)
);

AND2x4_ASAP7_75t_L g1873 ( 
.A(n_1834),
.B(n_1790),
.Y(n_1873)
);

HB1xp67_ASAP7_75t_L g1874 ( 
.A(n_1843),
.Y(n_1874)
);

AND2x2_ASAP7_75t_L g1875 ( 
.A(n_1837),
.B(n_1806),
.Y(n_1875)
);

NAND2xp5_ASAP7_75t_L g1876 ( 
.A(n_1837),
.B(n_1809),
.Y(n_1876)
);

HB1xp67_ASAP7_75t_L g1877 ( 
.A(n_1843),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1825),
.Y(n_1878)
);

HB1xp67_ASAP7_75t_L g1879 ( 
.A(n_1849),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1828),
.Y(n_1880)
);

BUFx2_ASAP7_75t_L g1881 ( 
.A(n_1828),
.Y(n_1881)
);

INVxp67_ASAP7_75t_L g1882 ( 
.A(n_1852),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1829),
.Y(n_1883)
);

HB1xp67_ASAP7_75t_L g1884 ( 
.A(n_1849),
.Y(n_1884)
);

NAND2xp5_ASAP7_75t_L g1885 ( 
.A(n_1837),
.B(n_1809),
.Y(n_1885)
);

NAND2xp5_ASAP7_75t_L g1886 ( 
.A(n_1838),
.B(n_1818),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1829),
.Y(n_1887)
);

OR2x2_ASAP7_75t_L g1888 ( 
.A(n_1827),
.B(n_1817),
.Y(n_1888)
);

OR2x2_ASAP7_75t_L g1889 ( 
.A(n_1827),
.B(n_1817),
.Y(n_1889)
);

INVx1_ASAP7_75t_SL g1890 ( 
.A(n_1844),
.Y(n_1890)
);

NOR2x1_ASAP7_75t_L g1891 ( 
.A(n_1831),
.B(n_1822),
.Y(n_1891)
);

CKINVDCx20_ASAP7_75t_R g1892 ( 
.A(n_1844),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1830),
.Y(n_1893)
);

AND2x2_ASAP7_75t_L g1894 ( 
.A(n_1838),
.B(n_1793),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1830),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1833),
.Y(n_1896)
);

NAND2xp5_ASAP7_75t_L g1897 ( 
.A(n_1838),
.B(n_1818),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_1833),
.Y(n_1898)
);

OR2x2_ASAP7_75t_L g1899 ( 
.A(n_1848),
.B(n_1793),
.Y(n_1899)
);

INVx2_ASAP7_75t_L g1900 ( 
.A(n_1836),
.Y(n_1900)
);

INVx2_ASAP7_75t_L g1901 ( 
.A(n_1836),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1835),
.Y(n_1902)
);

INVx1_ASAP7_75t_SL g1903 ( 
.A(n_1892),
.Y(n_1903)
);

AOI22xp5_ASAP7_75t_L g1904 ( 
.A1(n_1861),
.A2(n_1797),
.B1(n_1823),
.B2(n_1802),
.Y(n_1904)
);

NAND2xp5_ASAP7_75t_SL g1905 ( 
.A(n_1891),
.B(n_1844),
.Y(n_1905)
);

AND2x2_ASAP7_75t_L g1906 ( 
.A(n_1865),
.B(n_1834),
.Y(n_1906)
);

INVxp67_ASAP7_75t_L g1907 ( 
.A(n_1868),
.Y(n_1907)
);

AND2x2_ASAP7_75t_L g1908 ( 
.A(n_1865),
.B(n_1834),
.Y(n_1908)
);

OR2x2_ASAP7_75t_L g1909 ( 
.A(n_1888),
.B(n_1848),
.Y(n_1909)
);

OAI31xp33_ASAP7_75t_SL g1910 ( 
.A1(n_1891),
.A2(n_1831),
.A3(n_1789),
.B(n_1840),
.Y(n_1910)
);

NAND2xp5_ASAP7_75t_L g1911 ( 
.A(n_1869),
.B(n_1854),
.Y(n_1911)
);

AND2x2_ASAP7_75t_L g1912 ( 
.A(n_1869),
.B(n_1834),
.Y(n_1912)
);

INVx2_ASAP7_75t_L g1913 ( 
.A(n_1881),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1881),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1870),
.Y(n_1915)
);

AND2x2_ASAP7_75t_L g1916 ( 
.A(n_1861),
.B(n_1840),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1870),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1878),
.Y(n_1918)
);

AND2x2_ASAP7_75t_L g1919 ( 
.A(n_1861),
.B(n_1840),
.Y(n_1919)
);

AND2x2_ASAP7_75t_L g1920 ( 
.A(n_1861),
.B(n_1841),
.Y(n_1920)
);

OR2x2_ASAP7_75t_L g1921 ( 
.A(n_1888),
.B(n_1832),
.Y(n_1921)
);

INVx1_ASAP7_75t_SL g1922 ( 
.A(n_1857),
.Y(n_1922)
);

INVx2_ASAP7_75t_L g1923 ( 
.A(n_1900),
.Y(n_1923)
);

NOR2xp67_ASAP7_75t_L g1924 ( 
.A(n_1873),
.B(n_1791),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1878),
.Y(n_1925)
);

OR2x2_ASAP7_75t_L g1926 ( 
.A(n_1889),
.B(n_1832),
.Y(n_1926)
);

NAND2x1p5_ASAP7_75t_L g1927 ( 
.A(n_1872),
.B(n_1822),
.Y(n_1927)
);

OR2x6_ASAP7_75t_L g1928 ( 
.A(n_1861),
.B(n_1823),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1880),
.Y(n_1929)
);

NOR2xp33_ASAP7_75t_L g1930 ( 
.A(n_1882),
.B(n_1662),
.Y(n_1930)
);

INVx1_ASAP7_75t_L g1931 ( 
.A(n_1880),
.Y(n_1931)
);

AND2x2_ASAP7_75t_L g1932 ( 
.A(n_1864),
.B(n_1841),
.Y(n_1932)
);

NOR2xp33_ASAP7_75t_SL g1933 ( 
.A(n_1890),
.B(n_1791),
.Y(n_1933)
);

OR2x2_ASAP7_75t_L g1934 ( 
.A(n_1889),
.B(n_1832),
.Y(n_1934)
);

NAND2xp5_ASAP7_75t_L g1935 ( 
.A(n_1875),
.B(n_1845),
.Y(n_1935)
);

INVx2_ASAP7_75t_SL g1936 ( 
.A(n_1863),
.Y(n_1936)
);

INVx1_ASAP7_75t_L g1937 ( 
.A(n_1883),
.Y(n_1937)
);

AND2x2_ASAP7_75t_L g1938 ( 
.A(n_1864),
.B(n_1841),
.Y(n_1938)
);

INVx1_ASAP7_75t_L g1939 ( 
.A(n_1883),
.Y(n_1939)
);

NOR2xp33_ASAP7_75t_L g1940 ( 
.A(n_1857),
.B(n_1678),
.Y(n_1940)
);

NAND3xp33_ASAP7_75t_L g1941 ( 
.A(n_1904),
.B(n_1858),
.C(n_1859),
.Y(n_1941)
);

OAI31xp33_ASAP7_75t_L g1942 ( 
.A1(n_1907),
.A2(n_1789),
.A3(n_1800),
.B(n_1813),
.Y(n_1942)
);

INVx1_ASAP7_75t_L g1943 ( 
.A(n_1915),
.Y(n_1943)
);

INVx1_ASAP7_75t_SL g1944 ( 
.A(n_1903),
.Y(n_1944)
);

AOI32xp33_ASAP7_75t_L g1945 ( 
.A1(n_1916),
.A2(n_1919),
.A3(n_1920),
.B1(n_1922),
.B2(n_1928),
.Y(n_1945)
);

AOI22xp5_ASAP7_75t_L g1946 ( 
.A1(n_1928),
.A2(n_1800),
.B1(n_1805),
.B2(n_1860),
.Y(n_1946)
);

INVx3_ASAP7_75t_R g1947 ( 
.A(n_1913),
.Y(n_1947)
);

OR2x2_ASAP7_75t_L g1948 ( 
.A(n_1909),
.B(n_1876),
.Y(n_1948)
);

AOI22xp33_ASAP7_75t_L g1949 ( 
.A1(n_1928),
.A2(n_1805),
.B1(n_1860),
.B2(n_1798),
.Y(n_1949)
);

OAI22xp5_ASAP7_75t_L g1950 ( 
.A1(n_1928),
.A2(n_1799),
.B1(n_1873),
.B2(n_1885),
.Y(n_1950)
);

OAI22xp33_ASAP7_75t_L g1951 ( 
.A1(n_1933),
.A2(n_1799),
.B1(n_1798),
.B2(n_1886),
.Y(n_1951)
);

INVx1_ASAP7_75t_L g1952 ( 
.A(n_1915),
.Y(n_1952)
);

INVx2_ASAP7_75t_L g1953 ( 
.A(n_1906),
.Y(n_1953)
);

AOI22xp5_ASAP7_75t_L g1954 ( 
.A1(n_1916),
.A2(n_1805),
.B1(n_1798),
.B2(n_1900),
.Y(n_1954)
);

INVx1_ASAP7_75t_SL g1955 ( 
.A(n_1919),
.Y(n_1955)
);

OAI21xp33_ASAP7_75t_L g1956 ( 
.A1(n_1910),
.A2(n_1920),
.B(n_1909),
.Y(n_1956)
);

AOI222xp33_ASAP7_75t_L g1957 ( 
.A1(n_1923),
.A2(n_1867),
.B1(n_1758),
.B2(n_1759),
.C1(n_1757),
.C2(n_1901),
.Y(n_1957)
);

AOI22xp5_ASAP7_75t_L g1958 ( 
.A1(n_1940),
.A2(n_1805),
.B1(n_1798),
.B2(n_1901),
.Y(n_1958)
);

AND2x2_ASAP7_75t_L g1959 ( 
.A(n_1906),
.B(n_1863),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_1917),
.Y(n_1960)
);

NAND2xp5_ASAP7_75t_L g1961 ( 
.A(n_1913),
.B(n_1875),
.Y(n_1961)
);

AND2x2_ASAP7_75t_L g1962 ( 
.A(n_1908),
.B(n_1872),
.Y(n_1962)
);

AND2x4_ASAP7_75t_L g1963 ( 
.A(n_1936),
.B(n_1873),
.Y(n_1963)
);

O2A1O1Ixp33_ASAP7_75t_L g1964 ( 
.A1(n_1914),
.A2(n_1859),
.B(n_1862),
.C(n_1884),
.Y(n_1964)
);

AOI221xp5_ASAP7_75t_L g1965 ( 
.A1(n_1939),
.A2(n_1879),
.B1(n_1871),
.B2(n_1874),
.C(n_1877),
.Y(n_1965)
);

NAND2x1p5_ASAP7_75t_L g1966 ( 
.A(n_1905),
.B(n_1866),
.Y(n_1966)
);

HB1xp67_ASAP7_75t_L g1967 ( 
.A(n_1914),
.Y(n_1967)
);

NAND2xp5_ASAP7_75t_L g1968 ( 
.A(n_1944),
.B(n_1941),
.Y(n_1968)
);

AOI22xp5_ASAP7_75t_L g1969 ( 
.A1(n_1941),
.A2(n_1924),
.B1(n_1923),
.B2(n_1930),
.Y(n_1969)
);

NAND2xp5_ASAP7_75t_L g1970 ( 
.A(n_1967),
.B(n_1925),
.Y(n_1970)
);

AOI21xp5_ASAP7_75t_L g1971 ( 
.A1(n_1942),
.A2(n_1936),
.B(n_1866),
.Y(n_1971)
);

INVx2_ASAP7_75t_SL g1972 ( 
.A(n_1963),
.Y(n_1972)
);

XOR2x2_ASAP7_75t_L g1973 ( 
.A(n_1950),
.B(n_1697),
.Y(n_1973)
);

OR2x2_ASAP7_75t_L g1974 ( 
.A(n_1948),
.B(n_1921),
.Y(n_1974)
);

OAI22xp33_ASAP7_75t_L g1975 ( 
.A1(n_1946),
.A2(n_1798),
.B1(n_1934),
.B2(n_1926),
.Y(n_1975)
);

INVx1_ASAP7_75t_L g1976 ( 
.A(n_1943),
.Y(n_1976)
);

INVx2_ASAP7_75t_SL g1977 ( 
.A(n_1963),
.Y(n_1977)
);

NAND3xp33_ASAP7_75t_L g1978 ( 
.A(n_1942),
.B(n_1918),
.C(n_1917),
.Y(n_1978)
);

INVx1_ASAP7_75t_L g1979 ( 
.A(n_1952),
.Y(n_1979)
);

NAND2xp5_ASAP7_75t_L g1980 ( 
.A(n_1955),
.B(n_1921),
.Y(n_1980)
);

AND2x2_ASAP7_75t_L g1981 ( 
.A(n_1959),
.B(n_1908),
.Y(n_1981)
);

AND2x2_ASAP7_75t_SL g1982 ( 
.A(n_1961),
.B(n_1864),
.Y(n_1982)
);

AOI322xp5_ASAP7_75t_L g1983 ( 
.A1(n_1956),
.A2(n_1935),
.A3(n_1897),
.B1(n_1894),
.B2(n_1911),
.C1(n_1939),
.C2(n_1929),
.Y(n_1983)
);

NAND2xp5_ASAP7_75t_SL g1984 ( 
.A(n_1951),
.B(n_1873),
.Y(n_1984)
);

INVx2_ASAP7_75t_L g1985 ( 
.A(n_1953),
.Y(n_1985)
);

INVxp67_ASAP7_75t_SL g1986 ( 
.A(n_1966),
.Y(n_1986)
);

AOI221xp5_ASAP7_75t_L g1987 ( 
.A1(n_1949),
.A2(n_1918),
.B1(n_1929),
.B2(n_1937),
.C(n_1931),
.Y(n_1987)
);

AOI322xp5_ASAP7_75t_L g1988 ( 
.A1(n_1954),
.A2(n_1894),
.A3(n_1912),
.B1(n_1862),
.B2(n_1938),
.C1(n_1932),
.C2(n_1758),
.Y(n_1988)
);

INVx1_ASAP7_75t_SL g1989 ( 
.A(n_1968),
.Y(n_1989)
);

O2A1O1Ixp33_ASAP7_75t_SL g1990 ( 
.A1(n_1968),
.A2(n_1964),
.B(n_1965),
.C(n_1947),
.Y(n_1990)
);

INVxp67_ASAP7_75t_SL g1991 ( 
.A(n_1986),
.Y(n_1991)
);

XNOR2xp5_ASAP7_75t_L g1992 ( 
.A(n_1973),
.B(n_1966),
.Y(n_1992)
);

AOI211xp5_ASAP7_75t_L g1993 ( 
.A1(n_1978),
.A2(n_1960),
.B(n_1958),
.C(n_1962),
.Y(n_1993)
);

AOI221xp5_ASAP7_75t_L g1994 ( 
.A1(n_1978),
.A2(n_1987),
.B1(n_1971),
.B2(n_1975),
.C(n_1945),
.Y(n_1994)
);

OAI21xp5_ASAP7_75t_L g1995 ( 
.A1(n_1988),
.A2(n_1957),
.B(n_1938),
.Y(n_1995)
);

XNOR2xp5_ASAP7_75t_L g1996 ( 
.A(n_1972),
.B(n_1932),
.Y(n_1996)
);

NAND2xp5_ASAP7_75t_L g1997 ( 
.A(n_1977),
.B(n_1926),
.Y(n_1997)
);

INVx1_ASAP7_75t_L g1998 ( 
.A(n_1974),
.Y(n_1998)
);

OAI22xp33_ASAP7_75t_SL g1999 ( 
.A1(n_1984),
.A2(n_1934),
.B1(n_1927),
.B2(n_1899),
.Y(n_1999)
);

NAND3xp33_ASAP7_75t_SL g2000 ( 
.A(n_1989),
.B(n_1983),
.C(n_1969),
.Y(n_2000)
);

NOR2xp33_ASAP7_75t_L g2001 ( 
.A(n_1991),
.B(n_1980),
.Y(n_2001)
);

AOI21xp5_ASAP7_75t_L g2002 ( 
.A1(n_1990),
.A2(n_1970),
.B(n_1982),
.Y(n_2002)
);

AND2x2_ASAP7_75t_L g2003 ( 
.A(n_1998),
.B(n_1981),
.Y(n_2003)
);

NOR3xp33_ASAP7_75t_L g2004 ( 
.A(n_1991),
.B(n_1985),
.C(n_1970),
.Y(n_2004)
);

NAND2xp5_ASAP7_75t_SL g2005 ( 
.A(n_1999),
.B(n_1927),
.Y(n_2005)
);

OAI21xp5_ASAP7_75t_L g2006 ( 
.A1(n_1994),
.A2(n_1979),
.B(n_1976),
.Y(n_2006)
);

NOR3xp33_ASAP7_75t_L g2007 ( 
.A(n_1993),
.B(n_1997),
.C(n_1995),
.Y(n_2007)
);

NAND2xp5_ASAP7_75t_L g2008 ( 
.A(n_1996),
.B(n_1912),
.Y(n_2008)
);

BUFx2_ASAP7_75t_L g2009 ( 
.A(n_1992),
.Y(n_2009)
);

NAND2xp33_ASAP7_75t_SL g2010 ( 
.A(n_2003),
.B(n_2008),
.Y(n_2010)
);

INVx2_ASAP7_75t_SL g2011 ( 
.A(n_2005),
.Y(n_2011)
);

NOR3xp33_ASAP7_75t_SL g2012 ( 
.A(n_2000),
.B(n_2001),
.C(n_2006),
.Y(n_2012)
);

OAI21xp33_ASAP7_75t_L g2013 ( 
.A1(n_2007),
.A2(n_1927),
.B(n_1893),
.Y(n_2013)
);

NOR4xp25_ASAP7_75t_L g2014 ( 
.A(n_2004),
.B(n_1902),
.C(n_1898),
.D(n_1896),
.Y(n_2014)
);

NAND3xp33_ASAP7_75t_SL g2015 ( 
.A(n_2002),
.B(n_1899),
.C(n_1697),
.Y(n_2015)
);

NOR2x1_ASAP7_75t_L g2016 ( 
.A(n_2015),
.B(n_2009),
.Y(n_2016)
);

OAI321xp33_ASAP7_75t_L g2017 ( 
.A1(n_2011),
.A2(n_1798),
.A3(n_1898),
.B1(n_1896),
.B2(n_1895),
.C(n_1893),
.Y(n_2017)
);

AOI22xp5_ASAP7_75t_L g2018 ( 
.A1(n_2012),
.A2(n_2010),
.B1(n_2013),
.B2(n_2014),
.Y(n_2018)
);

INVx8_ASAP7_75t_L g2019 ( 
.A(n_2010),
.Y(n_2019)
);

NOR3xp33_ASAP7_75t_L g2020 ( 
.A(n_2015),
.B(n_1697),
.C(n_1698),
.Y(n_2020)
);

CKINVDCx11_ASAP7_75t_R g2021 ( 
.A(n_2010),
.Y(n_2021)
);

BUFx2_ASAP7_75t_L g2022 ( 
.A(n_2010),
.Y(n_2022)
);

NAND4xp75_ASAP7_75t_L g2023 ( 
.A(n_2018),
.B(n_1697),
.C(n_1895),
.D(n_1887),
.Y(n_2023)
);

INVx2_ASAP7_75t_L g2024 ( 
.A(n_2021),
.Y(n_2024)
);

NOR2x1_ASAP7_75t_L g2025 ( 
.A(n_2022),
.B(n_1887),
.Y(n_2025)
);

NOR2x1_ASAP7_75t_L g2026 ( 
.A(n_2016),
.B(n_2019),
.Y(n_2026)
);

INVx1_ASAP7_75t_L g2027 ( 
.A(n_2020),
.Y(n_2027)
);

NOR3xp33_ASAP7_75t_L g2028 ( 
.A(n_2017),
.B(n_1839),
.C(n_1836),
.Y(n_2028)
);

XNOR2xp5_ASAP7_75t_L g2029 ( 
.A(n_2026),
.B(n_1684),
.Y(n_2029)
);

NAND2x1_ASAP7_75t_SL g2030 ( 
.A(n_2024),
.B(n_1902),
.Y(n_2030)
);

NOR2xp33_ASAP7_75t_L g2031 ( 
.A(n_2023),
.B(n_1839),
.Y(n_2031)
);

INVx2_ASAP7_75t_L g2032 ( 
.A(n_2025),
.Y(n_2032)
);

INVx2_ASAP7_75t_L g2033 ( 
.A(n_2030),
.Y(n_2033)
);

OAI22x1_ASAP7_75t_L g2034 ( 
.A1(n_2033),
.A2(n_2029),
.B1(n_2032),
.B2(n_2027),
.Y(n_2034)
);

BUFx2_ASAP7_75t_L g2035 ( 
.A(n_2034),
.Y(n_2035)
);

AND3x2_ASAP7_75t_L g2036 ( 
.A(n_2034),
.B(n_2031),
.C(n_2028),
.Y(n_2036)
);

INVx1_ASAP7_75t_L g2037 ( 
.A(n_2035),
.Y(n_2037)
);

CKINVDCx20_ASAP7_75t_R g2038 ( 
.A(n_2036),
.Y(n_2038)
);

OAI22xp5_ASAP7_75t_SL g2039 ( 
.A1(n_2038),
.A2(n_1684),
.B1(n_1672),
.B2(n_1824),
.Y(n_2039)
);

AOI21xp33_ASAP7_75t_L g2040 ( 
.A1(n_2037),
.A2(n_1847),
.B(n_1839),
.Y(n_2040)
);

OR2x6_ASAP7_75t_L g2041 ( 
.A(n_2039),
.B(n_1684),
.Y(n_2041)
);

AOI22xp33_ASAP7_75t_L g2042 ( 
.A1(n_2041),
.A2(n_2040),
.B1(n_1853),
.B2(n_1847),
.Y(n_2042)
);

AOI221xp5_ASAP7_75t_L g2043 ( 
.A1(n_2042),
.A2(n_1847),
.B1(n_1853),
.B2(n_1820),
.C(n_1850),
.Y(n_2043)
);

AOI221xp5_ASAP7_75t_L g2044 ( 
.A1(n_2043),
.A2(n_1853),
.B1(n_1835),
.B2(n_1851),
.C(n_1850),
.Y(n_2044)
);

AOI211xp5_ASAP7_75t_L g2045 ( 
.A1(n_2044),
.A2(n_1674),
.B(n_1681),
.C(n_1745),
.Y(n_2045)
);


endmodule