module fake_jpeg_29496_n_297 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_297);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_297;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_127;
wire n_76;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_288;
wire n_272;
wire n_284;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_269;
wire n_122;
wire n_75;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_91;
wire n_54;
wire n_33;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_282;
wire n_96;

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_17),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_13),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_1),
.B(n_15),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_16),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_15),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_8),
.Y(n_34)
);

BUFx12_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_6),
.Y(n_38)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_11),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_43),
.Y(n_105)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_44),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_45),
.Y(n_77)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_46),
.Y(n_75)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_47),
.B(n_51),
.Y(n_76)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_48),
.Y(n_83)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_30),
.Y(n_49)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_49),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_26),
.Y(n_50)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_26),
.Y(n_52)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_52),
.Y(n_102)
);

INVx3_ASAP7_75t_SL g53 ( 
.A(n_20),
.Y(n_53)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_27),
.Y(n_54)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_54),
.Y(n_78)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_30),
.Y(n_55)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_55),
.Y(n_100)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_56),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_25),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_57),
.B(n_58),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_23),
.B(n_0),
.Y(n_58)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_25),
.Y(n_59)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_59),
.Y(n_89)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_27),
.Y(n_60)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_60),
.Y(n_108)
);

OR2x2_ASAP7_75t_L g61 ( 
.A(n_23),
.B(n_0),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_61),
.B(n_63),
.Y(n_74)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_27),
.Y(n_62)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_62),
.Y(n_90)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_31),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_64),
.B(n_65),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_25),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_24),
.B(n_18),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_66),
.B(n_67),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_31),
.Y(n_67)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_68),
.B(n_69),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_32),
.B(n_40),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_53),
.A2(n_32),
.B1(n_36),
.B2(n_40),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_73),
.A2(n_85),
.B1(n_88),
.B2(n_4),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_61),
.B(n_29),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_79),
.B(n_92),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_62),
.A2(n_40),
.B1(n_36),
.B2(n_31),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_80),
.A2(n_84),
.B1(n_94),
.B2(n_99),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_43),
.A2(n_36),
.B1(n_19),
.B2(n_28),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_49),
.A2(n_19),
.B1(n_28),
.B2(n_42),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_60),
.A2(n_19),
.B1(n_28),
.B2(n_42),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_46),
.B(n_38),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_91),
.B(n_97),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_69),
.B(n_29),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_50),
.A2(n_38),
.B1(n_34),
.B2(n_22),
.Y(n_94)
);

OAI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_48),
.A2(n_67),
.B1(n_52),
.B2(n_64),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_95),
.A2(n_63),
.B1(n_35),
.B2(n_3),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_44),
.B(n_33),
.Y(n_96)
);

OR2x2_ASAP7_75t_L g111 ( 
.A(n_96),
.B(n_98),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_59),
.B(n_34),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_45),
.B(n_33),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_68),
.A2(n_22),
.B1(n_21),
.B2(n_24),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_65),
.B(n_21),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_101),
.B(n_106),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_54),
.B(n_35),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_104),
.B(n_107),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_54),
.B(n_35),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_56),
.B(n_35),
.Y(n_107)
);

CKINVDCx14_ASAP7_75t_R g109 ( 
.A(n_101),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_109),
.B(n_123),
.Y(n_152)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_78),
.Y(n_110)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_110),
.Y(n_172)
);

INVx11_ASAP7_75t_L g113 ( 
.A(n_103),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_113),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_115),
.B(n_120),
.Y(n_160)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_87),
.Y(n_116)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_116),
.Y(n_149)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_87),
.Y(n_117)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_117),
.Y(n_154)
);

INVx1_ASAP7_75t_SL g120 ( 
.A(n_70),
.Y(n_120)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_105),
.Y(n_121)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_121),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_91),
.B(n_1),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_122),
.B(n_140),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_71),
.B(n_16),
.Y(n_123)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_89),
.Y(n_124)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_124),
.Y(n_167)
);

AND2x2_ASAP7_75t_SL g125 ( 
.A(n_97),
.B(n_2),
.Y(n_125)
);

AND2x2_ASAP7_75t_SL g158 ( 
.A(n_125),
.B(n_132),
.Y(n_158)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_89),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_126),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_93),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_127),
.A2(n_129),
.B1(n_133),
.B2(n_81),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_128),
.A2(n_104),
.B1(n_102),
.B2(n_72),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_93),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g130 ( 
.A(n_77),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_130),
.Y(n_157)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_75),
.Y(n_131)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_131),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_74),
.A2(n_5),
.B(n_7),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_82),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_71),
.B(n_9),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_134),
.B(n_138),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_70),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_135),
.Y(n_166)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_75),
.Y(n_136)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_136),
.Y(n_156)
);

AND2x2_ASAP7_75t_SL g137 ( 
.A(n_83),
.B(n_10),
.Y(n_137)
);

AND2x2_ASAP7_75t_SL g162 ( 
.A(n_137),
.B(n_100),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_74),
.B(n_10),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_82),
.B(n_96),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_139),
.B(n_106),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_76),
.B(n_12),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_99),
.B(n_12),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_141),
.B(n_98),
.Y(n_163)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_83),
.Y(n_143)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_143),
.Y(n_159)
);

OAI22x1_ASAP7_75t_L g147 ( 
.A1(n_118),
.A2(n_107),
.B1(n_81),
.B2(n_77),
.Y(n_147)
);

A2O1A1Ixp33_ASAP7_75t_SL g187 ( 
.A1(n_147),
.A2(n_129),
.B(n_127),
.C(n_133),
.Y(n_187)
);

O2A1O1Ixp33_ASAP7_75t_L g148 ( 
.A1(n_141),
.A2(n_100),
.B(n_107),
.C(n_104),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_148),
.A2(n_111),
.B(n_140),
.Y(n_190)
);

INVxp33_ASAP7_75t_L g150 ( 
.A(n_120),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_150),
.B(n_130),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_115),
.A2(n_90),
.B1(n_86),
.B2(n_89),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_153),
.A2(n_168),
.B1(n_170),
.B2(n_137),
.Y(n_179)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_131),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_161),
.B(n_163),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_162),
.B(n_125),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_165),
.B(n_119),
.Y(n_175)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_136),
.Y(n_169)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_169),
.Y(n_184)
);

MAJx2_ASAP7_75t_L g171 ( 
.A(n_112),
.B(n_86),
.C(n_108),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_171),
.B(n_125),
.C(n_137),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_112),
.A2(n_108),
.B1(n_102),
.B2(n_72),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_173),
.A2(n_142),
.B1(n_160),
.B2(n_118),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_174),
.B(n_175),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_176),
.A2(n_198),
.B1(n_90),
.B2(n_105),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_171),
.B(n_122),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_177),
.B(n_199),
.C(n_162),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_147),
.A2(n_132),
.B(n_139),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_178),
.A2(n_187),
.B(n_164),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_179),
.A2(n_172),
.B1(n_78),
.B2(n_103),
.Y(n_223)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_144),
.Y(n_180)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_180),
.Y(n_202)
);

BUFx2_ASAP7_75t_L g181 ( 
.A(n_144),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_181),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_160),
.A2(n_118),
.B(n_114),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_182),
.A2(n_166),
.B(n_164),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_183),
.B(n_170),
.Y(n_206)
);

OAI21xp33_ASAP7_75t_L g220 ( 
.A1(n_185),
.A2(n_191),
.B(n_150),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_163),
.B(n_114),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_186),
.B(n_197),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_151),
.B(n_138),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_188),
.B(n_201),
.Y(n_207)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_149),
.Y(n_189)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_189),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_190),
.A2(n_158),
.B(n_166),
.Y(n_208)
);

A2O1A1O1Ixp25_ASAP7_75t_L g191 ( 
.A1(n_151),
.A2(n_111),
.B(n_117),
.C(n_116),
.D(n_142),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_154),
.Y(n_192)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_192),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_152),
.B(n_110),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_193),
.B(n_194),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_159),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_145),
.B(n_126),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_195),
.B(n_196),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_157),
.B(n_158),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_162),
.B(n_143),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_160),
.A2(n_90),
.B1(n_105),
.B2(n_121),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_168),
.B(n_124),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_158),
.B(n_113),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_204),
.B(n_187),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_186),
.B(n_148),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_205),
.B(n_209),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_206),
.B(n_221),
.C(n_176),
.Y(n_229)
);

AOI221xp5_ASAP7_75t_L g230 ( 
.A1(n_208),
.A2(n_216),
.B1(n_220),
.B2(n_182),
.C(n_190),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_200),
.B(n_173),
.Y(n_209)
);

OAI21x1_ASAP7_75t_L g227 ( 
.A1(n_215),
.A2(n_197),
.B(n_185),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_177),
.B(n_156),
.Y(n_217)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_217),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_218),
.A2(n_146),
.B1(n_187),
.B2(n_215),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_183),
.B(n_155),
.C(n_167),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_178),
.A2(n_167),
.B(n_172),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_222),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_223),
.A2(n_198),
.B1(n_181),
.B2(n_180),
.Y(n_236)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_184),
.Y(n_224)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_224),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_227),
.A2(n_230),
.B(n_208),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_204),
.B(n_199),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_228),
.B(n_232),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_SL g245 ( 
.A(n_229),
.B(n_241),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_206),
.B(n_188),
.C(n_192),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_207),
.B(n_194),
.Y(n_233)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_233),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_210),
.Y(n_234)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_234),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_217),
.B(n_191),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_235),
.B(n_239),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_L g256 ( 
.A1(n_236),
.A2(n_211),
.B1(n_213),
.B2(n_224),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_209),
.A2(n_187),
.B1(n_184),
.B2(n_189),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_237),
.B(n_218),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_212),
.Y(n_238)
);

CKINVDCx14_ASAP7_75t_R g251 ( 
.A(n_238),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_240),
.A2(n_223),
.B1(n_225),
.B2(n_219),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_206),
.B(n_146),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_207),
.B(n_219),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_242),
.B(n_214),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_244),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_248),
.B(n_249),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_250),
.B(n_216),
.Y(n_259)
);

NOR3xp33_ASAP7_75t_SL g253 ( 
.A(n_243),
.B(n_205),
.C(n_210),
.Y(n_253)
);

NOR3xp33_ASAP7_75t_L g263 ( 
.A(n_253),
.B(n_203),
.C(n_232),
.Y(n_263)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_231),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_255),
.B(n_257),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_256),
.B(n_238),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_234),
.B(n_214),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_246),
.B(n_228),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_258),
.B(n_259),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_250),
.A2(n_225),
.B(n_239),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_260),
.A2(n_240),
.B(n_248),
.Y(n_271)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_262),
.Y(n_273)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_263),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_252),
.B(n_203),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_264),
.A2(n_266),
.B1(n_257),
.B2(n_251),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_253),
.B(n_212),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_245),
.B(n_229),
.C(n_241),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_268),
.B(n_246),
.C(n_254),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_258),
.B(n_245),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_269),
.B(n_274),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_270),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_271),
.B(n_276),
.Y(n_283)
);

INVx1_ASAP7_75t_SL g275 ( 
.A(n_267),
.Y(n_275)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_275),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_261),
.A2(n_247),
.B1(n_235),
.B2(n_226),
.Y(n_276)
);

AOI31xp33_ASAP7_75t_L g278 ( 
.A1(n_277),
.A2(n_260),
.A3(n_261),
.B(n_265),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_278),
.B(n_275),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_273),
.A2(n_247),
.B1(n_254),
.B2(n_255),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_279),
.B(n_280),
.Y(n_285)
);

CKINVDCx14_ASAP7_75t_R g280 ( 
.A(n_276),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_286),
.A2(n_288),
.B1(n_283),
.B2(n_221),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_281),
.B(n_274),
.C(n_272),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_287),
.B(n_289),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_282),
.A2(n_272),
.B1(n_271),
.B2(n_213),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_279),
.B(n_211),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_285),
.A2(n_284),
.B(n_281),
.Y(n_291)
);

NOR3xp33_ASAP7_75t_L g294 ( 
.A(n_291),
.B(n_287),
.C(n_221),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_292),
.A2(n_283),
.B(n_269),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_293),
.A2(n_294),
.B(n_290),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_295),
.A2(n_222),
.B(n_202),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_296),
.B(n_202),
.Y(n_297)
);


endmodule