module fake_netlist_1_4379_n_531 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_71, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_531);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_71;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_531;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_211;
wire n_334;
wire n_389;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_476;
wire n_105;
wire n_227;
wire n_384;
wire n_434;
wire n_231;
wire n_452;
wire n_518;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_73;
wire n_141;
wire n_119;
wire n_517;
wire n_479;
wire n_97;
wire n_167;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_502;
wire n_312;
wire n_455;
wire n_529;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_72;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_133;
wire n_149;
wire n_81;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_516;
wire n_254;
wire n_262;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_245;
wire n_357;
wire n_90;
wire n_260;
wire n_78;
wire n_201;
wire n_197;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_75;
wire n_376;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_520;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_497;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_74;
wire n_335;
wire n_272;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_418;
wire n_493;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_258;
wire n_253;
wire n_515;
wire n_266;
wire n_84;
wire n_213;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_494;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_109;
wire n_99;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx16_ASAP7_75t_R g72 ( .A(n_55), .Y(n_72) );
INVx1_ASAP7_75t_L g73 ( .A(n_22), .Y(n_73) );
INVx1_ASAP7_75t_L g74 ( .A(n_57), .Y(n_74) );
INVx1_ASAP7_75t_L g75 ( .A(n_36), .Y(n_75) );
INVx1_ASAP7_75t_L g76 ( .A(n_24), .Y(n_76) );
INVx2_ASAP7_75t_L g77 ( .A(n_53), .Y(n_77) );
INVxp67_ASAP7_75t_SL g78 ( .A(n_1), .Y(n_78) );
BUFx2_ASAP7_75t_L g79 ( .A(n_21), .Y(n_79) );
BUFx3_ASAP7_75t_L g80 ( .A(n_59), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_62), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_39), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_41), .Y(n_83) );
INVxp67_ASAP7_75t_SL g84 ( .A(n_71), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_45), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_48), .Y(n_86) );
HB1xp67_ASAP7_75t_L g87 ( .A(n_35), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_54), .Y(n_88) );
INVx2_ASAP7_75t_L g89 ( .A(n_56), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_25), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_33), .Y(n_91) );
CKINVDCx20_ASAP7_75t_R g92 ( .A(n_38), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_29), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_0), .Y(n_94) );
INVxp67_ASAP7_75t_SL g95 ( .A(n_65), .Y(n_95) );
INVxp67_ASAP7_75t_SL g96 ( .A(n_42), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_28), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_52), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_66), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_2), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_31), .Y(n_101) );
INVxp67_ASAP7_75t_L g102 ( .A(n_23), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_14), .Y(n_103) );
CKINVDCx20_ASAP7_75t_R g104 ( .A(n_30), .Y(n_104) );
AND3x2_ASAP7_75t_L g105 ( .A(n_79), .B(n_0), .C(n_1), .Y(n_105) );
BUFx6f_ASAP7_75t_L g106 ( .A(n_80), .Y(n_106) );
BUFx2_ASAP7_75t_L g107 ( .A(n_79), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_74), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_74), .Y(n_109) );
INVx2_ASAP7_75t_L g110 ( .A(n_77), .Y(n_110) );
HB1xp67_ASAP7_75t_L g111 ( .A(n_73), .Y(n_111) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_87), .B(n_2), .Y(n_112) );
INVx2_ASAP7_75t_L g113 ( .A(n_77), .Y(n_113) );
INVx2_ASAP7_75t_L g114 ( .A(n_77), .Y(n_114) );
BUFx6f_ASAP7_75t_L g115 ( .A(n_80), .Y(n_115) );
NAND2xp5_ASAP7_75t_L g116 ( .A(n_75), .B(n_76), .Y(n_116) );
NOR2xp33_ASAP7_75t_L g117 ( .A(n_75), .B(n_3), .Y(n_117) );
HB1xp67_ASAP7_75t_L g118 ( .A(n_73), .Y(n_118) );
INVx2_ASAP7_75t_L g119 ( .A(n_89), .Y(n_119) );
INVx2_ASAP7_75t_L g120 ( .A(n_89), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_76), .Y(n_121) );
CKINVDCx20_ASAP7_75t_R g122 ( .A(n_72), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_81), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_81), .Y(n_124) );
NAND2xp5_ASAP7_75t_L g125 ( .A(n_82), .B(n_3), .Y(n_125) );
BUFx6f_ASAP7_75t_L g126 ( .A(n_80), .Y(n_126) );
AND2x4_ASAP7_75t_L g127 ( .A(n_94), .B(n_4), .Y(n_127) );
AND2x2_ASAP7_75t_L g128 ( .A(n_72), .B(n_4), .Y(n_128) );
BUFx2_ASAP7_75t_L g129 ( .A(n_107), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_110), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_110), .Y(n_131) );
AND2x2_ASAP7_75t_L g132 ( .A(n_107), .B(n_103), .Y(n_132) );
AND2x4_ASAP7_75t_L g133 ( .A(n_127), .B(n_94), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_110), .Y(n_134) );
NAND2xp5_ASAP7_75t_SL g135 ( .A(n_108), .B(n_102), .Y(n_135) );
INVx2_ASAP7_75t_L g136 ( .A(n_106), .Y(n_136) );
INVx4_ASAP7_75t_L g137 ( .A(n_127), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_113), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_113), .Y(n_139) );
INVx1_ASAP7_75t_SL g140 ( .A(n_128), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_113), .Y(n_141) );
NAND2x1p5_ASAP7_75t_L g142 ( .A(n_127), .B(n_82), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_114), .Y(n_143) );
INVx6_ASAP7_75t_L g144 ( .A(n_106), .Y(n_144) );
AND2x4_ASAP7_75t_L g145 ( .A(n_127), .B(n_100), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g146 ( .A(n_108), .B(n_93), .Y(n_146) );
INVx1_ASAP7_75t_SL g147 ( .A(n_128), .Y(n_147) );
INVx5_ASAP7_75t_L g148 ( .A(n_106), .Y(n_148) );
INVxp67_ASAP7_75t_SL g149 ( .A(n_111), .Y(n_149) );
INVx5_ASAP7_75t_L g150 ( .A(n_106), .Y(n_150) );
INVx1_ASAP7_75t_SL g151 ( .A(n_122), .Y(n_151) );
NOR2xp33_ASAP7_75t_L g152 ( .A(n_116), .B(n_93), .Y(n_152) );
INVx4_ASAP7_75t_L g153 ( .A(n_106), .Y(n_153) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_126), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_114), .Y(n_155) );
AOI22x1_ASAP7_75t_L g156 ( .A1(n_109), .A2(n_89), .B1(n_85), .B2(n_101), .Y(n_156) );
BUFx2_ASAP7_75t_L g157 ( .A(n_149), .Y(n_157) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_154), .Y(n_158) );
INVx3_ASAP7_75t_L g159 ( .A(n_137), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_130), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_149), .B(n_118), .Y(n_161) );
AOI22xp33_ASAP7_75t_L g162 ( .A1(n_133), .A2(n_124), .B1(n_123), .B2(n_121), .Y(n_162) );
BUFx3_ASAP7_75t_L g163 ( .A(n_142), .Y(n_163) );
INVx1_ASAP7_75t_L g164 ( .A(n_130), .Y(n_164) );
BUFx2_ASAP7_75t_L g165 ( .A(n_129), .Y(n_165) );
OR2x2_ASAP7_75t_L g166 ( .A(n_129), .B(n_112), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_131), .Y(n_167) );
AOI22xp5_ASAP7_75t_L g168 ( .A1(n_140), .A2(n_92), .B1(n_104), .B2(n_117), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_131), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_134), .Y(n_170) );
BUFx3_ASAP7_75t_L g171 ( .A(n_142), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_134), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_138), .Y(n_173) );
INVx2_ASAP7_75t_SL g174 ( .A(n_142), .Y(n_174) );
BUFx2_ASAP7_75t_L g175 ( .A(n_140), .Y(n_175) );
CKINVDCx8_ASAP7_75t_R g176 ( .A(n_133), .Y(n_176) );
INVx2_ASAP7_75t_L g177 ( .A(n_136), .Y(n_177) );
NAND2x1p5_ASAP7_75t_L g178 ( .A(n_137), .B(n_109), .Y(n_178) );
BUFx6f_ASAP7_75t_L g179 ( .A(n_154), .Y(n_179) );
INVx2_ASAP7_75t_L g180 ( .A(n_136), .Y(n_180) );
AOI22xp5_ASAP7_75t_L g181 ( .A1(n_147), .A2(n_124), .B1(n_123), .B2(n_121), .Y(n_181) );
AND2x2_ASAP7_75t_SL g182 ( .A(n_137), .B(n_83), .Y(n_182) );
INVx1_ASAP7_75t_L g183 ( .A(n_138), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_139), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_139), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_141), .Y(n_186) );
BUFx6f_ASAP7_75t_L g187 ( .A(n_154), .Y(n_187) );
BUFx6f_ASAP7_75t_L g188 ( .A(n_154), .Y(n_188) );
NOR2xp33_ASAP7_75t_L g189 ( .A(n_135), .B(n_125), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_141), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_143), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_143), .Y(n_192) );
AOI21xp5_ASAP7_75t_L g193 ( .A1(n_160), .A2(n_133), .B(n_145), .Y(n_193) );
CKINVDCx20_ASAP7_75t_R g194 ( .A(n_165), .Y(n_194) );
INVx2_ASAP7_75t_SL g195 ( .A(n_174), .Y(n_195) );
INVx2_ASAP7_75t_L g196 ( .A(n_160), .Y(n_196) );
BUFx6f_ASAP7_75t_L g197 ( .A(n_163), .Y(n_197) );
AOI21xp5_ASAP7_75t_L g198 ( .A1(n_164), .A2(n_133), .B(n_145), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_164), .Y(n_199) );
BUFx2_ASAP7_75t_L g200 ( .A(n_163), .Y(n_200) );
AOI22xp5_ASAP7_75t_L g201 ( .A1(n_182), .A2(n_174), .B1(n_157), .B2(n_162), .Y(n_201) );
BUFx4f_ASAP7_75t_L g202 ( .A(n_178), .Y(n_202) );
INVx2_ASAP7_75t_L g203 ( .A(n_167), .Y(n_203) );
BUFx2_ASAP7_75t_L g204 ( .A(n_171), .Y(n_204) );
AND2x2_ASAP7_75t_L g205 ( .A(n_157), .B(n_147), .Y(n_205) );
OR2x6_ASAP7_75t_L g206 ( .A(n_171), .B(n_145), .Y(n_206) );
AND2x2_ASAP7_75t_L g207 ( .A(n_175), .B(n_132), .Y(n_207) );
BUFx2_ASAP7_75t_L g208 ( .A(n_165), .Y(n_208) );
AND2x2_ASAP7_75t_L g209 ( .A(n_175), .B(n_132), .Y(n_209) );
INVx2_ASAP7_75t_L g210 ( .A(n_167), .Y(n_210) );
AOI22xp33_ASAP7_75t_SL g211 ( .A1(n_182), .A2(n_156), .B1(n_145), .B2(n_78), .Y(n_211) );
AOI22xp5_ASAP7_75t_L g212 ( .A1(n_182), .A2(n_137), .B1(n_152), .B2(n_146), .Y(n_212) );
INVx2_ASAP7_75t_L g213 ( .A(n_169), .Y(n_213) );
BUFx12f_ASAP7_75t_L g214 ( .A(n_178), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_181), .B(n_146), .Y(n_215) );
INVx3_ASAP7_75t_L g216 ( .A(n_159), .Y(n_216) );
BUFx2_ASAP7_75t_L g217 ( .A(n_178), .Y(n_217) );
INVx2_ASAP7_75t_SL g218 ( .A(n_159), .Y(n_218) );
INVx1_ASAP7_75t_SL g219 ( .A(n_166), .Y(n_219) );
HB1xp67_ASAP7_75t_L g220 ( .A(n_176), .Y(n_220) );
AND2x2_ASAP7_75t_L g221 ( .A(n_161), .B(n_169), .Y(n_221) );
INVxp67_ASAP7_75t_SL g222 ( .A(n_181), .Y(n_222) );
AOI22xp33_ASAP7_75t_L g223 ( .A1(n_166), .A2(n_156), .B1(n_155), .B2(n_153), .Y(n_223) );
BUFx6f_ASAP7_75t_L g224 ( .A(n_176), .Y(n_224) );
AND2x2_ASAP7_75t_L g225 ( .A(n_170), .B(n_155), .Y(n_225) );
AOI221xp5_ASAP7_75t_L g226 ( .A1(n_189), .A2(n_100), .B1(n_103), .B2(n_119), .C(n_120), .Y(n_226) );
AOI22xp33_ASAP7_75t_L g227 ( .A1(n_219), .A2(n_168), .B1(n_159), .B2(n_151), .Y(n_227) );
INVx3_ASAP7_75t_L g228 ( .A(n_214), .Y(n_228) );
INVx8_ASAP7_75t_L g229 ( .A(n_214), .Y(n_229) );
INVx2_ASAP7_75t_L g230 ( .A(n_196), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_196), .Y(n_231) );
CKINVDCx11_ASAP7_75t_R g232 ( .A(n_194), .Y(n_232) );
OAI22xp33_ASAP7_75t_L g233 ( .A1(n_219), .A2(n_151), .B1(n_191), .B2(n_190), .Y(n_233) );
OAI22xp33_ASAP7_75t_L g234 ( .A1(n_214), .A2(n_192), .B1(n_191), .B2(n_190), .Y(n_234) );
AOI22xp33_ASAP7_75t_L g235 ( .A1(n_208), .A2(n_159), .B1(n_186), .B2(n_185), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_196), .Y(n_236) );
CKINVDCx14_ASAP7_75t_R g237 ( .A(n_208), .Y(n_237) );
AND2x2_ASAP7_75t_L g238 ( .A(n_221), .B(n_170), .Y(n_238) );
OAI22xp5_ASAP7_75t_L g239 ( .A1(n_222), .A2(n_192), .B1(n_184), .B2(n_183), .Y(n_239) );
A2O1A1Ixp33_ASAP7_75t_L g240 ( .A1(n_193), .A2(n_184), .B(n_172), .C(n_186), .Y(n_240) );
AOI22xp33_ASAP7_75t_L g241 ( .A1(n_207), .A2(n_172), .B1(n_173), .B2(n_185), .Y(n_241) );
INVx2_ASAP7_75t_SL g242 ( .A(n_202), .Y(n_242) );
OR2x2_ASAP7_75t_L g243 ( .A(n_205), .B(n_173), .Y(n_243) );
OAI22xp33_ASAP7_75t_L g244 ( .A1(n_201), .A2(n_183), .B1(n_105), .B2(n_85), .Y(n_244) );
OAI22xp33_ASAP7_75t_L g245 ( .A1(n_201), .A2(n_99), .B1(n_83), .B2(n_86), .Y(n_245) );
OR2x2_ASAP7_75t_L g246 ( .A(n_205), .B(n_114), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_203), .Y(n_247) );
INVx3_ASAP7_75t_L g248 ( .A(n_202), .Y(n_248) );
AND2x4_ASAP7_75t_L g249 ( .A(n_217), .B(n_86), .Y(n_249) );
BUFx6f_ASAP7_75t_L g250 ( .A(n_197), .Y(n_250) );
AOI221xp5_ASAP7_75t_L g251 ( .A1(n_207), .A2(n_119), .B1(n_120), .B2(n_90), .C(n_91), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_238), .B(n_221), .Y(n_252) );
AOI22xp33_ASAP7_75t_L g253 ( .A1(n_244), .A2(n_222), .B1(n_207), .B2(n_209), .Y(n_253) );
OAI22xp33_ASAP7_75t_L g254 ( .A1(n_229), .A2(n_202), .B1(n_212), .B2(n_206), .Y(n_254) );
AOI22xp33_ASAP7_75t_L g255 ( .A1(n_229), .A2(n_209), .B1(n_221), .B2(n_205), .Y(n_255) );
AOI22xp33_ASAP7_75t_L g256 ( .A1(n_229), .A2(n_209), .B1(n_211), .B2(n_220), .Y(n_256) );
CKINVDCx5p33_ASAP7_75t_R g257 ( .A(n_232), .Y(n_257) );
AOI22xp33_ASAP7_75t_L g258 ( .A1(n_229), .A2(n_211), .B1(n_224), .B2(n_202), .Y(n_258) );
HB1xp67_ASAP7_75t_L g259 ( .A(n_237), .Y(n_259) );
AOI221xp5_ASAP7_75t_L g260 ( .A1(n_245), .A2(n_226), .B1(n_215), .B2(n_212), .C(n_199), .Y(n_260) );
OAI22xp33_ASAP7_75t_L g261 ( .A1(n_229), .A2(n_206), .B1(n_224), .B2(n_217), .Y(n_261) );
OAI22xp5_ASAP7_75t_L g262 ( .A1(n_239), .A2(n_215), .B1(n_210), .B2(n_203), .Y(n_262) );
INVx2_ASAP7_75t_SL g263 ( .A(n_228), .Y(n_263) );
AOI221xp5_ASAP7_75t_L g264 ( .A1(n_233), .A2(n_226), .B1(n_199), .B2(n_193), .C(n_198), .Y(n_264) );
AOI221xp5_ASAP7_75t_L g265 ( .A1(n_239), .A2(n_198), .B1(n_223), .B2(n_225), .C(n_213), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_231), .Y(n_266) );
AOI22xp33_ASAP7_75t_SL g267 ( .A1(n_228), .A2(n_224), .B1(n_204), .B2(n_200), .Y(n_267) );
AO31x2_ASAP7_75t_L g268 ( .A1(n_240), .A2(n_203), .A3(n_210), .B(n_213), .Y(n_268) );
AND2x2_ASAP7_75t_L g269 ( .A(n_238), .B(n_225), .Y(n_269) );
AND2x2_ASAP7_75t_L g270 ( .A(n_231), .B(n_225), .Y(n_270) );
AOI22xp33_ASAP7_75t_L g271 ( .A1(n_249), .A2(n_224), .B1(n_206), .B2(n_210), .Y(n_271) );
AND2x4_ASAP7_75t_L g272 ( .A(n_248), .B(n_213), .Y(n_272) );
BUFx2_ASAP7_75t_L g273 ( .A(n_262), .Y(n_273) );
INVx1_ASAP7_75t_SL g274 ( .A(n_270), .Y(n_274) );
INVx2_ASAP7_75t_L g275 ( .A(n_268), .Y(n_275) );
AOI211xp5_ASAP7_75t_SL g276 ( .A1(n_254), .A2(n_234), .B(n_228), .C(n_248), .Y(n_276) );
INVx2_ASAP7_75t_L g277 ( .A(n_268), .Y(n_277) );
OAI211xp5_ASAP7_75t_L g278 ( .A1(n_253), .A2(n_227), .B(n_251), .C(n_241), .Y(n_278) );
AND2x2_ASAP7_75t_L g279 ( .A(n_270), .B(n_236), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_266), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_266), .Y(n_281) );
OAI22xp5_ASAP7_75t_L g282 ( .A1(n_262), .A2(n_243), .B1(n_247), .B2(n_236), .Y(n_282) );
OAI21x1_ASAP7_75t_L g283 ( .A1(n_265), .A2(n_230), .B(n_247), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_268), .Y(n_284) );
INVx2_ASAP7_75t_L g285 ( .A(n_268), .Y(n_285) );
NOR2xp33_ASAP7_75t_L g286 ( .A(n_259), .B(n_249), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_268), .Y(n_287) );
OAI33xp33_ASAP7_75t_L g288 ( .A1(n_261), .A2(n_88), .A3(n_90), .B1(n_91), .B2(n_97), .B3(n_98), .Y(n_288) );
INVx2_ASAP7_75t_L g289 ( .A(n_272), .Y(n_289) );
OAI211xp5_ASAP7_75t_L g290 ( .A1(n_255), .A2(n_235), .B(n_243), .C(n_204), .Y(n_290) );
NOR2xp33_ASAP7_75t_L g291 ( .A(n_252), .B(n_249), .Y(n_291) );
NAND4xp25_ASAP7_75t_SL g292 ( .A(n_256), .B(n_246), .C(n_230), .D(n_98), .Y(n_292) );
AOI21xp33_ASAP7_75t_L g293 ( .A1(n_264), .A2(n_249), .B(n_246), .Y(n_293) );
INVxp67_ASAP7_75t_SL g294 ( .A(n_252), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_269), .Y(n_295) );
OAI22xp5_ASAP7_75t_L g296 ( .A1(n_260), .A2(n_206), .B1(n_224), .B2(n_200), .Y(n_296) );
NOR2xp33_ASAP7_75t_L g297 ( .A(n_286), .B(n_257), .Y(n_297) );
AND2x4_ASAP7_75t_L g298 ( .A(n_289), .B(n_272), .Y(n_298) );
AND2x2_ASAP7_75t_L g299 ( .A(n_279), .B(n_269), .Y(n_299) );
AOI221xp5_ASAP7_75t_L g300 ( .A1(n_291), .A2(n_263), .B1(n_99), .B2(n_88), .C(n_101), .Y(n_300) );
AOI221xp5_ASAP7_75t_L g301 ( .A1(n_295), .A2(n_263), .B1(n_97), .B2(n_257), .C(n_258), .Y(n_301) );
AND2x2_ASAP7_75t_L g302 ( .A(n_279), .B(n_272), .Y(n_302) );
AO21x2_ASAP7_75t_L g303 ( .A1(n_282), .A2(n_272), .B(n_136), .Y(n_303) );
AND2x2_ASAP7_75t_L g304 ( .A(n_274), .B(n_271), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_280), .Y(n_305) );
INVx2_ASAP7_75t_L g306 ( .A(n_275), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_280), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_295), .B(n_267), .Y(n_308) );
AOI221xp5_ASAP7_75t_L g309 ( .A1(n_288), .A2(n_84), .B1(n_96), .B2(n_95), .C(n_126), .Y(n_309) );
NAND4xp25_ASAP7_75t_L g310 ( .A(n_276), .B(n_153), .C(n_248), .D(n_7), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_281), .Y(n_311) );
AOI31xp33_ASAP7_75t_SL g312 ( .A1(n_293), .A2(n_5), .A3(n_6), .B(n_7), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_281), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_284), .Y(n_314) );
NAND4xp25_ASAP7_75t_L g315 ( .A(n_276), .B(n_153), .C(n_6), .D(n_8), .Y(n_315) );
INVx2_ASAP7_75t_L g316 ( .A(n_275), .Y(n_316) );
NAND3xp33_ASAP7_75t_SL g317 ( .A(n_290), .B(n_5), .C(n_8), .Y(n_317) );
AOI31xp33_ASAP7_75t_L g318 ( .A1(n_290), .A2(n_242), .A3(n_195), .B(n_11), .Y(n_318) );
AND2x2_ASAP7_75t_L g319 ( .A(n_274), .B(n_250), .Y(n_319) );
AND2x2_ASAP7_75t_L g320 ( .A(n_289), .B(n_250), .Y(n_320) );
OAI222xp33_ASAP7_75t_L g321 ( .A1(n_296), .A2(n_242), .B1(n_206), .B2(n_195), .C1(n_12), .C2(n_13), .Y(n_321) );
AND2x2_ASAP7_75t_L g322 ( .A(n_289), .B(n_250), .Y(n_322) );
OAI33xp33_ASAP7_75t_L g323 ( .A1(n_282), .A2(n_9), .A3(n_10), .B1(n_11), .B2(n_12), .B3(n_13), .Y(n_323) );
AO21x2_ASAP7_75t_L g324 ( .A1(n_284), .A2(n_177), .B(n_180), .Y(n_324) );
OAI211xp5_ASAP7_75t_L g325 ( .A1(n_278), .A2(n_224), .B(n_106), .C(n_126), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_287), .Y(n_326) );
INVx2_ASAP7_75t_L g327 ( .A(n_275), .Y(n_327) );
INVx2_ASAP7_75t_SL g328 ( .A(n_283), .Y(n_328) );
OAI22xp5_ASAP7_75t_L g329 ( .A1(n_296), .A2(n_206), .B1(n_224), .B2(n_195), .Y(n_329) );
NAND2x1p5_ASAP7_75t_SL g330 ( .A(n_277), .B(n_218), .Y(n_330) );
OR2x2_ASAP7_75t_L g331 ( .A(n_294), .B(n_250), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_287), .Y(n_332) );
AND3x1_ASAP7_75t_L g333 ( .A(n_297), .B(n_292), .C(n_10), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_305), .Y(n_334) );
NAND3xp33_ASAP7_75t_L g335 ( .A(n_315), .B(n_115), .C(n_126), .Y(n_335) );
NAND4xp25_ASAP7_75t_L g336 ( .A(n_315), .B(n_273), .C(n_293), .D(n_278), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_299), .B(n_273), .Y(n_337) );
AND2x4_ASAP7_75t_L g338 ( .A(n_314), .B(n_285), .Y(n_338) );
AND2x2_ASAP7_75t_L g339 ( .A(n_305), .B(n_277), .Y(n_339) );
NOR2xp33_ASAP7_75t_L g340 ( .A(n_318), .B(n_292), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_307), .Y(n_341) );
INVx2_ASAP7_75t_L g342 ( .A(n_306), .Y(n_342) );
OR2x2_ASAP7_75t_L g343 ( .A(n_299), .B(n_277), .Y(n_343) );
OR2x2_ASAP7_75t_L g344 ( .A(n_302), .B(n_285), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_307), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_311), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_311), .Y(n_347) );
NAND4xp25_ASAP7_75t_L g348 ( .A(n_310), .B(n_285), .C(n_153), .D(n_15), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_313), .Y(n_349) );
INVx2_ASAP7_75t_SL g350 ( .A(n_331), .Y(n_350) );
OR2x2_ASAP7_75t_L g351 ( .A(n_302), .B(n_283), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_313), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_314), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_308), .B(n_283), .Y(n_354) );
OR2x6_ASAP7_75t_L g355 ( .A(n_329), .B(n_250), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_326), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_326), .Y(n_357) );
INVx2_ASAP7_75t_SL g358 ( .A(n_331), .Y(n_358) );
AND2x2_ASAP7_75t_L g359 ( .A(n_304), .B(n_9), .Y(n_359) );
OAI33xp33_ASAP7_75t_L g360 ( .A1(n_310), .A2(n_14), .A3(n_15), .B1(n_16), .B2(n_17), .B3(n_18), .Y(n_360) );
INVx2_ASAP7_75t_L g361 ( .A(n_306), .Y(n_361) );
INVx4_ASAP7_75t_L g362 ( .A(n_303), .Y(n_362) );
INVx1_ASAP7_75t_SL g363 ( .A(n_319), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_304), .B(n_16), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_332), .Y(n_365) );
AND2x2_ASAP7_75t_L g366 ( .A(n_298), .B(n_17), .Y(n_366) );
AND2x2_ASAP7_75t_L g367 ( .A(n_298), .B(n_18), .Y(n_367) );
OR2x2_ASAP7_75t_L g368 ( .A(n_330), .B(n_19), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_332), .Y(n_369) );
OR2x2_ASAP7_75t_L g370 ( .A(n_330), .B(n_19), .Y(n_370) );
BUFx2_ASAP7_75t_L g371 ( .A(n_330), .Y(n_371) );
INVxp67_ASAP7_75t_L g372 ( .A(n_303), .Y(n_372) );
AND2x2_ASAP7_75t_L g373 ( .A(n_306), .B(n_327), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_319), .B(n_20), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_298), .B(n_20), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_316), .Y(n_376) );
INVx2_ASAP7_75t_L g377 ( .A(n_316), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_298), .B(n_21), .Y(n_378) );
INVxp67_ASAP7_75t_L g379 ( .A(n_303), .Y(n_379) );
OAI21xp33_ASAP7_75t_L g380 ( .A1(n_317), .A2(n_126), .B(n_115), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_316), .Y(n_381) );
AND2x2_ASAP7_75t_L g382 ( .A(n_363), .B(n_322), .Y(n_382) );
OAI21xp33_ASAP7_75t_L g383 ( .A1(n_348), .A2(n_328), .B(n_325), .Y(n_383) );
INVx1_ASAP7_75t_SL g384 ( .A(n_343), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_337), .B(n_327), .Y(n_385) );
OR2x2_ASAP7_75t_L g386 ( .A(n_344), .B(n_327), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_334), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_341), .Y(n_388) );
NAND2xp5_ASAP7_75t_SL g389 ( .A(n_371), .B(n_328), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_359), .B(n_322), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_345), .Y(n_391) );
NOR2xp33_ASAP7_75t_SL g392 ( .A(n_340), .B(n_321), .Y(n_392) );
NAND4xp25_ASAP7_75t_L g393 ( .A(n_340), .B(n_336), .C(n_364), .D(n_335), .Y(n_393) );
AND2x2_ASAP7_75t_L g394 ( .A(n_350), .B(n_358), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_350), .B(n_320), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_358), .B(n_320), .Y(n_396) );
AO21x1_ASAP7_75t_L g397 ( .A1(n_362), .A2(n_312), .B(n_323), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_346), .B(n_324), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_347), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_349), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_352), .Y(n_401) );
NAND3xp33_ASAP7_75t_L g402 ( .A(n_372), .B(n_309), .C(n_300), .Y(n_402) );
AOI21xp33_ASAP7_75t_SL g403 ( .A1(n_368), .A2(n_22), .B(n_312), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_353), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_356), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_357), .Y(n_406) );
AND2x2_ASAP7_75t_L g407 ( .A(n_351), .B(n_339), .Y(n_407) );
INVx1_ASAP7_75t_SL g408 ( .A(n_366), .Y(n_408) );
INVxp67_ASAP7_75t_L g409 ( .A(n_370), .Y(n_409) );
INVx2_ASAP7_75t_L g410 ( .A(n_373), .Y(n_410) );
INVx1_ASAP7_75t_SL g411 ( .A(n_367), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_365), .Y(n_412) );
HB1xp67_ASAP7_75t_L g413 ( .A(n_373), .Y(n_413) );
OR2x2_ASAP7_75t_L g414 ( .A(n_369), .B(n_324), .Y(n_414) );
NOR2xp33_ASAP7_75t_L g415 ( .A(n_360), .B(n_288), .Y(n_415) );
INVx2_ASAP7_75t_SL g416 ( .A(n_339), .Y(n_416) );
NAND2xp33_ASAP7_75t_L g417 ( .A(n_380), .B(n_301), .Y(n_417) );
AND2x2_ASAP7_75t_L g418 ( .A(n_338), .B(n_324), .Y(n_418) );
INVx2_ASAP7_75t_L g419 ( .A(n_342), .Y(n_419) );
INVx2_ASAP7_75t_L g420 ( .A(n_342), .Y(n_420) );
NAND2x1p5_ASAP7_75t_L g421 ( .A(n_333), .B(n_197), .Y(n_421) );
INVx2_ASAP7_75t_L g422 ( .A(n_361), .Y(n_422) );
AOI221xp5_ASAP7_75t_L g423 ( .A1(n_360), .A2(n_115), .B1(n_126), .B2(n_154), .C(n_197), .Y(n_423) );
AOI22xp5_ASAP7_75t_L g424 ( .A1(n_375), .A2(n_197), .B1(n_115), .B2(n_218), .Y(n_424) );
OAI33xp33_ASAP7_75t_L g425 ( .A1(n_372), .A2(n_115), .A3(n_27), .B1(n_32), .B2(n_34), .B3(n_37), .Y(n_425) );
AOI211xp5_ASAP7_75t_L g426 ( .A1(n_374), .A2(n_115), .B(n_197), .C(n_154), .Y(n_426) );
OR2x2_ASAP7_75t_L g427 ( .A(n_376), .B(n_197), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_354), .B(n_197), .Y(n_428) );
NOR2xp33_ASAP7_75t_L g429 ( .A(n_378), .B(n_26), .Y(n_429) );
OR2x2_ASAP7_75t_L g430 ( .A(n_381), .B(n_40), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_338), .B(n_150), .Y(n_431) );
OR2x6_ASAP7_75t_L g432 ( .A(n_355), .B(n_218), .Y(n_432) );
OAI33xp33_ASAP7_75t_L g433 ( .A1(n_409), .A2(n_379), .A3(n_377), .B1(n_361), .B2(n_362), .B3(n_338), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_387), .Y(n_434) );
INVx2_ASAP7_75t_SL g435 ( .A(n_394), .Y(n_435) );
XOR2xp5_ASAP7_75t_L g436 ( .A(n_390), .B(n_377), .Y(n_436) );
XOR2xp5_ASAP7_75t_L g437 ( .A(n_393), .B(n_43), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_409), .B(n_379), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_388), .Y(n_439) );
NOR2xp33_ASAP7_75t_L g440 ( .A(n_392), .B(n_362), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_384), .B(n_355), .Y(n_441) );
HB1xp67_ASAP7_75t_L g442 ( .A(n_413), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_391), .Y(n_443) );
XNOR2xp5_ASAP7_75t_L g444 ( .A(n_408), .B(n_355), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_399), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_413), .B(n_150), .Y(n_446) );
NOR2x1_ASAP7_75t_L g447 ( .A(n_389), .B(n_216), .Y(n_447) );
INVxp67_ASAP7_75t_L g448 ( .A(n_389), .Y(n_448) );
AOI22xp5_ASAP7_75t_L g449 ( .A1(n_415), .A2(n_144), .B1(n_216), .B2(n_148), .Y(n_449) );
NAND2xp5_ASAP7_75t_SL g450 ( .A(n_423), .B(n_148), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_407), .B(n_150), .Y(n_451) );
NAND3xp33_ASAP7_75t_L g452 ( .A(n_423), .B(n_148), .C(n_150), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_400), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_401), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_404), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_405), .Y(n_456) );
AOI22xp5_ASAP7_75t_L g457 ( .A1(n_415), .A2(n_144), .B1(n_216), .B2(n_148), .Y(n_457) );
INVx1_ASAP7_75t_SL g458 ( .A(n_411), .Y(n_458) );
AO22x1_ASAP7_75t_L g459 ( .A1(n_416), .A2(n_216), .B1(n_150), .B2(n_148), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_385), .B(n_150), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_406), .Y(n_461) );
NOR2xp33_ASAP7_75t_L g462 ( .A(n_403), .B(n_44), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_412), .B(n_150), .Y(n_463) );
OR2x2_ASAP7_75t_L g464 ( .A(n_386), .B(n_46), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_395), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_410), .B(n_148), .Y(n_466) );
NOR2x1_ASAP7_75t_L g467 ( .A(n_432), .B(n_47), .Y(n_467) );
INVx1_ASAP7_75t_SL g468 ( .A(n_382), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_396), .Y(n_469) );
INVxp33_ASAP7_75t_L g470 ( .A(n_421), .Y(n_470) );
INVxp67_ASAP7_75t_L g471 ( .A(n_398), .Y(n_471) );
XNOR2x2_ASAP7_75t_SL g472 ( .A(n_418), .B(n_49), .Y(n_472) );
XOR2x2_ASAP7_75t_L g473 ( .A(n_421), .B(n_50), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_414), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_420), .B(n_148), .Y(n_475) );
AOI221xp5_ASAP7_75t_L g476 ( .A1(n_397), .A2(n_180), .B1(n_177), .B2(n_188), .C(n_179), .Y(n_476) );
AOI22x1_ASAP7_75t_L g477 ( .A1(n_430), .A2(n_51), .B1(n_58), .B2(n_60), .Y(n_477) );
NOR2x1_ASAP7_75t_L g478 ( .A(n_432), .B(n_61), .Y(n_478) );
INVxp67_ASAP7_75t_L g479 ( .A(n_425), .Y(n_479) );
INVxp67_ASAP7_75t_L g480 ( .A(n_425), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_420), .B(n_144), .Y(n_481) );
OAI211xp5_ASAP7_75t_L g482 ( .A1(n_383), .A2(n_63), .B(n_64), .C(n_67), .Y(n_482) );
A2O1A1Ixp33_ASAP7_75t_L g483 ( .A1(n_417), .A2(n_68), .B(n_69), .C(n_70), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_422), .Y(n_484) );
OAI21xp5_ASAP7_75t_L g485 ( .A1(n_417), .A2(n_144), .B(n_158), .Y(n_485) );
NAND2x1p5_ASAP7_75t_L g486 ( .A(n_427), .B(n_158), .Y(n_486) );
OR2x2_ASAP7_75t_L g487 ( .A(n_419), .B(n_158), .Y(n_487) );
INVx2_ASAP7_75t_L g488 ( .A(n_422), .Y(n_488) );
AOI22xp5_ASAP7_75t_SL g489 ( .A1(n_429), .A2(n_158), .B1(n_179), .B2(n_187), .Y(n_489) );
XNOR2xp5_ASAP7_75t_L g490 ( .A(n_402), .B(n_144), .Y(n_490) );
NOR2xp33_ASAP7_75t_L g491 ( .A(n_429), .B(n_158), .Y(n_491) );
INVx2_ASAP7_75t_L g492 ( .A(n_432), .Y(n_492) );
AOI22xp5_ASAP7_75t_L g493 ( .A1(n_426), .A2(n_179), .B1(n_187), .B2(n_188), .Y(n_493) );
AOI222xp33_ASAP7_75t_L g494 ( .A1(n_428), .A2(n_179), .B1(n_187), .B2(n_188), .C1(n_431), .C2(n_424), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_387), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_409), .B(n_188), .Y(n_496) );
A2O1A1Ixp33_ASAP7_75t_L g497 ( .A1(n_440), .A2(n_470), .B(n_480), .C(n_479), .Y(n_497) );
AOI321xp33_ASAP7_75t_L g498 ( .A1(n_462), .A2(n_438), .A3(n_469), .B1(n_465), .B2(n_492), .C(n_476), .Y(n_498) );
XNOR2x1_ASAP7_75t_L g499 ( .A(n_473), .B(n_458), .Y(n_499) );
AOI21xp33_ASAP7_75t_L g500 ( .A1(n_490), .A2(n_479), .B(n_480), .Y(n_500) );
OAI311xp33_ASAP7_75t_L g501 ( .A1(n_448), .A2(n_472), .A3(n_457), .B1(n_449), .C1(n_494), .Y(n_501) );
AOI22xp5_ASAP7_75t_L g502 ( .A1(n_448), .A2(n_435), .B1(n_436), .B2(n_437), .Y(n_502) );
OAI221xp5_ASAP7_75t_L g503 ( .A1(n_442), .A2(n_444), .B1(n_471), .B2(n_482), .C(n_462), .Y(n_503) );
XNOR2xp5_ASAP7_75t_L g504 ( .A(n_472), .B(n_468), .Y(n_504) );
OAI221xp5_ASAP7_75t_L g505 ( .A1(n_442), .A2(n_471), .B1(n_482), .B2(n_474), .C(n_467), .Y(n_505) );
AOI21xp5_ASAP7_75t_SL g506 ( .A1(n_450), .A2(n_452), .B(n_483), .Y(n_506) );
AOI22xp33_ASAP7_75t_L g507 ( .A1(n_433), .A2(n_451), .B1(n_441), .B2(n_445), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_443), .B(n_495), .Y(n_508) );
INVxp33_ASAP7_75t_SL g509 ( .A(n_478), .Y(n_509) );
OAI31xp33_ASAP7_75t_L g510 ( .A1(n_461), .A2(n_455), .A3(n_454), .B(n_453), .Y(n_510) );
OAI21xp5_ASAP7_75t_SL g511 ( .A1(n_447), .A2(n_493), .B(n_485), .Y(n_511) );
BUFx3_ASAP7_75t_L g512 ( .A(n_499), .Y(n_512) );
AO22x2_ASAP7_75t_L g513 ( .A1(n_508), .A2(n_434), .B1(n_439), .B2(n_456), .Y(n_513) );
AOI311xp33_ASAP7_75t_L g514 ( .A1(n_500), .A2(n_484), .A3(n_446), .B(n_463), .C(n_433), .Y(n_514) );
INVx2_ASAP7_75t_SL g515 ( .A(n_504), .Y(n_515) );
AO22x2_ASAP7_75t_L g516 ( .A1(n_507), .A2(n_464), .B1(n_488), .B2(n_496), .Y(n_516) );
AOI21xp5_ASAP7_75t_L g517 ( .A1(n_497), .A2(n_459), .B(n_489), .Y(n_517) );
AOI22xp33_ASAP7_75t_SL g518 ( .A1(n_509), .A2(n_477), .B1(n_460), .B2(n_491), .Y(n_518) );
AOI22xp5_ASAP7_75t_L g519 ( .A1(n_503), .A2(n_497), .B1(n_502), .B2(n_507), .Y(n_519) );
NAND5xp2_ASAP7_75t_L g520 ( .A(n_519), .B(n_498), .C(n_505), .D(n_511), .E(n_501), .Y(n_520) );
XOR2xp5_ASAP7_75t_L g521 ( .A(n_512), .B(n_466), .Y(n_521) );
NOR2xp67_ASAP7_75t_L g522 ( .A(n_517), .B(n_510), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_513), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_523), .Y(n_524) );
AOI22xp5_ASAP7_75t_L g525 ( .A1(n_522), .A2(n_515), .B1(n_516), .B2(n_513), .Y(n_525) );
NAND4xp75_ASAP7_75t_L g526 ( .A(n_525), .B(n_520), .C(n_514), .D(n_521), .Y(n_526) );
NAND2xp5_ASAP7_75t_SL g527 ( .A(n_524), .B(n_518), .Y(n_527) );
OAI22xp5_ASAP7_75t_SL g528 ( .A1(n_526), .A2(n_521), .B1(n_506), .B2(n_486), .Y(n_528) );
INVx2_ASAP7_75t_L g529 ( .A(n_528), .Y(n_529) );
AOI22xp5_ASAP7_75t_L g530 ( .A1(n_529), .A2(n_527), .B1(n_475), .B2(n_481), .Y(n_530) );
AOI221xp5_ASAP7_75t_L g531 ( .A1(n_530), .A2(n_486), .B1(n_487), .B2(n_188), .C(n_179), .Y(n_531) );
endmodule