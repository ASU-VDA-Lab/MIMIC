module fake_jpeg_2066_n_569 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_569);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_569;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx11_ASAP7_75t_R g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

CKINVDCx16_ASAP7_75t_R g27 ( 
.A(n_13),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_1),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_9),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_3),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_15),
.Y(n_40)
);

INVx13_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_4),
.Y(n_43)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_8),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_2),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_6),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_14),
.Y(n_47)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_9),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_10),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_7),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_9),
.Y(n_51)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_12),
.Y(n_52)
);

BUFx10_ASAP7_75t_L g53 ( 
.A(n_2),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_1),
.Y(n_54)
);

BUFx12_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g116 ( 
.A(n_55),
.Y(n_116)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

INVx11_ASAP7_75t_L g110 ( 
.A(n_56),
.Y(n_110)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_57),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_20),
.B(n_8),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_58),
.B(n_66),
.Y(n_163)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_59),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_19),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_60),
.Y(n_148)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_61),
.Y(n_121)
);

OR2x2_ASAP7_75t_L g62 ( 
.A(n_24),
.B(n_8),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_62),
.B(n_99),
.Y(n_130)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_18),
.Y(n_63)
);

INVx8_ASAP7_75t_L g132 ( 
.A(n_63),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_19),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_64),
.Y(n_153)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_65),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_20),
.B(n_8),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_24),
.Y(n_67)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_67),
.Y(n_139)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_24),
.Y(n_68)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_68),
.Y(n_169)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_69),
.Y(n_140)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_70),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_21),
.B(n_9),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_71),
.B(n_28),
.Y(n_113)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_72),
.Y(n_118)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_73),
.Y(n_129)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_52),
.Y(n_74)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_74),
.Y(n_146)
);

BUFx4f_ASAP7_75t_L g75 ( 
.A(n_52),
.Y(n_75)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_75),
.Y(n_147)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_19),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_76),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_19),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_77),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_26),
.A2(n_7),
.B1(n_16),
.B2(n_15),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_78),
.A2(n_25),
.B1(n_36),
.B2(n_47),
.Y(n_144)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_52),
.Y(n_79)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_79),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_26),
.Y(n_80)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_80),
.Y(n_123)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_22),
.Y(n_81)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_81),
.Y(n_167)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_22),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_82),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_37),
.B(n_28),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_83),
.B(n_106),
.Y(n_135)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_33),
.Y(n_84)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_84),
.Y(n_120)
);

BUFx2_ASAP7_75t_L g85 ( 
.A(n_22),
.Y(n_85)
);

INVx3_ASAP7_75t_SL g117 ( 
.A(n_85),
.Y(n_117)
);

INVx11_ASAP7_75t_L g86 ( 
.A(n_46),
.Y(n_86)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_86),
.Y(n_131)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_46),
.Y(n_87)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_87),
.Y(n_155)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_46),
.Y(n_88)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_88),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_26),
.Y(n_89)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_89),
.Y(n_124)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_33),
.Y(n_90)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_90),
.Y(n_157)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_46),
.Y(n_91)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_91),
.Y(n_159)
);

BUFx10_ASAP7_75t_L g92 ( 
.A(n_53),
.Y(n_92)
);

INVx5_ASAP7_75t_L g166 ( 
.A(n_92),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_26),
.Y(n_93)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_93),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_30),
.Y(n_94)
);

INVx6_ASAP7_75t_L g143 ( 
.A(n_94),
.Y(n_143)
);

INVx6_ASAP7_75t_SL g95 ( 
.A(n_41),
.Y(n_95)
);

INVx6_ASAP7_75t_SL g152 ( 
.A(n_95),
.Y(n_152)
);

BUFx5_ASAP7_75t_L g96 ( 
.A(n_49),
.Y(n_96)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_96),
.Y(n_170)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_23),
.Y(n_97)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_97),
.Y(n_174)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_54),
.Y(n_98)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_98),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_27),
.B(n_7),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_30),
.Y(n_100)
);

INVx6_ASAP7_75t_L g177 ( 
.A(n_100),
.Y(n_177)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_54),
.Y(n_101)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_101),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_53),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_102),
.B(n_34),
.Y(n_133)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_49),
.Y(n_103)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_103),
.Y(n_173)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_54),
.Y(n_104)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_104),
.Y(n_178)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_30),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_105),
.B(n_109),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_37),
.B(n_10),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_30),
.Y(n_107)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_107),
.Y(n_175)
);

BUFx5_ASAP7_75t_L g108 ( 
.A(n_27),
.Y(n_108)
);

INVx5_ASAP7_75t_SL g136 ( 
.A(n_108),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_38),
.Y(n_109)
);

OAI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_62),
.A2(n_50),
.B1(n_38),
.B2(n_54),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_111),
.A2(n_112),
.B1(n_115),
.B2(n_126),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_60),
.A2(n_34),
.B1(n_38),
.B2(n_50),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_113),
.B(n_128),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_99),
.A2(n_38),
.B1(n_50),
.B2(n_36),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_63),
.A2(n_44),
.B1(n_103),
.B2(n_84),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_125),
.A2(n_75),
.B1(n_86),
.B2(n_56),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_64),
.A2(n_34),
.B1(n_50),
.B2(n_51),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_81),
.B(n_18),
.C(n_21),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_127),
.B(n_133),
.Y(n_182)
);

OR2x2_ASAP7_75t_L g128 ( 
.A(n_73),
.B(n_23),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_74),
.A2(n_25),
.B1(n_29),
.B2(n_47),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_137),
.A2(n_144),
.B1(n_156),
.B2(n_171),
.Y(n_213)
);

OR2x2_ASAP7_75t_L g142 ( 
.A(n_63),
.B(n_23),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_142),
.B(n_150),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_85),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_82),
.B(n_29),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_151),
.B(n_158),
.Y(n_194)
);

OAI22xp33_ASAP7_75t_L g156 ( 
.A1(n_76),
.A2(n_44),
.B1(n_51),
.B2(n_32),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_57),
.B(n_40),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_90),
.B(n_40),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_160),
.B(n_165),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_88),
.B(n_105),
.C(n_55),
.Y(n_162)
);

NAND2x1_ASAP7_75t_L g235 ( 
.A(n_162),
.B(n_92),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_55),
.B(n_51),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_L g171 ( 
.A1(n_77),
.A2(n_32),
.B1(n_35),
.B2(n_44),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_L g172 ( 
.A1(n_80),
.A2(n_109),
.B1(n_107),
.B2(n_100),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_172),
.A2(n_94),
.B1(n_93),
.B2(n_89),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_148),
.Y(n_179)
);

INVx6_ASAP7_75t_L g264 ( 
.A(n_179),
.Y(n_264)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_147),
.Y(n_180)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_180),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_181),
.Y(n_244)
);

INVx6_ASAP7_75t_L g184 ( 
.A(n_148),
.Y(n_184)
);

BUFx2_ASAP7_75t_L g265 ( 
.A(n_184),
.Y(n_265)
);

BUFx12f_ASAP7_75t_L g185 ( 
.A(n_152),
.Y(n_185)
);

INVx1_ASAP7_75t_SL g298 ( 
.A(n_185),
.Y(n_298)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_161),
.Y(n_186)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_186),
.Y(n_259)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_132),
.Y(n_188)
);

INVx4_ASAP7_75t_L g288 ( 
.A(n_188),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_163),
.B(n_35),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_189),
.B(n_211),
.Y(n_249)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_174),
.Y(n_190)
);

BUFx2_ASAP7_75t_SL g292 ( 
.A(n_190),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_142),
.Y(n_191)
);

NAND3xp33_ASAP7_75t_L g262 ( 
.A(n_191),
.B(n_200),
.C(n_116),
.Y(n_262)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_149),
.Y(n_192)
);

INVx4_ASAP7_75t_L g293 ( 
.A(n_192),
.Y(n_293)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_176),
.Y(n_193)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_193),
.Y(n_260)
);

INVx5_ASAP7_75t_SL g195 ( 
.A(n_136),
.Y(n_195)
);

OR2x2_ASAP7_75t_L g268 ( 
.A(n_195),
.B(n_41),
.Y(n_268)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_169),
.Y(n_196)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_196),
.Y(n_248)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_178),
.Y(n_197)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_197),
.Y(n_270)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_139),
.Y(n_198)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_198),
.Y(n_263)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_140),
.Y(n_199)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_199),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_128),
.Y(n_200)
);

INVx4_ASAP7_75t_L g201 ( 
.A(n_149),
.Y(n_201)
);

INVx4_ASAP7_75t_L g295 ( 
.A(n_201),
.Y(n_295)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_117),
.Y(n_202)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_202),
.Y(n_300)
);

HB1xp67_ASAP7_75t_L g203 ( 
.A(n_117),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_203),
.Y(n_247)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_141),
.Y(n_204)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_204),
.Y(n_273)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_155),
.Y(n_205)
);

INVx3_ASAP7_75t_L g301 ( 
.A(n_205),
.Y(n_301)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_154),
.Y(n_207)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_207),
.Y(n_274)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_132),
.Y(n_208)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_208),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_125),
.A2(n_96),
.B(n_35),
.Y(n_209)
);

OA21x2_ASAP7_75t_L g250 ( 
.A1(n_209),
.A2(n_243),
.B(n_239),
.Y(n_250)
);

INVx4_ASAP7_75t_L g210 ( 
.A(n_118),
.Y(n_210)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_210),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_135),
.B(n_32),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_130),
.B(n_45),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_212),
.B(n_215),
.Y(n_255)
);

INVx4_ASAP7_75t_L g214 ( 
.A(n_118),
.Y(n_214)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_214),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_116),
.B(n_45),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_170),
.A2(n_72),
.B1(n_39),
.B2(n_45),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g284 ( 
.A1(n_216),
.A2(n_226),
.B1(n_230),
.B2(n_239),
.Y(n_284)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_159),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g246 ( 
.A(n_217),
.B(n_221),
.Y(n_246)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_119),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_218),
.B(n_220),
.Y(n_257)
);

INVx5_ASAP7_75t_L g219 ( 
.A(n_114),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_219),
.Y(n_269)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_121),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_167),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_175),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g275 ( 
.A(n_222),
.B(n_236),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_223),
.A2(n_232),
.B1(n_238),
.B2(n_136),
.Y(n_256)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_138),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_224),
.B(n_227),
.Y(n_258)
);

INVx8_ASAP7_75t_L g226 ( 
.A(n_153),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_129),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_111),
.B(n_31),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_228),
.B(n_234),
.Y(n_271)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_146),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_229),
.B(n_233),
.Y(n_266)
);

AOI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_170),
.A2(n_39),
.B1(n_31),
.B2(n_49),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_153),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_231),
.Y(n_279)
);

OAI22xp33_ASAP7_75t_L g232 ( 
.A1(n_112),
.A2(n_126),
.B1(n_156),
.B2(n_134),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_173),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_122),
.B(n_173),
.Y(n_234)
);

OAI21xp33_ASAP7_75t_L g297 ( 
.A1(n_235),
.A2(n_12),
.B(n_16),
.Y(n_297)
);

INVx4_ASAP7_75t_L g236 ( 
.A(n_131),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_168),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_237),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_172),
.A2(n_39),
.B1(n_31),
.B2(n_53),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_SL g239 ( 
.A1(n_120),
.A2(n_53),
.B1(n_41),
.B2(n_92),
.Y(n_239)
);

INVx4_ASAP7_75t_L g240 ( 
.A(n_131),
.Y(n_240)
);

AND2x2_ASAP7_75t_L g283 ( 
.A(n_240),
.B(n_241),
.Y(n_283)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_164),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_120),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_242),
.B(n_0),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_157),
.A2(n_41),
.B(n_53),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_182),
.B(n_145),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_245),
.B(n_290),
.Y(n_306)
);

OAI21xp33_ASAP7_75t_SL g342 ( 
.A1(n_250),
.A2(n_294),
.B(n_298),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_182),
.B(n_145),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_251),
.B(n_253),
.C(n_280),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_235),
.B(n_157),
.C(n_114),
.Y(n_253)
);

OAI22xp33_ASAP7_75t_SL g254 ( 
.A1(n_183),
.A2(n_171),
.B1(n_164),
.B2(n_168),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_254),
.A2(n_278),
.B1(n_0),
.B2(n_1),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_256),
.A2(n_276),
.B1(n_277),
.B2(n_281),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_206),
.A2(n_177),
.B1(n_123),
.B2(n_143),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_261),
.A2(n_237),
.B1(n_179),
.B2(n_226),
.Y(n_313)
);

NAND3xp33_ASAP7_75t_L g308 ( 
.A(n_262),
.B(n_201),
.C(n_202),
.Y(n_308)
);

CKINVDCx16_ASAP7_75t_R g330 ( 
.A(n_268),
.Y(n_330)
);

CKINVDCx16_ASAP7_75t_R g272 ( 
.A(n_243),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_272),
.B(n_302),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_213),
.A2(n_166),
.B1(n_177),
.B2(n_143),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_L g277 ( 
.A1(n_232),
.A2(n_110),
.B1(n_166),
.B2(n_124),
.Y(n_277)
);

OAI22x1_ASAP7_75t_L g278 ( 
.A1(n_225),
.A2(n_116),
.B1(n_124),
.B2(n_123),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_209),
.A2(n_134),
.B1(n_53),
.B2(n_110),
.Y(n_281)
);

INVx1_ASAP7_75t_SL g339 ( 
.A(n_282),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_187),
.A2(n_10),
.B1(n_16),
.B2(n_15),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g340 ( 
.A1(n_289),
.A2(n_299),
.B1(n_274),
.B2(n_273),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_194),
.B(n_0),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_186),
.B(n_0),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_291),
.B(n_0),
.Y(n_312)
);

AOI22xp33_ASAP7_75t_SL g294 ( 
.A1(n_188),
.A2(n_208),
.B1(n_222),
.B2(n_192),
.Y(n_294)
);

FAx1_ASAP7_75t_SL g296 ( 
.A(n_195),
.B(n_6),
.CI(n_16),
.CON(n_296),
.SN(n_296)
);

OAI21xp5_ASAP7_75t_SL g317 ( 
.A1(n_296),
.A2(n_180),
.B(n_5),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_297),
.B(n_216),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_241),
.A2(n_5),
.B1(n_15),
.B2(n_14),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_185),
.B(n_17),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_185),
.B(n_17),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_303),
.B(n_298),
.Y(n_335)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_263),
.Y(n_304)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_304),
.Y(n_355)
);

AOI22xp33_ASAP7_75t_L g305 ( 
.A1(n_271),
.A2(n_197),
.B1(n_193),
.B2(n_231),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g380 ( 
.A1(n_305),
.A2(n_323),
.B1(n_327),
.B2(n_328),
.Y(n_380)
);

INVxp67_ASAP7_75t_L g362 ( 
.A(n_308),
.Y(n_362)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_268),
.A2(n_181),
.B(n_230),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g360 ( 
.A1(n_309),
.A2(n_316),
.B(n_334),
.Y(n_360)
);

INVxp67_ASAP7_75t_L g396 ( 
.A(n_310),
.Y(n_396)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_300),
.Y(n_311)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_311),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_312),
.B(n_319),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_313),
.A2(n_320),
.B1(n_333),
.B2(n_337),
.Y(n_370)
);

O2A1O1Ixp33_ASAP7_75t_SL g314 ( 
.A1(n_250),
.A2(n_219),
.B(n_236),
.C(n_240),
.Y(n_314)
);

A2O1A1Ixp33_ASAP7_75t_L g383 ( 
.A1(n_314),
.A2(n_322),
.B(n_324),
.C(n_349),
.Y(n_383)
);

INVx2_ASAP7_75t_SL g315 ( 
.A(n_265),
.Y(n_315)
);

INVx1_ASAP7_75t_SL g367 ( 
.A(n_315),
.Y(n_367)
);

AOI21xp5_ASAP7_75t_L g316 ( 
.A1(n_250),
.A2(n_214),
.B(n_210),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_SL g385 ( 
.A(n_317),
.B(n_335),
.Y(n_385)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_263),
.Y(n_318)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_318),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_291),
.B(n_184),
.Y(n_319)
);

OAI22xp33_ASAP7_75t_SL g320 ( 
.A1(n_276),
.A2(n_17),
.B1(n_13),
.B2(n_5),
.Y(n_320)
);

BUFx6f_ASAP7_75t_L g321 ( 
.A(n_264),
.Y(n_321)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_321),
.Y(n_361)
);

AND2x2_ASAP7_75t_L g373 ( 
.A(n_322),
.B(n_340),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_261),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_SL g324 ( 
.A1(n_245),
.A2(n_4),
.B(n_2),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_L g356 ( 
.A1(n_324),
.A2(n_247),
.B(n_286),
.Y(n_356)
);

BUFx6f_ASAP7_75t_L g325 ( 
.A(n_264),
.Y(n_325)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_325),
.Y(n_371)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_267),
.Y(n_326)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_326),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_256),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_327)
);

AOI22xp33_ASAP7_75t_L g328 ( 
.A1(n_244),
.A2(n_3),
.B1(n_279),
.B2(n_285),
.Y(n_328)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_267),
.Y(n_331)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_331),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_332),
.B(n_341),
.C(n_252),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_281),
.A2(n_284),
.B1(n_244),
.B2(n_290),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_L g334 ( 
.A1(n_253),
.A2(n_278),
.B(n_251),
.Y(n_334)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_273),
.Y(n_336)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_336),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_255),
.A2(n_249),
.B1(n_248),
.B2(n_289),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_279),
.A2(n_285),
.B1(n_248),
.B2(n_280),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_L g387 ( 
.A1(n_338),
.A2(n_348),
.B1(n_350),
.B2(n_354),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_274),
.B(n_257),
.C(n_258),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_342),
.A2(n_345),
.B1(n_346),
.B2(n_333),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_296),
.B(n_269),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_343),
.B(n_349),
.Y(n_366)
);

INVx2_ASAP7_75t_SL g344 ( 
.A(n_265),
.Y(n_344)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_344),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_L g345 ( 
.A1(n_296),
.A2(n_299),
.B1(n_269),
.B2(n_288),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_L g346 ( 
.A1(n_288),
.A2(n_266),
.B1(n_283),
.B2(n_246),
.Y(n_346)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_300),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_347),
.B(n_351),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_292),
.A2(n_283),
.B1(n_246),
.B2(n_275),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_275),
.B(n_246),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_283),
.A2(n_275),
.B1(n_270),
.B2(n_259),
.Y(n_350)
);

INVx3_ASAP7_75t_L g351 ( 
.A(n_293),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_259),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_352),
.B(n_354),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_260),
.B(n_270),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_353),
.B(n_304),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_260),
.A2(n_301),
.B1(n_286),
.B2(n_287),
.Y(n_354)
);

OAI21x1_ASAP7_75t_L g423 ( 
.A1(n_356),
.A2(n_378),
.B(n_393),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_334),
.A2(n_301),
.B1(n_287),
.B2(n_252),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_357),
.A2(n_397),
.B1(n_380),
.B2(n_387),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g409 ( 
.A(n_359),
.B(n_325),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_SL g364 ( 
.A(n_306),
.B(n_247),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_364),
.B(n_379),
.Y(n_417)
);

AOI21xp5_ASAP7_75t_L g368 ( 
.A1(n_316),
.A2(n_293),
.B(n_295),
.Y(n_368)
);

OAI21xp5_ASAP7_75t_L g408 ( 
.A1(n_368),
.A2(n_374),
.B(n_383),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_SL g369 ( 
.A(n_332),
.B(n_295),
.Y(n_369)
);

XOR2xp5_ASAP7_75t_L g425 ( 
.A(n_369),
.B(n_357),
.Y(n_425)
);

NAND2x1_ASAP7_75t_SL g374 ( 
.A(n_343),
.B(n_330),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_306),
.B(n_341),
.C(n_329),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_375),
.B(n_386),
.C(n_311),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_L g424 ( 
.A1(n_376),
.A2(n_394),
.B1(n_386),
.B2(n_380),
.Y(n_424)
);

OAI21xp5_ASAP7_75t_L g378 ( 
.A1(n_309),
.A2(n_314),
.B(n_317),
.Y(n_378)
);

CKINVDCx16_ASAP7_75t_R g382 ( 
.A(n_353),
.Y(n_382)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_382),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_319),
.B(n_312),
.Y(n_384)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_384),
.Y(n_413)
);

XOR2xp5_ASAP7_75t_L g386 ( 
.A(n_337),
.B(n_310),
.Y(n_386)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_389),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_339),
.B(n_336),
.Y(n_390)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_390),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_338),
.Y(n_391)
);

CKINVDCx14_ASAP7_75t_R g419 ( 
.A(n_391),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_SL g393 ( 
.A(n_339),
.B(n_326),
.Y(n_393)
);

NAND3xp33_ASAP7_75t_L g410 ( 
.A(n_393),
.B(n_395),
.C(n_374),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_307),
.A2(n_327),
.B1(n_313),
.B2(n_314),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_SL g395 ( 
.A(n_318),
.B(n_331),
.Y(n_395)
);

CKINVDCx16_ASAP7_75t_R g397 ( 
.A(n_350),
.Y(n_397)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_397),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_L g398 ( 
.A1(n_394),
.A2(n_323),
.B1(n_348),
.B2(n_321),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_L g461 ( 
.A1(n_398),
.A2(n_416),
.B1(n_404),
.B2(n_431),
.Y(n_461)
);

OAI32xp33_ASAP7_75t_L g399 ( 
.A1(n_366),
.A2(n_352),
.A3(n_315),
.B1(n_344),
.B2(n_347),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_399),
.B(n_401),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_L g437 ( 
.A(n_400),
.B(n_358),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_395),
.Y(n_401)
);

BUFx6f_ASAP7_75t_L g402 ( 
.A(n_361),
.Y(n_402)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_402),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_375),
.B(n_351),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_SL g443 ( 
.A(n_403),
.B(n_405),
.Y(n_443)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_404),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_385),
.B(n_321),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_369),
.B(n_344),
.C(n_315),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_406),
.B(n_409),
.C(n_427),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_385),
.B(n_325),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_SL g450 ( 
.A(n_407),
.B(n_414),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_410),
.B(n_381),
.Y(n_446)
);

OAI21xp5_ASAP7_75t_L g411 ( 
.A1(n_360),
.A2(n_374),
.B(n_378),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_411),
.B(n_415),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_359),
.B(n_390),
.Y(n_414)
);

OAI21xp5_ASAP7_75t_L g415 ( 
.A1(n_360),
.A2(n_396),
.B(n_366),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_L g416 ( 
.A1(n_376),
.A2(n_391),
.B1(n_370),
.B2(n_382),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_373),
.A2(n_370),
.B1(n_383),
.B2(n_387),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_SL g441 ( 
.A1(n_418),
.A2(n_377),
.B1(n_388),
.B2(n_381),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_SL g420 ( 
.A1(n_373),
.A2(n_368),
.B1(n_365),
.B2(n_384),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_L g447 ( 
.A1(n_420),
.A2(n_422),
.B1(n_424),
.B2(n_392),
.Y(n_447)
);

INVx1_ASAP7_75t_SL g421 ( 
.A(n_356),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_421),
.B(n_426),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_SL g422 ( 
.A1(n_373),
.A2(n_365),
.B1(n_364),
.B2(n_379),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_SL g440 ( 
.A(n_423),
.B(n_362),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_SL g454 ( 
.A(n_425),
.B(n_367),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_363),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_355),
.B(n_358),
.C(n_388),
.Y(n_427)
);

HB1xp67_ASAP7_75t_L g428 ( 
.A(n_363),
.Y(n_428)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_428),
.Y(n_451)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_389),
.Y(n_432)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_432),
.Y(n_464)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_355),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_433),
.B(n_392),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_437),
.B(n_462),
.C(n_463),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_419),
.Y(n_439)
);

AOI22xp33_ASAP7_75t_L g478 ( 
.A1(n_439),
.A2(n_445),
.B1(n_453),
.B2(n_402),
.Y(n_478)
);

AOI21xp33_ASAP7_75t_L g465 ( 
.A1(n_440),
.A2(n_446),
.B(n_411),
.Y(n_465)
);

AOI22xp5_ASAP7_75t_L g480 ( 
.A1(n_441),
.A2(n_461),
.B1(n_464),
.B2(n_453),
.Y(n_480)
);

XOR2xp5_ASAP7_75t_L g444 ( 
.A(n_409),
.B(n_377),
.Y(n_444)
);

XOR2xp5_ASAP7_75t_L g471 ( 
.A(n_444),
.B(n_454),
.Y(n_471)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_417),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_L g473 ( 
.A1(n_447),
.A2(n_457),
.B1(n_398),
.B2(n_412),
.Y(n_473)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_448),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_401),
.B(n_372),
.Y(n_449)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_449),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_417),
.B(n_372),
.Y(n_452)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_452),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_SL g453 ( 
.A(n_429),
.B(n_367),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_427),
.B(n_361),
.Y(n_455)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_455),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_426),
.B(n_371),
.Y(n_456)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_456),
.Y(n_484)
);

AOI22xp5_ASAP7_75t_L g457 ( 
.A1(n_416),
.A2(n_371),
.B1(n_432),
.B2(n_429),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_413),
.B(n_422),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_458),
.B(n_433),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_430),
.B(n_413),
.Y(n_460)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_460),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_400),
.B(n_425),
.C(n_406),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_415),
.B(n_430),
.C(n_431),
.Y(n_463)
);

AOI21xp5_ASAP7_75t_L g510 ( 
.A1(n_465),
.A2(n_474),
.B(n_467),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_439),
.B(n_412),
.Y(n_467)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_467),
.Y(n_496)
);

OAI22xp5_ASAP7_75t_SL g468 ( 
.A1(n_457),
.A2(n_418),
.B1(n_408),
.B2(n_421),
.Y(n_468)
);

AOI22xp5_ASAP7_75t_L g491 ( 
.A1(n_468),
.A2(n_473),
.B1(n_477),
.B2(n_485),
.Y(n_491)
);

AOI21xp5_ASAP7_75t_L g474 ( 
.A1(n_435),
.A2(n_408),
.B(n_436),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_462),
.B(n_423),
.C(n_420),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_475),
.B(n_435),
.C(n_463),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_476),
.B(n_479),
.Y(n_498)
);

OAI22xp5_ASAP7_75t_SL g477 ( 
.A1(n_447),
.A2(n_399),
.B1(n_402),
.B2(n_434),
.Y(n_477)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_478),
.Y(n_501)
);

CKINVDCx20_ASAP7_75t_R g479 ( 
.A(n_448),
.Y(n_479)
);

AOI22xp5_ASAP7_75t_L g500 ( 
.A1(n_480),
.A2(n_442),
.B1(n_436),
.B2(n_460),
.Y(n_500)
);

XOR2xp5_ASAP7_75t_L g482 ( 
.A(n_459),
.B(n_437),
.Y(n_482)
);

XOR2xp5_ASAP7_75t_L g492 ( 
.A(n_482),
.B(n_488),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_450),
.B(n_443),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_483),
.B(n_490),
.Y(n_512)
);

AOI22xp5_ASAP7_75t_L g485 ( 
.A1(n_461),
.A2(n_434),
.B1(n_441),
.B2(n_464),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_445),
.B(n_455),
.Y(n_486)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_486),
.Y(n_502)
);

BUFx6f_ASAP7_75t_L g487 ( 
.A(n_438),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_487),
.B(n_438),
.Y(n_494)
);

XNOR2xp5_ASAP7_75t_L g488 ( 
.A(n_459),
.B(n_444),
.Y(n_488)
);

XNOR2xp5_ASAP7_75t_L g495 ( 
.A(n_488),
.B(n_450),
.Y(n_495)
);

CKINVDCx20_ASAP7_75t_R g490 ( 
.A(n_449),
.Y(n_490)
);

MAJx2_ASAP7_75t_L g517 ( 
.A(n_492),
.B(n_493),
.C(n_497),
.Y(n_517)
);

XOR2xp5_ASAP7_75t_L g493 ( 
.A(n_472),
.B(n_454),
.Y(n_493)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_494),
.Y(n_514)
);

XNOR2xp5_ASAP7_75t_L g521 ( 
.A(n_495),
.B(n_504),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_472),
.B(n_443),
.Y(n_499)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_499),
.Y(n_515)
);

OAI22xp5_ASAP7_75t_L g528 ( 
.A1(n_500),
.A2(n_510),
.B1(n_466),
.B2(n_469),
.Y(n_528)
);

XOR2xp5_ASAP7_75t_L g503 ( 
.A(n_471),
.B(n_440),
.Y(n_503)
);

XOR2xp5_ASAP7_75t_L g526 ( 
.A(n_503),
.B(n_480),
.Y(n_526)
);

XNOR2xp5_ASAP7_75t_L g504 ( 
.A(n_482),
.B(n_442),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_475),
.B(n_456),
.C(n_452),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_505),
.B(n_506),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_481),
.B(n_451),
.C(n_471),
.Y(n_506)
);

XNOR2xp5_ASAP7_75t_L g507 ( 
.A(n_481),
.B(n_451),
.Y(n_507)
);

XNOR2xp5_ASAP7_75t_L g525 ( 
.A(n_507),
.B(n_485),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_486),
.B(n_468),
.C(n_474),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_508),
.B(n_509),
.Y(n_529)
);

MAJIxp5_ASAP7_75t_L g509 ( 
.A(n_466),
.B(n_484),
.C(n_489),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_489),
.B(n_479),
.Y(n_511)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_511),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_507),
.B(n_490),
.Y(n_513)
);

OR2x2_ASAP7_75t_L g540 ( 
.A(n_513),
.B(n_518),
.Y(n_540)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_500),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_498),
.B(n_512),
.Y(n_520)
);

CKINVDCx20_ASAP7_75t_R g537 ( 
.A(n_520),
.Y(n_537)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_496),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_522),
.B(n_523),
.Y(n_530)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_509),
.Y(n_523)
);

CKINVDCx20_ASAP7_75t_R g524 ( 
.A(n_502),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_SL g536 ( 
.A(n_524),
.B(n_470),
.Y(n_536)
);

HB1xp67_ASAP7_75t_L g541 ( 
.A(n_525),
.Y(n_541)
);

XOR2xp5_ASAP7_75t_L g539 ( 
.A(n_526),
.B(n_506),
.Y(n_539)
);

AOI21xp5_ASAP7_75t_L g527 ( 
.A1(n_508),
.A2(n_484),
.B(n_469),
.Y(n_527)
);

OAI21xp5_ASAP7_75t_SL g535 ( 
.A1(n_527),
.A2(n_529),
.B(n_513),
.Y(n_535)
);

AND2x2_ASAP7_75t_SL g543 ( 
.A(n_528),
.B(n_503),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_515),
.B(n_495),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_531),
.B(n_532),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_SL g532 ( 
.A(n_520),
.B(n_505),
.Y(n_532)
);

MAJIxp5_ASAP7_75t_L g533 ( 
.A(n_519),
.B(n_492),
.C(n_497),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_533),
.B(n_534),
.Y(n_553)
);

OAI22xp5_ASAP7_75t_L g534 ( 
.A1(n_516),
.A2(n_501),
.B1(n_491),
.B2(n_470),
.Y(n_534)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_535),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_536),
.B(n_538),
.Y(n_549)
);

OAI21xp5_ASAP7_75t_L g538 ( 
.A1(n_518),
.A2(n_477),
.B(n_504),
.Y(n_538)
);

XNOR2xp5_ASAP7_75t_L g547 ( 
.A(n_539),
.B(n_521),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_SL g542 ( 
.A(n_514),
.B(n_493),
.Y(n_542)
);

CKINVDCx16_ASAP7_75t_R g548 ( 
.A(n_542),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_543),
.B(n_521),
.Y(n_551)
);

MAJIxp5_ASAP7_75t_L g544 ( 
.A(n_539),
.B(n_527),
.C(n_517),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_544),
.B(n_546),
.Y(n_555)
);

AOI22xp5_ASAP7_75t_L g546 ( 
.A1(n_537),
.A2(n_525),
.B1(n_526),
.B2(n_514),
.Y(n_546)
);

XOR2xp5_ASAP7_75t_L g557 ( 
.A(n_547),
.B(n_543),
.Y(n_557)
);

AO21x1_ASAP7_75t_L g554 ( 
.A1(n_551),
.A2(n_552),
.B(n_535),
.Y(n_554)
);

AOI22xp5_ASAP7_75t_L g552 ( 
.A1(n_538),
.A2(n_487),
.B1(n_517),
.B2(n_540),
.Y(n_552)
);

XOR2xp5_ASAP7_75t_L g560 ( 
.A(n_554),
.B(n_556),
.Y(n_560)
);

OAI21xp5_ASAP7_75t_L g556 ( 
.A1(n_550),
.A2(n_530),
.B(n_533),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_L g562 ( 
.A(n_557),
.B(n_558),
.Y(n_562)
);

XNOR2xp5_ASAP7_75t_SL g558 ( 
.A(n_545),
.B(n_541),
.Y(n_558)
);

OAI21xp5_ASAP7_75t_SL g559 ( 
.A1(n_553),
.A2(n_540),
.B(n_543),
.Y(n_559)
);

AND2x2_ASAP7_75t_SL g561 ( 
.A(n_559),
.B(n_552),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_561),
.B(n_555),
.Y(n_564)
);

AO21x2_ASAP7_75t_L g563 ( 
.A1(n_560),
.A2(n_549),
.B(n_546),
.Y(n_563)
);

MAJIxp5_ASAP7_75t_L g565 ( 
.A(n_563),
.B(n_564),
.C(n_555),
.Y(n_565)
);

XOR2xp5_ASAP7_75t_L g566 ( 
.A(n_565),
.B(n_562),
.Y(n_566)
);

OAI21xp5_ASAP7_75t_L g567 ( 
.A1(n_566),
.A2(n_548),
.B(n_549),
.Y(n_567)
);

AOI21xp5_ASAP7_75t_SL g568 ( 
.A1(n_567),
.A2(n_544),
.B(n_551),
.Y(n_568)
);

AOI21xp5_ASAP7_75t_L g569 ( 
.A1(n_568),
.A2(n_547),
.B(n_487),
.Y(n_569)
);


endmodule