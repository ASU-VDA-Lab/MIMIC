module fake_jpeg_20360_n_104 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_8, n_15, n_7, n_104);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_8;
input n_15;
input n_7;

output n_104;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_8),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_13),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_29),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_25),
.B(n_30),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_21),
.B(n_15),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_12),
.B(n_31),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_26),
.B(n_2),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_46),
.B(n_0),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_50),
.B(n_53),
.Y(n_57)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_51),
.B(n_54),
.Y(n_61)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_52),
.B(n_37),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_46),
.B(n_0),
.Y(n_53)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

OAI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_48),
.A2(n_45),
.B1(n_40),
.B2(n_36),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_55),
.A2(n_41),
.B1(n_39),
.B2(n_1),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_53),
.Y(n_56)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_58),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

BUFx2_ASAP7_75t_L g67 ( 
.A(n_59),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_62),
.B(n_65),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_53),
.B(n_44),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_53),
.B(n_42),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_66),
.B(n_2),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_57),
.B(n_32),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_68),
.B(n_70),
.Y(n_83)
);

AO21x1_ASAP7_75t_L g82 ( 
.A1(n_72),
.A2(n_78),
.B(n_17),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_61),
.A2(n_64),
.B1(n_60),
.B2(n_6),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_73),
.B(n_18),
.Y(n_84)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_63),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_74),
.B(n_77),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_SL g76 ( 
.A1(n_57),
.A2(n_3),
.B(n_5),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_L g80 ( 
.A(n_76),
.B(n_14),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_59),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_64),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_61),
.Y(n_79)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_79),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_80),
.B(n_84),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_82),
.B(n_86),
.Y(n_91)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_75),
.Y(n_85)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_85),
.Y(n_90)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_67),
.Y(n_86)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_69),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_88),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_87),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_93),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_92),
.A2(n_71),
.B1(n_83),
.B2(n_84),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_95),
.Y(n_96)
);

XOR2xp5_ASAP7_75t_L g97 ( 
.A(n_96),
.B(n_89),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_97),
.B(n_94),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_98),
.A2(n_90),
.B(n_91),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_99),
.B(n_81),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_100),
.A2(n_69),
.B(n_72),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_101),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_102),
.A2(n_19),
.B(n_20),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_103),
.B(n_24),
.Y(n_104)
);


endmodule