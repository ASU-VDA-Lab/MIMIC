module fake_jpeg_19542_n_38 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_38);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_38;

wire n_13;
wire n_21;
wire n_33;
wire n_23;
wire n_10;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_36;
wire n_11;
wire n_25;
wire n_31;
wire n_17;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_15;

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_3),
.Y(n_10)
);

INVx13_ASAP7_75t_L g11 ( 
.A(n_9),
.Y(n_11)
);

INVx8_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

INVx6_ASAP7_75t_SL g14 ( 
.A(n_7),
.Y(n_14)
);

INVx3_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_2),
.B(n_5),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_16),
.B(n_0),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_19),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_L g20 ( 
.A1(n_18),
.A2(n_8),
.B1(n_4),
.B2(n_5),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_SL g27 ( 
.A1(n_20),
.A2(n_23),
.B1(n_24),
.B2(n_18),
.Y(n_27)
);

OR2x4_ASAP7_75t_L g21 ( 
.A(n_13),
.B(n_1),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_21),
.B(n_22),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_11),
.Y(n_23)
);

INVx1_ASAP7_75t_SL g24 ( 
.A(n_10),
.Y(n_24)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_27),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_25),
.A2(n_24),
.B1(n_20),
.B2(n_22),
.Y(n_28)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_28),
.Y(n_30)
);

A2O1A1Ixp33_ASAP7_75t_SL g31 ( 
.A1(n_30),
.A2(n_29),
.B(n_28),
.C(n_27),
.Y(n_31)
);

OAI21xp5_ASAP7_75t_L g34 ( 
.A1(n_31),
.A2(n_32),
.B(n_17),
.Y(n_34)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_30),
.Y(n_32)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g33 ( 
.A1(n_31),
.A2(n_25),
.B(n_26),
.C(n_11),
.D(n_17),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_33),
.B(n_34),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g35 ( 
.A(n_34),
.B(n_14),
.C(n_15),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_35),
.B(n_12),
.C(n_15),
.Y(n_37)
);

XOR2xp5_ASAP7_75t_L g38 ( 
.A(n_37),
.B(n_36),
.Y(n_38)
);


endmodule