module fake_jpeg_17447_n_47 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_47);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_47;

wire n_21;
wire n_33;
wire n_45;
wire n_23;
wire n_27;
wire n_22;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_25;
wire n_17;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_32;

INVx3_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx24_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_18),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_22),
.B(n_24),
.Y(n_32)
);

BUFx2_ASAP7_75t_L g23 ( 
.A(n_18),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_23),
.Y(n_30)
);

INVx5_ASAP7_75t_L g24 ( 
.A(n_18),
.Y(n_24)
);

NOR4xp25_ASAP7_75t_SL g25 ( 
.A(n_20),
.B(n_16),
.C(n_15),
.D(n_14),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_25),
.B(n_21),
.C(n_17),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_19),
.B(n_20),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_26),
.B(n_17),
.Y(n_28)
);

OAI21x1_ASAP7_75t_L g36 ( 
.A1(n_27),
.A2(n_28),
.B(n_0),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

A2O1A1Ixp33_ASAP7_75t_SL g35 ( 
.A1(n_29),
.A2(n_24),
.B(n_1),
.C(n_2),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_25),
.A2(n_13),
.B1(n_12),
.B2(n_11),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_31),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_33),
.A2(n_37),
.B1(n_3),
.B2(n_5),
.Y(n_39)
);

A2O1A1O1Ixp25_ASAP7_75t_L g34 ( 
.A1(n_27),
.A2(n_21),
.B(n_10),
.C(n_23),
.D(n_22),
.Y(n_34)
);

OAI21xp5_ASAP7_75t_SL g41 ( 
.A1(n_34),
.A2(n_35),
.B(n_36),
.Y(n_41)
);

AOI21xp5_ASAP7_75t_L g37 ( 
.A1(n_31),
.A2(n_3),
.B(n_5),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_35),
.B(n_30),
.C(n_32),
.Y(n_38)
);

XOR2xp5_ASAP7_75t_L g43 ( 
.A(n_38),
.B(n_29),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_39),
.A2(n_40),
.B1(n_30),
.B2(n_7),
.Y(n_42)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_42),
.A2(n_43),
.B1(n_44),
.B2(n_38),
.Y(n_45)
);

A2O1A1Ixp33_ASAP7_75t_L g44 ( 
.A1(n_41),
.A2(n_6),
.B(n_8),
.C(n_9),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_45),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_46),
.B(n_44),
.Y(n_47)
);


endmodule