module fake_jpeg_15947_n_121 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_121);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_121;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

INVx3_ASAP7_75t_SL g13 ( 
.A(n_12),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

HB1xp67_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_3),
.B(n_2),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_6),
.B(n_11),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_23),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_26),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g27 ( 
.A(n_24),
.B(n_0),
.Y(n_27)
);

OAI21xp5_ASAP7_75t_SL g51 ( 
.A1(n_27),
.A2(n_28),
.B(n_19),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_24),
.B(n_0),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_14),
.B(n_0),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_29),
.B(n_39),
.Y(n_42)
);

INVx1_ASAP7_75t_SL g30 ( 
.A(n_25),
.Y(n_30)
);

OR2x2_ASAP7_75t_L g46 ( 
.A(n_30),
.B(n_31),
.Y(n_46)
);

CKINVDCx16_ASAP7_75t_R g31 ( 
.A(n_18),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_33),
.Y(n_61)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_34),
.Y(n_50)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_35),
.B(n_37),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_13),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_36),
.A2(n_38),
.B1(n_39),
.B2(n_29),
.Y(n_48)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_14),
.B(n_1),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_38),
.B(n_4),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_17),
.B(n_2),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_27),
.B(n_20),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_40),
.B(n_51),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_34),
.A2(n_17),
.B1(n_5),
.B2(n_6),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_44),
.A2(n_22),
.B1(n_10),
.B2(n_12),
.Y(n_70)
);

INVx13_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_45),
.B(n_47),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_31),
.B(n_18),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_48),
.A2(n_8),
.B1(n_51),
.B2(n_42),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_52),
.B(n_53),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_27),
.B(n_4),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_33),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_54),
.B(n_62),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_L g56 ( 
.A(n_28),
.B(n_15),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_56),
.B(n_58),
.C(n_8),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_32),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_57),
.B(n_59),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_30),
.B(n_16),
.C(n_22),
.Y(n_58)
);

INVx13_ASAP7_75t_L g59 ( 
.A(n_26),
.Y(n_59)
);

INVx13_ASAP7_75t_L g60 ( 
.A(n_26),
.Y(n_60)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_60),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_28),
.B(n_22),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_SL g63 ( 
.A1(n_62),
.A2(n_52),
.B(n_53),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_63),
.B(n_50),
.C(n_46),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_52),
.A2(n_35),
.B1(n_30),
.B2(n_5),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_65),
.A2(n_68),
.B1(n_69),
.B2(n_70),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_49),
.A2(n_35),
.B1(n_6),
.B2(n_16),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_44),
.A2(n_56),
.B1(n_42),
.B2(n_48),
.Y(n_69)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_71),
.B(n_74),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_SL g84 ( 
.A(n_72),
.B(n_43),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_49),
.A2(n_57),
.B1(n_45),
.B2(n_41),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_50),
.A2(n_58),
.B1(n_54),
.B2(n_61),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_78),
.B(n_46),
.Y(n_80)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_67),
.Y(n_79)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_79),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_80),
.A2(n_65),
.B1(n_73),
.B2(n_66),
.Y(n_98)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_64),
.Y(n_81)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_81),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_82),
.B(n_84),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_77),
.B(n_46),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_83),
.B(n_87),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_SL g85 ( 
.A(n_63),
.B(n_61),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_85),
.B(n_82),
.C(n_72),
.Y(n_93)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_64),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_86),
.B(n_88),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_71),
.B(n_55),
.Y(n_87)
);

BUFx2_ASAP7_75t_L g88 ( 
.A(n_77),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_66),
.B(n_75),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_90),
.B(n_91),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_76),
.B(n_59),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_93),
.B(n_94),
.C(n_97),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_84),
.B(n_73),
.C(n_74),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g97 ( 
.A(n_85),
.B(n_66),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_98),
.B(n_97),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g100 ( 
.A(n_92),
.B(n_89),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_100),
.A2(n_55),
.B(n_88),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_95),
.A2(n_87),
.B1(n_89),
.B2(n_92),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_104),
.B(n_105),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_100),
.A2(n_70),
.B1(n_68),
.B2(n_60),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_106),
.B(n_108),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_94),
.A2(n_55),
.B1(n_93),
.B2(n_99),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_107),
.A2(n_106),
.B1(n_105),
.B2(n_104),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_101),
.A2(n_102),
.B1(n_103),
.B2(n_96),
.Y(n_108)
);

AOI31xp33_ASAP7_75t_L g112 ( 
.A1(n_110),
.A2(n_101),
.A3(n_109),
.B(n_107),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_111),
.B(n_112),
.Y(n_118)
);

OR2x2_ASAP7_75t_L g114 ( 
.A(n_109),
.B(n_95),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_114),
.B(n_113),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_115),
.Y(n_116)
);

AO21x1_ASAP7_75t_L g120 ( 
.A1(n_116),
.A2(n_117),
.B(n_111),
.Y(n_120)
);

HB1xp67_ASAP7_75t_L g119 ( 
.A(n_117),
.Y(n_119)
);

AOI21x1_ASAP7_75t_SL g121 ( 
.A1(n_119),
.A2(n_120),
.B(n_118),
.Y(n_121)
);


endmodule