module fake_jpeg_6434_n_96 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_96);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_96;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_62;
wire n_43;
wire n_82;

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_11),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_3),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_2),
.Y(n_47)
);

HB1xp67_ASAP7_75t_L g48 ( 
.A(n_23),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_33),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_8),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_0),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_26),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_16),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_14),
.B(n_6),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_21),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_41),
.B(n_1),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_57),
.B(n_62),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_45),
.B(n_51),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_58),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_49),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_59),
.B(n_60),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_48),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_61),
.Y(n_63)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_57),
.A2(n_53),
.B1(n_52),
.B2(n_42),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_65),
.A2(n_44),
.B1(n_55),
.B2(n_54),
.Y(n_70)
);

CKINVDCx12_ASAP7_75t_R g66 ( 
.A(n_58),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_66),
.B(n_67),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_57),
.B(n_46),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_70),
.A2(n_69),
.B1(n_56),
.B2(n_50),
.Y(n_75)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_63),
.Y(n_71)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_71),
.Y(n_76)
);

BUFx2_ASAP7_75t_SL g73 ( 
.A(n_68),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_73),
.B(n_5),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_72),
.B(n_64),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_74),
.B(n_75),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_77),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_73),
.A2(n_47),
.B(n_43),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_78),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_73),
.A2(n_38),
.B1(n_10),
.B2(n_12),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_79),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_72),
.B(n_9),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_83),
.A2(n_80),
.B1(n_76),
.B2(n_17),
.Y(n_85)
);

OAI21xp33_ASAP7_75t_L g87 ( 
.A1(n_85),
.A2(n_86),
.B(n_18),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_82),
.A2(n_13),
.B(n_15),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_87),
.B(n_81),
.C(n_84),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_88),
.B(n_19),
.C(n_22),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_SL g90 ( 
.A(n_89),
.B(n_24),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_90),
.B(n_25),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_91),
.B(n_27),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_92),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_93),
.Y(n_94)
);

OAI31xp67_ASAP7_75t_L g95 ( 
.A1(n_94),
.A2(n_28),
.A3(n_29),
.B(n_30),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_95),
.B(n_32),
.Y(n_96)
);


endmodule