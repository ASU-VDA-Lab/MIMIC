module fake_jpeg_15485_n_392 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_392);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_392;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

BUFx16f_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx16f_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_11),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_11),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_6),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_8),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_3),
.Y(n_34)
);

INVx11_ASAP7_75t_SL g35 ( 
.A(n_2),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_8),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_40),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_41),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_20),
.B(n_7),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_42),
.B(n_52),
.Y(n_99)
);

INVx6_ASAP7_75t_SL g43 ( 
.A(n_16),
.Y(n_43)
);

INVx2_ASAP7_75t_SL g100 ( 
.A(n_43),
.Y(n_100)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_44),
.Y(n_85)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_45),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_21),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_46),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_27),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_47),
.B(n_54),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_21),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_48),
.Y(n_83)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_49),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_16),
.Y(n_50)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_50),
.Y(n_118)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_27),
.Y(n_51)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_51),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_20),
.B(n_7),
.Y(n_52)
);

INVx8_ASAP7_75t_SL g53 ( 
.A(n_35),
.Y(n_53)
);

BUFx2_ASAP7_75t_L g80 ( 
.A(n_53),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_16),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_27),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_55),
.B(n_63),
.Y(n_82)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_27),
.Y(n_56)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_21),
.Y(n_57)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_57),
.Y(n_110)
);

BUFx12f_ASAP7_75t_SL g58 ( 
.A(n_35),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_58),
.B(n_69),
.Y(n_76)
);

BUFx24_ASAP7_75t_L g59 ( 
.A(n_27),
.Y(n_59)
);

BUFx2_ASAP7_75t_L g109 ( 
.A(n_59),
.Y(n_109)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_60),
.Y(n_112)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_21),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g122 ( 
.A(n_61),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_62),
.Y(n_73)
);

INVx1_ASAP7_75t_SL g63 ( 
.A(n_16),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_18),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_64),
.B(n_30),
.Y(n_107)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_18),
.Y(n_65)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_65),
.Y(n_104)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_18),
.Y(n_66)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_66),
.Y(n_113)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_15),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_67),
.B(n_25),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_37),
.Y(n_68)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_68),
.Y(n_77)
);

INVx2_ASAP7_75t_R g69 ( 
.A(n_18),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_37),
.Y(n_70)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_70),
.Y(n_119)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_37),
.Y(n_71)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_71),
.Y(n_114)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_18),
.Y(n_72)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_72),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_45),
.A2(n_17),
.B1(n_29),
.B2(n_28),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_81),
.A2(n_92),
.B1(n_97),
.B2(n_115),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_58),
.A2(n_17),
.B1(n_26),
.B2(n_28),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_87),
.A2(n_88),
.B1(n_91),
.B2(n_105),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_69),
.A2(n_17),
.B1(n_26),
.B2(n_28),
.Y(n_88)
);

BUFx12f_ASAP7_75t_L g89 ( 
.A(n_61),
.Y(n_89)
);

INVx5_ASAP7_75t_L g146 ( 
.A(n_89),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_40),
.B(n_14),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_90),
.A2(n_100),
.B1(n_86),
.B2(n_77),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_49),
.A2(n_26),
.B1(n_29),
.B2(n_32),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_60),
.A2(n_29),
.B1(n_34),
.B2(n_31),
.Y(n_92)
);

BUFx8_ASAP7_75t_L g93 ( 
.A(n_72),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_93),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_94),
.B(n_98),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_70),
.A2(n_38),
.B1(n_34),
.B2(n_22),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_67),
.B(n_38),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_71),
.B(n_22),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_101),
.B(n_8),
.Y(n_126)
);

OAI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_51),
.A2(n_31),
.B1(n_30),
.B2(n_23),
.Y(n_102)
);

OAI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_102),
.A2(n_9),
.B1(n_1),
.B2(n_3),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_65),
.A2(n_24),
.B1(n_33),
.B2(n_32),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_66),
.A2(n_24),
.B1(n_33),
.B2(n_32),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_106),
.A2(n_123),
.B1(n_125),
.B2(n_111),
.Y(n_164)
);

CKINVDCx14_ASAP7_75t_R g171 ( 
.A(n_107),
.Y(n_171)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_61),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g152 ( 
.A(n_108),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_59),
.B(n_33),
.C(n_25),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_111),
.B(n_8),
.C(n_1),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_56),
.A2(n_44),
.B1(n_46),
.B2(n_57),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_41),
.B(n_23),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_116),
.B(n_117),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_62),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_63),
.A2(n_25),
.B1(n_24),
.B2(n_19),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_120),
.A2(n_86),
.B1(n_79),
.B2(n_108),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_48),
.A2(n_19),
.B1(n_15),
.B2(n_36),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_121),
.A2(n_12),
.B1(n_13),
.B2(n_0),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_43),
.A2(n_19),
.B1(n_36),
.B2(n_14),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_68),
.B(n_36),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_124),
.B(n_0),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_59),
.A2(n_14),
.B1(n_1),
.B2(n_2),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_126),
.B(n_142),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_124),
.A2(n_54),
.B1(n_50),
.B2(n_2),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_127),
.A2(n_147),
.B1(n_122),
.B2(n_155),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g201 ( 
.A(n_128),
.B(n_130),
.Y(n_201)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_95),
.Y(n_129)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_129),
.Y(n_176)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_119),
.Y(n_131)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_131),
.Y(n_184)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_119),
.Y(n_132)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_132),
.Y(n_196)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_74),
.Y(n_133)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_133),
.Y(n_181)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_74),
.Y(n_134)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_134),
.Y(n_188)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_104),
.Y(n_137)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_137),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_103),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_138),
.B(n_141),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_99),
.B(n_7),
.Y(n_139)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_139),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_76),
.A2(n_7),
.B1(n_1),
.B2(n_3),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_140),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_118),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_82),
.B(n_9),
.Y(n_142)
);

OAI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_143),
.A2(n_150),
.B1(n_151),
.B2(n_156),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_120),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_144),
.B(n_145),
.Y(n_199)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_89),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_110),
.A2(n_4),
.B1(n_6),
.B2(n_10),
.Y(n_147)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_104),
.Y(n_148)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_148),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_76),
.A2(n_6),
.B1(n_11),
.B2(n_12),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_149),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_76),
.A2(n_6),
.B1(n_11),
.B2(n_12),
.Y(n_150)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_84),
.Y(n_153)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_153),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_78),
.Y(n_154)
);

INVx1_ASAP7_75t_SL g205 ( 
.A(n_154),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_90),
.B(n_12),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_155),
.B(n_170),
.Y(n_183)
);

INVx3_ASAP7_75t_SL g156 ( 
.A(n_78),
.Y(n_156)
);

OAI22xp33_ASAP7_75t_L g157 ( 
.A1(n_110),
.A2(n_13),
.B1(n_73),
.B2(n_77),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_157),
.A2(n_166),
.B1(n_79),
.B2(n_83),
.Y(n_187)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_113),
.Y(n_159)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_159),
.Y(n_180)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_89),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_160),
.B(n_162),
.Y(n_202)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_113),
.Y(n_161)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_161),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_75),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_84),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_163),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g214 ( 
.A(n_164),
.B(n_174),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_90),
.A2(n_114),
.B1(n_96),
.B2(n_112),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_93),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_167),
.B(n_168),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_100),
.B(n_85),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_114),
.B(n_96),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_112),
.B(n_73),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_172),
.B(n_170),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_173),
.A2(n_163),
.B(n_153),
.Y(n_209)
);

INVx2_ASAP7_75t_SL g175 ( 
.A(n_80),
.Y(n_175)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_175),
.Y(n_206)
);

BUFx24_ASAP7_75t_SL g179 ( 
.A(n_165),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_179),
.B(n_186),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_135),
.B(n_115),
.C(n_85),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_185),
.B(n_204),
.C(n_221),
.Y(n_241)
);

INVx5_ASAP7_75t_L g186 ( 
.A(n_146),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_L g231 ( 
.A1(n_187),
.A2(n_194),
.B1(n_204),
.B2(n_186),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_174),
.A2(n_83),
.B1(n_93),
.B2(n_109),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_189),
.A2(n_190),
.B1(n_156),
.B2(n_157),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_128),
.A2(n_109),
.B1(n_122),
.B2(n_80),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g228 ( 
.A(n_191),
.B(n_183),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_131),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_195),
.B(n_208),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_129),
.B(n_165),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_197),
.B(n_203),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_127),
.B(n_130),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_173),
.B(n_166),
.C(n_172),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_132),
.Y(n_208)
);

AO21x1_ASAP7_75t_L g230 ( 
.A1(n_209),
.A2(n_199),
.B(n_189),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_158),
.B(n_136),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_210),
.B(n_216),
.Y(n_242)
);

AOI32xp33_ASAP7_75t_L g212 ( 
.A1(n_146),
.A2(n_158),
.A3(n_169),
.B1(n_151),
.B2(n_147),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_SL g233 ( 
.A1(n_212),
.A2(n_214),
.B(n_193),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_134),
.B(n_133),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_154),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_217),
.B(n_177),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_137),
.B(n_159),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_218),
.B(n_220),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_148),
.B(n_161),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_169),
.B(n_152),
.C(n_171),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_201),
.B(n_145),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_222),
.B(n_247),
.C(n_248),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_197),
.B(n_152),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_223),
.B(n_226),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_224),
.A2(n_225),
.B1(n_227),
.B2(n_238),
.Y(n_274)
);

OAI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_178),
.A2(n_156),
.B1(n_160),
.B2(n_175),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_207),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_214),
.A2(n_175),
.B1(n_185),
.B2(n_210),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_228),
.B(n_249),
.Y(n_271)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_218),
.Y(n_229)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_229),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_230),
.A2(n_233),
.B(n_255),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_231),
.A2(n_247),
.B1(n_248),
.B2(n_249),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_202),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_232),
.B(n_238),
.Y(n_286)
);

AOI22xp33_ASAP7_75t_L g235 ( 
.A1(n_187),
.A2(n_209),
.B1(n_182),
.B2(n_194),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_L g266 ( 
.A1(n_235),
.A2(n_244),
.B1(n_224),
.B2(n_230),
.Y(n_266)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_216),
.Y(n_236)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_236),
.Y(n_295)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_176),
.Y(n_238)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_239),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_220),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_240),
.B(n_254),
.Y(n_291)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_184),
.Y(n_243)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_243),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_L g244 ( 
.A1(n_178),
.A2(n_193),
.B(n_214),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_244),
.A2(n_252),
.B(n_253),
.Y(n_283)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_184),
.Y(n_245)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_245),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_203),
.A2(n_191),
.B1(n_183),
.B2(n_221),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_176),
.A2(n_201),
.B1(n_190),
.B2(n_196),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_201),
.B(n_213),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_196),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g273 ( 
.A(n_250),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_211),
.B(n_215),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_213),
.B(n_219),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g254 ( 
.A(n_181),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_188),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_200),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_256),
.Y(n_270)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_180),
.Y(n_257)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_257),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_200),
.B(n_192),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_258),
.B(n_262),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_198),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_259),
.Y(n_272)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_180),
.Y(n_260)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_260),
.Y(n_293)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_177),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_261),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_206),
.B(n_205),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_242),
.A2(n_205),
.B1(n_206),
.B2(n_228),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_264),
.A2(n_265),
.B1(n_275),
.B2(n_285),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_242),
.A2(n_228),
.B1(n_241),
.B2(n_233),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_266),
.A2(n_251),
.B1(n_254),
.B2(n_283),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_269),
.B(n_265),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_274),
.A2(n_267),
.B1(n_295),
.B2(n_279),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_241),
.A2(n_230),
.B1(n_240),
.B2(n_227),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_278),
.B(n_280),
.C(n_284),
.Y(n_300)
);

OR2x6_ASAP7_75t_L g279 ( 
.A(n_223),
.B(n_246),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_279),
.A2(n_252),
.B(n_260),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_222),
.B(n_237),
.C(n_229),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_237),
.B(n_236),
.C(n_246),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_243),
.A2(n_245),
.B1(n_250),
.B2(n_258),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_257),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_287),
.B(n_270),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_234),
.B(n_253),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_288),
.B(n_294),
.C(n_280),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_262),
.A2(n_256),
.B1(n_234),
.B2(n_259),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_290),
.A2(n_279),
.B1(n_264),
.B2(n_285),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_261),
.B(n_239),
.C(n_255),
.Y(n_294)
);

CKINVDCx14_ASAP7_75t_R g338 ( 
.A(n_296),
.Y(n_338)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_292),
.Y(n_297)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_297),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_298),
.A2(n_301),
.B1(n_302),
.B2(n_310),
.Y(n_324)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_292),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_299),
.B(n_304),
.Y(n_328)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_293),
.Y(n_304)
);

BUFx5_ASAP7_75t_L g305 ( 
.A(n_279),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_305),
.B(n_311),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_263),
.B(n_288),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_306),
.B(n_307),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_263),
.B(n_279),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_308),
.B(n_309),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_277),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_275),
.A2(n_271),
.B1(n_295),
.B2(n_278),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_271),
.A2(n_267),
.B1(n_282),
.B2(n_269),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_293),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_312),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_282),
.A2(n_284),
.B1(n_280),
.B2(n_283),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_313),
.B(n_315),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_314),
.Y(n_337)
);

AOI21xp5_ASAP7_75t_L g315 ( 
.A1(n_268),
.A2(n_291),
.B(n_281),
.Y(n_315)
);

OA21x2_ASAP7_75t_L g316 ( 
.A1(n_290),
.A2(n_289),
.B(n_276),
.Y(n_316)
);

BUFx2_ASAP7_75t_L g331 ( 
.A(n_316),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_L g317 ( 
.A1(n_294),
.A2(n_286),
.B(n_273),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_317),
.B(n_320),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_272),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_318),
.B(n_319),
.C(n_300),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_263),
.B(n_246),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_L g321 ( 
.A1(n_279),
.A2(n_271),
.B(n_244),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_321),
.B(n_322),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_L g322 ( 
.A1(n_282),
.A2(n_279),
.B(n_275),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_310),
.B(n_313),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_326),
.B(n_327),
.C(n_329),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_300),
.B(n_319),
.C(n_301),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_300),
.B(n_319),
.C(n_306),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_332),
.B(n_333),
.C(n_339),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_303),
.B(n_320),
.C(n_317),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_303),
.B(n_311),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_322),
.B(n_298),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_342),
.B(n_343),
.C(n_297),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_308),
.B(n_302),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_340),
.A2(n_296),
.B1(n_321),
.B2(n_307),
.Y(n_344)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_344),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_328),
.B(n_296),
.Y(n_345)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_345),
.Y(n_366)
);

MAJx2_ASAP7_75t_L g346 ( 
.A(n_329),
.B(n_321),
.C(n_316),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_334),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_347),
.B(n_350),
.Y(n_360)
);

AND2x2_ASAP7_75t_L g348 ( 
.A(n_325),
.B(n_314),
.Y(n_348)
);

AOI21xp5_ASAP7_75t_L g363 ( 
.A1(n_348),
.A2(n_356),
.B(n_359),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_338),
.A2(n_316),
.B1(n_305),
.B2(n_317),
.Y(n_349)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_349),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_341),
.A2(n_316),
.B1(n_305),
.B2(n_309),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_343),
.Y(n_351)
);

AOI21xp33_ASAP7_75t_L g367 ( 
.A1(n_351),
.A2(n_353),
.B(n_354),
.Y(n_367)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_335),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_L g354 ( 
.A1(n_337),
.A2(n_318),
.B1(n_315),
.B2(n_304),
.Y(n_354)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_336),
.Y(n_356)
);

XOR2xp5_ASAP7_75t_L g370 ( 
.A(n_357),
.B(n_330),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_324),
.A2(n_299),
.B1(n_312),
.B2(n_331),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_358),
.B(n_323),
.Y(n_364)
);

OAI21xp5_ASAP7_75t_L g359 ( 
.A1(n_331),
.A2(n_342),
.B(n_325),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_352),
.B(n_327),
.C(n_332),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_361),
.B(n_365),
.C(n_369),
.Y(n_371)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_364),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_352),
.B(n_333),
.C(n_323),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_355),
.B(n_357),
.C(n_351),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_370),
.B(n_359),
.C(n_344),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_364),
.B(n_355),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_372),
.B(n_373),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_360),
.B(n_358),
.Y(n_373)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_374),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_365),
.B(n_350),
.Y(n_375)
);

INVx6_ASAP7_75t_L g381 ( 
.A(n_375),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_366),
.B(n_356),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_376),
.A2(n_345),
.B1(n_360),
.B2(n_347),
.Y(n_378)
);

XOR2xp5_ASAP7_75t_L g384 ( 
.A(n_378),
.B(n_363),
.Y(n_384)
);

OR2x2_ASAP7_75t_L g382 ( 
.A(n_379),
.B(n_377),
.Y(n_382)
);

AO221x1_ASAP7_75t_L g386 ( 
.A1(n_382),
.A2(n_384),
.B1(n_367),
.B2(n_363),
.C(n_346),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_378),
.B(n_353),
.Y(n_383)
);

INVxp67_ASAP7_75t_L g385 ( 
.A(n_383),
.Y(n_385)
);

AOI21xp5_ASAP7_75t_L g387 ( 
.A1(n_386),
.A2(n_379),
.B(n_383),
.Y(n_387)
);

OAI21xp5_ASAP7_75t_SL g388 ( 
.A1(n_387),
.A2(n_385),
.B(n_380),
.Y(n_388)
);

AOI321xp33_ASAP7_75t_L g389 ( 
.A1(n_388),
.A2(n_381),
.A3(n_371),
.B1(n_362),
.B2(n_368),
.C(n_361),
.Y(n_389)
);

BUFx24_ASAP7_75t_SL g390 ( 
.A(n_389),
.Y(n_390)
);

AOI21xp5_ASAP7_75t_L g391 ( 
.A1(n_390),
.A2(n_381),
.B(n_370),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_391),
.B(n_371),
.Y(n_392)
);


endmodule